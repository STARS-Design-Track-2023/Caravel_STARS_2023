magic
tech sky130A
magscale 1 2
timestamp 1693187644
<< viali >>
rect 1501 39049 1535 39083
rect 4905 39049 4939 39083
rect 9321 39049 9355 39083
rect 11621 39049 11655 39083
rect 13185 39049 13219 39083
rect 17785 39049 17819 39083
rect 22109 39049 22143 39083
rect 27169 39049 27203 39083
rect 33149 39049 33183 39083
rect 35725 39049 35759 39083
rect 11897 38981 11931 39015
rect 15761 38981 15795 39015
rect 31217 38981 31251 39015
rect 1777 38913 1811 38947
rect 5089 38913 5123 38947
rect 9229 38913 9263 38947
rect 12081 38913 12115 38947
rect 13001 38913 13035 38947
rect 17969 38913 18003 38947
rect 19441 38913 19475 38947
rect 20085 38913 20119 38947
rect 22385 38913 22419 38947
rect 27077 38913 27111 38947
rect 27721 38913 27755 38947
rect 33057 38913 33091 38947
rect 35633 38913 35667 38947
rect 37473 38913 37507 38947
rect 20361 38845 20395 38879
rect 15577 38777 15611 38811
rect 31033 38777 31067 38811
rect 37657 38777 37691 38811
rect 12265 38709 12299 38743
rect 19625 38709 19659 38743
rect 27629 38709 27663 38743
rect 4997 38505 5031 38539
rect 8769 38505 8803 38539
rect 18337 38505 18371 38539
rect 32229 38505 32263 38539
rect 34897 38505 34931 38539
rect 37841 38505 37875 38539
rect 19533 38369 19567 38403
rect 27261 38369 27295 38403
rect 29653 38369 29687 38403
rect 5181 38301 5215 38335
rect 8585 38301 8619 38335
rect 9045 38301 9079 38335
rect 9137 38301 9171 38335
rect 9321 38301 9355 38335
rect 13093 38301 13127 38335
rect 13277 38301 13311 38335
rect 13369 38301 13403 38335
rect 18521 38301 18555 38335
rect 18889 38301 18923 38335
rect 18981 38301 19015 38335
rect 19257 38301 19291 38335
rect 21281 38301 21315 38335
rect 21557 38301 21591 38335
rect 21649 38301 21683 38335
rect 21833 38301 21867 38335
rect 25053 38301 25087 38335
rect 25145 38301 25179 38335
rect 25329 38301 25363 38335
rect 29561 38301 29595 38335
rect 32045 38301 32079 38335
rect 34713 38301 34747 38335
rect 9597 38233 9631 38267
rect 12817 38233 12851 38267
rect 22109 38233 22143 38267
rect 25605 38233 25639 38267
rect 27537 38233 27571 38267
rect 29285 38233 29319 38267
rect 37565 38233 37599 38267
rect 11069 38165 11103 38199
rect 11345 38165 11379 38199
rect 21005 38165 21039 38199
rect 21465 38165 21499 38199
rect 23581 38165 23615 38199
rect 27077 38165 27111 38199
rect 9781 37961 9815 37995
rect 10241 37961 10275 37995
rect 11897 37961 11931 37995
rect 12265 37961 12299 37995
rect 12357 37961 12391 37995
rect 19441 37961 19475 37995
rect 19809 37961 19843 37995
rect 22017 37961 22051 37995
rect 22385 37961 22419 37995
rect 26249 37961 26283 37995
rect 26801 37961 26835 37995
rect 28365 37961 28399 37995
rect 13921 37893 13955 37927
rect 17049 37893 17083 37927
rect 17417 37893 17451 37927
rect 23581 37893 23615 37927
rect 24409 37893 24443 37927
rect 25789 37893 25823 37927
rect 9965 37825 9999 37859
rect 10609 37825 10643 37859
rect 12541 37825 12575 37859
rect 13277 37825 13311 37859
rect 13737 37825 13771 37859
rect 13829 37825 13863 37859
rect 14059 37825 14093 37859
rect 14376 37825 14410 37859
rect 14473 37825 14507 37859
rect 14565 37825 14599 37859
rect 14749 37825 14783 37859
rect 15945 37825 15979 37859
rect 16129 37825 16163 37859
rect 16221 37825 16255 37859
rect 16313 37825 16347 37859
rect 16681 37825 16715 37859
rect 16865 37825 16899 37859
rect 17233 37825 17267 37859
rect 17509 37825 17543 37859
rect 17601 37825 17635 37859
rect 20361 37825 20395 37859
rect 23397 37825 23431 37859
rect 23673 37825 23707 37859
rect 23765 37825 23799 37859
rect 24041 37825 24075 37859
rect 24225 37825 24259 37859
rect 25053 37825 25087 37859
rect 25329 37825 25363 37859
rect 25513 37825 25547 37859
rect 25973 37825 26007 37859
rect 26065 37825 26099 37859
rect 26433 37825 26467 37859
rect 26617 37825 26651 37859
rect 27721 37825 27755 37859
rect 28181 37825 28215 37859
rect 28825 37825 28859 37859
rect 29101 37825 29135 37859
rect 31217 37825 31251 37859
rect 10701 37757 10735 37791
rect 10793 37757 10827 37791
rect 11713 37757 11747 37791
rect 11805 37757 11839 37791
rect 13369 37757 13403 37791
rect 14197 37757 14231 37791
rect 14657 37757 14691 37791
rect 19901 37757 19935 37791
rect 19993 37757 20027 37791
rect 20913 37757 20947 37791
rect 22477 37757 22511 37791
rect 22569 37757 22603 37791
rect 25237 37757 25271 37791
rect 25697 37757 25731 37791
rect 27537 37757 27571 37791
rect 27997 37757 28031 37791
rect 29377 37757 29411 37791
rect 30849 37757 30883 37791
rect 24869 37689 24903 37723
rect 29009 37689 29043 37723
rect 13553 37621 13587 37655
rect 16497 37621 16531 37655
rect 17785 37621 17819 37655
rect 23949 37621 23983 37655
rect 27905 37621 27939 37655
rect 31033 37621 31067 37655
rect 17785 37417 17819 37451
rect 23857 37417 23891 37451
rect 26065 37417 26099 37451
rect 27353 37417 27387 37451
rect 1685 37281 1719 37315
rect 17877 37281 17911 37315
rect 22201 37281 22235 37315
rect 22845 37281 22879 37315
rect 22937 37281 22971 37315
rect 26617 37281 26651 37315
rect 27997 37281 28031 37315
rect 30205 37281 30239 37315
rect 8309 37213 8343 37247
rect 8585 37213 8619 37247
rect 8677 37213 8711 37247
rect 8953 37213 8987 37247
rect 18061 37213 18095 37247
rect 18337 37213 18371 37247
rect 18521 37213 18555 37247
rect 18613 37213 18647 37247
rect 20177 37213 20211 37247
rect 20269 37213 20303 37247
rect 20453 37213 20487 37247
rect 22753 37213 22787 37247
rect 23305 37213 23339 37247
rect 23673 37213 23707 37247
rect 26433 37213 26467 37247
rect 27813 37213 27847 37247
rect 29653 37213 29687 37247
rect 29745 37213 29779 37247
rect 29929 37213 29963 37247
rect 32597 37213 32631 37247
rect 37657 37213 37691 37247
rect 1501 37145 1535 37179
rect 9229 37145 9263 37179
rect 17785 37145 17819 37179
rect 20729 37145 20763 37179
rect 23489 37145 23523 37179
rect 23581 37145 23615 37179
rect 8493 37077 8527 37111
rect 10701 37077 10735 37111
rect 18245 37077 18279 37111
rect 22385 37077 22419 37111
rect 26525 37077 26559 37111
rect 27721 37077 27755 37111
rect 31677 37077 31711 37111
rect 32505 37077 32539 37111
rect 37841 37077 37875 37111
rect 9321 36873 9355 36907
rect 9781 36873 9815 36907
rect 20913 36873 20947 36907
rect 28089 36873 28123 36907
rect 29193 36873 29227 36907
rect 30941 36873 30975 36907
rect 31309 36873 31343 36907
rect 8769 36805 8803 36839
rect 24041 36805 24075 36839
rect 7297 36737 7331 36771
rect 9689 36737 9723 36771
rect 21097 36737 21131 36771
rect 23857 36737 23891 36771
rect 24501 36737 24535 36771
rect 24685 36737 24719 36771
rect 24777 36737 24811 36771
rect 27721 36737 27755 36771
rect 27997 36737 28031 36771
rect 28273 36737 28307 36771
rect 29561 36737 29595 36771
rect 30849 36737 30883 36771
rect 32321 36737 32355 36771
rect 8033 36669 8067 36703
rect 9873 36669 9907 36703
rect 23673 36669 23707 36703
rect 29653 36669 29687 36703
rect 29837 36669 29871 36703
rect 30665 36669 30699 36703
rect 32597 36669 32631 36703
rect 7573 36533 7607 36567
rect 24685 36533 24719 36567
rect 24961 36533 24995 36567
rect 27629 36533 27663 36567
rect 28457 36533 28491 36567
rect 34069 36533 34103 36567
rect 14289 36329 14323 36363
rect 18061 36329 18095 36363
rect 24133 36329 24167 36363
rect 27905 36329 27939 36363
rect 32229 36329 32263 36363
rect 11805 36261 11839 36295
rect 12541 36261 12575 36295
rect 12725 36261 12759 36295
rect 16497 36261 16531 36295
rect 32597 36261 32631 36295
rect 12633 36193 12667 36227
rect 19809 36193 19843 36227
rect 28733 36193 28767 36227
rect 33149 36193 33183 36227
rect 5733 36125 5767 36159
rect 5825 36125 5859 36159
rect 6009 36125 6043 36159
rect 9505 36125 9539 36159
rect 9781 36125 9815 36159
rect 11253 36125 11287 36159
rect 11529 36125 11563 36159
rect 11621 36125 11655 36159
rect 12111 36125 12145 36159
rect 12904 36125 12938 36159
rect 13276 36125 13310 36159
rect 13369 36125 13403 36159
rect 14289 36125 14323 36159
rect 14381 36125 14415 36159
rect 14657 36125 14691 36159
rect 14749 36125 14783 36159
rect 15301 36125 15335 36159
rect 15393 36125 15427 36159
rect 15669 36125 15703 36159
rect 15761 36125 15795 36159
rect 15945 36125 15979 36159
rect 16221 36125 16255 36159
rect 16313 36125 16347 36159
rect 16773 36125 16807 36159
rect 16866 36125 16900 36159
rect 17141 36125 17175 36159
rect 17279 36125 17313 36159
rect 17509 36125 17543 36159
rect 17877 36125 17911 36159
rect 18521 36125 18555 36159
rect 18705 36125 18739 36159
rect 20213 36125 20247 36159
rect 23581 36125 23615 36159
rect 23949 36125 23983 36159
rect 25513 36125 25547 36159
rect 25881 36125 25915 36159
rect 27261 36125 27295 36159
rect 27354 36125 27388 36159
rect 27537 36125 27571 36159
rect 27767 36125 27801 36159
rect 28549 36125 28583 36159
rect 32045 36125 32079 36159
rect 33057 36125 33091 36159
rect 6285 36057 6319 36091
rect 11437 36057 11471 36091
rect 13001 36057 13035 36091
rect 13093 36057 13127 36091
rect 14565 36057 14599 36091
rect 15577 36057 15611 36091
rect 16129 36057 16163 36091
rect 17049 36057 17083 36091
rect 17693 36057 17727 36091
rect 17785 36057 17819 36091
rect 19809 36057 19843 36091
rect 19993 36057 20027 36091
rect 20085 36057 20119 36091
rect 23765 36057 23799 36091
rect 23857 36057 23891 36091
rect 25697 36057 25731 36091
rect 25789 36057 25823 36091
rect 27629 36057 27663 36091
rect 7757 35989 7791 36023
rect 9413 35989 9447 36023
rect 9597 35989 9631 36023
rect 11989 35989 12023 36023
rect 12173 35989 12207 36023
rect 15301 35989 15335 36023
rect 17417 35989 17451 36023
rect 18613 35989 18647 36023
rect 26065 35989 26099 36023
rect 32965 35989 32999 36023
rect 6561 35785 6595 35819
rect 7665 35785 7699 35819
rect 13645 35785 13679 35819
rect 13921 35785 13955 35819
rect 29193 35785 29227 35819
rect 30757 35785 30791 35819
rect 9505 35717 9539 35751
rect 13277 35717 13311 35751
rect 14013 35717 14047 35751
rect 19074 35717 19108 35751
rect 19211 35717 19245 35751
rect 20821 35717 20855 35751
rect 25053 35717 25087 35751
rect 6745 35649 6779 35683
rect 7757 35649 7791 35683
rect 9137 35649 9171 35683
rect 13093 35649 13127 35683
rect 13553 35649 13587 35683
rect 13737 35649 13771 35683
rect 14841 35649 14875 35683
rect 18889 35649 18923 35683
rect 18981 35649 19015 35683
rect 21005 35649 21039 35683
rect 21097 35649 21131 35683
rect 21189 35649 21223 35683
rect 21373 35649 21407 35683
rect 21925 35649 21959 35683
rect 22073 35649 22107 35683
rect 22201 35649 22235 35683
rect 22293 35649 22327 35683
rect 22390 35649 22424 35683
rect 22845 35649 22879 35683
rect 22993 35649 23027 35683
rect 23121 35649 23155 35683
rect 23213 35649 23247 35683
rect 23310 35649 23344 35683
rect 23765 35649 23799 35683
rect 23857 35649 23891 35683
rect 23949 35649 23983 35683
rect 24133 35649 24167 35683
rect 24869 35649 24903 35683
rect 25145 35649 25179 35683
rect 25237 35649 25271 35683
rect 25697 35649 25731 35683
rect 25789 35649 25823 35683
rect 25973 35649 26007 35683
rect 26065 35649 26099 35683
rect 26157 35649 26191 35683
rect 26249 35649 26283 35683
rect 26433 35649 26467 35683
rect 26525 35649 26559 35683
rect 29653 35649 29687 35683
rect 29746 35649 29780 35683
rect 29929 35649 29963 35683
rect 30021 35649 30055 35683
rect 30159 35649 30193 35683
rect 30573 35649 30607 35683
rect 30849 35649 30883 35683
rect 31401 35649 31435 35683
rect 32965 35649 32999 35683
rect 33517 35649 33551 35683
rect 7849 35581 7883 35615
rect 8309 35581 8343 35615
rect 9229 35581 9263 35615
rect 12909 35581 12943 35615
rect 19349 35581 19383 35615
rect 25513 35581 25547 35615
rect 27445 35581 27479 35615
rect 27721 35581 27755 35615
rect 7297 35513 7331 35547
rect 13369 35513 13403 35547
rect 22569 35513 22603 35547
rect 30297 35513 30331 35547
rect 10977 35445 11011 35479
rect 18705 35445 18739 35479
rect 23489 35445 23523 35479
rect 23581 35445 23615 35479
rect 25421 35445 25455 35479
rect 26709 35445 26743 35479
rect 30389 35445 30423 35479
rect 31217 35445 31251 35479
rect 32873 35445 32907 35479
rect 33333 35445 33367 35479
rect 9505 35241 9539 35275
rect 17509 35241 17543 35275
rect 28181 35173 28215 35207
rect 10149 35105 10183 35139
rect 23581 35105 23615 35139
rect 23673 35105 23707 35139
rect 27537 35105 27571 35139
rect 30941 35105 30975 35139
rect 32689 35105 32723 35139
rect 32965 35105 32999 35139
rect 6653 35037 6687 35071
rect 6745 35037 6779 35071
rect 6929 35037 6963 35071
rect 9965 35037 9999 35071
rect 17325 35037 17359 35071
rect 23305 35037 23339 35071
rect 23489 35037 23523 35071
rect 23765 35037 23799 35071
rect 25329 35037 25363 35071
rect 25513 35037 25547 35071
rect 25605 35037 25639 35071
rect 25697 35037 25731 35071
rect 26341 35037 26375 35071
rect 26433 35037 26467 35071
rect 26525 35037 26559 35071
rect 26709 35037 26743 35071
rect 28365 35037 28399 35071
rect 28917 35037 28951 35071
rect 30389 35037 30423 35071
rect 30481 35037 30515 35071
rect 30665 35037 30699 35071
rect 7205 34969 7239 35003
rect 9873 34969 9907 35003
rect 26065 34969 26099 35003
rect 27721 34969 27755 35003
rect 8677 34901 8711 34935
rect 23949 34901 23983 34935
rect 25973 34901 26007 34935
rect 27629 34901 27663 34935
rect 28089 34901 28123 34935
rect 28825 34901 28859 34935
rect 32413 34901 32447 34935
rect 34437 34901 34471 34935
rect 7665 34697 7699 34731
rect 7941 34697 7975 34731
rect 16865 34697 16899 34731
rect 31217 34697 31251 34731
rect 33333 34697 33367 34731
rect 33701 34697 33735 34731
rect 11897 34629 11931 34663
rect 21005 34629 21039 34663
rect 21221 34629 21255 34663
rect 22293 34629 22327 34663
rect 23673 34629 23707 34663
rect 31677 34629 31711 34663
rect 5641 34561 5675 34595
rect 7849 34561 7883 34595
rect 8309 34561 8343 34595
rect 8401 34561 8435 34595
rect 11667 34561 11701 34595
rect 11805 34561 11839 34595
rect 12080 34561 12114 34595
rect 12173 34561 12207 34595
rect 17141 34561 17175 34595
rect 17325 34561 17359 34595
rect 21925 34561 21959 34595
rect 22073 34561 22107 34595
rect 22201 34561 22235 34595
rect 22390 34561 22424 34595
rect 23397 34561 23431 34595
rect 23581 34561 23615 34595
rect 23765 34561 23799 34595
rect 28641 34561 28675 34595
rect 31585 34561 31619 34595
rect 33241 34561 33275 34595
rect 37565 34561 37599 34595
rect 8585 34493 8619 34527
rect 31861 34493 31895 34527
rect 33149 34493 33183 34527
rect 37841 34493 37875 34527
rect 21373 34425 21407 34459
rect 5457 34357 5491 34391
rect 11529 34357 11563 34391
rect 16865 34357 16899 34391
rect 16957 34357 16991 34391
rect 17049 34357 17083 34391
rect 21189 34357 21223 34391
rect 22569 34357 22603 34391
rect 23949 34357 23983 34391
rect 28898 34357 28932 34391
rect 30389 34357 30423 34391
rect 6745 34153 6779 34187
rect 14657 34153 14691 34187
rect 14841 34153 14875 34187
rect 16681 34153 16715 34187
rect 28089 34153 28123 34187
rect 11621 34085 11655 34119
rect 15945 34085 15979 34119
rect 17417 34085 17451 34119
rect 19441 34085 19475 34119
rect 19901 34085 19935 34119
rect 26065 34085 26099 34119
rect 28457 34085 28491 34119
rect 31125 34085 31159 34119
rect 34069 34085 34103 34119
rect 5273 34017 5307 34051
rect 13185 34017 13219 34051
rect 13737 34017 13771 34051
rect 14749 34017 14783 34051
rect 15117 34017 15151 34051
rect 16865 34017 16899 34051
rect 19257 34017 19291 34051
rect 29009 34017 29043 34051
rect 34989 34017 35023 34051
rect 4721 33949 4755 33983
rect 4813 33949 4847 33983
rect 4997 33949 5031 33983
rect 7297 33949 7331 33983
rect 8585 33949 8619 33983
rect 9505 33949 9539 33983
rect 9873 33949 9907 33983
rect 11621 33949 11655 33983
rect 11897 33949 11931 33983
rect 14381 33949 14415 33983
rect 14565 33949 14599 33983
rect 15761 33949 15795 33983
rect 16037 33949 16071 33983
rect 16221 33949 16255 33983
rect 16313 33949 16347 33983
rect 16405 33949 16439 33983
rect 17693 33949 17727 33983
rect 17786 33949 17820 33983
rect 18061 33949 18095 33983
rect 18158 33949 18192 33983
rect 18429 33949 18463 33983
rect 18797 33949 18831 33983
rect 19533 33949 19567 33983
rect 20085 33949 20119 33983
rect 20269 33949 20303 33983
rect 20453 33949 20487 33983
rect 20821 33949 20855 33983
rect 21925 33949 21959 33983
rect 22569 33949 22603 33983
rect 22661 33949 22695 33983
rect 22845 33949 22879 33983
rect 22937 33949 22971 33983
rect 23213 33949 23247 33983
rect 23306 33949 23340 33983
rect 23581 33949 23615 33983
rect 23678 33949 23712 33983
rect 25605 33949 25639 33983
rect 25697 33949 25731 33983
rect 25881 33949 25915 33983
rect 25973 33949 26007 33983
rect 26249 33949 26283 33983
rect 26341 33949 26375 33983
rect 26433 33949 26467 33983
rect 26617 33949 26651 33983
rect 27261 33949 27295 33983
rect 27905 33949 27939 33983
rect 28917 33949 28951 33983
rect 30481 33949 30515 33983
rect 30601 33949 30635 33983
rect 30946 33949 30980 33983
rect 31493 33949 31527 33983
rect 31769 33949 31803 33983
rect 33885 33949 33919 33983
rect 34345 33949 34379 33983
rect 34437 33949 34471 33983
rect 34713 33949 34747 33983
rect 13461 33881 13495 33915
rect 15393 33881 15427 33915
rect 15577 33881 15611 33915
rect 17233 33881 17267 33915
rect 17969 33881 18003 33915
rect 18613 33881 18647 33915
rect 18705 33881 18739 33915
rect 20177 33881 20211 33915
rect 23489 33881 23523 33915
rect 30757 33881 30791 33915
rect 30849 33881 30883 33915
rect 36737 33881 36771 33915
rect 7205 33813 7239 33847
rect 8677 33813 8711 33847
rect 8953 33813 8987 33847
rect 9689 33813 9723 33847
rect 11805 33813 11839 33847
rect 13369 33813 13403 33847
rect 13553 33813 13587 33847
rect 15669 33813 15703 33847
rect 17049 33813 17083 33847
rect 17141 33813 17175 33847
rect 18337 33813 18371 33847
rect 18981 33813 19015 33847
rect 19533 33813 19567 33847
rect 21833 33813 21867 33847
rect 23121 33813 23155 33847
rect 23857 33813 23891 33847
rect 25421 33813 25455 33847
rect 27169 33813 27203 33847
rect 28825 33813 28859 33847
rect 31585 33813 31619 33847
rect 31953 33813 31987 33847
rect 5457 33609 5491 33643
rect 5825 33609 5859 33643
rect 14289 33609 14323 33643
rect 14565 33609 14599 33643
rect 17433 33609 17467 33643
rect 17601 33609 17635 33643
rect 21097 33609 21131 33643
rect 21281 33609 21315 33643
rect 33333 33609 33367 33643
rect 33793 33609 33827 33643
rect 34161 33609 34195 33643
rect 34621 33609 34655 33643
rect 36921 33609 36955 33643
rect 9229 33541 9263 33575
rect 14197 33541 14231 33575
rect 17233 33541 17267 33575
rect 20821 33541 20855 33575
rect 21465 33541 21499 33575
rect 25237 33541 25271 33575
rect 34253 33541 34287 33575
rect 7021 33473 7055 33507
rect 8953 33473 8987 33507
rect 14013 33473 14047 33507
rect 14381 33473 14415 33507
rect 19708 33473 19742 33507
rect 19901 33473 19935 33507
rect 20269 33473 20303 33507
rect 20361 33473 20395 33507
rect 20637 33473 20671 33507
rect 20729 33473 20763 33507
rect 20913 33473 20947 33507
rect 21833 33473 21867 33507
rect 22017 33473 22051 33507
rect 23765 33473 23799 33507
rect 23857 33473 23891 33507
rect 26617 33473 26651 33507
rect 26985 33473 27019 33507
rect 33425 33473 33459 33507
rect 34713 33473 34747 33507
rect 36737 33473 36771 33507
rect 5917 33405 5951 33439
rect 6101 33405 6135 33439
rect 7297 33405 7331 33439
rect 8769 33405 8803 33439
rect 19073 33405 19107 33439
rect 23489 33405 23523 33439
rect 23581 33405 23615 33439
rect 27261 33405 27295 33439
rect 29009 33405 29043 33439
rect 33241 33405 33275 33439
rect 34069 33405 34103 33439
rect 21833 33337 21867 33371
rect 24869 33337 24903 33371
rect 26801 33337 26835 33371
rect 10701 33269 10735 33303
rect 17417 33269 17451 33303
rect 21281 33269 21315 33303
rect 24041 33269 24075 33303
rect 25237 33269 25271 33303
rect 25421 33269 25455 33303
rect 34897 33269 34931 33303
rect 7665 33065 7699 33099
rect 10149 33065 10183 33099
rect 18613 33065 18647 33099
rect 26617 33065 26651 33099
rect 19717 32997 19751 33031
rect 19809 32997 19843 33031
rect 20729 32997 20763 33031
rect 6101 32929 6135 32963
rect 6745 32929 6779 32963
rect 6837 32929 6871 32963
rect 8125 32929 8159 32963
rect 8401 32929 8435 32963
rect 9597 32929 9631 32963
rect 16957 32929 16991 32963
rect 19625 32929 19659 32963
rect 27261 32929 27295 32963
rect 34989 32929 35023 32963
rect 4077 32861 4111 32895
rect 4169 32861 4203 32895
rect 4353 32861 4387 32895
rect 6653 32861 6687 32895
rect 7849 32861 7883 32895
rect 7941 32861 7975 32895
rect 8217 32861 8251 32895
rect 8493 32861 8527 32895
rect 9781 32861 9815 32895
rect 11713 32861 11747 32895
rect 11806 32861 11840 32895
rect 11989 32861 12023 32895
rect 12178 32861 12212 32895
rect 16221 32861 16255 32895
rect 17325 32861 17359 32895
rect 18337 32861 18371 32895
rect 18429 32861 18463 32895
rect 18705 32861 18739 32895
rect 19901 32861 19935 32895
rect 20177 32861 20211 32895
rect 20453 32861 20487 32895
rect 20545 32861 20579 32895
rect 21465 32861 21499 32895
rect 22109 32861 22143 32895
rect 23397 32861 23431 32895
rect 27537 32861 27571 32895
rect 30389 32861 30423 32895
rect 30941 32861 30975 32895
rect 31217 32861 31251 32895
rect 34345 32861 34379 32895
rect 34437 32861 34471 32895
rect 34713 32861 34747 32895
rect 4629 32793 4663 32827
rect 12081 32793 12115 32827
rect 18797 32793 18831 32827
rect 20361 32793 20395 32827
rect 23213 32793 23247 32827
rect 27813 32793 27847 32827
rect 31493 32793 31527 32827
rect 36737 32793 36771 32827
rect 6285 32725 6319 32759
rect 9689 32725 9723 32759
rect 12357 32725 12391 32759
rect 21005 32725 21039 32759
rect 23581 32725 23615 32759
rect 26985 32725 27019 32759
rect 27077 32725 27111 32759
rect 29285 32725 29319 32759
rect 30205 32725 30239 32759
rect 31125 32725 31159 32759
rect 32965 32725 32999 32759
rect 4997 32521 5031 32555
rect 12081 32521 12115 32555
rect 17693 32521 17727 32555
rect 19993 32521 20027 32555
rect 27813 32521 27847 32555
rect 29009 32521 29043 32555
rect 31401 32521 31435 32555
rect 36001 32521 36035 32555
rect 11713 32453 11747 32487
rect 12265 32453 12299 32487
rect 12449 32453 12483 32487
rect 16681 32453 16715 32487
rect 16865 32453 16899 32487
rect 17325 32453 17359 32487
rect 17509 32453 17543 32487
rect 23121 32453 23155 32487
rect 23213 32453 23247 32487
rect 5181 32385 5215 32419
rect 11529 32385 11563 32419
rect 11805 32385 11839 32419
rect 11897 32385 11931 32419
rect 18429 32385 18463 32419
rect 18613 32385 18647 32419
rect 18705 32385 18739 32419
rect 18889 32385 18923 32419
rect 18981 32385 19015 32419
rect 21281 32385 21315 32419
rect 21925 32385 21959 32419
rect 23029 32385 23063 32419
rect 23397 32385 23431 32419
rect 23765 32385 23799 32419
rect 23903 32385 23937 32419
rect 24041 32385 24075 32419
rect 24133 32385 24167 32419
rect 27905 32385 27939 32419
rect 28549 32385 28583 32419
rect 29193 32385 29227 32419
rect 30849 32385 30883 32419
rect 31493 32385 31527 32419
rect 32413 32385 32447 32419
rect 33149 32385 33183 32419
rect 33425 32385 33459 32419
rect 35633 32385 35667 32419
rect 35817 32385 35851 32419
rect 28273 32317 28307 32351
rect 28457 32317 28491 32351
rect 30665 32317 30699 32351
rect 30757 32317 30791 32351
rect 32689 32317 32723 32351
rect 12633 32249 12667 32283
rect 17049 32249 17083 32283
rect 28917 32249 28951 32283
rect 31217 32249 31251 32283
rect 32137 32249 32171 32283
rect 16865 32181 16899 32215
rect 17475 32181 17509 32215
rect 22201 32181 22235 32215
rect 22845 32181 22879 32215
rect 24317 32181 24351 32215
rect 19073 31977 19107 32011
rect 18705 31909 18739 31943
rect 19993 31909 20027 31943
rect 24961 31909 24995 31943
rect 25329 31909 25363 31943
rect 26801 31909 26835 31943
rect 7205 31841 7239 31875
rect 3985 31773 4019 31807
rect 4077 31773 4111 31807
rect 4261 31773 4295 31807
rect 6285 31773 6319 31807
rect 6561 31773 6595 31807
rect 7481 31773 7515 31807
rect 7573 31773 7607 31807
rect 7665 31773 7699 31807
rect 7849 31773 7883 31807
rect 8125 31773 8159 31807
rect 8493 31773 8527 31807
rect 9229 31773 9263 31807
rect 9321 31773 9355 31807
rect 9505 31773 9539 31807
rect 13645 31773 13679 31807
rect 18889 31773 18923 31807
rect 19073 31773 19107 31807
rect 21281 31773 21315 31807
rect 21925 31773 21959 31807
rect 22018 31773 22052 31807
rect 22201 31773 22235 31807
rect 22293 31773 22327 31807
rect 22390 31773 22424 31807
rect 22661 31773 22695 31807
rect 22809 31773 22843 31807
rect 23167 31773 23201 31807
rect 23397 31773 23431 31807
rect 23490 31773 23524 31807
rect 23903 31773 23937 31807
rect 24409 31773 24443 31807
rect 24777 31773 24811 31807
rect 25145 31773 25179 31807
rect 25237 31773 25271 31807
rect 25421 31773 25455 31807
rect 26157 31773 26191 31807
rect 26249 31773 26283 31807
rect 26525 31773 26559 31807
rect 26985 31773 27019 31807
rect 27997 31773 28031 31807
rect 28273 31773 28307 31807
rect 29561 31773 29595 31807
rect 29699 31773 29733 31807
rect 29837 31773 29871 31807
rect 29929 31773 29963 31807
rect 30067 31773 30101 31807
rect 30481 31773 30515 31807
rect 31493 31773 31527 31807
rect 31769 31773 31803 31807
rect 31953 31773 31987 31807
rect 34897 31773 34931 31807
rect 34989 31773 35023 31807
rect 35449 31773 35483 31807
rect 4537 31705 4571 31739
rect 9781 31705 9815 31739
rect 13093 31705 13127 31739
rect 13369 31705 13403 31739
rect 22937 31705 22971 31739
rect 23029 31705 23063 31739
rect 23673 31705 23707 31739
rect 23765 31705 23799 31739
rect 24593 31705 24627 31739
rect 24685 31705 24719 31739
rect 26341 31705 26375 31739
rect 31585 31705 31619 31739
rect 35081 31705 35115 31739
rect 7297 31637 7331 31671
rect 8033 31637 8067 31671
rect 8309 31637 8343 31671
rect 11253 31637 11287 31671
rect 13277 31637 13311 31671
rect 13461 31637 13495 31671
rect 22569 31637 22603 31671
rect 23305 31637 23339 31671
rect 24041 31637 24075 31671
rect 25605 31637 25639 31671
rect 25973 31637 26007 31671
rect 27905 31637 27939 31671
rect 28089 31637 28123 31671
rect 30205 31637 30239 31671
rect 30389 31637 30423 31671
rect 34805 31637 34839 31671
rect 35265 31637 35299 31671
rect 9873 31433 9907 31467
rect 10149 31433 10183 31467
rect 10609 31433 10643 31467
rect 13461 31433 13495 31467
rect 18705 31433 18739 31467
rect 19901 31433 19935 31467
rect 21005 31433 21039 31467
rect 22109 31433 22143 31467
rect 22201 31433 22235 31467
rect 22385 31433 22419 31467
rect 8125 31365 8159 31399
rect 11805 31365 11839 31399
rect 14749 31365 14783 31399
rect 16957 31365 16991 31399
rect 21833 31365 21867 31399
rect 23397 31365 23431 31399
rect 25145 31365 25179 31399
rect 27997 31365 28031 31399
rect 10057 31297 10091 31331
rect 10517 31297 10551 31331
rect 11529 31297 11563 31331
rect 11713 31297 11747 31331
rect 11897 31297 11931 31331
rect 15485 31297 15519 31331
rect 15669 31297 15703 31331
rect 15945 31297 15979 31331
rect 16129 31297 16163 31331
rect 16221 31297 16255 31331
rect 16313 31297 16347 31331
rect 16681 31297 16715 31331
rect 16774 31297 16808 31331
rect 17049 31297 17083 31331
rect 17187 31297 17221 31331
rect 17417 31297 17451 31331
rect 17601 31297 17635 31331
rect 17693 31297 17727 31331
rect 17785 31297 17819 31331
rect 18521 31297 18555 31331
rect 18797 31297 18831 31331
rect 19441 31297 19475 31331
rect 19717 31297 19751 31331
rect 20545 31297 20579 31331
rect 20637 31297 20671 31331
rect 20821 31297 20855 31331
rect 20913 31297 20947 31331
rect 21189 31297 21223 31331
rect 21281 31297 21315 31331
rect 22017 31297 22051 31331
rect 22845 31297 22879 31331
rect 23029 31297 23063 31331
rect 23305 31297 23339 31331
rect 25421 31297 25455 31331
rect 25605 31297 25639 31331
rect 25973 31297 26007 31331
rect 26341 31297 26375 31331
rect 26985 31297 27019 31331
rect 27169 31297 27203 31331
rect 27261 31297 27295 31331
rect 27353 31297 27387 31331
rect 29653 31297 29687 31331
rect 29929 31297 29963 31331
rect 32413 31297 32447 31331
rect 34437 31297 34471 31331
rect 34529 31297 34563 31331
rect 7849 31229 7883 31263
rect 9597 31229 9631 31263
rect 10793 31229 10827 31263
rect 15393 31229 15427 31263
rect 15853 31229 15887 31263
rect 21373 31229 21407 31263
rect 21465 31229 21499 31263
rect 22937 31229 22971 31263
rect 23121 31229 23155 31263
rect 27721 31229 27755 31263
rect 30205 31229 30239 31263
rect 31953 31229 31987 31263
rect 34161 31229 34195 31263
rect 34805 31229 34839 31263
rect 36553 31229 36587 31263
rect 17325 31161 17359 31195
rect 26709 31161 26743 31195
rect 29837 31161 29871 31195
rect 12081 31093 12115 31127
rect 16497 31093 16531 31127
rect 17969 31093 18003 31127
rect 18337 31093 18371 31127
rect 20361 31093 20395 31127
rect 22661 31093 22695 31127
rect 27629 31093 27663 31127
rect 29469 31093 29503 31127
rect 7849 30889 7883 30923
rect 8953 30889 8987 30923
rect 14473 30889 14507 30923
rect 16497 30889 16531 30923
rect 19349 30889 19383 30923
rect 21281 30889 21315 30923
rect 24501 30889 24535 30923
rect 24869 30889 24903 30923
rect 26617 30889 26651 30923
rect 28089 30889 28123 30923
rect 30113 30889 30147 30923
rect 34069 30889 34103 30923
rect 35449 30889 35483 30923
rect 20729 30821 20763 30855
rect 33793 30821 33827 30855
rect 8401 30753 8435 30787
rect 9413 30753 9447 30787
rect 9505 30753 9539 30787
rect 13369 30753 13403 30787
rect 13921 30753 13955 30787
rect 14565 30753 14599 30787
rect 21741 30753 21775 30787
rect 24593 30753 24627 30787
rect 28641 30753 28675 30787
rect 30757 30753 30791 30787
rect 33149 30753 33183 30787
rect 34805 30753 34839 30787
rect 4537 30685 4571 30719
rect 5641 30685 5675 30719
rect 5733 30685 5767 30719
rect 5917 30685 5951 30719
rect 14381 30685 14415 30719
rect 14657 30685 14691 30719
rect 14841 30685 14875 30719
rect 16313 30685 16347 30719
rect 16589 30685 16623 30719
rect 16682 30685 16716 30719
rect 16865 30685 16899 30719
rect 17095 30685 17129 30719
rect 19349 30685 19383 30719
rect 20361 30685 20395 30719
rect 21373 30685 21407 30719
rect 24501 30685 24535 30719
rect 26065 30685 26099 30719
rect 26157 30685 26191 30719
rect 26341 30685 26375 30719
rect 26433 30685 26467 30719
rect 30481 30685 30515 30719
rect 33425 30685 33459 30719
rect 33885 30685 33919 30719
rect 6193 30617 6227 30651
rect 8217 30617 8251 30651
rect 13737 30617 13771 30651
rect 16129 30617 16163 30651
rect 16957 30617 16991 30651
rect 19073 30617 19107 30651
rect 21557 30617 21591 30651
rect 28549 30617 28583 30651
rect 30941 30617 30975 30651
rect 34989 30617 35023 30651
rect 4445 30549 4479 30583
rect 7665 30549 7699 30583
rect 8309 30549 8343 30583
rect 9321 30549 9355 30583
rect 13553 30549 13587 30583
rect 13645 30549 13679 30583
rect 14105 30549 14139 30583
rect 17233 30549 17267 30583
rect 17785 30549 17819 30583
rect 20913 30549 20947 30583
rect 21005 30549 21039 30583
rect 21097 30549 21131 30583
rect 28457 30549 28491 30583
rect 30573 30549 30607 30583
rect 32229 30549 32263 30583
rect 33333 30549 33367 30583
rect 35081 30549 35115 30583
rect 6009 30345 6043 30379
rect 6469 30345 6503 30379
rect 7389 30277 7423 30311
rect 13001 30277 13035 30311
rect 19901 30277 19935 30311
rect 20085 30277 20119 30311
rect 20453 30277 20487 30311
rect 20637 30277 20671 30311
rect 25881 30277 25915 30311
rect 6653 30209 6687 30243
rect 7665 30209 7699 30243
rect 7757 30209 7791 30243
rect 7849 30209 7883 30243
rect 8033 30209 8067 30243
rect 8585 30209 8619 30243
rect 11621 30209 11655 30243
rect 11714 30209 11748 30243
rect 11897 30209 11931 30243
rect 11989 30209 12023 30243
rect 12127 30209 12161 30243
rect 14749 30209 14783 30243
rect 17693 30209 17727 30243
rect 18429 30209 18463 30243
rect 18521 30209 18555 30243
rect 18613 30209 18647 30243
rect 18797 30209 18831 30243
rect 23397 30209 23431 30243
rect 25697 30209 25731 30243
rect 25969 30209 26003 30243
rect 26065 30209 26099 30243
rect 30389 30209 30423 30243
rect 32137 30209 32171 30243
rect 32321 30209 32355 30243
rect 32413 30209 32447 30243
rect 32505 30209 32539 30243
rect 4261 30141 4295 30175
rect 4537 30141 4571 30175
rect 6745 30141 6779 30175
rect 17785 30141 17819 30175
rect 25145 30141 25179 30175
rect 7481 30073 7515 30107
rect 20269 30073 20303 30107
rect 29101 30073 29135 30107
rect 8677 30005 8711 30039
rect 12265 30005 12299 30039
rect 17785 30005 17819 30039
rect 18061 30005 18095 30039
rect 18153 30005 18187 30039
rect 20085 30005 20119 30039
rect 20637 30005 20671 30039
rect 20821 30005 20855 30039
rect 26249 30005 26283 30039
rect 32781 30005 32815 30039
rect 15761 29801 15795 29835
rect 16681 29801 16715 29835
rect 24593 29801 24627 29835
rect 8493 29733 8527 29767
rect 13737 29733 13771 29767
rect 14105 29733 14139 29767
rect 14381 29733 14415 29767
rect 15117 29733 15151 29767
rect 6101 29665 6135 29699
rect 9229 29665 9263 29699
rect 14473 29665 14507 29699
rect 27629 29665 27663 29699
rect 33977 29665 34011 29699
rect 36829 29665 36863 29699
rect 4169 29597 4203 29631
rect 8309 29597 8343 29631
rect 8585 29597 8619 29631
rect 8677 29597 8711 29631
rect 8953 29597 8987 29631
rect 12541 29597 12575 29631
rect 12725 29597 12759 29631
rect 12909 29597 12943 29631
rect 13461 29597 13495 29631
rect 13553 29597 13587 29631
rect 13829 29597 13863 29631
rect 14289 29597 14323 29631
rect 14565 29597 14599 29631
rect 14749 29597 14783 29631
rect 15301 29597 15335 29631
rect 15393 29597 15427 29631
rect 15485 29597 15519 29631
rect 15669 29597 15703 29631
rect 15945 29597 15979 29631
rect 16045 29597 16079 29631
rect 16313 29597 16347 29631
rect 16865 29597 16899 29631
rect 18245 29597 18279 29631
rect 18337 29597 18371 29631
rect 18613 29597 18647 29631
rect 18705 29597 18739 29631
rect 20637 29597 20671 29631
rect 20913 29597 20947 29631
rect 22891 29597 22925 29631
rect 23304 29597 23338 29631
rect 23397 29597 23431 29631
rect 23765 29597 23799 29631
rect 24041 29597 24075 29631
rect 24685 29597 24719 29631
rect 24777 29597 24811 29631
rect 25769 29597 25803 29631
rect 25881 29597 25915 29631
rect 25973 29597 26007 29631
rect 26157 29597 26191 29631
rect 26433 29597 26467 29631
rect 26525 29597 26559 29631
rect 26709 29597 26743 29631
rect 26801 29597 26835 29631
rect 27445 29597 27479 29631
rect 27813 29597 27847 29631
rect 28549 29597 28583 29631
rect 29377 29597 29411 29631
rect 29837 29597 29871 29631
rect 29929 29597 29963 29631
rect 30021 29597 30055 29631
rect 30205 29597 30239 29631
rect 30297 29597 30331 29631
rect 30390 29597 30424 29631
rect 30665 29597 30699 29631
rect 30803 29597 30837 29631
rect 31217 29597 31251 29631
rect 34161 29597 34195 29631
rect 34805 29597 34839 29631
rect 5825 29529 5859 29563
rect 16129 29529 16163 29563
rect 17233 29529 17267 29563
rect 18521 29529 18555 29563
rect 23009 29529 23043 29563
rect 23121 29529 23155 29563
rect 26249 29529 26283 29563
rect 30573 29529 30607 29563
rect 32965 29529 32999 29563
rect 35081 29529 35115 29563
rect 4077 29461 4111 29495
rect 5457 29461 5491 29495
rect 5917 29461 5951 29495
rect 10701 29461 10735 29495
rect 13277 29461 13311 29495
rect 16957 29461 16991 29495
rect 17049 29461 17083 29495
rect 18889 29461 18923 29495
rect 20821 29461 20855 29495
rect 21005 29461 21039 29495
rect 21189 29461 21223 29495
rect 22753 29461 22787 29495
rect 23581 29461 23615 29495
rect 23949 29461 23983 29495
rect 24409 29461 24443 29495
rect 25513 29461 25547 29495
rect 27353 29461 27387 29495
rect 27905 29461 27939 29495
rect 28273 29461 28307 29495
rect 28365 29461 28399 29495
rect 29285 29461 29319 29495
rect 29561 29461 29595 29495
rect 30941 29461 30975 29495
rect 34069 29461 34103 29495
rect 34529 29461 34563 29495
rect 9873 29257 9907 29291
rect 18889 29257 18923 29291
rect 21281 29257 21315 29291
rect 29009 29257 29043 29291
rect 34989 29257 35023 29291
rect 7113 29189 7147 29223
rect 9137 29189 9171 29223
rect 11345 29189 11379 29223
rect 22109 29189 22143 29223
rect 23673 29189 23707 29223
rect 23765 29189 23799 29223
rect 26065 29189 26099 29223
rect 27537 29189 27571 29223
rect 31585 29189 31619 29223
rect 3893 29121 3927 29155
rect 5917 29121 5951 29155
rect 6929 29121 6963 29155
rect 7021 29121 7055 29155
rect 7297 29121 7331 29155
rect 7665 29121 7699 29155
rect 13093 29121 13127 29155
rect 13277 29121 13311 29155
rect 18521 29121 18555 29155
rect 18705 29121 18739 29155
rect 20729 29121 20763 29155
rect 20913 29121 20947 29155
rect 21005 29121 21039 29155
rect 21097 29121 21131 29155
rect 21833 29121 21867 29155
rect 21981 29121 22015 29155
rect 22201 29121 22235 29155
rect 22298 29121 22332 29155
rect 22569 29121 22603 29155
rect 22845 29121 22879 29155
rect 23029 29121 23063 29155
rect 23489 29121 23523 29155
rect 23857 29121 23891 29155
rect 25513 29121 25547 29155
rect 25605 29121 25639 29155
rect 25789 29121 25823 29155
rect 25881 29121 25915 29155
rect 26157 29121 26191 29155
rect 26341 29121 26375 29155
rect 26433 29121 26467 29155
rect 26525 29121 26559 29155
rect 27261 29121 27295 29155
rect 29193 29121 29227 29155
rect 31496 29143 31530 29177
rect 31769 29121 31803 29155
rect 31953 29121 31987 29155
rect 32137 29121 32171 29155
rect 32321 29121 32355 29155
rect 32413 29121 32447 29155
rect 32506 29143 32540 29177
rect 33057 29121 33091 29155
rect 34621 29121 34655 29155
rect 35081 29121 35115 29155
rect 36645 29121 36679 29155
rect 36829 29121 36863 29155
rect 8217 29053 8251 29087
rect 9229 29053 9263 29087
rect 9413 29053 9447 29087
rect 22753 29053 22787 29087
rect 30941 29053 30975 29087
rect 8769 28985 8803 29019
rect 12909 28985 12943 29019
rect 22477 28985 22511 29019
rect 22937 28985 22971 29019
rect 24041 28985 24075 29019
rect 26801 28985 26835 29019
rect 32781 28985 32815 29019
rect 34805 28985 34839 29019
rect 37013 28985 37047 29019
rect 4156 28917 4190 28951
rect 6745 28917 6779 28951
rect 18613 28917 18647 28951
rect 23213 28917 23247 28951
rect 29456 28917 29490 28951
rect 32873 28917 32907 28951
rect 4537 28713 4571 28747
rect 25789 28713 25823 28747
rect 7941 28645 7975 28679
rect 29285 28645 29319 28679
rect 6009 28577 6043 28611
rect 6193 28577 6227 28611
rect 6469 28577 6503 28611
rect 30021 28577 30055 28611
rect 30205 28577 30239 28611
rect 32045 28577 32079 28611
rect 33885 28577 33919 28611
rect 34069 28577 34103 28611
rect 36461 28577 36495 28611
rect 4353 28509 4387 28543
rect 4721 28509 4755 28543
rect 6101 28509 6135 28543
rect 8309 28509 8343 28543
rect 9965 28509 9999 28543
rect 10057 28509 10091 28543
rect 10241 28509 10275 28543
rect 16129 28509 16163 28543
rect 16313 28509 16347 28543
rect 16497 28509 16531 28543
rect 19717 28509 19751 28543
rect 19809 28509 19843 28543
rect 20085 28509 20119 28543
rect 20821 28509 20855 28543
rect 22569 28509 22603 28543
rect 24593 28509 24627 28543
rect 24685 28509 24719 28543
rect 24961 28509 24995 28543
rect 25973 28509 26007 28543
rect 26065 28509 26099 28543
rect 26341 28509 26375 28543
rect 29101 28509 29135 28543
rect 30389 28509 30423 28543
rect 30482 28509 30516 28543
rect 30757 28509 30791 28543
rect 30854 28509 30888 28543
rect 31309 28509 31343 28543
rect 31569 28519 31603 28553
rect 31769 28509 31803 28543
rect 34713 28509 34747 28543
rect 10517 28441 10551 28475
rect 16405 28441 16439 28475
rect 19901 28441 19935 28475
rect 24777 28441 24811 28475
rect 26157 28441 26191 28475
rect 30665 28441 30699 28475
rect 31493 28441 31527 28475
rect 34989 28441 35023 28475
rect 4261 28373 4295 28407
rect 8217 28373 8251 28407
rect 11989 28373 12023 28407
rect 16681 28373 16715 28407
rect 19533 28373 19567 28407
rect 24409 28373 24443 28407
rect 29561 28373 29595 28407
rect 29929 28373 29963 28407
rect 31033 28373 31067 28407
rect 31125 28373 31159 28407
rect 33517 28373 33551 28407
rect 34161 28373 34195 28407
rect 34529 28373 34563 28407
rect 5825 28169 5859 28203
rect 6745 28169 6779 28203
rect 10609 28169 10643 28203
rect 11529 28169 11563 28203
rect 13737 28169 13771 28203
rect 13921 28169 13955 28203
rect 17325 28169 17359 28203
rect 23121 28169 23155 28203
rect 23857 28169 23891 28203
rect 31861 28169 31895 28203
rect 32597 28169 32631 28203
rect 32965 28169 32999 28203
rect 34437 28169 34471 28203
rect 34897 28169 34931 28203
rect 6837 28101 6871 28135
rect 11897 28101 11931 28135
rect 17049 28101 17083 28135
rect 19073 28101 19107 28135
rect 19273 28101 19307 28135
rect 21097 28101 21131 28135
rect 21189 28101 21223 28135
rect 4077 28033 4111 28067
rect 7665 28033 7699 28067
rect 9965 28033 9999 28067
rect 10793 28033 10827 28067
rect 12449 28033 12483 28067
rect 12633 28033 12667 28067
rect 12725 28033 12759 28067
rect 12817 28033 12851 28067
rect 13829 28033 13863 28067
rect 14657 28033 14691 28067
rect 14749 28033 14783 28067
rect 14933 28033 14967 28067
rect 16681 28033 16715 28067
rect 16774 28033 16808 28067
rect 16957 28033 16991 28067
rect 17187 28033 17221 28067
rect 19625 28033 19659 28067
rect 19809 28033 19843 28067
rect 19901 28033 19935 28067
rect 20545 28033 20579 28067
rect 20637 28033 20671 28067
rect 20821 28033 20855 28067
rect 20914 28033 20948 28067
rect 21327 28033 21361 28067
rect 22477 28033 22511 28067
rect 22845 28033 22879 28067
rect 23305 28033 23339 28067
rect 23397 28033 23431 28067
rect 23489 28033 23523 28067
rect 23673 28033 23707 28067
rect 23765 28033 23799 28067
rect 24133 28033 24167 28067
rect 31953 28033 31987 28067
rect 32505 28033 32539 28067
rect 34253 28033 34287 28067
rect 34989 28033 35023 28067
rect 37381 28033 37415 28067
rect 4353 27965 4387 27999
rect 7021 27965 7055 27999
rect 7941 27965 7975 27999
rect 10057 27965 10091 27999
rect 10149 27965 10183 27999
rect 11989 27965 12023 27999
rect 12081 27965 12115 27999
rect 13553 27965 13587 27999
rect 20177 27965 20211 27999
rect 20361 27965 20395 27999
rect 20453 27965 20487 27999
rect 21925 27965 21959 27999
rect 22293 27965 22327 27999
rect 22753 27965 22787 27999
rect 32413 27965 32447 27999
rect 9413 27897 9447 27931
rect 14105 27897 14139 27931
rect 14565 27897 14599 27931
rect 19441 27897 19475 27931
rect 19717 27897 19751 27931
rect 20085 27897 20119 27931
rect 21465 27897 21499 27931
rect 24041 27897 24075 27931
rect 6377 27829 6411 27863
rect 9597 27829 9631 27863
rect 13001 27829 13035 27863
rect 14197 27829 14231 27863
rect 14473 27829 14507 27863
rect 19257 27829 19291 27863
rect 24225 27829 24259 27863
rect 24501 27829 24535 27863
rect 37565 27829 37599 27863
rect 4629 27625 4663 27659
rect 8309 27625 8343 27659
rect 14657 27625 14691 27659
rect 23765 27625 23799 27659
rect 14105 27557 14139 27591
rect 16037 27557 16071 27591
rect 33793 27557 33827 27591
rect 12081 27489 12115 27523
rect 12173 27489 12207 27523
rect 13093 27489 13127 27523
rect 27537 27489 27571 27523
rect 4813 27421 4847 27455
rect 6929 27421 6963 27455
rect 8493 27421 8527 27455
rect 9505 27421 9539 27455
rect 9597 27421 9631 27455
rect 9781 27421 9815 27455
rect 13277 27421 13311 27455
rect 14473 27421 14507 27455
rect 15577 27421 15611 27455
rect 15669 27421 15703 27455
rect 15853 27421 15887 27455
rect 16681 27421 16715 27455
rect 16774 27421 16808 27455
rect 16957 27421 16991 27455
rect 17146 27421 17180 27455
rect 17417 27421 17451 27455
rect 17601 27421 17635 27455
rect 17693 27421 17727 27455
rect 17785 27421 17819 27455
rect 18153 27421 18187 27455
rect 18337 27421 18371 27455
rect 18429 27421 18463 27455
rect 18613 27421 18647 27455
rect 22937 27421 22971 27455
rect 23213 27421 23247 27455
rect 23581 27421 23615 27455
rect 25513 27421 25547 27455
rect 25605 27421 25639 27455
rect 25789 27421 25823 27455
rect 27905 27421 27939 27455
rect 28181 27421 28215 27455
rect 29561 27421 29595 27455
rect 30021 27421 30055 27455
rect 30389 27421 30423 27455
rect 30482 27421 30516 27455
rect 30665 27421 30699 27455
rect 30757 27421 30791 27455
rect 30895 27421 30929 27455
rect 33701 27421 33735 27455
rect 33977 27421 34011 27455
rect 10057 27353 10091 27387
rect 11989 27353 12023 27387
rect 17049 27353 17083 27387
rect 18061 27353 18095 27387
rect 18521 27353 18555 27387
rect 22753 27353 22787 27387
rect 23121 27353 23155 27387
rect 23397 27353 23431 27387
rect 23489 27353 23523 27387
rect 26065 27353 26099 27387
rect 6837 27285 6871 27319
rect 11529 27285 11563 27319
rect 11621 27285 11655 27319
rect 14289 27285 14323 27319
rect 14381 27285 14415 27319
rect 17325 27285 17359 27319
rect 18797 27285 18831 27319
rect 27813 27285 27847 27319
rect 27997 27285 28031 27319
rect 29653 27285 29687 27319
rect 29837 27285 29871 27319
rect 31033 27285 31067 27319
rect 33609 27285 33643 27319
rect 10241 27081 10275 27115
rect 16681 27081 16715 27115
rect 16957 27081 16991 27115
rect 18061 27081 18095 27115
rect 18797 27081 18831 27115
rect 26985 27081 27019 27115
rect 15485 27013 15519 27047
rect 22477 27013 22511 27047
rect 26433 27013 26467 27047
rect 29745 27013 29779 27047
rect 6653 26945 6687 26979
rect 10425 26945 10459 26979
rect 12254 26945 12288 26979
rect 12358 26945 12392 26979
rect 12541 26945 12575 26979
rect 12633 26945 12667 26979
rect 12771 26945 12805 26979
rect 14461 26967 14495 27001
rect 14933 26945 14967 26979
rect 15669 26945 15703 26979
rect 16865 26945 16899 26979
rect 17049 26945 17083 26979
rect 17693 26945 17727 26979
rect 17785 26945 17819 26979
rect 19165 26945 19199 26979
rect 22385 26945 22419 26979
rect 22569 26945 22603 26979
rect 22753 26945 22787 26979
rect 27169 26945 27203 26979
rect 27537 26945 27571 26979
rect 29469 26945 29503 26979
rect 31677 26945 31711 26979
rect 33149 26945 33183 26979
rect 33425 26945 33459 26979
rect 6929 26877 6963 26911
rect 14657 26877 14691 26911
rect 14749 26877 14783 26911
rect 19073 26877 19107 26911
rect 26157 26877 26191 26911
rect 26341 26877 26375 26911
rect 27813 26877 27847 26911
rect 33701 26877 33735 26911
rect 35449 26877 35483 26911
rect 14565 26809 14599 26843
rect 17233 26809 17267 26843
rect 26801 26809 26835 26843
rect 33333 26809 33367 26843
rect 8401 26741 8435 26775
rect 12909 26741 12943 26775
rect 14289 26741 14323 26775
rect 17693 26741 17727 26775
rect 18981 26741 19015 26775
rect 22201 26741 22235 26775
rect 29285 26741 29319 26775
rect 31217 26741 31251 26775
rect 31493 26741 31527 26775
rect 7757 26537 7791 26571
rect 13829 26537 13863 26571
rect 14473 26537 14507 26571
rect 15117 26537 15151 26571
rect 17417 26537 17451 26571
rect 27813 26537 27847 26571
rect 30297 26537 30331 26571
rect 33241 26537 33275 26571
rect 8033 26469 8067 26503
rect 21373 26469 21407 26503
rect 25973 26469 26007 26503
rect 34897 26469 34931 26503
rect 7573 26401 7607 26435
rect 8585 26401 8619 26435
rect 28365 26401 28399 26435
rect 29653 26401 29687 26435
rect 31309 26401 31343 26435
rect 33057 26401 33091 26435
rect 33885 26401 33919 26435
rect 35265 26401 35299 26435
rect 4537 26333 4571 26367
rect 4629 26333 4663 26367
rect 4813 26333 4847 26367
rect 6837 26333 6871 26367
rect 7297 26333 7331 26367
rect 7941 26333 7975 26367
rect 8401 26333 8435 26367
rect 9137 26333 9171 26367
rect 13553 26333 13587 26367
rect 13645 26333 13679 26367
rect 13921 26333 13955 26367
rect 14657 26333 14691 26367
rect 14749 26333 14783 26367
rect 15025 26333 15059 26367
rect 15301 26333 15335 26367
rect 15485 26333 15519 26367
rect 15669 26333 15703 26367
rect 16221 26333 16255 26367
rect 16865 26333 16899 26367
rect 17141 26333 17175 26367
rect 17233 26333 17267 26367
rect 20821 26333 20855 26367
rect 21189 26333 21223 26367
rect 23581 26333 23615 26367
rect 23857 26333 23891 26367
rect 25421 26333 25455 26367
rect 25697 26333 25731 26367
rect 25789 26333 25823 26367
rect 26252 26311 26286 26345
rect 26341 26333 26375 26367
rect 26525 26333 26559 26367
rect 26617 26333 26651 26367
rect 29837 26333 29871 26367
rect 30757 26333 30791 26367
rect 30849 26333 30883 26367
rect 31033 26333 31067 26367
rect 33609 26333 33643 26367
rect 34713 26333 34747 26367
rect 34989 26333 35023 26367
rect 5089 26265 5123 26299
rect 7389 26265 7423 26299
rect 8493 26265 8527 26299
rect 13369 26265 13403 26299
rect 14841 26265 14875 26299
rect 15393 26265 15427 26299
rect 16037 26265 16071 26299
rect 16405 26265 16439 26299
rect 17049 26265 17083 26299
rect 20269 26265 20303 26299
rect 20453 26265 20487 26299
rect 20637 26265 20671 26299
rect 21005 26265 21039 26299
rect 21097 26265 21131 26299
rect 23397 26265 23431 26299
rect 25605 26265 25639 26299
rect 28273 26265 28307 26299
rect 29929 26265 29963 26299
rect 37013 26265 37047 26299
rect 6929 26197 6963 26231
rect 9045 26197 9079 26231
rect 23765 26197 23799 26231
rect 26065 26197 26099 26231
rect 28181 26197 28215 26231
rect 33701 26197 33735 26231
rect 5457 25993 5491 26027
rect 16405 25993 16439 26027
rect 19073 25993 19107 26027
rect 23949 25993 23983 26027
rect 25237 25993 25271 26027
rect 32137 25993 32171 26027
rect 34805 25993 34839 26027
rect 35265 25993 35299 26027
rect 18797 25925 18831 25959
rect 18889 25925 18923 25959
rect 19533 25925 19567 25959
rect 20637 25925 20671 25959
rect 31953 25925 31987 25959
rect 1777 25857 1811 25891
rect 3065 25857 3099 25891
rect 5641 25857 5675 25891
rect 16221 25857 16255 25891
rect 18705 25857 18739 25891
rect 19303 25857 19337 25891
rect 19441 25857 19475 25891
rect 19661 25857 19695 25891
rect 19809 25857 19843 25891
rect 20453 25857 20487 25891
rect 20729 25857 20763 25891
rect 20821 25857 20855 25891
rect 22477 25857 22511 25891
rect 22661 25857 22695 25891
rect 22753 25857 22787 25891
rect 23121 25857 23155 25891
rect 23397 25857 23431 25891
rect 23857 25857 23891 25891
rect 24317 25857 24351 25891
rect 24593 25857 24627 25891
rect 24777 25857 24811 25891
rect 24869 25857 24903 25891
rect 24961 25857 24995 25891
rect 25513 25857 25547 25891
rect 25605 25857 25639 25891
rect 25697 25857 25731 25891
rect 25881 25857 25915 25891
rect 25973 25857 26007 25891
rect 26157 25857 26191 25891
rect 26249 25857 26283 25891
rect 26341 25857 26375 25891
rect 31493 25857 31527 25891
rect 31585 25857 31619 25891
rect 31769 25857 31803 25891
rect 32505 25857 32539 25891
rect 32965 25857 32999 25891
rect 33149 25857 33183 25891
rect 33241 25857 33275 25891
rect 33333 25857 33367 25891
rect 34345 25857 34379 25891
rect 34437 25857 34471 25891
rect 35081 25857 35115 25891
rect 35173 25857 35207 25891
rect 3341 25789 3375 25823
rect 3617 25789 3651 25823
rect 8677 25789 8711 25823
rect 8953 25789 8987 25823
rect 23765 25789 23799 25823
rect 24225 25789 24259 25823
rect 32597 25789 32631 25823
rect 32689 25789 32723 25823
rect 34161 25789 34195 25823
rect 18521 25721 18555 25755
rect 22569 25721 22603 25755
rect 23489 25721 23523 25755
rect 34989 25721 35023 25755
rect 1501 25653 1535 25687
rect 2881 25653 2915 25687
rect 5089 25653 5123 25687
rect 10425 25653 10459 25687
rect 19165 25653 19199 25687
rect 21005 25653 21039 25687
rect 22293 25653 22327 25687
rect 23857 25653 23891 25687
rect 24133 25653 24167 25687
rect 25329 25653 25363 25687
rect 26617 25653 26651 25687
rect 33609 25653 33643 25687
rect 3893 25449 3927 25483
rect 9045 25449 9079 25483
rect 18797 25449 18831 25483
rect 22845 25449 22879 25483
rect 20913 25381 20947 25415
rect 21097 25381 21131 25415
rect 27813 25381 27847 25415
rect 2145 25313 2179 25347
rect 9873 25313 9907 25347
rect 11897 25313 11931 25347
rect 12541 25313 12575 25347
rect 14841 25313 14875 25347
rect 17417 25313 17451 25347
rect 21005 25313 21039 25347
rect 23673 25313 23707 25347
rect 28917 25313 28951 25347
rect 1869 25245 1903 25279
rect 4077 25245 4111 25279
rect 7573 25245 7607 25279
rect 9229 25245 9263 25279
rect 9689 25245 9723 25279
rect 10149 25245 10183 25279
rect 12357 25245 12391 25279
rect 12955 25245 12989 25279
rect 13093 25245 13127 25279
rect 13185 25245 13219 25279
rect 13368 25245 13402 25279
rect 13461 25245 13495 25279
rect 14565 25245 14599 25279
rect 15945 25245 15979 25279
rect 16680 25223 16714 25257
rect 16773 25245 16807 25279
rect 16865 25245 16899 25279
rect 17049 25245 17083 25279
rect 17233 25245 17267 25279
rect 18429 25245 18463 25279
rect 18521 25245 18555 25279
rect 18613 25245 18647 25279
rect 20729 25245 20763 25279
rect 21276 25245 21310 25279
rect 21465 25245 21499 25279
rect 21593 25245 21627 25279
rect 21741 25245 21775 25279
rect 22201 25245 22235 25279
rect 22294 25245 22328 25279
rect 22666 25245 22700 25279
rect 23029 25245 23063 25279
rect 24777 25245 24811 25279
rect 24961 25245 24995 25279
rect 25053 25245 25087 25279
rect 25237 25245 25271 25279
rect 25329 25245 25363 25279
rect 27169 25245 27203 25279
rect 27262 25245 27296 25279
rect 27445 25245 27479 25279
rect 27634 25245 27668 25279
rect 28457 25245 28491 25279
rect 28733 25245 28767 25279
rect 29193 25245 29227 25279
rect 30021 25245 30055 25279
rect 30205 25245 30239 25279
rect 30297 25245 30331 25279
rect 30389 25245 30423 25279
rect 34345 25245 34379 25279
rect 34713 25245 34747 25279
rect 10425 25177 10459 25211
rect 12449 25177 12483 25211
rect 16405 25177 16439 25211
rect 21373 25177 21407 25211
rect 22477 25177 22511 25211
rect 22569 25177 22603 25211
rect 27537 25177 27571 25211
rect 34989 25177 35023 25211
rect 36737 25177 36771 25211
rect 3617 25109 3651 25143
rect 7481 25109 7515 25143
rect 9321 25109 9355 25143
rect 9781 25109 9815 25143
rect 11989 25109 12023 25143
rect 12817 25109 12851 25143
rect 16129 25109 16163 25143
rect 20545 25109 20579 25143
rect 28549 25109 28583 25143
rect 29101 25109 29135 25143
rect 30665 25109 30699 25143
rect 34529 25109 34563 25143
rect 4353 24905 4387 24939
rect 4721 24905 4755 24939
rect 9597 24905 9631 24939
rect 10333 24905 10367 24939
rect 10609 24905 10643 24939
rect 14289 24905 14323 24939
rect 21465 24905 21499 24939
rect 23397 24905 23431 24939
rect 26985 24905 27019 24939
rect 34253 24905 34287 24939
rect 34621 24905 34655 24939
rect 12357 24837 12391 24871
rect 13001 24837 13035 24871
rect 18521 24837 18555 24871
rect 21097 24837 21131 24871
rect 21373 24837 21407 24871
rect 27353 24837 27387 24871
rect 30941 24837 30975 24871
rect 5917 24769 5951 24803
rect 10425 24769 10459 24803
rect 10793 24769 10827 24803
rect 12173 24769 12207 24803
rect 12449 24769 12483 24803
rect 12541 24769 12575 24803
rect 12817 24769 12851 24803
rect 14289 24769 14323 24803
rect 14933 24769 14967 24803
rect 15393 24769 15427 24803
rect 16221 24769 16255 24803
rect 16865 24769 16899 24803
rect 17233 24769 17267 24803
rect 17877 24769 17911 24803
rect 18613 24769 18647 24803
rect 19073 24769 19107 24803
rect 21281 24769 21315 24803
rect 23489 24769 23523 24803
rect 23857 24769 23891 24803
rect 25881 24769 25915 24803
rect 26157 24769 26191 24803
rect 28641 24769 28675 24803
rect 28917 24769 28951 24803
rect 31125 24769 31159 24803
rect 31309 24769 31343 24803
rect 31585 24769 31619 24803
rect 31953 24769 31987 24803
rect 33057 24769 33091 24803
rect 33241 24769 33275 24803
rect 33517 24769 33551 24803
rect 1409 24701 1443 24735
rect 1685 24701 1719 24735
rect 4813 24701 4847 24735
rect 4997 24701 5031 24735
rect 7297 24701 7331 24735
rect 7573 24701 7607 24735
rect 9045 24701 9079 24735
rect 9689 24701 9723 24735
rect 9873 24701 9907 24735
rect 15025 24701 15059 24735
rect 16681 24701 16715 24735
rect 17325 24701 17359 24735
rect 24133 24701 24167 24735
rect 27445 24701 27479 24735
rect 27537 24701 27571 24735
rect 29193 24701 29227 24735
rect 34713 24701 34747 24735
rect 34805 24701 34839 24735
rect 12725 24633 12759 24667
rect 28825 24633 28859 24667
rect 33425 24633 33459 24667
rect 3157 24565 3191 24599
rect 5733 24565 5767 24599
rect 9229 24565 9263 24599
rect 13185 24565 13219 24599
rect 18337 24565 18371 24599
rect 21649 24565 21683 24599
rect 25789 24565 25823 24599
rect 25973 24565 26007 24599
rect 31217 24565 31251 24599
rect 33149 24565 33183 24599
rect 1777 24361 1811 24395
rect 3801 24361 3835 24395
rect 7941 24361 7975 24395
rect 13737 24361 13771 24395
rect 13921 24361 13955 24395
rect 18613 24361 18647 24395
rect 18797 24361 18831 24395
rect 19901 24361 19935 24395
rect 22109 24361 22143 24395
rect 27353 24361 27387 24395
rect 31769 24361 31803 24395
rect 7021 24293 7055 24327
rect 15209 24293 15243 24327
rect 16405 24293 16439 24327
rect 20729 24293 20763 24327
rect 24041 24293 24075 24327
rect 33057 24293 33091 24327
rect 33517 24293 33551 24327
rect 33701 24293 33735 24327
rect 34437 24293 34471 24327
rect 2973 24225 3007 24259
rect 4353 24225 4387 24259
rect 5273 24225 5307 24259
rect 5549 24225 5583 24259
rect 13001 24225 13035 24259
rect 19993 24225 20027 24259
rect 23305 24225 23339 24259
rect 24869 24225 24903 24259
rect 25605 24225 25639 24259
rect 25881 24225 25915 24259
rect 28273 24225 28307 24259
rect 1961 24157 1995 24191
rect 4169 24157 4203 24191
rect 8125 24157 8159 24191
rect 9137 24157 9171 24191
rect 12817 24157 12851 24191
rect 14381 24157 14415 24191
rect 14749 24157 14783 24191
rect 15117 24157 15151 24191
rect 15761 24157 15795 24191
rect 15945 24157 15979 24191
rect 16037 24157 16071 24191
rect 16163 24157 16197 24191
rect 17107 24157 17141 24191
rect 17233 24157 17267 24191
rect 17325 24157 17359 24191
rect 17509 24157 17543 24191
rect 17877 24157 17911 24191
rect 18153 24157 18187 24191
rect 18705 24157 18739 24191
rect 18889 24157 18923 24191
rect 19073 24157 19107 24191
rect 19533 24157 19567 24191
rect 19717 24157 19751 24191
rect 20361 24157 20395 24191
rect 20821 24157 20855 24191
rect 22109 24157 22143 24191
rect 22937 24157 22971 24191
rect 23673 24157 23707 24191
rect 23949 24157 23983 24191
rect 24777 24157 24811 24191
rect 25329 24157 25363 24191
rect 28181 24157 28215 24191
rect 28457 24157 28491 24191
rect 29561 24157 29595 24191
rect 29740 24157 29774 24191
rect 29837 24157 29871 24191
rect 29929 24157 29963 24191
rect 31401 24157 31435 24191
rect 31585 24157 31619 24191
rect 31677 24157 31711 24191
rect 32229 24157 32263 24191
rect 32413 24157 32447 24191
rect 32781 24157 32815 24191
rect 32873 24157 32907 24191
rect 33149 24157 33183 24191
rect 33241 24157 33275 24191
rect 33333 24157 33367 24191
rect 33609 24157 33643 24191
rect 33885 24157 33919 24191
rect 34069 24157 34103 24191
rect 34161 24157 34195 24191
rect 34345 24157 34379 24191
rect 13783 24123 13817 24157
rect 13553 24089 13587 24123
rect 16865 24089 16899 24123
rect 20085 24089 20119 24123
rect 20453 24089 20487 24123
rect 33517 24089 33551 24123
rect 33977 24089 34011 24123
rect 2329 24021 2363 24055
rect 2697 24021 2731 24055
rect 2789 24021 2823 24055
rect 4261 24021 4295 24055
rect 9045 24021 9079 24055
rect 12633 24021 12667 24055
rect 18153 24021 18187 24055
rect 18337 24021 18371 24055
rect 19257 24021 19291 24055
rect 19625 24021 19659 24055
rect 20545 24021 20579 24055
rect 30205 24021 30239 24055
rect 31493 24021 31527 24055
rect 32137 24021 32171 24055
rect 32413 24021 32447 24055
rect 32597 24021 32631 24055
rect 6377 23817 6411 23851
rect 12725 23817 12759 23851
rect 15761 23817 15795 23851
rect 18705 23817 18739 23851
rect 19901 23817 19935 23851
rect 29101 23817 29135 23851
rect 32229 23817 32263 23851
rect 13461 23749 13495 23783
rect 14289 23749 14323 23783
rect 14657 23749 14691 23783
rect 15025 23749 15059 23783
rect 18521 23749 18555 23783
rect 19815 23749 19849 23783
rect 21097 23749 21131 23783
rect 25881 23749 25915 23783
rect 27261 23749 27295 23783
rect 27905 23749 27939 23783
rect 27997 23749 28031 23783
rect 28733 23749 28767 23783
rect 5641 23681 5675 23715
rect 6745 23681 6779 23715
rect 6837 23681 6871 23715
rect 8677 23681 8711 23715
rect 11253 23681 11287 23715
rect 12909 23681 12943 23715
rect 13093 23681 13127 23715
rect 14197 23681 14231 23715
rect 14749 23681 14783 23715
rect 14841 23681 14875 23715
rect 15301 23681 15335 23715
rect 15485 23681 15519 23715
rect 15669 23681 15703 23715
rect 17325 23681 17359 23715
rect 17417 23681 17451 23715
rect 17969 23681 18003 23715
rect 18061 23681 18095 23715
rect 19073 23681 19107 23715
rect 19165 23681 19199 23715
rect 19257 23681 19291 23715
rect 19441 23681 19475 23715
rect 19993 23681 20027 23715
rect 20269 23681 20303 23715
rect 20821 23681 20855 23715
rect 22385 23681 22419 23715
rect 22569 23681 22603 23715
rect 23305 23681 23339 23715
rect 23673 23681 23707 23715
rect 23857 23681 23891 23715
rect 24685 23681 24719 23715
rect 25053 23681 25087 23715
rect 25145 23681 25179 23715
rect 26065 23681 26099 23715
rect 27077 23681 27111 23715
rect 27353 23681 27387 23715
rect 27445 23681 27479 23715
rect 27721 23681 27755 23715
rect 28089 23681 28123 23715
rect 28641 23681 28675 23715
rect 32137 23681 32171 23715
rect 33149 23681 33183 23715
rect 35541 23681 35575 23715
rect 6929 23613 6963 23647
rect 8953 23613 8987 23647
rect 10425 23613 10459 23647
rect 16037 23613 16071 23647
rect 17233 23613 17267 23647
rect 17509 23613 17543 23647
rect 22661 23613 22695 23647
rect 23213 23613 23247 23647
rect 26249 23613 26283 23647
rect 28457 23613 28491 23647
rect 34897 23613 34931 23647
rect 35633 23613 35667 23647
rect 15853 23545 15887 23579
rect 18981 23545 19015 23579
rect 19533 23545 19567 23579
rect 20177 23545 20211 23579
rect 22201 23545 22235 23579
rect 24317 23545 24351 23579
rect 27629 23545 27663 23579
rect 28273 23545 28307 23579
rect 5549 23477 5583 23511
rect 10609 23477 10643 23511
rect 15117 23477 15151 23511
rect 15945 23477 15979 23511
rect 17693 23477 17727 23511
rect 17785 23477 17819 23511
rect 33241 23477 33275 23511
rect 2237 23273 2271 23307
rect 2973 23273 3007 23307
rect 4261 23273 4295 23307
rect 4997 23273 5031 23307
rect 6285 23273 6319 23307
rect 6478 23273 6512 23307
rect 7021 23273 7055 23307
rect 9321 23273 9355 23307
rect 14105 23273 14139 23307
rect 20637 23273 20671 23307
rect 20821 23273 20855 23307
rect 23857 23273 23891 23307
rect 35725 23273 35759 23307
rect 23489 23205 23523 23239
rect 34805 23205 34839 23239
rect 35541 23205 35575 23239
rect 5733 23137 5767 23171
rect 8125 23137 8159 23171
rect 12817 23137 12851 23171
rect 14749 23137 14783 23171
rect 15485 23137 15519 23171
rect 16221 23137 16255 23171
rect 18705 23137 18739 23171
rect 20545 23137 20579 23171
rect 22017 23137 22051 23171
rect 35633 23137 35667 23171
rect 36277 23137 36311 23171
rect 1961 23069 1995 23103
rect 2513 23069 2547 23103
rect 2605 23069 2639 23103
rect 2697 23069 2731 23103
rect 2881 23069 2915 23103
rect 3157 23069 3191 23103
rect 3617 23069 3651 23103
rect 4445 23069 4479 23103
rect 4905 23069 4939 23103
rect 5198 23079 5232 23113
rect 5365 23069 5399 23103
rect 5641 23069 5675 23103
rect 5917 23069 5951 23103
rect 6101 23069 6135 23103
rect 6193 23069 6227 23103
rect 6745 23069 6779 23103
rect 6929 23069 6963 23103
rect 7205 23069 7239 23103
rect 7665 23069 7699 23103
rect 9505 23069 9539 23103
rect 9597 23069 9631 23103
rect 9873 23069 9907 23103
rect 10517 23069 10551 23103
rect 10609 23069 10643 23103
rect 10793 23069 10827 23103
rect 15393 23069 15427 23103
rect 15761 23069 15795 23103
rect 15853 23069 15887 23103
rect 16681 23069 16715 23103
rect 17049 23069 17083 23103
rect 17141 23069 17175 23103
rect 17325 23069 17359 23103
rect 17693 23069 17727 23103
rect 18061 23069 18095 23103
rect 18613 23069 18647 23103
rect 20453 23069 20487 23103
rect 21189 23069 21223 23103
rect 21741 23069 21775 23103
rect 22753 23069 22787 23103
rect 22937 23069 22971 23103
rect 23397 23069 23431 23103
rect 23765 23069 23799 23103
rect 23949 23069 23983 23103
rect 24961 23069 24995 23103
rect 25237 23069 25271 23103
rect 25697 23069 25731 23103
rect 26065 23069 26099 23103
rect 29745 23069 29779 23103
rect 29929 23069 29963 23103
rect 32505 23069 32539 23103
rect 32781 23069 32815 23103
rect 32873 23069 32907 23103
rect 33057 23069 33091 23103
rect 34713 23069 34747 23103
rect 34989 23069 35023 23103
rect 35357 23069 35391 23103
rect 35909 23069 35943 23103
rect 36185 23069 36219 23103
rect 36369 23069 36403 23103
rect 3249 23001 3283 23035
rect 3341 23001 3375 23035
rect 3479 23001 3513 23035
rect 4537 23001 4571 23035
rect 4629 23001 4663 23035
rect 4747 23001 4781 23035
rect 5273 23001 5307 23035
rect 5483 23001 5517 23035
rect 6437 23001 6471 23035
rect 6653 23001 6687 23035
rect 6837 23001 6871 23035
rect 7297 23001 7331 23035
rect 7389 23001 7423 23035
rect 7507 23001 7541 23035
rect 7757 23001 7791 23035
rect 7941 23001 7975 23035
rect 9689 23001 9723 23035
rect 11069 23001 11103 23035
rect 14289 23001 14323 23035
rect 14473 23001 14507 23035
rect 21005 23001 21039 23035
rect 25881 23001 25915 23035
rect 25973 23001 26007 23035
rect 30021 23001 30055 23035
rect 33241 23001 33275 23035
rect 35173 23001 35207 23035
rect 35265 23001 35299 23035
rect 1777 22933 1811 22967
rect 25421 22933 25455 22967
rect 26249 22933 26283 22967
rect 32321 22933 32355 22967
rect 32689 22933 32723 22967
rect 36093 22933 36127 22967
rect 2881 22729 2915 22763
rect 3433 22729 3467 22763
rect 3985 22729 4019 22763
rect 5089 22729 5123 22763
rect 5549 22729 5583 22763
rect 9505 22729 9539 22763
rect 11069 22729 11103 22763
rect 11897 22729 11931 22763
rect 13001 22729 13035 22763
rect 15485 22729 15519 22763
rect 17969 22729 18003 22763
rect 22109 22729 22143 22763
rect 24409 22729 24443 22763
rect 27537 22729 27571 22763
rect 27997 22729 28031 22763
rect 30297 22729 30331 22763
rect 32229 22729 32263 22763
rect 35357 22729 35391 22763
rect 37381 22729 37415 22763
rect 5457 22661 5491 22695
rect 6377 22661 6411 22695
rect 7849 22661 7883 22695
rect 13645 22661 13679 22695
rect 20361 22661 20395 22695
rect 33701 22661 33735 22695
rect 35173 22661 35207 22695
rect 36829 22661 36863 22695
rect 2789 22593 2823 22627
rect 2973 22593 3007 22627
rect 3617 22593 3651 22627
rect 3801 22593 3835 22627
rect 3893 22593 3927 22627
rect 4077 22593 4111 22627
rect 5273 22593 5307 22627
rect 5549 22593 5583 22627
rect 5733 22593 5767 22627
rect 6561 22593 6595 22627
rect 6745 22593 6779 22627
rect 8033 22593 8067 22627
rect 9689 22593 9723 22627
rect 11253 22593 11287 22627
rect 12357 22593 12391 22627
rect 12541 22593 12575 22627
rect 12633 22593 12667 22627
rect 12725 22593 12759 22627
rect 13369 22593 13403 22627
rect 13553 22593 13587 22627
rect 14197 22593 14231 22627
rect 14565 22593 14599 22627
rect 15423 22593 15457 22627
rect 16129 22593 16163 22627
rect 16313 22593 16347 22627
rect 17141 22593 17175 22627
rect 17325 22593 17359 22627
rect 17877 22593 17911 22627
rect 20729 22593 20763 22627
rect 22017 22593 22051 22627
rect 22201 22593 22235 22627
rect 22569 22593 22603 22627
rect 22661 22593 22695 22627
rect 22937 22593 22971 22627
rect 23305 22593 23339 22627
rect 23673 22593 23707 22627
rect 24041 22593 24075 22627
rect 24317 22593 24351 22627
rect 24501 22593 24535 22627
rect 25605 22593 25639 22627
rect 26985 22593 27019 22627
rect 27169 22593 27203 22627
rect 27261 22593 27295 22627
rect 27353 22593 27387 22627
rect 27721 22593 27755 22627
rect 29653 22593 29687 22627
rect 29837 22593 29871 22627
rect 29929 22593 29963 22627
rect 30205 22593 30239 22627
rect 30389 22593 30423 22627
rect 30481 22593 30515 22627
rect 30665 22593 30699 22627
rect 32137 22593 32171 22627
rect 32321 22593 32355 22627
rect 32781 22593 32815 22627
rect 32873 22593 32907 22627
rect 33149 22593 33183 22627
rect 33241 22593 33275 22627
rect 33425 22593 33459 22627
rect 33517 22593 33551 22627
rect 35449 22593 35483 22627
rect 36093 22593 36127 22627
rect 36277 22593 36311 22627
rect 36369 22593 36403 22627
rect 36553 22593 36587 22627
rect 36645 22593 36679 22627
rect 37289 22593 37323 22627
rect 37657 22593 37691 22627
rect 9965 22525 9999 22559
rect 11989 22525 12023 22559
rect 12081 22525 12115 22559
rect 14657 22525 14691 22559
rect 15945 22525 15979 22559
rect 16497 22525 16531 22559
rect 25789 22525 25823 22559
rect 30021 22525 30055 22559
rect 32689 22525 32723 22559
rect 32965 22525 32999 22559
rect 8217 22457 8251 22491
rect 11529 22457 11563 22491
rect 15853 22457 15887 22491
rect 23949 22457 23983 22491
rect 37841 22457 37875 22491
rect 9873 22389 9907 22423
rect 15301 22389 15335 22423
rect 25421 22389 25455 22423
rect 29469 22389 29503 22423
rect 30665 22389 30699 22423
rect 32505 22389 32539 22423
rect 35173 22389 35207 22423
rect 36093 22389 36127 22423
rect 36461 22389 36495 22423
rect 37013 22389 37047 22423
rect 3985 22185 4019 22219
rect 10333 22185 10367 22219
rect 12173 22185 12207 22219
rect 29193 22185 29227 22219
rect 14565 22117 14599 22151
rect 17049 22117 17083 22151
rect 19349 22117 19383 22151
rect 22661 22117 22695 22151
rect 30757 22117 30791 22151
rect 32229 22117 32263 22151
rect 32505 22117 32539 22151
rect 10057 22049 10091 22083
rect 11621 22049 11655 22083
rect 12265 22049 12299 22083
rect 23673 22049 23707 22083
rect 25329 22049 25363 22083
rect 27261 22049 27295 22083
rect 30389 22049 30423 22083
rect 31217 22049 31251 22083
rect 31401 22049 31435 22083
rect 32873 22049 32907 22083
rect 33057 22049 33091 22083
rect 33149 22049 33183 22083
rect 33241 22049 33275 22083
rect 35265 22049 35299 22083
rect 35725 22049 35759 22083
rect 35817 22049 35851 22083
rect 36001 22049 36035 22083
rect 37013 22049 37047 22083
rect 1961 21981 1995 22015
rect 4261 21981 4295 22015
rect 7757 21981 7791 22015
rect 10241 21981 10275 22015
rect 10425 21981 10459 22015
rect 12817 21981 12851 22015
rect 14841 21981 14875 22015
rect 15025 21981 15059 22015
rect 15577 21981 15611 22015
rect 15761 21981 15795 22015
rect 15853 21981 15887 22015
rect 16037 21981 16071 22015
rect 16405 21981 16439 22015
rect 16589 21981 16623 22015
rect 16865 21981 16899 22015
rect 17049 21981 17083 22015
rect 17509 21981 17543 22015
rect 19441 21981 19475 22015
rect 19717 21981 19751 22015
rect 19993 21981 20027 22015
rect 20085 21981 20119 22015
rect 22201 21981 22235 22015
rect 22385 21981 22419 22015
rect 22753 21981 22787 22015
rect 22937 21981 22971 22015
rect 23581 21981 23615 22015
rect 23857 21981 23891 22015
rect 24685 21981 24719 22015
rect 24869 21981 24903 22015
rect 24961 21981 24995 22015
rect 25053 21981 25087 22015
rect 25789 21981 25823 22015
rect 26065 21981 26099 22015
rect 26209 21981 26243 22015
rect 27445 21981 27479 22015
rect 27721 21981 27755 22015
rect 27997 21981 28031 22015
rect 28365 21981 28399 22015
rect 28641 21981 28675 22015
rect 28825 21981 28859 22015
rect 28917 21981 28951 22015
rect 29009 21981 29043 22015
rect 31125 21981 31159 22015
rect 31861 21981 31895 22015
rect 31953 21981 31987 22015
rect 32413 21981 32447 22015
rect 32597 21981 32631 22015
rect 32689 21981 32723 22015
rect 33333 21981 33367 22015
rect 35081 21981 35115 22015
rect 35909 21981 35943 22015
rect 36829 21981 36863 22015
rect 32137 21947 32171 21981
rect 3801 21913 3835 21947
rect 12449 21913 12483 21947
rect 16681 21913 16715 21947
rect 25973 21913 26007 21947
rect 27813 21913 27847 21947
rect 28181 21913 28215 21947
rect 28273 21913 28307 21947
rect 29561 21913 29595 21947
rect 35173 21913 35207 21947
rect 1777 21845 1811 21879
rect 4001 21845 4035 21879
rect 4169 21845 4203 21879
rect 4353 21845 4387 21879
rect 8217 21845 8251 21879
rect 9413 21845 9447 21879
rect 9781 21845 9815 21879
rect 9873 21845 9907 21879
rect 11713 21845 11747 21879
rect 11805 21845 11839 21879
rect 12541 21845 12575 21879
rect 12633 21845 12667 21879
rect 26358 21845 26392 21879
rect 27629 21845 27663 21879
rect 28549 21845 28583 21879
rect 32038 21845 32072 21879
rect 34713 21845 34747 21879
rect 35541 21845 35575 21879
rect 36645 21845 36679 21879
rect 3249 21641 3283 21675
rect 9137 21641 9171 21675
rect 9781 21641 9815 21675
rect 11529 21641 11563 21675
rect 14933 21641 14967 21675
rect 17325 21641 17359 21675
rect 22937 21641 22971 21675
rect 25421 21641 25455 21675
rect 32597 21641 32631 21675
rect 35265 21641 35299 21675
rect 35909 21641 35943 21675
rect 36461 21641 36495 21675
rect 1685 21573 1719 21607
rect 4583 21573 4617 21607
rect 5181 21573 5215 21607
rect 18889 21573 18923 21607
rect 25053 21573 25087 21607
rect 25605 21573 25639 21607
rect 27445 21573 27479 21607
rect 29745 21573 29779 21607
rect 29929 21573 29963 21607
rect 3617 21505 3651 21539
rect 3709 21505 3743 21539
rect 4077 21505 4111 21539
rect 4261 21505 4295 21539
rect 4353 21505 4387 21539
rect 4445 21505 4479 21539
rect 4721 21505 4755 21539
rect 4997 21505 5031 21539
rect 5733 21505 5767 21539
rect 5825 21505 5859 21539
rect 5917 21505 5951 21539
rect 6101 21505 6135 21539
rect 9321 21505 9355 21539
rect 9413 21505 9447 21539
rect 9505 21505 9539 21539
rect 9689 21505 9723 21539
rect 9965 21505 9999 21539
rect 10057 21505 10091 21539
rect 10149 21505 10183 21539
rect 10333 21505 10367 21539
rect 11897 21505 11931 21539
rect 13369 21505 13403 21539
rect 15112 21505 15146 21539
rect 15209 21505 15243 21539
rect 15301 21505 15335 21539
rect 15484 21505 15518 21539
rect 15577 21505 15611 21539
rect 17509 21505 17543 21539
rect 17693 21505 17727 21539
rect 17785 21505 17819 21539
rect 17877 21505 17911 21539
rect 18061 21505 18095 21539
rect 19533 21505 19567 21539
rect 19901 21505 19935 21539
rect 20177 21505 20211 21539
rect 20361 21505 20395 21539
rect 23029 21505 23063 21539
rect 23121 21505 23155 21539
rect 23397 21505 23431 21539
rect 24869 21505 24903 21539
rect 25145 21505 25179 21539
rect 25237 21505 25271 21539
rect 25697 21505 25731 21539
rect 27629 21505 27663 21539
rect 27721 21505 27755 21539
rect 30021 21505 30055 21539
rect 30757 21505 30791 21539
rect 30941 21505 30975 21539
rect 32505 21505 32539 21539
rect 32689 21505 32723 21539
rect 33333 21505 33367 21539
rect 33425 21505 33459 21539
rect 33517 21505 33551 21539
rect 33701 21505 33735 21539
rect 33793 21505 33827 21539
rect 33977 21505 34011 21539
rect 35173 21505 35207 21539
rect 35817 21505 35851 21539
rect 36277 21505 36311 21539
rect 36369 21505 36403 21539
rect 36737 21505 36771 21539
rect 1409 21437 1443 21471
rect 3157 21437 3191 21471
rect 3893 21437 3927 21471
rect 5365 21437 5399 21471
rect 6561 21437 6595 21471
rect 6837 21437 6871 21471
rect 11989 21437 12023 21471
rect 12173 21437 12207 21471
rect 13093 21437 13127 21471
rect 14289 21437 14323 21471
rect 18153 21437 18187 21471
rect 18521 21437 18555 21471
rect 19625 21437 19659 21471
rect 19809 21437 19843 21471
rect 23213 21437 23247 21471
rect 36001 21437 36035 21471
rect 8309 21369 8343 21403
rect 13829 21369 13863 21403
rect 23581 21369 23615 21403
rect 5457 21301 5491 21335
rect 20269 21301 20303 21335
rect 23121 21301 23155 21335
rect 27537 21301 27571 21335
rect 29745 21301 29779 21335
rect 30941 21301 30975 21335
rect 33057 21301 33091 21335
rect 33885 21301 33919 21335
rect 35449 21301 35483 21335
rect 4353 21097 4387 21131
rect 6929 21097 6963 21131
rect 9505 21097 9539 21131
rect 10149 21097 10183 21131
rect 16957 21097 16991 21131
rect 18429 21097 18463 21131
rect 21189 21097 21223 21131
rect 22017 21097 22051 21131
rect 22845 21097 22879 21131
rect 25053 21097 25087 21131
rect 26801 21097 26835 21131
rect 30573 21097 30607 21131
rect 7205 21029 7239 21063
rect 15485 21029 15519 21063
rect 16313 21029 16347 21063
rect 4077 20961 4111 20995
rect 4169 20961 4203 20995
rect 7757 20961 7791 20995
rect 14381 20961 14415 20995
rect 18981 20961 19015 20995
rect 20269 20961 20303 20995
rect 25145 20961 25179 20995
rect 30665 20961 30699 20995
rect 1777 20893 1811 20927
rect 3893 20893 3927 20927
rect 3985 20893 4019 20927
rect 5457 20893 5491 20927
rect 7113 20893 7147 20927
rect 7573 20893 7607 20927
rect 8953 20893 8987 20927
rect 9321 20893 9355 20927
rect 9597 20893 9631 20927
rect 9873 20893 9907 20927
rect 9965 20893 9999 20927
rect 14565 20893 14599 20927
rect 14749 20893 14783 20927
rect 14841 20893 14875 20927
rect 14933 20893 14967 20927
rect 15209 20893 15243 20927
rect 15306 20893 15340 20927
rect 16129 20893 16163 20927
rect 16221 20893 16255 20927
rect 16405 20893 16439 20927
rect 17136 20893 17170 20927
rect 17509 20893 17543 20927
rect 18554 20893 18588 20927
rect 19073 20893 19107 20927
rect 19349 20893 19383 20927
rect 19533 20893 19567 20927
rect 20177 20893 20211 20927
rect 20361 20893 20395 20927
rect 20545 20893 20579 20927
rect 20693 20893 20727 20927
rect 21010 20893 21044 20927
rect 21373 20893 21407 20927
rect 21466 20893 21500 20927
rect 21741 20893 21775 20927
rect 21838 20893 21872 20927
rect 22201 20893 22235 20927
rect 22385 20893 22419 20927
rect 22477 20893 22511 20927
rect 22569 20893 22603 20927
rect 25053 20893 25087 20927
rect 25329 20893 25363 20927
rect 26985 20893 27019 20927
rect 27077 20893 27111 20927
rect 27353 20893 27387 20927
rect 27629 20893 27663 20927
rect 27813 20893 27847 20927
rect 30389 20893 30423 20927
rect 34988 20893 35022 20927
rect 35081 20893 35115 20927
rect 35173 20893 35207 20927
rect 35357 20893 35391 20927
rect 35449 20893 35483 20927
rect 35633 20893 35667 20927
rect 37197 20893 37231 20927
rect 5273 20825 5307 20859
rect 5641 20825 5675 20859
rect 7665 20825 7699 20859
rect 9137 20825 9171 20859
rect 9229 20825 9263 20859
rect 9781 20825 9815 20859
rect 15117 20825 15151 20859
rect 15761 20825 15795 20859
rect 17233 20825 17267 20859
rect 17325 20825 17359 20859
rect 20821 20825 20855 20859
rect 20913 20825 20947 20859
rect 21649 20825 21683 20859
rect 27169 20825 27203 20859
rect 27445 20825 27479 20859
rect 34713 20825 34747 20859
rect 35541 20825 35575 20859
rect 37565 20825 37599 20859
rect 1501 20757 1535 20791
rect 18613 20757 18647 20791
rect 19441 20757 19475 20791
rect 24869 20757 24903 20791
rect 30205 20757 30239 20791
rect 37381 20757 37415 20791
rect 37841 20757 37875 20791
rect 3709 20553 3743 20587
rect 14841 20553 14875 20587
rect 15853 20553 15887 20587
rect 20177 20553 20211 20587
rect 21281 20553 21315 20587
rect 27813 20553 27847 20587
rect 35449 20553 35483 20587
rect 7573 20485 7607 20519
rect 14657 20485 14691 20519
rect 19809 20485 19843 20519
rect 20545 20485 20579 20519
rect 27537 20485 27571 20519
rect 2789 20417 2823 20451
rect 3525 20417 3559 20451
rect 3801 20417 3835 20451
rect 7665 20417 7699 20451
rect 11713 20417 11747 20451
rect 15945 20417 15979 20451
rect 18061 20417 18095 20451
rect 18153 20417 18187 20451
rect 18521 20417 18555 20451
rect 19257 20417 19291 20451
rect 19993 20417 20027 20451
rect 20085 20417 20119 20451
rect 20361 20417 20395 20451
rect 20637 20417 20671 20451
rect 20730 20417 20764 20451
rect 20913 20417 20947 20451
rect 21005 20417 21039 20451
rect 21102 20417 21136 20451
rect 24317 20417 24351 20451
rect 24409 20417 24443 20451
rect 24593 20417 24627 20451
rect 25145 20417 25179 20451
rect 25237 20417 25271 20451
rect 25789 20417 25823 20451
rect 25973 20417 26007 20451
rect 26065 20417 26099 20451
rect 26157 20417 26191 20451
rect 27261 20417 27295 20451
rect 27445 20417 27479 20451
rect 27629 20417 27663 20451
rect 28917 20417 28951 20451
rect 29101 20417 29135 20451
rect 29745 20417 29779 20451
rect 30297 20417 30331 20451
rect 30573 20417 30607 20451
rect 30757 20417 30791 20451
rect 31033 20417 31067 20451
rect 33149 20417 33183 20451
rect 35909 20417 35943 20451
rect 2881 20349 2915 20383
rect 3065 20349 3099 20383
rect 3341 20349 3375 20383
rect 7757 20349 7791 20383
rect 11621 20349 11655 20383
rect 14289 20349 14323 20383
rect 15485 20349 15519 20383
rect 17601 20349 17635 20383
rect 18613 20349 18647 20383
rect 18797 20349 18831 20383
rect 19165 20349 19199 20383
rect 24501 20349 24535 20383
rect 29653 20349 29687 20383
rect 33241 20349 33275 20383
rect 35633 20349 35667 20383
rect 35725 20349 35759 20383
rect 35817 20349 35851 20383
rect 15669 20281 15703 20315
rect 30665 20281 30699 20315
rect 33517 20281 33551 20315
rect 2421 20213 2455 20247
rect 3893 20213 3927 20247
rect 7205 20213 7239 20247
rect 11989 20213 12023 20247
rect 14657 20213 14691 20247
rect 19441 20213 19475 20247
rect 19717 20213 19751 20247
rect 24133 20213 24167 20247
rect 24961 20213 24995 20247
rect 26341 20213 26375 20247
rect 28917 20213 28951 20247
rect 30021 20213 30055 20247
rect 3801 20009 3835 20043
rect 9781 20009 9815 20043
rect 11621 20009 11655 20043
rect 12173 20009 12207 20043
rect 13829 20009 13863 20043
rect 15669 20009 15703 20043
rect 16405 20009 16439 20043
rect 16865 20009 16899 20043
rect 20177 20009 20211 20043
rect 22845 20009 22879 20043
rect 23489 20009 23523 20043
rect 23949 20009 23983 20043
rect 25605 20009 25639 20043
rect 26341 20009 26375 20043
rect 26433 20009 26467 20043
rect 36737 20009 36771 20043
rect 5089 19941 5123 19975
rect 10425 19941 10459 19975
rect 11989 19941 12023 19975
rect 12909 19941 12943 19975
rect 16681 19941 16715 19975
rect 24133 19941 24167 19975
rect 31677 19941 31711 19975
rect 2881 19873 2915 19907
rect 4445 19873 4479 19907
rect 4813 19873 4847 19907
rect 5733 19873 5767 19907
rect 13277 19873 13311 19907
rect 19533 19873 19567 19907
rect 20269 19873 20303 19907
rect 23029 19873 23063 19907
rect 23857 19873 23891 19907
rect 24869 19873 24903 19907
rect 25697 19873 25731 19907
rect 26157 19873 26191 19907
rect 31217 19873 31251 19907
rect 32045 19873 32079 19907
rect 32321 19873 32355 19907
rect 36093 19873 36127 19907
rect 36461 19873 36495 19907
rect 1961 19805 1995 19839
rect 3341 19805 3375 19839
rect 3985 19805 4019 19839
rect 4077 19805 4111 19839
rect 4721 19805 4755 19839
rect 5549 19805 5583 19839
rect 6193 19805 6227 19839
rect 6285 19805 6319 19839
rect 6561 19805 6595 19839
rect 6653 19805 6687 19839
rect 9229 19805 9263 19839
rect 9505 19805 9539 19839
rect 9597 19805 9631 19839
rect 9873 19805 9907 19839
rect 10057 19805 10091 19839
rect 10149 19805 10183 19839
rect 10241 19805 10275 19839
rect 12265 19805 12299 19839
rect 13185 19805 13219 19839
rect 13553 19805 13587 19839
rect 13645 19805 13679 19839
rect 14105 19805 14139 19839
rect 14473 19805 14507 19839
rect 14565 19805 14599 19839
rect 15209 19805 15243 19839
rect 15301 19805 15335 19839
rect 15708 19805 15742 19839
rect 16313 19805 16347 19839
rect 16497 19805 16531 19839
rect 16957 19805 16991 19839
rect 17417 19805 17451 19839
rect 17877 19805 17911 19839
rect 18153 19805 18187 19839
rect 18705 19805 18739 19839
rect 18889 19805 18923 19839
rect 18981 19805 19015 19839
rect 19625 19805 19659 19839
rect 19901 19805 19935 19839
rect 19993 19805 20027 19839
rect 20545 19805 20579 19839
rect 20637 19805 20671 19839
rect 20729 19805 20763 19839
rect 20913 19805 20947 19839
rect 23121 19805 23155 19839
rect 23673 19805 23707 19839
rect 24041 19805 24075 19839
rect 24225 19805 24259 19839
rect 24409 19805 24443 19839
rect 24593 19805 24627 19839
rect 24777 19805 24811 19839
rect 24961 19805 24995 19839
rect 25053 19805 25087 19839
rect 25421 19805 25455 19839
rect 26065 19805 26099 19839
rect 26617 19805 26651 19839
rect 26709 19805 26743 19839
rect 26985 19805 27019 19839
rect 28457 19805 28491 19839
rect 28641 19805 28675 19839
rect 28825 19805 28859 19839
rect 28917 19805 28951 19839
rect 29009 19805 29043 19839
rect 29193 19805 29227 19839
rect 29745 19805 29779 19839
rect 29837 19805 29871 19839
rect 30021 19805 30055 19839
rect 30113 19805 30147 19839
rect 30389 19805 30423 19839
rect 30665 19805 30699 19839
rect 31493 19805 31527 19839
rect 31953 19805 31987 19839
rect 33425 19805 33459 19839
rect 33609 19805 33643 19839
rect 35081 19805 35115 19839
rect 35173 19805 35207 19839
rect 35357 19805 35391 19839
rect 35449 19805 35483 19839
rect 36001 19805 36035 19839
rect 36369 19805 36403 19839
rect 36553 19805 36587 19839
rect 36645 19805 36679 19839
rect 4169 19737 4203 19771
rect 4307 19737 4341 19771
rect 6377 19737 6411 19771
rect 6929 19737 6963 19771
rect 9413 19737 9447 19771
rect 11621 19737 11655 19771
rect 13461 19737 13495 19771
rect 22845 19737 22879 19771
rect 23949 19737 23983 19771
rect 25237 19737 25271 19771
rect 25329 19737 25363 19771
rect 26801 19737 26835 19771
rect 28549 19737 28583 19771
rect 34897 19737 34931 19771
rect 1777 19669 1811 19703
rect 5181 19669 5215 19703
rect 5641 19669 5675 19703
rect 6009 19669 6043 19703
rect 8401 19669 8435 19703
rect 11437 19669 11471 19703
rect 12725 19669 12759 19703
rect 15853 19669 15887 19703
rect 23305 19669 23339 19703
rect 24409 19669 24443 19703
rect 29193 19669 29227 19703
rect 29561 19669 29595 19703
rect 33517 19669 33551 19703
rect 35541 19669 35575 19703
rect 35909 19669 35943 19703
rect 5917 19465 5951 19499
rect 7021 19465 7055 19499
rect 9321 19465 9355 19499
rect 12357 19465 12391 19499
rect 13185 19465 13219 19499
rect 19809 19465 19843 19499
rect 22661 19465 22695 19499
rect 27813 19465 27847 19499
rect 30205 19465 30239 19499
rect 33793 19465 33827 19499
rect 33977 19465 34011 19499
rect 36001 19465 36035 19499
rect 1685 19397 1719 19431
rect 8953 19397 8987 19431
rect 13001 19397 13035 19431
rect 22201 19397 22235 19431
rect 33333 19397 33367 19431
rect 1409 19329 1443 19363
rect 3525 19329 3559 19363
rect 3709 19329 3743 19363
rect 4169 19329 4203 19363
rect 7205 19329 7239 19363
rect 7941 19329 7975 19363
rect 8769 19329 8803 19363
rect 9045 19329 9079 19363
rect 9137 19329 9171 19363
rect 9597 19329 9631 19363
rect 9781 19329 9815 19363
rect 11161 19329 11195 19363
rect 11345 19329 11379 19363
rect 11529 19329 11563 19363
rect 11989 19329 12023 19363
rect 12541 19329 12575 19363
rect 12633 19329 12667 19363
rect 13369 19329 13403 19363
rect 14381 19329 14415 19363
rect 14565 19329 14599 19363
rect 14749 19329 14783 19363
rect 16681 19329 16715 19363
rect 17141 19329 17175 19363
rect 17601 19329 17635 19363
rect 18153 19329 18187 19363
rect 19717 19329 19751 19363
rect 19901 19329 19935 19363
rect 22385 19329 22419 19363
rect 22477 19329 22511 19363
rect 22753 19329 22787 19363
rect 23581 19329 23615 19363
rect 24041 19329 24075 19363
rect 27261 19329 27295 19363
rect 27445 19329 27479 19363
rect 27537 19329 27571 19363
rect 27629 19329 27663 19363
rect 27905 19329 27939 19363
rect 28181 19329 28215 19363
rect 28273 19329 28307 19363
rect 29009 19329 29043 19363
rect 29193 19329 29227 19363
rect 29285 19329 29319 19363
rect 29469 19329 29503 19363
rect 29745 19329 29779 19363
rect 29837 19329 29871 19363
rect 30021 19329 30055 19363
rect 30205 19329 30239 19363
rect 32965 19329 32999 19363
rect 33149 19329 33183 19363
rect 33885 19329 33919 19363
rect 34161 19329 34195 19363
rect 34253 19329 34287 19363
rect 34437 19329 34471 19363
rect 34713 19329 34747 19363
rect 34897 19329 34931 19363
rect 35817 19329 35851 19363
rect 36001 19329 36035 19363
rect 3893 19261 3927 19295
rect 4445 19261 4479 19295
rect 8309 19261 8343 19295
rect 9413 19261 9447 19295
rect 11897 19261 11931 19295
rect 13553 19261 13587 19295
rect 16773 19261 16807 19295
rect 18245 19261 18279 19295
rect 23857 19261 23891 19295
rect 24317 19261 24351 19295
rect 29377 19261 29411 19295
rect 34805 19261 34839 19295
rect 3157 19193 3191 19227
rect 11713 19193 11747 19227
rect 14657 19193 14691 19227
rect 33609 19193 33643 19227
rect 11345 19125 11379 19159
rect 11805 19125 11839 19159
rect 12265 19125 12299 19159
rect 12909 19125 12943 19159
rect 22201 19125 22235 19159
rect 24225 19125 24259 19159
rect 29653 19125 29687 19159
rect 33149 19125 33183 19159
rect 34621 19125 34655 19159
rect 4721 18921 4755 18955
rect 19809 18921 19843 18955
rect 20821 18921 20855 18955
rect 21005 18921 21039 18955
rect 22569 18921 22603 18955
rect 32965 18921 32999 18955
rect 17877 18853 17911 18887
rect 18337 18853 18371 18887
rect 22017 18853 22051 18887
rect 33609 18853 33643 18887
rect 3341 18785 3375 18819
rect 5733 18785 5767 18819
rect 10885 18785 10919 18819
rect 19349 18785 19383 18819
rect 20177 18785 20211 18819
rect 20453 18785 20487 18819
rect 21833 18785 21867 18819
rect 22661 18785 22695 18819
rect 36737 18785 36771 18819
rect 3065 18717 3099 18751
rect 4905 18717 4939 18751
rect 6009 18717 6043 18751
rect 6101 18717 6135 18751
rect 10793 18717 10827 18751
rect 11805 18717 11839 18751
rect 11897 18717 11931 18751
rect 11989 18717 12023 18751
rect 12173 18717 12207 18751
rect 17693 18717 17727 18751
rect 17969 18717 18003 18751
rect 18061 18717 18095 18751
rect 18245 18717 18279 18751
rect 18521 18717 18555 18751
rect 18613 18717 18647 18751
rect 19257 18717 19291 18751
rect 19533 18717 19567 18751
rect 19625 18717 19659 18751
rect 19998 18717 20032 18751
rect 20545 18717 20579 18751
rect 21557 18717 21591 18751
rect 21649 18717 21683 18751
rect 22385 18717 22419 18751
rect 31033 18717 31067 18751
rect 31217 18717 31251 18751
rect 31401 18717 31435 18751
rect 31585 18717 31619 18751
rect 32413 18717 32447 18751
rect 32505 18717 32539 18751
rect 32689 18717 32723 18751
rect 32781 18717 32815 18751
rect 33701 18717 33735 18751
rect 34989 18717 35023 18751
rect 36921 18717 36955 18751
rect 1409 18649 1443 18683
rect 1777 18649 1811 18683
rect 5641 18649 5675 18683
rect 10701 18649 10735 18683
rect 11529 18649 11563 18683
rect 14381 18649 14415 18683
rect 14565 18649 14599 18683
rect 18337 18649 18371 18683
rect 21189 18649 21223 18683
rect 31493 18649 31527 18683
rect 34713 18649 34747 18683
rect 2697 18581 2731 18615
rect 3157 18581 3191 18615
rect 6285 18581 6319 18615
rect 10333 18581 10367 18615
rect 14197 18581 14231 18615
rect 17509 18581 17543 18615
rect 18061 18581 18095 18615
rect 20979 18581 21013 18615
rect 22201 18581 22235 18615
rect 31217 18581 31251 18615
rect 34811 18581 34845 18615
rect 34897 18581 34931 18615
rect 37105 18581 37139 18615
rect 13921 18377 13955 18411
rect 15393 18377 15427 18411
rect 19901 18377 19935 18411
rect 25605 18377 25639 18411
rect 32781 18377 32815 18411
rect 34253 18377 34287 18411
rect 4353 18309 4387 18343
rect 9505 18309 9539 18343
rect 12081 18309 12115 18343
rect 15025 18309 15059 18343
rect 25237 18309 25271 18343
rect 31033 18309 31067 18343
rect 32137 18309 32171 18343
rect 32965 18309 32999 18343
rect 33149 18309 33183 18343
rect 37565 18309 37599 18343
rect 1869 18241 1903 18275
rect 2329 18241 2363 18275
rect 6193 18241 6227 18275
rect 11529 18241 11563 18275
rect 11713 18241 11747 18275
rect 12357 18241 12391 18275
rect 12541 18241 12575 18275
rect 14105 18241 14139 18275
rect 14289 18241 14323 18275
rect 14473 18241 14507 18275
rect 15669 18241 15703 18275
rect 16773 18241 16807 18275
rect 17141 18241 17175 18275
rect 18797 18241 18831 18275
rect 18889 18241 18923 18275
rect 19199 18241 19233 18275
rect 19533 18241 19567 18275
rect 19687 18241 19721 18275
rect 22477 18241 22511 18275
rect 22753 18241 22787 18275
rect 23305 18241 23339 18275
rect 25053 18241 25087 18275
rect 25329 18241 25363 18275
rect 25421 18241 25455 18275
rect 25881 18241 25915 18275
rect 27997 18241 28031 18275
rect 28181 18241 28215 18275
rect 29561 18241 29595 18275
rect 29745 18241 29779 18275
rect 30389 18241 30423 18275
rect 30665 18241 30699 18275
rect 31217 18241 31251 18275
rect 31401 18241 31435 18275
rect 31493 18241 31527 18275
rect 31677 18241 31711 18275
rect 32873 18241 32907 18275
rect 34345 18241 34379 18275
rect 34805 18241 34839 18275
rect 34989 18241 35023 18275
rect 35173 18241 35207 18275
rect 36921 18241 36955 18275
rect 1685 18173 1719 18207
rect 2145 18173 2179 18207
rect 5917 18173 5951 18207
rect 7573 18173 7607 18207
rect 7849 18173 7883 18207
rect 9321 18173 9355 18207
rect 12173 18173 12207 18207
rect 15577 18173 15611 18207
rect 16037 18173 16071 18207
rect 22937 18173 22971 18207
rect 25789 18173 25823 18207
rect 30481 18173 30515 18207
rect 31861 18173 31895 18207
rect 32505 18173 32539 18207
rect 32597 18173 32631 18207
rect 34069 18173 34103 18207
rect 10793 18105 10827 18139
rect 11713 18105 11747 18139
rect 19441 18105 19475 18139
rect 23581 18105 23615 18139
rect 26249 18105 26283 18139
rect 33149 18105 33183 18139
rect 34713 18105 34747 18139
rect 2053 18037 2087 18071
rect 2513 18037 2547 18071
rect 3065 18037 3099 18071
rect 18429 18037 18463 18071
rect 19257 18037 19291 18071
rect 28089 18037 28123 18071
rect 29561 18037 29595 18071
rect 34897 18037 34931 18071
rect 37105 18037 37139 18071
rect 37841 18037 37875 18071
rect 2053 17833 2087 17867
rect 2973 17833 3007 17867
rect 7849 17833 7883 17867
rect 8033 17833 8067 17867
rect 11345 17833 11379 17867
rect 12449 17833 12483 17867
rect 12817 17833 12851 17867
rect 13093 17833 13127 17867
rect 15301 17833 15335 17867
rect 17693 17833 17727 17867
rect 20637 17833 20671 17867
rect 22937 17833 22971 17867
rect 27353 17833 27387 17867
rect 31309 17833 31343 17867
rect 32137 17833 32171 17867
rect 8953 17765 8987 17799
rect 11253 17765 11287 17799
rect 16037 17765 16071 17799
rect 23949 17765 23983 17799
rect 25605 17765 25639 17799
rect 26617 17765 26651 17799
rect 34069 17765 34103 17799
rect 1593 17697 1627 17731
rect 3985 17697 4019 17731
rect 9413 17697 9447 17731
rect 9505 17697 9539 17731
rect 10057 17697 10091 17731
rect 10885 17697 10919 17731
rect 11989 17697 12023 17731
rect 15485 17697 15519 17731
rect 23489 17697 23523 17731
rect 24685 17697 24719 17731
rect 24961 17697 24995 17731
rect 25145 17697 25179 17731
rect 26341 17697 26375 17731
rect 26985 17697 27019 17731
rect 27721 17697 27755 17731
rect 1777 17629 1811 17663
rect 2237 17629 2271 17663
rect 3249 17629 3283 17663
rect 3341 17629 3375 17663
rect 3433 17629 3467 17663
rect 3617 17629 3651 17663
rect 6101 17629 6135 17663
rect 8217 17629 8251 17663
rect 10149 17629 10183 17663
rect 10425 17629 10459 17663
rect 11069 17629 11103 17663
rect 11253 17629 11287 17663
rect 11805 17629 11839 17663
rect 12449 17629 12483 17663
rect 12633 17629 12667 17663
rect 12725 17629 12759 17663
rect 12902 17629 12936 17663
rect 13001 17631 13035 17665
rect 13185 17629 13219 17663
rect 13737 17629 13771 17663
rect 13921 17629 13955 17663
rect 14289 17629 14323 17663
rect 15577 17629 15611 17663
rect 15853 17629 15887 17663
rect 16313 17629 16347 17663
rect 16405 17629 16439 17663
rect 16497 17629 16531 17663
rect 16681 17629 16715 17663
rect 17417 17629 17451 17663
rect 17509 17629 17543 17663
rect 17877 17629 17911 17663
rect 18061 17629 18095 17663
rect 18153 17629 18187 17663
rect 18245 17629 18279 17663
rect 18429 17629 18463 17663
rect 18797 17629 18831 17663
rect 18981 17629 19015 17663
rect 20361 17629 20395 17663
rect 22293 17629 22327 17663
rect 22477 17629 22511 17663
rect 22569 17629 22603 17663
rect 22661 17629 22695 17663
rect 23581 17629 23615 17663
rect 24593 17629 24627 17663
rect 25237 17629 25271 17663
rect 26249 17629 26283 17663
rect 27077 17629 27111 17663
rect 27905 17629 27939 17663
rect 28365 17629 28399 17663
rect 28549 17629 28583 17663
rect 29009 17629 29043 17663
rect 29561 17629 29595 17663
rect 29745 17629 29779 17663
rect 29837 17629 29871 17663
rect 29929 17629 29963 17663
rect 30297 17629 30331 17663
rect 30481 17629 30515 17663
rect 31217 17629 31251 17663
rect 32045 17629 32079 17663
rect 33793 17629 33827 17663
rect 34069 17629 34103 17663
rect 4261 17561 4295 17595
rect 6377 17561 6411 17595
rect 11713 17561 11747 17595
rect 14657 17561 14691 17595
rect 15945 17561 15979 17595
rect 20545 17561 20579 17595
rect 1961 17493 1995 17527
rect 5733 17493 5767 17527
rect 9321 17493 9355 17527
rect 12265 17493 12299 17527
rect 13645 17493 13679 17527
rect 18613 17493 18647 17527
rect 18889 17493 18923 17527
rect 30205 17493 30239 17527
rect 30389 17493 30423 17527
rect 33885 17493 33919 17527
rect 3433 17289 3467 17323
rect 4261 17289 4295 17323
rect 4537 17289 4571 17323
rect 6561 17289 6595 17323
rect 6929 17289 6963 17323
rect 7389 17289 7423 17323
rect 11989 17289 12023 17323
rect 12357 17289 12391 17323
rect 14013 17289 14047 17323
rect 28174 17289 28208 17323
rect 28365 17289 28399 17323
rect 28533 17289 28567 17323
rect 29193 17289 29227 17323
rect 33149 17289 33183 17323
rect 33993 17289 34027 17323
rect 34161 17289 34195 17323
rect 3065 17221 3099 17255
rect 4905 17221 4939 17255
rect 5917 17221 5951 17255
rect 9965 17221 9999 17255
rect 19901 17221 19935 17255
rect 28733 17221 28767 17255
rect 31677 17221 31711 17255
rect 31861 17221 31895 17255
rect 33793 17221 33827 17255
rect 3249 17153 3283 17187
rect 4445 17153 4479 17187
rect 4997 17153 5031 17187
rect 5733 17153 5767 17187
rect 6745 17153 6779 17187
rect 7297 17153 7331 17187
rect 8953 17153 8987 17187
rect 9137 17153 9171 17187
rect 10240 17153 10274 17187
rect 10333 17153 10367 17187
rect 10425 17153 10459 17187
rect 10609 17153 10643 17187
rect 11989 17153 12023 17187
rect 12173 17153 12207 17187
rect 12265 17153 12299 17187
rect 12449 17153 12483 17187
rect 16681 17153 16715 17187
rect 16865 17153 16899 17187
rect 19625 17153 19659 17187
rect 19718 17153 19752 17187
rect 19993 17153 20027 17187
rect 20090 17153 20124 17187
rect 20637 17153 20671 17187
rect 20729 17153 20763 17187
rect 20821 17153 20855 17187
rect 21005 17153 21039 17187
rect 22385 17153 22419 17187
rect 22937 17153 22971 17187
rect 23489 17153 23523 17187
rect 27997 17153 28031 17187
rect 28089 17153 28123 17187
rect 28273 17153 28307 17187
rect 29009 17153 29043 17187
rect 29193 17153 29227 17187
rect 29561 17153 29595 17187
rect 31953 17153 31987 17187
rect 32873 17153 32907 17187
rect 33057 17153 33091 17187
rect 34437 17153 34471 17187
rect 34897 17153 34931 17187
rect 5089 17085 5123 17119
rect 7573 17085 7607 17119
rect 14473 17085 14507 17119
rect 20361 17085 20395 17119
rect 22477 17085 22511 17119
rect 32321 17085 32355 17119
rect 32413 17085 32447 17119
rect 32505 17085 32539 17119
rect 32597 17085 32631 17119
rect 32781 17085 32815 17119
rect 34529 17085 34563 17119
rect 34989 17085 35023 17119
rect 35173 17085 35207 17119
rect 14197 17017 14231 17051
rect 31677 17017 31711 17051
rect 6101 16949 6135 16983
rect 9321 16949 9355 16983
rect 16681 16949 16715 16983
rect 17049 16949 17083 16983
rect 20269 16949 20303 16983
rect 22753 16949 22787 16983
rect 28549 16949 28583 16983
rect 33977 16949 34011 16983
rect 34437 16949 34471 16983
rect 34805 16949 34839 16983
rect 35081 16949 35115 16983
rect 16497 16745 16531 16779
rect 16681 16745 16715 16779
rect 30113 16745 30147 16779
rect 31217 16745 31251 16779
rect 32137 16745 32171 16779
rect 35173 16745 35207 16779
rect 35449 16745 35483 16779
rect 3801 16677 3835 16711
rect 8401 16677 8435 16711
rect 34345 16677 34379 16711
rect 34437 16677 34471 16711
rect 35357 16677 35391 16711
rect 2789 16609 2823 16643
rect 2973 16609 3007 16643
rect 4445 16609 4479 16643
rect 9137 16609 9171 16643
rect 16129 16609 16163 16643
rect 16773 16609 16807 16643
rect 17693 16609 17727 16643
rect 23213 16609 23247 16643
rect 23505 16609 23539 16643
rect 23949 16609 23983 16643
rect 25605 16609 25639 16643
rect 34253 16609 34287 16643
rect 35541 16609 35575 16643
rect 1961 16541 1995 16575
rect 2237 16541 2271 16575
rect 3985 16541 4019 16575
rect 4169 16541 4203 16575
rect 4537 16541 4571 16575
rect 8585 16541 8619 16575
rect 8769 16541 8803 16575
rect 14197 16541 14231 16575
rect 15025 16541 15059 16575
rect 16957 16541 16991 16575
rect 17233 16541 17267 16575
rect 17969 16541 18003 16575
rect 18153 16541 18187 16575
rect 18337 16541 18371 16575
rect 18613 16541 18647 16575
rect 20269 16541 20303 16575
rect 20362 16541 20396 16575
rect 20775 16541 20809 16575
rect 21005 16541 21039 16575
rect 21373 16541 21407 16575
rect 21833 16541 21867 16575
rect 22293 16541 22327 16575
rect 23421 16541 23455 16575
rect 25237 16541 25271 16575
rect 25421 16541 25455 16575
rect 26065 16541 26099 16575
rect 30021 16541 30055 16575
rect 30205 16541 30239 16575
rect 30573 16541 30607 16575
rect 30757 16541 30791 16575
rect 31401 16541 31435 16575
rect 32321 16541 32355 16575
rect 34529 16541 34563 16575
rect 35449 16541 35483 16575
rect 4077 16473 4111 16507
rect 4307 16473 4341 16507
rect 9413 16473 9447 16507
rect 19073 16473 19107 16507
rect 20545 16473 20579 16507
rect 20637 16473 20671 16507
rect 22109 16473 22143 16507
rect 22845 16473 22879 16507
rect 23765 16473 23799 16507
rect 26249 16473 26283 16507
rect 32505 16473 32539 16507
rect 34989 16473 35023 16507
rect 1777 16405 1811 16439
rect 2053 16405 2087 16439
rect 2329 16405 2363 16439
rect 2697 16405 2731 16439
rect 4629 16405 4663 16439
rect 10885 16405 10919 16439
rect 16497 16405 16531 16439
rect 17141 16405 17175 16439
rect 20913 16405 20947 16439
rect 23305 16405 23339 16439
rect 26433 16405 26467 16439
rect 30757 16405 30791 16439
rect 35189 16405 35223 16439
rect 35817 16405 35851 16439
rect 3893 16201 3927 16235
rect 4061 16201 4095 16235
rect 5181 16201 5215 16235
rect 9505 16201 9539 16235
rect 9781 16201 9815 16235
rect 10149 16201 10183 16235
rect 14289 16201 14323 16235
rect 16865 16201 16899 16235
rect 17049 16201 17083 16235
rect 20729 16201 20763 16235
rect 21465 16201 21499 16235
rect 29285 16201 29319 16235
rect 30481 16201 30515 16235
rect 30849 16201 30883 16235
rect 34989 16201 35023 16235
rect 1685 16133 1719 16167
rect 4261 16133 4295 16167
rect 10241 16133 10275 16167
rect 17233 16133 17267 16167
rect 17509 16133 17543 16167
rect 17709 16133 17743 16167
rect 18797 16133 18831 16167
rect 20177 16133 20211 16167
rect 20361 16133 20395 16167
rect 20561 16133 20595 16167
rect 23029 16133 23063 16167
rect 29377 16133 29411 16167
rect 31033 16133 31067 16167
rect 31217 16133 31251 16167
rect 5549 16065 5583 16099
rect 9689 16065 9723 16099
rect 12265 16065 12299 16099
rect 12357 16065 12391 16099
rect 14473 16065 14507 16099
rect 14749 16065 14783 16099
rect 16957 16065 16991 16099
rect 17969 16065 18003 16099
rect 18153 16065 18187 16099
rect 18245 16065 18279 16099
rect 18337 16065 18371 16099
rect 20269 16065 20303 16099
rect 21281 16065 21315 16099
rect 22845 16065 22879 16099
rect 23121 16065 23155 16099
rect 23213 16065 23247 16099
rect 24685 16065 24719 16099
rect 25237 16065 25271 16099
rect 26249 16065 26283 16099
rect 26341 16065 26375 16099
rect 27077 16065 27111 16099
rect 27169 16065 27203 16099
rect 27353 16065 27387 16099
rect 29101 16065 29135 16099
rect 29285 16065 29319 16099
rect 29561 16065 29595 16099
rect 30113 16065 30147 16099
rect 30665 16065 30699 16099
rect 30941 16065 30975 16099
rect 34897 16065 34931 16099
rect 35173 16065 35207 16099
rect 37657 16065 37691 16099
rect 1409 15997 1443 16031
rect 5641 15997 5675 16031
rect 5825 15997 5859 16031
rect 10333 15997 10367 16031
rect 12541 15997 12575 16031
rect 14657 15997 14691 16031
rect 21005 15997 21039 16031
rect 26525 15997 26559 16031
rect 27261 15997 27295 16031
rect 29745 15997 29779 16031
rect 29929 15997 29963 16031
rect 11897 15929 11931 15963
rect 17877 15929 17911 15963
rect 35173 15929 35207 15963
rect 3157 15861 3191 15895
rect 4077 15861 4111 15895
rect 16681 15861 16715 15895
rect 17693 15861 17727 15895
rect 18613 15861 18647 15895
rect 18889 15861 18923 15895
rect 20545 15861 20579 15895
rect 21097 15861 21131 15895
rect 23397 15861 23431 15895
rect 26065 15861 26099 15895
rect 27537 15861 27571 15895
rect 30297 15861 30331 15895
rect 31401 15861 31435 15895
rect 37841 15861 37875 15895
rect 1501 15657 1535 15691
rect 3801 15657 3835 15691
rect 4997 15657 5031 15691
rect 7941 15657 7975 15691
rect 10241 15657 10275 15691
rect 14289 15657 14323 15691
rect 14749 15657 14783 15691
rect 18153 15657 18187 15691
rect 20821 15657 20855 15691
rect 26341 15657 26375 15691
rect 32321 15657 32355 15691
rect 32781 15657 32815 15691
rect 33241 15657 33275 15691
rect 35173 15657 35207 15691
rect 35449 15657 35483 15691
rect 18981 15589 19015 15623
rect 32413 15589 32447 15623
rect 4077 15521 4111 15555
rect 4537 15521 4571 15555
rect 6193 15521 6227 15555
rect 11529 15521 11563 15555
rect 15485 15521 15519 15555
rect 15669 15521 15703 15555
rect 16221 15521 16255 15555
rect 18797 15521 18831 15555
rect 20637 15521 20671 15555
rect 27721 15521 27755 15555
rect 27997 15521 28031 15555
rect 31861 15521 31895 15555
rect 32229 15521 32263 15555
rect 33333 15521 33367 15555
rect 34805 15521 34839 15555
rect 35633 15521 35667 15555
rect 1777 15453 1811 15487
rect 3985 15453 4019 15487
rect 4169 15453 4203 15487
rect 4261 15453 4295 15487
rect 4629 15453 4663 15487
rect 8953 15453 8987 15487
rect 11437 15453 11471 15487
rect 11897 15453 11931 15487
rect 13921 15453 13955 15487
rect 14197 15453 14231 15487
rect 14565 15453 14599 15487
rect 15761 15453 15795 15487
rect 15853 15453 15887 15487
rect 15945 15453 15979 15487
rect 16129 15453 16163 15487
rect 16313 15453 16347 15487
rect 18245 15453 18279 15487
rect 19074 15453 19108 15487
rect 19349 15453 19383 15487
rect 19993 15453 20027 15487
rect 20729 15453 20763 15487
rect 22937 15453 22971 15487
rect 23121 15453 23155 15487
rect 23397 15453 23431 15487
rect 23673 15453 23707 15487
rect 23765 15453 23799 15487
rect 24501 15453 24535 15487
rect 24777 15453 24811 15487
rect 24961 15453 24995 15487
rect 25237 15453 25271 15487
rect 25421 15453 25455 15487
rect 25973 15453 26007 15487
rect 26157 15453 26191 15487
rect 26433 15453 26467 15487
rect 27629 15453 27663 15487
rect 28181 15453 28215 15487
rect 28457 15453 28491 15487
rect 28641 15453 28675 15487
rect 28733 15453 28767 15487
rect 29653 15453 29687 15487
rect 29837 15453 29871 15487
rect 31493 15453 31527 15487
rect 31677 15453 31711 15487
rect 32505 15453 32539 15487
rect 33425 15453 33459 15487
rect 34897 15453 34931 15487
rect 35725 15453 35759 15487
rect 6469 15385 6503 15419
rect 11345 15385 11379 15419
rect 12173 15385 12207 15419
rect 18429 15385 18463 15419
rect 32749 15385 32783 15419
rect 32965 15385 32999 15419
rect 10977 15317 11011 15351
rect 18613 15317 18647 15351
rect 25605 15317 25639 15351
rect 26617 15317 26651 15351
rect 27261 15317 27295 15351
rect 28365 15317 28399 15351
rect 30665 15317 30699 15351
rect 32597 15317 32631 15351
rect 33057 15317 33091 15351
rect 2973 15113 3007 15147
rect 3709 15113 3743 15147
rect 4077 15113 4111 15147
rect 6653 15113 6687 15147
rect 7573 15113 7607 15147
rect 13921 15113 13955 15147
rect 15761 15113 15795 15147
rect 20177 15113 20211 15147
rect 27077 15113 27111 15147
rect 34345 15113 34379 15147
rect 4905 15045 4939 15079
rect 9045 15045 9079 15079
rect 11897 15045 11931 15079
rect 11989 15045 12023 15079
rect 14749 15045 14783 15079
rect 15025 15045 15059 15079
rect 29009 15045 29043 15079
rect 2881 14977 2915 15011
rect 3433 14977 3467 15011
rect 3617 14977 3651 15011
rect 4721 14977 4755 15011
rect 6837 14977 6871 15011
rect 7481 14977 7515 15011
rect 8033 14977 8067 15011
rect 8125 14977 8159 15011
rect 8401 14977 8435 15011
rect 10517 14977 10551 15011
rect 13001 14977 13035 15011
rect 13369 14977 13403 15011
rect 14105 14977 14139 15011
rect 14197 14977 14231 15011
rect 14289 14977 14323 15011
rect 14473 14977 14507 15011
rect 14565 14977 14599 15011
rect 14841 14977 14875 15011
rect 15117 14977 15151 15011
rect 15393 14977 15427 15011
rect 15577 14977 15611 15011
rect 16221 14977 16255 15011
rect 16497 14977 16531 15011
rect 16773 14977 16807 15011
rect 17049 14977 17083 15011
rect 17141 14977 17175 15011
rect 17601 14977 17635 15011
rect 17693 14977 17727 15011
rect 18245 14977 18279 15011
rect 18797 14977 18831 15011
rect 19165 14977 19199 15011
rect 19625 14977 19659 15011
rect 20085 14977 20119 15011
rect 20361 14977 20395 15011
rect 22017 14977 22051 15011
rect 22201 14977 22235 15011
rect 22661 14977 22695 15011
rect 25513 14977 25547 15011
rect 25697 14977 25731 15011
rect 25789 14977 25823 15011
rect 25973 14977 26007 15011
rect 26985 14977 27019 15011
rect 27261 14977 27295 15011
rect 27813 14977 27847 15011
rect 27905 14977 27939 15011
rect 28089 14977 28123 15011
rect 28273 14977 28307 15011
rect 28457 14977 28491 15011
rect 28549 14977 28583 15011
rect 28825 14977 28859 15011
rect 30665 14977 30699 15011
rect 30757 14977 30791 15011
rect 30849 14977 30883 15011
rect 30941 14977 30975 15011
rect 31125 14977 31159 15011
rect 33057 14977 33091 15011
rect 33977 14977 34011 15011
rect 3157 14909 3191 14943
rect 4169 14909 4203 14943
rect 4261 14909 4295 14943
rect 4537 14909 4571 14943
rect 7665 14909 7699 14943
rect 9505 14909 9539 14943
rect 9597 14909 9631 14943
rect 12173 14909 12207 14943
rect 18705 14909 18739 14943
rect 21833 14909 21867 14943
rect 23213 14909 23247 14943
rect 28641 14909 28675 14943
rect 32965 14909 32999 14943
rect 33885 14909 33919 14943
rect 7113 14841 7147 14875
rect 9045 14841 9079 14875
rect 11529 14841 11563 14875
rect 14841 14841 14875 14875
rect 15945 14841 15979 14875
rect 27445 14841 27479 14875
rect 27997 14841 28031 14875
rect 33425 14841 33459 14875
rect 2513 14773 2547 14807
rect 3617 14773 3651 14807
rect 8309 14773 8343 14807
rect 8677 14773 8711 14807
rect 8861 14773 8895 14807
rect 9781 14773 9815 14807
rect 10333 14773 10367 14807
rect 13553 14773 13587 14807
rect 16405 14773 16439 14807
rect 20545 14773 20579 14807
rect 25605 14773 25639 14807
rect 25973 14773 26007 14807
rect 27629 14773 27663 14807
rect 31033 14773 31067 14807
rect 3157 14569 3191 14603
rect 4077 14569 4111 14603
rect 7389 14569 7423 14603
rect 13461 14569 13495 14603
rect 16589 14569 16623 14603
rect 17049 14569 17083 14603
rect 17417 14569 17451 14603
rect 19625 14569 19659 14603
rect 31953 14569 31987 14603
rect 23121 14501 23155 14535
rect 10149 14433 10183 14467
rect 11897 14433 11931 14467
rect 12817 14433 12851 14467
rect 13001 14433 13035 14467
rect 15485 14433 15519 14467
rect 21005 14433 21039 14467
rect 21649 14433 21683 14467
rect 23305 14433 23339 14467
rect 23397 14433 23431 14467
rect 31585 14433 31619 14467
rect 1409 14365 1443 14399
rect 4077 14365 4111 14399
rect 4261 14365 4295 14399
rect 5641 14365 5675 14399
rect 8953 14365 8987 14399
rect 9137 14365 9171 14399
rect 9229 14365 9263 14399
rect 9321 14365 9355 14399
rect 9873 14365 9907 14399
rect 15301 14365 15335 14399
rect 16589 14365 16623 14399
rect 16773 14365 16807 14399
rect 17049 14365 17083 14399
rect 17233 14365 17267 14399
rect 17325 14365 17359 14399
rect 17969 14365 18003 14399
rect 18153 14365 18187 14399
rect 19257 14365 19291 14399
rect 19901 14365 19935 14399
rect 20545 14365 20579 14399
rect 20821 14365 20855 14399
rect 21281 14365 21315 14399
rect 22017 14365 22051 14399
rect 22661 14365 22695 14399
rect 23581 14365 23615 14399
rect 30297 14365 30331 14399
rect 30389 14365 30423 14399
rect 31217 14365 31251 14399
rect 31401 14365 31435 14399
rect 31493 14365 31527 14399
rect 31769 14365 31803 14399
rect 1685 14297 1719 14331
rect 5917 14297 5951 14331
rect 9597 14297 9631 14331
rect 18061 14297 18095 14331
rect 30573 14297 30607 14331
rect 30665 14297 30699 14331
rect 30849 14297 30883 14331
rect 13093 14229 13127 14263
rect 19634 14229 19668 14263
rect 23765 14229 23799 14263
rect 31033 14229 31067 14263
rect 1961 14025 1995 14059
rect 6377 14025 6411 14059
rect 6653 14025 6687 14059
rect 7021 14025 7055 14059
rect 8677 14025 8711 14059
rect 17785 14025 17819 14059
rect 17877 14025 17911 14059
rect 19809 14025 19843 14059
rect 23489 14025 23523 14059
rect 29101 14025 29135 14059
rect 31401 14025 31435 14059
rect 32873 14025 32907 14059
rect 7113 13957 7147 13991
rect 17233 13957 17267 13991
rect 22845 13957 22879 13991
rect 25421 13957 25455 13991
rect 26433 13957 26467 13991
rect 1777 13889 1811 13923
rect 2145 13889 2179 13923
rect 6561 13889 6595 13923
rect 8401 13889 8435 13923
rect 8493 13889 8527 13923
rect 14657 13889 14691 13923
rect 15301 13889 15335 13923
rect 16221 13889 16255 13923
rect 16681 13889 16715 13923
rect 16773 13889 16807 13923
rect 19717 13889 19751 13923
rect 20269 13889 20303 13923
rect 20637 13889 20671 13923
rect 20913 13889 20947 13923
rect 21097 13889 21131 13923
rect 21189 13889 21223 13923
rect 21282 13879 21316 13913
rect 22109 13889 22143 13923
rect 22293 13889 22327 13923
rect 22661 13889 22695 13923
rect 24133 13889 24167 13923
rect 24501 13889 24535 13923
rect 24777 13889 24811 13923
rect 24869 13889 24903 13923
rect 25053 13889 25087 13923
rect 25145 13889 25179 13923
rect 25605 13889 25639 13923
rect 25697 13889 25731 13923
rect 25881 13889 25915 13923
rect 25973 13889 26007 13923
rect 26065 13889 26099 13923
rect 26249 13889 26283 13923
rect 26341 13889 26375 13923
rect 26525 13889 26559 13923
rect 26617 13889 26651 13923
rect 26801 13889 26835 13923
rect 27077 13879 27111 13913
rect 27261 13889 27295 13923
rect 28825 13889 28859 13923
rect 29101 13889 29135 13923
rect 29285 13889 29319 13923
rect 30205 13889 30239 13923
rect 30389 13889 30423 13923
rect 30481 13889 30515 13923
rect 30757 13889 30791 13923
rect 30941 13889 30975 13923
rect 31953 13889 31987 13923
rect 32781 13889 32815 13923
rect 32965 13889 32999 13923
rect 33057 13889 33091 13923
rect 33241 13889 33275 13923
rect 1501 13821 1535 13855
rect 7205 13821 7239 13855
rect 15577 13821 15611 13855
rect 17969 13821 18003 13855
rect 21925 13821 21959 13855
rect 22477 13821 22511 13855
rect 23029 13821 23063 13855
rect 23121 13821 23155 13855
rect 23213 13821 23247 13855
rect 23305 13821 23339 13855
rect 23673 13821 23707 13855
rect 28917 13821 28951 13855
rect 30573 13821 30607 13855
rect 31677 13821 31711 13855
rect 21557 13753 21591 13787
rect 24409 13753 24443 13787
rect 25329 13753 25363 13787
rect 15025 13685 15059 13719
rect 17417 13685 17451 13719
rect 26157 13685 26191 13719
rect 26801 13685 26835 13719
rect 27169 13685 27203 13719
rect 28549 13685 28583 13719
rect 31861 13685 31895 13719
rect 33241 13685 33275 13719
rect 4261 13481 4295 13515
rect 10517 13481 10551 13515
rect 15393 13481 15427 13515
rect 16681 13481 16715 13515
rect 17877 13481 17911 13515
rect 18429 13481 18463 13515
rect 18889 13481 18923 13515
rect 19717 13481 19751 13515
rect 20637 13481 20671 13515
rect 27445 13481 27479 13515
rect 28089 13481 28123 13515
rect 28365 13481 28399 13515
rect 29101 13481 29135 13515
rect 29193 13481 29227 13515
rect 33149 13481 33183 13515
rect 33241 13481 33275 13515
rect 33701 13481 33735 13515
rect 9137 13413 9171 13447
rect 13553 13413 13587 13447
rect 22661 13413 22695 13447
rect 22937 13413 22971 13447
rect 28273 13413 28307 13447
rect 4353 13345 4387 13379
rect 6377 13345 6411 13379
rect 7113 13345 7147 13379
rect 9781 13345 9815 13379
rect 10977 13345 11011 13379
rect 12909 13345 12943 13379
rect 21005 13345 21039 13379
rect 24777 13345 24811 13379
rect 26249 13345 26283 13379
rect 26341 13345 26375 13379
rect 26709 13345 26743 13379
rect 29009 13345 29043 13379
rect 32965 13345 32999 13379
rect 34069 13345 34103 13379
rect 3893 13277 3927 13311
rect 8769 13277 8803 13311
rect 10149 13277 10183 13311
rect 10241 13277 10275 13311
rect 10609 13277 10643 13311
rect 10701 13277 10735 13311
rect 13185 13277 13219 13311
rect 13829 13277 13863 13311
rect 15025 13277 15059 13311
rect 17785 13277 17819 13311
rect 19993 13277 20027 13311
rect 20085 13277 20119 13311
rect 20177 13277 20211 13311
rect 20361 13277 20395 13311
rect 21097 13277 21131 13311
rect 21373 13277 21407 13311
rect 21741 13277 21775 13311
rect 22385 13277 22419 13311
rect 22569 13277 22603 13311
rect 22937 13277 22971 13311
rect 23213 13277 23247 13311
rect 23489 13277 23523 13311
rect 24409 13277 24443 13311
rect 24593 13277 24627 13311
rect 25697 13277 25731 13311
rect 25881 13277 25915 13311
rect 25973 13277 26007 13311
rect 26157 13277 26191 13311
rect 26525 13277 26559 13311
rect 26801 13277 26835 13311
rect 26985 13277 27019 13311
rect 27077 13277 27111 13311
rect 27189 13277 27223 13311
rect 28457 13277 28491 13311
rect 28549 13277 28583 13311
rect 28733 13277 28767 13311
rect 29285 13277 29319 13311
rect 29561 13277 29595 13311
rect 29745 13277 29779 13311
rect 32873 13277 32907 13311
rect 33425 13277 33459 13311
rect 33517 13277 33551 13311
rect 33885 13277 33919 13311
rect 4077 13209 4111 13243
rect 4629 13209 4663 13243
rect 6929 13209 6963 13243
rect 9965 13209 9999 13243
rect 11253 13209 11287 13243
rect 15209 13209 15243 13243
rect 16681 13209 16715 13243
rect 16865 13209 16899 13243
rect 18245 13209 18279 13243
rect 18873 13209 18907 13243
rect 19073 13209 19107 13243
rect 20453 13209 20487 13243
rect 20653 13209 20687 13243
rect 23305 13209 23339 13243
rect 23673 13209 23707 13243
rect 32505 13209 32539 13243
rect 32597 13209 32631 13243
rect 6561 13141 6595 13175
rect 7021 13141 7055 13175
rect 8585 13141 8619 13175
rect 9505 13141 9539 13175
rect 9597 13141 9631 13175
rect 10885 13141 10919 13175
rect 12725 13141 12759 13175
rect 13093 13141 13127 13175
rect 13645 13141 13679 13175
rect 16497 13141 16531 13175
rect 18445 13141 18479 13175
rect 18613 13141 18647 13175
rect 18705 13141 18739 13175
rect 20821 13141 20855 13175
rect 21557 13141 21591 13175
rect 25789 13141 25823 13175
rect 29653 13141 29687 13175
rect 3157 12937 3191 12971
rect 4997 12937 5031 12971
rect 8125 12937 8159 12971
rect 10517 12937 10551 12971
rect 14933 12937 14967 12971
rect 15577 12937 15611 12971
rect 19743 12937 19777 12971
rect 20361 12937 20395 12971
rect 21649 12937 21683 12971
rect 22017 12937 22051 12971
rect 26249 12937 26283 12971
rect 31217 12937 31251 12971
rect 31861 12937 31895 12971
rect 32873 12937 32907 12971
rect 4077 12869 4111 12903
rect 4537 12869 4571 12903
rect 8585 12869 8619 12903
rect 13461 12869 13495 12903
rect 17601 12869 17635 12903
rect 19533 12869 19567 12903
rect 31493 12869 31527 12903
rect 31709 12869 31743 12903
rect 32505 12869 32539 12903
rect 1409 12801 1443 12835
rect 3985 12801 4019 12835
rect 4445 12801 4479 12835
rect 4629 12801 4663 12835
rect 5181 12801 5215 12835
rect 6009 12801 6043 12835
rect 6377 12801 6411 12835
rect 8309 12801 8343 12835
rect 10333 12801 10367 12835
rect 10609 12801 10643 12835
rect 13093 12801 13127 12835
rect 13185 12801 13219 12835
rect 15485 12801 15519 12835
rect 16865 12801 16899 12835
rect 20545 12801 20579 12835
rect 21119 12801 21153 12835
rect 21465 12801 21499 12835
rect 21833 12801 21867 12835
rect 24685 12801 24719 12835
rect 24961 12801 24995 12835
rect 25053 12801 25087 12835
rect 26433 12801 26467 12835
rect 26525 12801 26559 12835
rect 26709 12801 26743 12835
rect 26801 12801 26835 12835
rect 29101 12801 29135 12835
rect 30665 12801 30699 12835
rect 31217 12801 31251 12835
rect 31401 12801 31435 12835
rect 32137 12801 32171 12835
rect 32321 12801 32355 12835
rect 33149 12801 33183 12835
rect 1685 12733 1719 12767
rect 4169 12733 4203 12767
rect 6653 12733 6687 12767
rect 12265 12733 12299 12767
rect 15669 12733 15703 12767
rect 20177 12733 20211 12767
rect 22293 12733 22327 12767
rect 22385 12733 22419 12767
rect 24409 12733 24443 12767
rect 24501 12733 24535 12767
rect 24593 12733 24627 12767
rect 25237 12733 25271 12767
rect 29377 12733 29411 12767
rect 30573 12733 30607 12767
rect 32873 12733 32907 12767
rect 33057 12733 33091 12767
rect 6193 12665 6227 12699
rect 10057 12665 10091 12699
rect 19901 12665 19935 12699
rect 29193 12665 29227 12699
rect 31033 12665 31067 12699
rect 3617 12597 3651 12631
rect 10149 12597 10183 12631
rect 15117 12597 15151 12631
rect 19717 12597 19751 12631
rect 19993 12597 20027 12631
rect 21465 12597 21499 12631
rect 24869 12597 24903 12631
rect 25145 12597 25179 12631
rect 29285 12597 29319 12631
rect 31677 12597 31711 12631
rect 1961 12393 1995 12427
rect 3801 12393 3835 12427
rect 3985 12393 4019 12427
rect 4261 12393 4295 12427
rect 6469 12393 6503 12427
rect 8585 12393 8619 12427
rect 11529 12393 11563 12427
rect 16865 12393 16899 12427
rect 21741 12393 21775 12427
rect 25237 12393 25271 12427
rect 26893 12393 26927 12427
rect 29561 12393 29595 12427
rect 30205 12393 30239 12427
rect 17601 12325 17635 12359
rect 3065 12257 3099 12291
rect 3249 12257 3283 12291
rect 6929 12257 6963 12291
rect 7113 12257 7147 12291
rect 9781 12257 9815 12291
rect 12173 12257 12207 12291
rect 18061 12257 18095 12291
rect 18245 12257 18279 12291
rect 18429 12257 18463 12291
rect 23029 12257 23063 12291
rect 23121 12257 23155 12291
rect 23213 12257 23247 12291
rect 23397 12257 23431 12291
rect 23765 12257 23799 12291
rect 25789 12257 25823 12291
rect 26249 12257 26283 12291
rect 2145 12189 2179 12223
rect 2973 12189 3007 12223
rect 4261 12189 4295 12223
rect 4537 12189 4571 12223
rect 6837 12189 6871 12223
rect 8217 12189 8251 12223
rect 8401 12189 8435 12223
rect 9965 12189 9999 12223
rect 10149 12189 10183 12223
rect 11989 12189 12023 12223
rect 14749 12189 14783 12223
rect 15117 12189 15151 12223
rect 18613 12189 18647 12223
rect 18981 12189 19015 12223
rect 19349 12189 19383 12223
rect 22937 12189 22971 12223
rect 23489 12189 23523 12223
rect 23581 12189 23615 12223
rect 25605 12189 25639 12223
rect 26433 12189 26467 12223
rect 29837 12189 29871 12223
rect 30021 12189 30055 12223
rect 30297 12189 30331 12223
rect 30389 12189 30423 12223
rect 30573 12189 30607 12223
rect 33149 12189 33183 12223
rect 33517 12189 33551 12223
rect 4169 12121 4203 12155
rect 4445 12121 4479 12155
rect 8677 12121 8711 12155
rect 11897 12121 11931 12155
rect 15393 12121 15427 12155
rect 18889 12121 18923 12155
rect 21557 12121 21591 12155
rect 21773 12121 21807 12155
rect 29929 12121 29963 12155
rect 2605 12053 2639 12087
rect 3959 12053 3993 12087
rect 8033 12053 8067 12087
rect 14933 12053 14967 12087
rect 17969 12053 18003 12087
rect 19533 12053 19567 12087
rect 21925 12053 21959 12087
rect 23765 12053 23799 12087
rect 25697 12053 25731 12087
rect 26525 12053 26559 12087
rect 30481 12053 30515 12087
rect 33149 12053 33183 12087
rect 1593 11849 1627 11883
rect 12173 11849 12207 11883
rect 24402 11849 24436 11883
rect 29285 11849 29319 11883
rect 29745 11849 29779 11883
rect 30205 11849 30239 11883
rect 32413 11849 32447 11883
rect 12541 11781 12575 11815
rect 27905 11781 27939 11815
rect 27675 11747 27709 11781
rect 1501 11713 1535 11747
rect 10701 11713 10735 11747
rect 10793 11713 10827 11747
rect 11989 11713 12023 11747
rect 15945 11713 15979 11747
rect 18613 11713 18647 11747
rect 18797 11713 18831 11747
rect 23489 11713 23523 11747
rect 23765 11713 23799 11747
rect 24225 11713 24259 11747
rect 24317 11713 24351 11747
rect 24501 11713 24535 11747
rect 24593 11713 24627 11747
rect 24777 11713 24811 11747
rect 24869 11713 24903 11747
rect 25053 11713 25087 11747
rect 27169 11713 27203 11747
rect 27353 11713 27387 11747
rect 27445 11713 27479 11747
rect 29469 11713 29503 11747
rect 29929 11713 29963 11747
rect 30573 11713 30607 11747
rect 32597 11713 32631 11747
rect 32689 11713 32723 11747
rect 10885 11645 10919 11679
rect 12265 11645 12299 11679
rect 14289 11645 14323 11679
rect 16037 11645 16071 11679
rect 16129 11645 16163 11679
rect 24961 11645 24995 11679
rect 29561 11645 29595 11679
rect 29837 11645 29871 11679
rect 30665 11645 30699 11679
rect 18705 11577 18739 11611
rect 24593 11577 24627 11611
rect 27537 11577 27571 11611
rect 10333 11509 10367 11543
rect 15577 11509 15611 11543
rect 23581 11509 23615 11543
rect 26985 11509 27019 11543
rect 27721 11509 27755 11543
rect 30849 11509 30883 11543
rect 3157 11305 3191 11339
rect 5733 11305 5767 11339
rect 8493 11305 8527 11339
rect 12449 11305 12483 11339
rect 17601 11305 17635 11339
rect 28917 11305 28951 11339
rect 29285 11305 29319 11339
rect 31401 11305 31435 11339
rect 32137 11305 32171 11339
rect 8033 11237 8067 11271
rect 9321 11237 9355 11271
rect 9965 11237 9999 11271
rect 14105 11237 14139 11271
rect 15761 11237 15795 11271
rect 21925 11237 21959 11271
rect 30573 11237 30607 11271
rect 1409 11169 1443 11203
rect 4353 11169 4387 11203
rect 8309 11169 8343 11203
rect 9229 11169 9263 11203
rect 10057 11169 10091 11203
rect 10333 11169 10367 11203
rect 11805 11169 11839 11203
rect 13001 11169 13035 11203
rect 14657 11169 14691 11203
rect 16129 11169 16163 11203
rect 19441 11169 19475 11203
rect 23765 11169 23799 11203
rect 26249 11169 26283 11203
rect 27169 11169 27203 11203
rect 30113 11169 30147 11203
rect 30389 11169 30423 11203
rect 5917 11101 5951 11135
rect 6101 11101 6135 11135
rect 7389 11101 7423 11135
rect 7481 11101 7515 11135
rect 7665 11101 7699 11135
rect 7757 11101 7791 11135
rect 8585 11101 8619 11135
rect 9137 11101 9171 11135
rect 9413 11101 9447 11135
rect 9781 11101 9815 11135
rect 12817 11101 12851 11135
rect 13737 11101 13771 11135
rect 14473 11101 14507 11135
rect 15577 11101 15611 11135
rect 15853 11101 15887 11135
rect 18613 11101 18647 11135
rect 18797 11101 18831 11135
rect 19257 11101 19291 11135
rect 19901 11101 19935 11135
rect 19993 11101 20027 11135
rect 20085 11101 20119 11135
rect 21373 11101 21407 11135
rect 21649 11101 21683 11135
rect 21741 11101 21775 11135
rect 22017 11101 22051 11135
rect 22201 11101 22235 11135
rect 22477 11101 22511 11135
rect 23581 11101 23615 11135
rect 25421 11101 25455 11135
rect 25605 11101 25639 11135
rect 26433 11101 26467 11135
rect 26893 11101 26927 11135
rect 27077 11101 27111 11135
rect 27261 11101 27295 11135
rect 27445 11101 27479 11135
rect 27721 11101 27755 11135
rect 27905 11101 27939 11135
rect 28181 11101 28215 11135
rect 28273 11101 28307 11135
rect 28457 11101 28491 11135
rect 29101 11101 29135 11135
rect 29377 11101 29411 11135
rect 30205 11101 30239 11135
rect 30297 11101 30331 11135
rect 31585 11101 31619 11135
rect 31861 11101 31895 11135
rect 32045 11101 32079 11135
rect 32321 11101 32355 11135
rect 32597 11101 32631 11135
rect 32781 11101 32815 11135
rect 32873 11101 32907 11135
rect 33057 11101 33091 11135
rect 37565 11101 37599 11135
rect 1685 11033 1719 11067
rect 4169 11033 4203 11067
rect 7941 11033 7975 11067
rect 8953 11033 8987 11067
rect 12909 11033 12943 11067
rect 14565 11033 14599 11067
rect 18429 11033 18463 11067
rect 20269 11033 20303 11067
rect 21557 11033 21591 11067
rect 25513 11033 25547 11067
rect 28089 11033 28123 11067
rect 28365 11033 28399 11067
rect 37933 11033 37967 11067
rect 3801 10965 3835 10999
rect 4261 10965 4295 10999
rect 13921 10965 13955 10999
rect 22385 10965 22419 10999
rect 23397 10965 23431 10999
rect 26341 10965 26375 10999
rect 26801 10965 26835 10999
rect 27629 10965 27663 10999
rect 32965 10965 32999 10999
rect 1777 10761 1811 10795
rect 2789 10761 2823 10795
rect 5825 10761 5859 10795
rect 8677 10761 8711 10795
rect 9045 10761 9079 10795
rect 19165 10761 19199 10795
rect 24133 10761 24167 10795
rect 32229 10761 32263 10795
rect 33701 10761 33735 10795
rect 35081 10761 35115 10795
rect 7389 10693 7423 10727
rect 7573 10693 7607 10727
rect 14197 10693 14231 10727
rect 15945 10693 15979 10727
rect 20821 10693 20855 10727
rect 21021 10693 21055 10727
rect 23029 10693 23063 10727
rect 23121 10693 23155 10727
rect 23259 10693 23293 10727
rect 1961 10625 1995 10659
rect 2697 10625 2731 10659
rect 3341 10625 3375 10659
rect 6009 10625 6043 10659
rect 6193 10625 6227 10659
rect 6745 10625 6779 10659
rect 7205 10625 7239 10659
rect 8585 10625 8619 10659
rect 8861 10625 8895 10659
rect 9597 10625 9631 10659
rect 10977 10625 11011 10659
rect 13921 10625 13955 10659
rect 16865 10625 16899 10659
rect 17049 10625 17083 10659
rect 17141 10625 17175 10659
rect 17233 10625 17267 10659
rect 18153 10625 18187 10659
rect 18337 10625 18371 10659
rect 18981 10625 19015 10659
rect 20269 10625 20303 10659
rect 21465 10625 21499 10659
rect 22100 10625 22134 10659
rect 22201 10625 22235 10659
rect 22385 10625 22419 10659
rect 22477 10625 22511 10659
rect 22937 10625 22971 10659
rect 24225 10625 24259 10659
rect 26985 10625 27019 10659
rect 27169 10625 27203 10659
rect 27261 10625 27295 10659
rect 27353 10625 27387 10659
rect 28181 10625 28215 10659
rect 28365 10625 28399 10659
rect 28733 10625 28767 10659
rect 28917 10625 28951 10659
rect 30297 10625 30331 10659
rect 30481 10625 30515 10659
rect 32137 10625 32171 10659
rect 32321 10625 32355 10659
rect 32597 10625 32631 10659
rect 33517 10625 33551 10659
rect 33793 10625 33827 10659
rect 34069 10625 34103 10659
rect 34713 10625 34747 10659
rect 2973 10557 3007 10591
rect 3433 10557 3467 10591
rect 3709 10557 3743 10591
rect 4077 10557 4111 10591
rect 4353 10557 4387 10591
rect 6101 10557 6135 10591
rect 6837 10557 6871 10591
rect 6929 10557 6963 10591
rect 9137 10557 9171 10591
rect 11069 10557 11103 10591
rect 11253 10557 11287 10591
rect 21281 10557 21315 10591
rect 21649 10557 21683 10591
rect 23397 10557 23431 10591
rect 23949 10557 23983 10591
rect 30389 10557 30423 10591
rect 32505 10557 32539 10591
rect 33977 10557 34011 10591
rect 34621 10557 34655 10591
rect 2329 10489 2363 10523
rect 10609 10489 10643 10523
rect 17509 10489 17543 10523
rect 24593 10489 24627 10523
rect 28457 10489 28491 10523
rect 28733 10489 28767 10523
rect 34437 10489 34471 10523
rect 6377 10421 6411 10455
rect 9321 10421 9355 10455
rect 18061 10421 18095 10455
rect 20177 10421 20211 10455
rect 21005 10421 21039 10455
rect 21189 10421 21223 10455
rect 21925 10421 21959 10455
rect 22753 10421 22787 10455
rect 27629 10421 27663 10455
rect 32873 10421 32907 10455
rect 33517 10421 33551 10455
rect 4629 10217 4663 10251
rect 6193 10217 6227 10251
rect 7573 10217 7607 10251
rect 20453 10217 20487 10251
rect 20913 10217 20947 10251
rect 22385 10217 22419 10251
rect 22661 10217 22695 10251
rect 32689 10217 32723 10251
rect 33517 10217 33551 10251
rect 8493 10149 8527 10183
rect 20821 10149 20855 10183
rect 21189 10149 21223 10183
rect 21649 10149 21683 10183
rect 29009 10149 29043 10183
rect 5641 10081 5675 10115
rect 5825 10081 5859 10115
rect 7757 10081 7791 10115
rect 9045 10081 9079 10115
rect 9321 10081 9355 10115
rect 13737 10081 13771 10115
rect 21281 10081 21315 10115
rect 21373 10081 21407 10115
rect 22385 10081 22419 10115
rect 30481 10081 30515 10115
rect 2973 10013 3007 10047
rect 4813 10013 4847 10047
rect 5549 10013 5583 10047
rect 6009 10013 6043 10047
rect 6193 10013 6227 10047
rect 7481 10013 7515 10047
rect 7849 10013 7883 10047
rect 8334 10013 8368 10047
rect 9137 10013 9171 10047
rect 9229 10013 9263 10047
rect 11437 10013 11471 10047
rect 11713 10013 11747 10047
rect 17693 10013 17727 10047
rect 17785 10013 17819 10047
rect 18061 10013 18095 10047
rect 18245 10013 18279 10047
rect 18337 10013 18371 10047
rect 18429 10013 18463 10047
rect 20269 10013 20303 10047
rect 20453 10013 20487 10047
rect 20545 10013 20579 10047
rect 21097 10013 21131 10047
rect 21557 10013 21591 10047
rect 21925 10013 21959 10047
rect 22293 10013 22327 10047
rect 28641 10013 28675 10047
rect 28733 10013 28767 10047
rect 28917 10013 28951 10047
rect 30113 10013 30147 10047
rect 30297 10013 30331 10047
rect 30389 10013 30423 10047
rect 30665 10013 30699 10047
rect 32597 10013 32631 10047
rect 33793 10013 33827 10047
rect 33885 10013 33919 10047
rect 33977 10013 34011 10047
rect 34161 10013 34195 10047
rect 2789 9945 2823 9979
rect 11989 9945 12023 9979
rect 17969 9945 18003 9979
rect 19349 9945 19383 9979
rect 19717 9945 19751 9979
rect 20821 9945 20855 9979
rect 21649 9945 21683 9979
rect 28457 9945 28491 9979
rect 3157 9877 3191 9911
rect 5181 9877 5215 9911
rect 7757 9877 7791 9911
rect 8125 9877 8159 9911
rect 8217 9877 8251 9911
rect 9505 9877 9539 9911
rect 11621 9877 11655 9911
rect 18705 9877 18739 9911
rect 20637 9877 20671 9911
rect 21833 9877 21867 9911
rect 28273 9877 28307 9911
rect 30849 9877 30883 9911
rect 11805 9673 11839 9707
rect 13553 9673 13587 9707
rect 16037 9673 16071 9707
rect 22477 9673 22511 9707
rect 33241 9673 33275 9707
rect 6377 9605 6411 9639
rect 8309 9605 8343 9639
rect 8585 9605 8619 9639
rect 15485 9605 15519 9639
rect 24593 9605 24627 9639
rect 24685 9605 24719 9639
rect 26341 9605 26375 9639
rect 33057 9605 33091 9639
rect 3249 9537 3283 9571
rect 3341 9537 3375 9571
rect 3433 9537 3467 9571
rect 3617 9537 3651 9571
rect 6653 9537 6687 9571
rect 6745 9537 6779 9571
rect 6837 9537 6871 9571
rect 7021 9537 7055 9571
rect 7757 9537 7791 9571
rect 8033 9537 8067 9571
rect 8493 9537 8527 9571
rect 8677 9537 8711 9571
rect 10241 9537 10275 9571
rect 10701 9537 10735 9571
rect 10793 9537 10827 9571
rect 12173 9537 12207 9571
rect 12265 9537 12299 9571
rect 13461 9537 13495 9571
rect 15577 9537 15611 9571
rect 16221 9537 16255 9571
rect 16773 9537 16807 9571
rect 18429 9537 18463 9571
rect 18797 9537 18831 9571
rect 19809 9537 19843 9571
rect 20085 9537 20119 9571
rect 22661 9537 22695 9571
rect 22753 9537 22787 9571
rect 23029 9537 23063 9571
rect 24133 9537 24167 9571
rect 24317 9537 24351 9571
rect 24409 9537 24443 9571
rect 24777 9537 24811 9571
rect 26157 9537 26191 9571
rect 26433 9537 26467 9571
rect 26617 9537 26651 9571
rect 26985 9537 27019 9571
rect 27169 9537 27203 9571
rect 27445 9537 27479 9571
rect 29009 9537 29043 9571
rect 29653 9537 29687 9571
rect 29837 9537 29871 9571
rect 29937 9537 29971 9571
rect 30113 9527 30147 9561
rect 30757 9537 30791 9571
rect 31033 9537 31067 9571
rect 31309 9537 31343 9571
rect 31585 9537 31619 9571
rect 32505 9537 32539 9571
rect 32873 9537 32907 9571
rect 10885 9469 10919 9503
rect 12449 9469 12483 9503
rect 13645 9469 13679 9503
rect 15301 9469 15335 9503
rect 17141 9469 17175 9503
rect 18245 9469 18279 9503
rect 18889 9469 18923 9503
rect 19441 9469 19475 9503
rect 19901 9469 19935 9503
rect 19993 9469 20027 9503
rect 23121 9469 23155 9503
rect 25973 9469 26007 9503
rect 28825 9469 28859 9503
rect 29745 9469 29779 9503
rect 32413 9469 32447 9503
rect 7481 9401 7515 9435
rect 8033 9401 8067 9435
rect 10333 9401 10367 9435
rect 15945 9401 15979 9435
rect 24961 9401 24995 9435
rect 31217 9401 31251 9435
rect 32137 9401 32171 9435
rect 2973 9333 3007 9367
rect 10057 9333 10091 9367
rect 13093 9333 13127 9367
rect 19625 9333 19659 9367
rect 24317 9333 24351 9367
rect 26525 9333 26559 9367
rect 27629 9333 27663 9367
rect 29193 9333 29227 9367
rect 30021 9333 30055 9367
rect 11529 9129 11563 9163
rect 17509 9129 17543 9163
rect 20913 9129 20947 9163
rect 23949 9129 23983 9163
rect 29377 9129 29411 9163
rect 29745 9129 29779 9163
rect 31769 9129 31803 9163
rect 32873 9129 32907 9163
rect 33241 9129 33275 9163
rect 22845 9061 22879 9095
rect 29929 9061 29963 9095
rect 32413 9061 32447 9095
rect 4629 8993 4663 9027
rect 8677 8993 8711 9027
rect 9781 8993 9815 9027
rect 10057 8993 10091 9027
rect 13645 8993 13679 9027
rect 15393 8993 15427 9027
rect 15577 8993 15611 9027
rect 18337 8993 18371 9027
rect 20729 8993 20763 9027
rect 22201 8993 22235 9027
rect 22661 8993 22695 9027
rect 25329 8993 25363 9027
rect 25789 8993 25823 9027
rect 27997 8993 28031 9027
rect 31493 8993 31527 9027
rect 1777 8925 1811 8959
rect 4169 8925 4203 8959
rect 4261 8925 4295 8959
rect 4353 8925 4387 8959
rect 4537 8925 4571 8959
rect 4997 8925 5031 8959
rect 5825 8925 5859 8959
rect 12725 8925 12759 8959
rect 12909 8925 12943 8959
rect 13369 8925 13403 8959
rect 14105 8925 14139 8959
rect 14289 8925 14323 8959
rect 14381 8925 14415 8959
rect 14473 8925 14507 8959
rect 15301 8925 15335 8959
rect 15761 8925 15795 8959
rect 17969 8925 18003 8959
rect 18521 8925 18555 8959
rect 19717 8925 19751 8959
rect 19993 8925 20027 8959
rect 20637 8925 20671 8959
rect 22569 8925 22603 8959
rect 22937 8925 22971 8959
rect 23030 8925 23064 8959
rect 23213 8925 23247 8959
rect 23402 8925 23436 8959
rect 23857 8925 23891 8959
rect 24409 8925 24443 8959
rect 24502 8925 24536 8959
rect 24893 8925 24927 8959
rect 25237 8925 25271 8959
rect 25513 8925 25547 8959
rect 25605 8925 25639 8959
rect 25881 8925 25915 8959
rect 26065 8925 26099 8959
rect 26157 8925 26191 8959
rect 26249 8925 26283 8959
rect 26801 8925 26835 8959
rect 26985 8925 27019 8959
rect 27077 8925 27111 8959
rect 27169 8925 27203 8959
rect 27353 8925 27387 8959
rect 27629 8925 27663 8959
rect 28181 8925 28215 8959
rect 28365 8925 28399 8959
rect 28457 8925 28491 8959
rect 28549 8925 28583 8959
rect 28917 8925 28951 8959
rect 29101 8925 29135 8959
rect 29193 8925 29227 8959
rect 29377 8925 29411 8959
rect 29561 8925 29595 8959
rect 29653 8925 29687 8959
rect 30021 8925 30055 8959
rect 30205 8925 30239 8959
rect 31585 8925 31619 8959
rect 31861 8925 31895 8959
rect 32137 8925 32171 8959
rect 32597 8925 32631 8959
rect 32689 8925 32723 8959
rect 32965 8925 32999 8959
rect 33057 8925 33091 8959
rect 33241 8925 33275 8959
rect 33517 8925 33551 8959
rect 37933 8925 37967 8959
rect 1409 8857 1443 8891
rect 4813 8857 4847 8891
rect 6009 8857 6043 8891
rect 6193 8857 6227 8891
rect 8401 8857 8435 8891
rect 12817 8857 12851 8891
rect 16037 8857 16071 8891
rect 19901 8857 19935 8891
rect 20269 8857 20303 8891
rect 22293 8857 22327 8891
rect 23305 8857 23339 8891
rect 24685 8857 24719 8891
rect 24777 8857 24811 8891
rect 27813 8857 27847 8891
rect 30389 8857 30423 8891
rect 37657 8857 37691 8891
rect 3893 8789 3927 8823
rect 8033 8789 8067 8823
rect 8493 8789 8527 8823
rect 13001 8789 13035 8823
rect 13461 8789 13495 8823
rect 14749 8789 14783 8823
rect 14933 8789 14967 8823
rect 19533 8789 19567 8823
rect 23581 8789 23615 8823
rect 25053 8789 25087 8823
rect 26525 8789 26559 8823
rect 27537 8789 27571 8823
rect 28825 8789 28859 8823
rect 29009 8789 29043 8823
rect 31125 8789 31159 8823
rect 31953 8789 31987 8823
rect 4261 8585 4295 8619
rect 5089 8585 5123 8619
rect 9321 8585 9355 8619
rect 10057 8585 10091 8619
rect 10609 8585 10643 8619
rect 13369 8585 13403 8619
rect 15209 8585 15243 8619
rect 18889 8585 18923 8619
rect 24961 8585 24995 8619
rect 29285 8585 29319 8619
rect 31309 8585 31343 8619
rect 5917 8517 5951 8551
rect 6545 8517 6579 8551
rect 6745 8517 6779 8551
rect 7849 8517 7883 8551
rect 12449 8517 12483 8551
rect 12633 8517 12667 8551
rect 13737 8517 13771 8551
rect 19533 8517 19567 8551
rect 19717 8517 19751 8551
rect 22109 8517 22143 8551
rect 24869 8517 24903 8551
rect 3433 8449 3467 8483
rect 4169 8449 4203 8483
rect 5457 8449 5491 8483
rect 6101 8449 6135 8483
rect 6193 8449 6227 8483
rect 10149 8449 10183 8483
rect 10517 8449 10551 8483
rect 11529 8449 11563 8483
rect 11989 8449 12023 8483
rect 12357 8449 12391 8483
rect 12541 8449 12575 8483
rect 13001 8449 13035 8483
rect 13185 8449 13219 8483
rect 17417 8449 17451 8483
rect 18797 8449 18831 8483
rect 18981 8449 19015 8483
rect 19809 8449 19843 8483
rect 21925 8449 21959 8483
rect 23213 8449 23247 8483
rect 23489 8449 23523 8483
rect 23673 8449 23707 8483
rect 26985 8449 27019 8483
rect 27169 8449 27203 8483
rect 27261 8449 27295 8483
rect 27353 8449 27387 8483
rect 27537 8449 27571 8483
rect 28917 8449 28951 8483
rect 29101 8449 29135 8483
rect 31585 8449 31619 8483
rect 31861 8449 31895 8483
rect 33149 8449 33183 8483
rect 4445 8381 4479 8415
rect 5549 8381 5583 8415
rect 5733 8381 5767 8415
rect 10333 8381 10367 8415
rect 11897 8381 11931 8415
rect 13461 8381 13495 8415
rect 17601 8381 17635 8415
rect 24777 8381 24811 8415
rect 31401 8381 31435 8415
rect 33241 8381 33275 8415
rect 3801 8313 3835 8347
rect 5917 8313 5951 8347
rect 6377 8313 6411 8347
rect 9689 8313 9723 8347
rect 17233 8313 17267 8347
rect 27721 8313 27755 8347
rect 32781 8313 32815 8347
rect 3249 8245 3283 8279
rect 6561 8245 6595 8279
rect 19533 8245 19567 8279
rect 22293 8245 22327 8279
rect 23029 8245 23063 8279
rect 25329 8245 25363 8279
rect 29009 8245 29043 8279
rect 5641 8041 5675 8075
rect 8677 8041 8711 8075
rect 12817 8041 12851 8075
rect 13553 8041 13587 8075
rect 13737 8041 13771 8075
rect 20177 8041 20211 8075
rect 31861 8041 31895 8075
rect 17509 7973 17543 8007
rect 21649 7973 21683 8007
rect 23305 7973 23339 8007
rect 30757 7973 30791 8007
rect 6653 7905 6687 7939
rect 6929 7905 6963 7939
rect 12173 7905 12207 7939
rect 12633 7905 12667 7939
rect 15945 7905 15979 7939
rect 22385 7905 22419 7939
rect 30297 7905 30331 7939
rect 5641 7837 5675 7871
rect 5825 7837 5859 7871
rect 6469 7837 6503 7871
rect 9689 7837 9723 7871
rect 9873 7837 9907 7871
rect 13369 7837 13403 7871
rect 13737 7837 13771 7871
rect 13921 7837 13955 7871
rect 15761 7837 15795 7871
rect 15853 7837 15887 7871
rect 17233 7837 17267 7871
rect 17601 7837 17635 7871
rect 17785 7837 17819 7871
rect 19717 7837 19751 7871
rect 19901 7837 19935 7871
rect 20085 7837 20119 7871
rect 20269 7837 20303 7871
rect 21557 7837 21591 7871
rect 21741 7837 21775 7871
rect 21833 7837 21867 7871
rect 21925 7837 21959 7871
rect 22109 7837 22143 7871
rect 22201 7837 22235 7871
rect 22661 7837 22695 7871
rect 30021 7837 30055 7871
rect 30205 7837 30239 7871
rect 30389 7837 30423 7871
rect 30573 7837 30607 7871
rect 30941 7837 30975 7871
rect 31401 7837 31435 7871
rect 31493 7837 31527 7871
rect 7205 7769 7239 7803
rect 10425 7769 10459 7803
rect 12357 7769 12391 7803
rect 17509 7769 17543 7803
rect 17693 7769 17727 7803
rect 19809 7769 19843 7803
rect 22753 7769 22787 7803
rect 23121 7769 23155 7803
rect 31309 7769 31343 7803
rect 31677 7769 31711 7803
rect 6101 7701 6135 7735
rect 6561 7701 6595 7735
rect 9781 7701 9815 7735
rect 15393 7701 15427 7735
rect 17325 7701 17359 7735
rect 22293 7701 22327 7735
rect 31217 7701 31251 7735
rect 5641 7497 5675 7531
rect 7665 7497 7699 7531
rect 22385 7497 22419 7531
rect 23213 7497 23247 7531
rect 26617 7497 26651 7531
rect 30113 7497 30147 7531
rect 2881 7429 2915 7463
rect 9689 7429 9723 7463
rect 11805 7429 11839 7463
rect 19349 7429 19383 7463
rect 20177 7429 20211 7463
rect 22937 7429 22971 7463
rect 23949 7429 23983 7463
rect 25605 7429 25639 7463
rect 1501 7361 1535 7395
rect 2605 7361 2639 7395
rect 5549 7361 5583 7395
rect 6745 7361 6779 7395
rect 7849 7361 7883 7395
rect 9413 7361 9447 7395
rect 14289 7361 14323 7395
rect 14565 7361 14599 7395
rect 14841 7361 14875 7395
rect 15485 7361 15519 7395
rect 17785 7361 17819 7395
rect 17969 7361 18003 7395
rect 19165 7361 19199 7395
rect 19533 7361 19567 7395
rect 19625 7361 19659 7395
rect 19809 7361 19843 7395
rect 20361 7361 20395 7395
rect 20821 7361 20855 7395
rect 21833 7361 21867 7395
rect 22109 7361 22143 7395
rect 22201 7361 22235 7395
rect 22569 7361 22603 7395
rect 22717 7361 22751 7395
rect 22845 7361 22879 7395
rect 23075 7361 23109 7395
rect 23857 7361 23891 7395
rect 24041 7361 24075 7395
rect 24133 7361 24167 7395
rect 24317 7361 24351 7395
rect 24501 7361 24535 7395
rect 24685 7361 24719 7395
rect 25145 7361 25179 7395
rect 26433 7361 26467 7395
rect 26617 7361 26651 7395
rect 27629 7361 27663 7395
rect 27813 7361 27847 7395
rect 27905 7361 27939 7395
rect 27997 7361 28031 7395
rect 28457 7361 28491 7395
rect 29009 7361 29043 7395
rect 29101 7361 29135 7395
rect 29377 7361 29411 7395
rect 29653 7361 29687 7395
rect 30113 7361 30147 7395
rect 30297 7361 30331 7395
rect 30757 7361 30791 7395
rect 31401 7361 31435 7395
rect 31769 7361 31803 7395
rect 31861 7361 31895 7395
rect 1685 7293 1719 7327
rect 4353 7293 4387 7327
rect 5733 7293 5767 7327
rect 6377 7293 6411 7327
rect 6837 7293 6871 7327
rect 11529 7293 11563 7327
rect 13829 7293 13863 7327
rect 14657 7293 14691 7327
rect 15025 7293 15059 7327
rect 18981 7293 19015 7327
rect 20913 7293 20947 7327
rect 24409 7293 24443 7327
rect 25329 7293 25363 7327
rect 27721 7293 27755 7327
rect 28641 7293 28675 7327
rect 31309 7293 31343 7327
rect 14473 7225 14507 7259
rect 19993 7225 20027 7259
rect 21189 7225 21223 7259
rect 5181 7157 5215 7191
rect 11161 7157 11195 7191
rect 13277 7157 13311 7191
rect 15669 7157 15703 7191
rect 17877 7157 17911 7191
rect 21925 7157 21959 7191
rect 24869 7157 24903 7191
rect 24961 7157 24995 7191
rect 25145 7157 25179 7191
rect 6009 6953 6043 6987
rect 12357 6953 12391 6987
rect 12817 6953 12851 6987
rect 15742 6953 15776 6987
rect 17233 6953 17267 6987
rect 18061 6953 18095 6987
rect 25421 6953 25455 6987
rect 31493 6953 31527 6987
rect 17693 6885 17727 6919
rect 30665 6885 30699 6919
rect 4261 6817 4295 6851
rect 12633 6817 12667 6851
rect 15485 6817 15519 6851
rect 17877 6817 17911 6851
rect 19993 6817 20027 6851
rect 20453 6817 20487 6851
rect 24869 6817 24903 6851
rect 27077 6817 27111 6851
rect 27261 6817 27295 6851
rect 28549 6817 28583 6851
rect 32781 6817 32815 6851
rect 32965 6817 32999 6851
rect 33149 6817 33183 6851
rect 8953 6749 8987 6783
rect 9137 6749 9171 6783
rect 12909 6749 12943 6783
rect 15209 6749 15243 6783
rect 17601 6749 17635 6783
rect 17969 6749 18003 6783
rect 18153 6749 18187 6783
rect 18337 6749 18371 6783
rect 18429 6749 18463 6783
rect 18521 6749 18555 6783
rect 20085 6749 20119 6783
rect 21189 6749 21223 6783
rect 21281 6749 21315 6783
rect 21465 6749 21499 6783
rect 24961 6749 24995 6783
rect 25697 6749 25731 6783
rect 25973 6749 26007 6783
rect 26157 6749 26191 6783
rect 26249 6749 26283 6783
rect 26341 6749 26375 6783
rect 26985 6749 27019 6783
rect 27537 6749 27571 6783
rect 27630 6749 27664 6783
rect 27905 6749 27939 6783
rect 28002 6749 28036 6783
rect 28273 6749 28307 6783
rect 28365 6749 28399 6783
rect 29929 6749 29963 6783
rect 30113 6749 30147 6783
rect 30389 6749 30423 6783
rect 30757 6749 30791 6783
rect 30849 6749 30883 6783
rect 31769 6749 31803 6783
rect 31861 6749 31895 6783
rect 31953 6749 31987 6783
rect 32137 6749 32171 6783
rect 32505 6749 32539 6783
rect 32597 6749 32631 6783
rect 32689 6749 32723 6783
rect 33241 6749 33275 6783
rect 4537 6681 4571 6715
rect 18797 6681 18831 6715
rect 25421 6681 25455 6715
rect 27261 6681 27295 6715
rect 27813 6681 27847 6715
rect 9045 6613 9079 6647
rect 14565 6613 14599 6647
rect 21649 6613 21683 6647
rect 25329 6613 25363 6647
rect 25605 6613 25639 6647
rect 26617 6613 26651 6647
rect 28181 6613 28215 6647
rect 28733 6613 28767 6647
rect 33609 6613 33643 6647
rect 4721 6409 4755 6443
rect 7849 6409 7883 6443
rect 15301 6409 15335 6443
rect 18705 6409 18739 6443
rect 19901 6409 19935 6443
rect 22385 6409 22419 6443
rect 23765 6409 23799 6443
rect 24231 6409 24265 6443
rect 25513 6409 25547 6443
rect 27997 6409 28031 6443
rect 28181 6409 28215 6443
rect 7757 6341 7791 6375
rect 9965 6341 9999 6375
rect 13369 6341 13403 6375
rect 19073 6341 19107 6375
rect 23397 6341 23431 6375
rect 23489 6341 23523 6375
rect 24133 6341 24167 6375
rect 32781 6341 32815 6375
rect 4905 6273 4939 6307
rect 8401 6273 8435 6307
rect 9505 6273 9539 6307
rect 9689 6273 9723 6307
rect 10057 6273 10091 6307
rect 12265 6273 12299 6307
rect 12449 6273 12483 6307
rect 12541 6273 12575 6307
rect 12817 6273 12851 6307
rect 14013 6273 14047 6307
rect 14105 6273 14139 6307
rect 15025 6273 15059 6307
rect 15577 6273 15611 6307
rect 18061 6273 18095 6307
rect 18245 6273 18279 6307
rect 18337 6273 18371 6307
rect 18429 6273 18463 6307
rect 18889 6273 18923 6307
rect 19717 6273 19751 6307
rect 19901 6273 19935 6307
rect 22753 6273 22787 6307
rect 23213 6273 23247 6307
rect 23581 6273 23615 6307
rect 24317 6273 24351 6307
rect 24409 6273 24443 6307
rect 25421 6273 25455 6307
rect 25605 6273 25639 6307
rect 27813 6273 27847 6307
rect 28089 6273 28123 6307
rect 28273 6273 28307 6307
rect 32505 6273 32539 6307
rect 32597 6273 32631 6307
rect 7941 6205 7975 6239
rect 8585 6205 8619 6239
rect 8677 6205 8711 6239
rect 8769 6205 8803 6239
rect 9321 6205 9355 6239
rect 12081 6205 12115 6239
rect 14841 6205 14875 6239
rect 15393 6205 15427 6239
rect 22845 6205 22879 6239
rect 27537 6205 27571 6239
rect 9689 6137 9723 6171
rect 18153 6137 18187 6171
rect 32781 6137 32815 6171
rect 7389 6069 7423 6103
rect 8217 6069 8251 6103
rect 15669 6069 15703 6103
rect 18521 6069 18555 6103
rect 19257 6069 19291 6103
rect 23029 6069 23063 6103
rect 27629 6069 27663 6103
rect 12817 5865 12851 5899
rect 15715 5865 15749 5899
rect 22661 5865 22695 5899
rect 30481 5865 30515 5899
rect 32045 5865 32079 5899
rect 32229 5865 32263 5899
rect 9137 5797 9171 5831
rect 22201 5797 22235 5831
rect 29837 5797 29871 5831
rect 5089 5729 5123 5763
rect 6929 5729 6963 5763
rect 7205 5729 7239 5763
rect 8677 5729 8711 5763
rect 9321 5729 9355 5763
rect 12541 5729 12575 5763
rect 14933 5729 14967 5763
rect 17509 5729 17543 5763
rect 19257 5729 19291 5763
rect 19717 5729 19751 5763
rect 29561 5729 29595 5763
rect 9045 5661 9079 5695
rect 9413 5661 9447 5695
rect 9506 5661 9540 5695
rect 9781 5661 9815 5695
rect 9919 5661 9953 5695
rect 10149 5661 10183 5695
rect 10297 5661 10331 5695
rect 10653 5661 10687 5695
rect 12725 5661 12759 5695
rect 12909 5661 12943 5695
rect 13645 5661 13679 5695
rect 13921 5661 13955 5695
rect 14749 5661 14783 5695
rect 15393 5661 15427 5695
rect 17141 5661 17175 5695
rect 19625 5661 19659 5695
rect 20085 5661 20119 5695
rect 20453 5661 20487 5695
rect 20637 5661 20671 5695
rect 22201 5661 22235 5695
rect 22385 5661 22419 5695
rect 22937 5661 22971 5695
rect 23121 5661 23155 5695
rect 23581 5661 23615 5695
rect 23673 5661 23707 5695
rect 24593 5661 24627 5695
rect 24869 5661 24903 5695
rect 25053 5661 25087 5695
rect 32137 5661 32171 5695
rect 32321 5661 32355 5695
rect 5365 5593 5399 5627
rect 9689 5593 9723 5627
rect 10425 5593 10459 5627
rect 10517 5593 10551 5627
rect 11989 5593 12023 5627
rect 15485 5593 15519 5627
rect 19349 5593 19383 5627
rect 30113 5593 30147 5627
rect 30297 5593 30331 5627
rect 31677 5593 31711 5627
rect 31861 5593 31895 5627
rect 6837 5525 6871 5559
rect 9045 5525 9079 5559
rect 10057 5525 10091 5559
rect 10793 5525 10827 5559
rect 13461 5525 13495 5559
rect 13829 5525 13863 5559
rect 14381 5525 14415 5559
rect 14841 5525 14875 5559
rect 19901 5525 19935 5559
rect 20453 5525 20487 5559
rect 24409 5525 24443 5559
rect 30021 5525 30055 5559
rect 6469 5321 6503 5355
rect 8861 5321 8895 5355
rect 15209 5321 15243 5355
rect 17325 5321 17359 5355
rect 19717 5321 19751 5355
rect 23121 5321 23155 5355
rect 23673 5321 23707 5355
rect 27537 5321 27571 5355
rect 29469 5321 29503 5355
rect 30205 5321 30239 5355
rect 31493 5321 31527 5355
rect 9505 5253 9539 5287
rect 9689 5253 9723 5287
rect 11805 5253 11839 5287
rect 13737 5253 13771 5287
rect 19349 5253 19383 5287
rect 19533 5253 19567 5287
rect 21097 5253 21131 5287
rect 22937 5253 22971 5287
rect 25881 5253 25915 5287
rect 6653 5185 6687 5219
rect 8217 5185 8251 5219
rect 9321 5185 9355 5219
rect 9597 5185 9631 5219
rect 10517 5185 10551 5219
rect 11529 5185 11563 5219
rect 13461 5185 13495 5219
rect 19809 5185 19843 5219
rect 19993 5185 20027 5219
rect 20913 5185 20947 5219
rect 22293 5185 22327 5219
rect 23029 5185 23063 5219
rect 23213 5185 23247 5219
rect 23397 5185 23431 5219
rect 25605 5185 25639 5219
rect 25697 5185 25731 5219
rect 27169 5185 27203 5219
rect 27629 5185 27663 5219
rect 27721 5185 27755 5219
rect 27905 5185 27939 5219
rect 28549 5185 28583 5219
rect 28733 5185 28767 5219
rect 28917 5185 28951 5219
rect 29009 5185 29043 5219
rect 29561 5185 29595 5219
rect 29745 5185 29779 5219
rect 29929 5185 29963 5219
rect 30021 5185 30055 5219
rect 30481 5185 30515 5219
rect 30757 5185 30791 5219
rect 31125 5185 31159 5219
rect 10241 5117 10275 5151
rect 15853 5117 15887 5151
rect 16681 5117 16715 5151
rect 22385 5117 22419 5151
rect 23673 5117 23707 5151
rect 25881 5117 25915 5151
rect 27077 5117 27111 5151
rect 30573 5117 30607 5151
rect 31033 5117 31067 5151
rect 13277 5049 13311 5083
rect 21281 5049 21315 5083
rect 27905 5049 27939 5083
rect 29285 5049 29319 5083
rect 29837 5049 29871 5083
rect 30665 5049 30699 5083
rect 9137 4981 9171 5015
rect 11161 4981 11195 5015
rect 16405 4981 16439 5015
rect 19901 4981 19935 5015
rect 23489 4981 23523 5015
rect 30297 4981 30331 5015
rect 9873 4777 9907 4811
rect 10964 4777 10998 4811
rect 12449 4777 12483 4811
rect 15945 4777 15979 4811
rect 16589 4777 16623 4811
rect 20177 4777 20211 4811
rect 20361 4777 20395 4811
rect 23489 4777 23523 4811
rect 24409 4777 24443 4811
rect 25697 4777 25731 4811
rect 26065 4777 26099 4811
rect 27537 4777 27571 4811
rect 29653 4777 29687 4811
rect 30021 4777 30055 4811
rect 10701 4641 10735 4675
rect 14197 4641 14231 4675
rect 19533 4641 19567 4675
rect 24593 4641 24627 4675
rect 26617 4641 26651 4675
rect 27077 4641 27111 4675
rect 27997 4641 28031 4675
rect 28641 4641 28675 4675
rect 1777 4573 1811 4607
rect 10057 4573 10091 4607
rect 10241 4573 10275 4607
rect 16037 4573 16071 4607
rect 16313 4573 16347 4607
rect 16405 4573 16439 4607
rect 19441 4573 19475 4607
rect 21281 4573 21315 4607
rect 21833 4573 21867 4607
rect 23204 4573 23238 4607
rect 24685 4573 24719 4607
rect 24777 4573 24811 4607
rect 24869 4573 24903 4607
rect 25053 4573 25087 4607
rect 25329 4573 25363 4607
rect 25605 4573 25639 4607
rect 26157 4573 26191 4607
rect 26341 4573 26375 4607
rect 26709 4573 26743 4607
rect 27353 4573 27387 4607
rect 27905 4573 27939 4607
rect 29561 4573 29595 4607
rect 30113 4573 30147 4607
rect 30205 4573 30239 4607
rect 30297 4573 30331 4607
rect 1409 4505 1443 4539
rect 14473 4505 14507 4539
rect 16221 4505 16255 4539
rect 19993 4505 20027 4539
rect 20209 4505 20243 4539
rect 23489 4505 23523 4539
rect 25145 4505 25179 4539
rect 25513 4505 25547 4539
rect 26249 4505 26283 4539
rect 27169 4505 27203 4539
rect 19809 4437 19843 4471
rect 23305 4437 23339 4471
rect 26433 4437 26467 4471
rect 9781 4233 9815 4267
rect 14565 4233 14599 4267
rect 25421 4233 25455 4267
rect 27905 4233 27939 4267
rect 8309 4165 8343 4199
rect 8033 4097 8067 4131
rect 14381 4097 14415 4131
rect 24961 4097 24995 4131
rect 25145 4097 25179 4131
rect 25237 4097 25271 4131
rect 25421 4097 25455 4131
rect 27813 4097 27847 4131
rect 27997 4097 28031 4131
rect 25145 3961 25179 3995
rect 37565 3077 37599 3111
rect 1961 3009 1995 3043
rect 2421 3009 2455 3043
rect 12541 3009 12575 3043
rect 13185 3009 13219 3043
rect 15117 3009 15151 3043
rect 17233 3009 17267 3043
rect 19993 3009 20027 3043
rect 1777 2805 1811 2839
rect 2237 2805 2271 2839
rect 12357 2805 12391 2839
rect 13001 2805 13035 2839
rect 14933 2805 14967 2839
rect 17417 2805 17451 2839
rect 19809 2805 19843 2839
rect 37657 2805 37691 2839
rect 8677 2601 8711 2635
rect 11161 2601 11195 2635
rect 37657 2533 37691 2567
rect 1777 2397 1811 2431
rect 2421 2397 2455 2431
rect 4353 2397 4387 2431
rect 6929 2397 6963 2431
rect 8493 2397 8527 2431
rect 13093 2397 13127 2431
rect 15025 2397 15059 2431
rect 17601 2397 17635 2431
rect 19809 2397 19843 2431
rect 37473 2397 37507 2431
rect 1409 2329 1443 2363
rect 2053 2329 2087 2363
rect 3985 2329 4019 2363
rect 6561 2329 6595 2363
rect 11253 2329 11287 2363
rect 19441 2329 19475 2363
rect 27077 2329 27111 2363
rect 13185 2261 13219 2295
rect 15301 2261 15335 2295
rect 17693 2261 17727 2295
rect 27169 2261 27203 2295
<< metal1 >>
rect 1104 39194 38272 39216
rect 1104 39142 4874 39194
rect 4926 39142 4938 39194
rect 4990 39142 5002 39194
rect 5054 39142 5066 39194
rect 5118 39142 5130 39194
rect 5182 39142 35594 39194
rect 35646 39142 35658 39194
rect 35710 39142 35722 39194
rect 35774 39142 35786 39194
rect 35838 39142 35850 39194
rect 35902 39142 38272 39194
rect 1104 39120 38272 39142
rect 14 39040 20 39092
rect 72 39080 78 39092
rect 1489 39083 1547 39089
rect 1489 39080 1501 39083
rect 72 39052 1501 39080
rect 72 39040 78 39052
rect 1489 39049 1501 39052
rect 1535 39049 1547 39083
rect 1489 39043 1547 39049
rect 4522 39040 4528 39092
rect 4580 39080 4586 39092
rect 4893 39083 4951 39089
rect 4893 39080 4905 39083
rect 4580 39052 4905 39080
rect 4580 39040 4586 39052
rect 4893 39049 4905 39052
rect 4939 39049 4951 39083
rect 4893 39043 4951 39049
rect 9030 39040 9036 39092
rect 9088 39080 9094 39092
rect 9309 39083 9367 39089
rect 9309 39080 9321 39083
rect 9088 39052 9321 39080
rect 9088 39040 9094 39052
rect 9309 39049 9321 39052
rect 9355 39049 9367 39083
rect 9309 39043 9367 39049
rect 11054 39040 11060 39092
rect 11112 39080 11118 39092
rect 11609 39083 11667 39089
rect 11609 39080 11621 39083
rect 11112 39052 11621 39080
rect 11112 39040 11118 39052
rect 11609 39049 11621 39052
rect 11655 39049 11667 39083
rect 11609 39043 11667 39049
rect 13170 39040 13176 39092
rect 13228 39040 13234 39092
rect 17402 39040 17408 39092
rect 17460 39080 17466 39092
rect 17773 39083 17831 39089
rect 17773 39080 17785 39083
rect 17460 39052 17785 39080
rect 17460 39040 17466 39052
rect 17773 39049 17785 39052
rect 17819 39049 17831 39083
rect 17773 39043 17831 39049
rect 21910 39040 21916 39092
rect 21968 39080 21974 39092
rect 22097 39083 22155 39089
rect 22097 39080 22109 39083
rect 21968 39052 22109 39080
rect 21968 39040 21974 39052
rect 22097 39049 22109 39052
rect 22143 39049 22155 39083
rect 22097 39043 22155 39049
rect 26418 39040 26424 39092
rect 26476 39080 26482 39092
rect 27157 39083 27215 39089
rect 27157 39080 27169 39083
rect 26476 39052 27169 39080
rect 26476 39040 26482 39052
rect 27157 39049 27169 39052
rect 27203 39049 27215 39083
rect 27157 39043 27215 39049
rect 33134 39040 33140 39092
rect 33192 39040 33198 39092
rect 35434 39040 35440 39092
rect 35492 39080 35498 39092
rect 35713 39083 35771 39089
rect 35713 39080 35725 39083
rect 35492 39052 35725 39080
rect 35492 39040 35498 39052
rect 35713 39049 35725 39052
rect 35759 39049 35771 39083
rect 35713 39043 35771 39049
rect 11885 39015 11943 39021
rect 11885 38981 11897 39015
rect 11931 39012 11943 39015
rect 12342 39012 12348 39024
rect 11931 38984 12348 39012
rect 11931 38981 11943 38984
rect 11885 38975 11943 38981
rect 12342 38972 12348 38984
rect 12400 38972 12406 39024
rect 15470 38972 15476 39024
rect 15528 39012 15534 39024
rect 15749 39015 15807 39021
rect 15749 39012 15761 39015
rect 15528 38984 15761 39012
rect 15528 38972 15534 38984
rect 15749 38981 15761 38984
rect 15795 38981 15807 39015
rect 15749 38975 15807 38981
rect 30926 38972 30932 39024
rect 30984 39012 30990 39024
rect 31205 39015 31263 39021
rect 31205 39012 31217 39015
rect 30984 38984 31217 39012
rect 30984 38972 30990 38984
rect 31205 38981 31217 38984
rect 31251 38981 31263 39015
rect 31205 38975 31263 38981
rect 1762 38904 1768 38956
rect 1820 38904 1826 38956
rect 5074 38904 5080 38956
rect 5132 38904 5138 38956
rect 9214 38904 9220 38956
rect 9272 38904 9278 38956
rect 12066 38904 12072 38956
rect 12124 38904 12130 38956
rect 12526 38904 12532 38956
rect 12584 38944 12590 38956
rect 12989 38947 13047 38953
rect 12989 38944 13001 38947
rect 12584 38916 13001 38944
rect 12584 38904 12590 38916
rect 12989 38913 13001 38916
rect 13035 38913 13047 38947
rect 12989 38907 13047 38913
rect 17954 38904 17960 38956
rect 18012 38904 18018 38956
rect 19426 38904 19432 38956
rect 19484 38904 19490 38956
rect 20070 38904 20076 38956
rect 20128 38904 20134 38956
rect 22370 38904 22376 38956
rect 22428 38904 22434 38956
rect 27062 38904 27068 38956
rect 27120 38904 27126 38956
rect 27706 38904 27712 38956
rect 27764 38904 27770 38956
rect 33042 38904 33048 38956
rect 33100 38904 33106 38956
rect 35618 38904 35624 38956
rect 35676 38904 35682 38956
rect 37366 38904 37372 38956
rect 37424 38944 37430 38956
rect 37461 38947 37519 38953
rect 37461 38944 37473 38947
rect 37424 38916 37473 38944
rect 37424 38904 37430 38916
rect 37461 38913 37473 38916
rect 37507 38913 37519 38947
rect 37461 38907 37519 38913
rect 13998 38836 14004 38888
rect 14056 38876 14062 38888
rect 20349 38879 20407 38885
rect 20349 38876 20361 38879
rect 14056 38848 20361 38876
rect 14056 38836 14062 38848
rect 20349 38845 20361 38848
rect 20395 38845 20407 38879
rect 20349 38839 20407 38845
rect 15562 38768 15568 38820
rect 15620 38768 15626 38820
rect 29730 38768 29736 38820
rect 29788 38808 29794 38820
rect 31021 38811 31079 38817
rect 31021 38808 31033 38811
rect 29788 38780 31033 38808
rect 29788 38768 29794 38780
rect 31021 38777 31033 38780
rect 31067 38777 31079 38811
rect 31021 38771 31079 38777
rect 37642 38768 37648 38820
rect 37700 38768 37706 38820
rect 12253 38743 12311 38749
rect 12253 38709 12265 38743
rect 12299 38740 12311 38743
rect 12802 38740 12808 38752
rect 12299 38712 12808 38740
rect 12299 38709 12311 38712
rect 12253 38703 12311 38709
rect 12802 38700 12808 38712
rect 12860 38700 12866 38752
rect 19610 38700 19616 38752
rect 19668 38700 19674 38752
rect 27614 38700 27620 38752
rect 27672 38700 27678 38752
rect 1104 38650 38272 38672
rect 1104 38598 4214 38650
rect 4266 38598 4278 38650
rect 4330 38598 4342 38650
rect 4394 38598 4406 38650
rect 4458 38598 4470 38650
rect 4522 38598 34934 38650
rect 34986 38598 34998 38650
rect 35050 38598 35062 38650
rect 35114 38598 35126 38650
rect 35178 38598 35190 38650
rect 35242 38598 38272 38650
rect 1104 38576 38272 38598
rect 4985 38539 5043 38545
rect 4985 38505 4997 38539
rect 5031 38536 5043 38539
rect 5074 38536 5080 38548
rect 5031 38508 5080 38536
rect 5031 38505 5043 38508
rect 4985 38499 5043 38505
rect 5074 38496 5080 38508
rect 5132 38496 5138 38548
rect 8757 38539 8815 38545
rect 8757 38505 8769 38539
rect 8803 38536 8815 38539
rect 9214 38536 9220 38548
rect 8803 38508 9220 38536
rect 8803 38505 8815 38508
rect 8757 38499 8815 38505
rect 9214 38496 9220 38508
rect 9272 38496 9278 38548
rect 17954 38496 17960 38548
rect 18012 38536 18018 38548
rect 18325 38539 18383 38545
rect 18325 38536 18337 38539
rect 18012 38508 18337 38536
rect 18012 38496 18018 38508
rect 18325 38505 18337 38508
rect 18371 38505 18383 38539
rect 22462 38536 22468 38548
rect 18325 38499 18383 38505
rect 18432 38508 22468 38536
rect 13630 38428 13636 38480
rect 13688 38468 13694 38480
rect 18432 38468 18460 38508
rect 22462 38496 22468 38508
rect 22520 38496 22526 38548
rect 27706 38536 27712 38548
rect 25056 38508 27712 38536
rect 13688 38440 18460 38468
rect 13688 38428 13694 38440
rect 12710 38360 12716 38412
rect 12768 38400 12774 38412
rect 19521 38403 19579 38409
rect 12768 38372 18920 38400
rect 12768 38360 12774 38372
rect 5166 38292 5172 38344
rect 5224 38292 5230 38344
rect 8570 38292 8576 38344
rect 8628 38292 8634 38344
rect 9030 38292 9036 38344
rect 9088 38292 9094 38344
rect 9125 38335 9183 38341
rect 9125 38301 9137 38335
rect 9171 38332 9183 38335
rect 9309 38335 9367 38341
rect 9309 38332 9321 38335
rect 9171 38304 9321 38332
rect 9171 38301 9183 38304
rect 9125 38295 9183 38301
rect 9309 38301 9321 38304
rect 9355 38301 9367 38335
rect 9309 38295 9367 38301
rect 13081 38335 13139 38341
rect 13081 38301 13093 38335
rect 13127 38332 13139 38335
rect 13265 38335 13323 38341
rect 13265 38332 13277 38335
rect 13127 38304 13277 38332
rect 13127 38301 13139 38304
rect 13081 38295 13139 38301
rect 13265 38301 13277 38304
rect 13311 38301 13323 38335
rect 13265 38295 13323 38301
rect 13357 38335 13415 38341
rect 13357 38301 13369 38335
rect 13403 38332 13415 38335
rect 13446 38332 13452 38344
rect 13403 38304 13452 38332
rect 13403 38301 13415 38304
rect 13357 38295 13415 38301
rect 13446 38292 13452 38304
rect 13504 38332 13510 38344
rect 13504 38304 18460 38332
rect 13504 38292 13510 38304
rect 9582 38224 9588 38276
rect 9640 38224 9646 38276
rect 10226 38224 10232 38276
rect 10284 38224 10290 38276
rect 10888 38236 11638 38264
rect 9122 38156 9128 38208
rect 9180 38196 9186 38208
rect 10888 38196 10916 38236
rect 12802 38224 12808 38276
rect 12860 38224 12866 38276
rect 9180 38168 10916 38196
rect 11057 38199 11115 38205
rect 9180 38156 9186 38168
rect 11057 38165 11069 38199
rect 11103 38196 11115 38199
rect 11238 38196 11244 38208
rect 11103 38168 11244 38196
rect 11103 38165 11115 38168
rect 11057 38159 11115 38165
rect 11238 38156 11244 38168
rect 11296 38156 11302 38208
rect 11330 38156 11336 38208
rect 11388 38156 11394 38208
rect 18432 38196 18460 38304
rect 18506 38292 18512 38344
rect 18564 38292 18570 38344
rect 18892 38341 18920 38372
rect 19521 38369 19533 38403
rect 19567 38400 19579 38403
rect 19610 38400 19616 38412
rect 19567 38372 19616 38400
rect 19567 38369 19579 38372
rect 19521 38363 19579 38369
rect 19610 38360 19616 38372
rect 19668 38360 19674 38412
rect 21192 38372 23244 38400
rect 21192 38344 21220 38372
rect 18877 38335 18935 38341
rect 18877 38301 18889 38335
rect 18923 38301 18935 38335
rect 18877 38295 18935 38301
rect 18969 38335 19027 38341
rect 18969 38301 18981 38335
rect 19015 38332 19027 38335
rect 19245 38335 19303 38341
rect 19245 38332 19257 38335
rect 19015 38304 19257 38332
rect 19015 38301 19027 38304
rect 18969 38295 19027 38301
rect 19245 38301 19257 38304
rect 19291 38301 19303 38335
rect 21174 38332 21180 38344
rect 20654 38304 21180 38332
rect 19245 38295 19303 38301
rect 21174 38292 21180 38304
rect 21232 38292 21238 38344
rect 21266 38292 21272 38344
rect 21324 38292 21330 38344
rect 21545 38335 21603 38341
rect 21545 38301 21557 38335
rect 21591 38301 21603 38335
rect 21545 38295 21603 38301
rect 21637 38335 21695 38341
rect 21637 38301 21649 38335
rect 21683 38332 21695 38335
rect 21821 38335 21879 38341
rect 21821 38332 21833 38335
rect 21683 38304 21833 38332
rect 21683 38301 21695 38304
rect 21637 38295 21695 38301
rect 21821 38301 21833 38304
rect 21867 38301 21879 38335
rect 23216 38332 23244 38372
rect 25056 38341 25084 38508
rect 27706 38496 27712 38508
rect 27764 38536 27770 38548
rect 32217 38539 32275 38545
rect 27764 38508 29592 38536
rect 27764 38496 27770 38508
rect 26050 38360 26056 38412
rect 26108 38400 26114 38412
rect 27249 38403 27307 38409
rect 26108 38372 27200 38400
rect 26108 38360 26114 38372
rect 25041 38335 25099 38341
rect 23216 38318 24992 38332
rect 23230 38304 24992 38318
rect 21821 38295 21879 38301
rect 21560 38264 21588 38295
rect 20824 38236 21588 38264
rect 22097 38267 22155 38273
rect 20824 38196 20852 38236
rect 22097 38233 22109 38267
rect 22143 38233 22155 38267
rect 22097 38227 22155 38233
rect 18432 38168 20852 38196
rect 20990 38156 20996 38208
rect 21048 38156 21054 38208
rect 21453 38199 21511 38205
rect 21453 38165 21465 38199
rect 21499 38196 21511 38199
rect 22112 38196 22140 38227
rect 21499 38168 22140 38196
rect 21499 38165 21511 38168
rect 21453 38159 21511 38165
rect 23474 38156 23480 38208
rect 23532 38196 23538 38208
rect 23569 38199 23627 38205
rect 23569 38196 23581 38199
rect 23532 38168 23581 38196
rect 23532 38156 23538 38168
rect 23569 38165 23581 38168
rect 23615 38165 23627 38199
rect 24964 38196 24992 38304
rect 25041 38301 25053 38335
rect 25087 38301 25099 38335
rect 25041 38295 25099 38301
rect 25133 38335 25191 38341
rect 25133 38301 25145 38335
rect 25179 38332 25191 38335
rect 25317 38335 25375 38341
rect 25317 38332 25329 38335
rect 25179 38304 25329 38332
rect 25179 38301 25191 38304
rect 25133 38295 25191 38301
rect 25317 38301 25329 38304
rect 25363 38301 25375 38335
rect 25317 38295 25375 38301
rect 25590 38224 25596 38276
rect 25648 38224 25654 38276
rect 26050 38264 26056 38276
rect 25976 38236 26056 38264
rect 25976 38196 26004 38236
rect 26050 38224 26056 38236
rect 26108 38224 26114 38276
rect 24964 38168 26004 38196
rect 23569 38159 23627 38165
rect 26510 38156 26516 38208
rect 26568 38196 26574 38208
rect 27065 38199 27123 38205
rect 27065 38196 27077 38199
rect 26568 38168 27077 38196
rect 26568 38156 26574 38168
rect 27065 38165 27077 38168
rect 27111 38165 27123 38199
rect 27172 38196 27200 38372
rect 27249 38369 27261 38403
rect 27295 38400 27307 38403
rect 27614 38400 27620 38412
rect 27295 38372 27620 38400
rect 27295 38369 27307 38372
rect 27249 38363 27307 38369
rect 27614 38360 27620 38372
rect 27672 38360 27678 38412
rect 29564 38344 29592 38508
rect 32217 38505 32229 38539
rect 32263 38536 32275 38539
rect 33042 38536 33048 38548
rect 32263 38508 33048 38536
rect 32263 38505 32275 38508
rect 32217 38499 32275 38505
rect 33042 38496 33048 38508
rect 33100 38496 33106 38548
rect 34885 38539 34943 38545
rect 34885 38505 34897 38539
rect 34931 38536 34943 38539
rect 35618 38536 35624 38548
rect 34931 38508 35624 38536
rect 34931 38505 34943 38508
rect 34885 38499 34943 38505
rect 35618 38496 35624 38508
rect 35676 38496 35682 38548
rect 37829 38539 37887 38545
rect 37829 38505 37841 38539
rect 37875 38536 37887 38539
rect 37918 38536 37924 38548
rect 37875 38508 37924 38536
rect 37875 38505 37887 38508
rect 37829 38499 37887 38505
rect 37918 38496 37924 38508
rect 37976 38496 37982 38548
rect 29638 38360 29644 38412
rect 29696 38360 29702 38412
rect 29546 38292 29552 38344
rect 29604 38292 29610 38344
rect 32033 38335 32091 38341
rect 32033 38332 32045 38335
rect 29656 38304 32045 38332
rect 27522 38224 27528 38276
rect 27580 38224 27586 38276
rect 27908 38236 28014 38264
rect 27908 38196 27936 38236
rect 29270 38224 29276 38276
rect 29328 38224 29334 38276
rect 29454 38224 29460 38276
rect 29512 38264 29518 38276
rect 29656 38264 29684 38304
rect 32033 38301 32045 38304
rect 32079 38301 32091 38335
rect 32033 38295 32091 38301
rect 34701 38335 34759 38341
rect 34701 38301 34713 38335
rect 34747 38301 34759 38335
rect 34701 38295 34759 38301
rect 29512 38236 29684 38264
rect 29512 38224 29518 38236
rect 31662 38224 31668 38276
rect 31720 38264 31726 38276
rect 34716 38264 34744 38295
rect 31720 38236 34744 38264
rect 37553 38267 37611 38273
rect 31720 38224 31726 38236
rect 37553 38233 37565 38267
rect 37599 38233 37611 38267
rect 37553 38227 37611 38233
rect 28534 38196 28540 38208
rect 27172 38168 28540 38196
rect 27065 38159 27123 38165
rect 28534 38156 28540 38168
rect 28592 38196 28598 38208
rect 30374 38196 30380 38208
rect 28592 38168 30380 38196
rect 28592 38156 28598 38168
rect 30374 38156 30380 38168
rect 30432 38156 30438 38208
rect 31110 38156 31116 38208
rect 31168 38196 31174 38208
rect 37568 38196 37596 38227
rect 31168 38168 37596 38196
rect 31168 38156 31174 38168
rect 1104 38106 38272 38128
rect 1104 38054 4874 38106
rect 4926 38054 4938 38106
rect 4990 38054 5002 38106
rect 5054 38054 5066 38106
rect 5118 38054 5130 38106
rect 5182 38054 35594 38106
rect 35646 38054 35658 38106
rect 35710 38054 35722 38106
rect 35774 38054 35786 38106
rect 35838 38054 35850 38106
rect 35902 38054 38272 38106
rect 1104 38032 38272 38054
rect 9582 37952 9588 38004
rect 9640 37992 9646 38004
rect 9769 37995 9827 38001
rect 9769 37992 9781 37995
rect 9640 37964 9781 37992
rect 9640 37952 9646 37964
rect 9769 37961 9781 37964
rect 9815 37961 9827 37995
rect 9769 37955 9827 37961
rect 10229 37995 10287 38001
rect 10229 37961 10241 37995
rect 10275 37961 10287 37995
rect 10229 37955 10287 37961
rect 9953 37859 10011 37865
rect 9953 37825 9965 37859
rect 9999 37856 10011 37859
rect 10244 37856 10272 37955
rect 11330 37952 11336 38004
rect 11388 37992 11394 38004
rect 11882 37992 11888 38004
rect 11388 37964 11888 37992
rect 11388 37952 11394 37964
rect 11882 37952 11888 37964
rect 11940 37952 11946 38004
rect 12066 37952 12072 38004
rect 12124 37992 12130 38004
rect 12253 37995 12311 38001
rect 12253 37992 12265 37995
rect 12124 37964 12265 37992
rect 12124 37952 12130 37964
rect 12253 37961 12265 37964
rect 12299 37961 12311 37995
rect 12253 37955 12311 37961
rect 12342 37952 12348 38004
rect 12400 37952 12406 38004
rect 13630 37952 13636 38004
rect 13688 37952 13694 38004
rect 13740 37964 15332 37992
rect 13648 37924 13676 37952
rect 11716 37896 13676 37924
rect 9999 37828 10272 37856
rect 10597 37859 10655 37865
rect 9999 37825 10011 37828
rect 9953 37819 10011 37825
rect 10597 37825 10609 37859
rect 10643 37856 10655 37859
rect 11238 37856 11244 37868
rect 10643 37828 11244 37856
rect 10643 37825 10655 37828
rect 10597 37819 10655 37825
rect 11238 37816 11244 37828
rect 11296 37816 11302 37868
rect 10689 37791 10747 37797
rect 10689 37788 10701 37791
rect 10612 37760 10701 37788
rect 10612 37664 10640 37760
rect 10689 37757 10701 37760
rect 10735 37757 10747 37791
rect 10689 37751 10747 37757
rect 10778 37748 10784 37800
rect 10836 37748 10842 37800
rect 11716 37797 11744 37896
rect 12529 37859 12587 37865
rect 12529 37825 12541 37859
rect 12575 37856 12587 37859
rect 13170 37856 13176 37868
rect 12575 37828 13176 37856
rect 12575 37825 12587 37828
rect 12529 37819 12587 37825
rect 13170 37816 13176 37828
rect 13228 37816 13234 37868
rect 13740 37865 13768 37964
rect 13909 37927 13967 37933
rect 13909 37893 13921 37927
rect 13955 37924 13967 37927
rect 13955 37896 14688 37924
rect 13955 37893 13967 37896
rect 13909 37887 13967 37893
rect 13265 37859 13323 37865
rect 13265 37825 13277 37859
rect 13311 37825 13323 37859
rect 13265 37819 13323 37825
rect 13725 37859 13783 37865
rect 13725 37825 13737 37859
rect 13771 37825 13783 37859
rect 13725 37819 13783 37825
rect 11701 37791 11759 37797
rect 11701 37757 11713 37791
rect 11747 37757 11759 37791
rect 11701 37751 11759 37757
rect 11793 37791 11851 37797
rect 11793 37757 11805 37791
rect 11839 37757 11851 37791
rect 11793 37751 11851 37757
rect 10594 37612 10600 37664
rect 10652 37652 10658 37664
rect 11808 37652 11836 37751
rect 11882 37748 11888 37800
rect 11940 37748 11946 37800
rect 13078 37748 13084 37800
rect 13136 37788 13142 37800
rect 13280 37788 13308 37819
rect 13814 37816 13820 37868
rect 13872 37816 13878 37868
rect 14090 37865 14096 37868
rect 14047 37859 14096 37865
rect 14047 37825 14059 37859
rect 14093 37825 14096 37859
rect 14047 37819 14096 37825
rect 14090 37816 14096 37819
rect 14148 37816 14154 37868
rect 14366 37865 14372 37868
rect 14364 37819 14372 37865
rect 14366 37816 14372 37819
rect 14424 37816 14430 37868
rect 14461 37859 14519 37865
rect 14461 37825 14473 37859
rect 14507 37825 14519 37859
rect 14461 37819 14519 37825
rect 14553 37859 14611 37865
rect 14553 37825 14565 37859
rect 14599 37825 14611 37859
rect 14553 37819 14611 37825
rect 13136 37760 13308 37788
rect 13357 37791 13415 37797
rect 13136 37748 13142 37760
rect 13357 37757 13369 37791
rect 13403 37788 13415 37791
rect 14185 37791 14243 37797
rect 14185 37788 14197 37791
rect 13403 37760 14197 37788
rect 13403 37757 13415 37760
rect 13357 37751 13415 37757
rect 14185 37757 14197 37760
rect 14231 37757 14243 37791
rect 14185 37751 14243 37757
rect 11900 37720 11928 37748
rect 13262 37720 13268 37732
rect 11900 37692 13268 37720
rect 13262 37680 13268 37692
rect 13320 37720 13326 37732
rect 14476 37720 14504 37819
rect 13320 37692 14504 37720
rect 14568 37720 14596 37819
rect 14660 37797 14688 37896
rect 15304 37868 15332 37964
rect 15948 37964 18000 37992
rect 15948 37868 15976 37964
rect 16942 37924 16948 37936
rect 16316 37896 16948 37924
rect 14737 37859 14795 37865
rect 14737 37825 14749 37859
rect 14783 37825 14795 37859
rect 14737 37819 14795 37825
rect 14645 37791 14703 37797
rect 14645 37757 14657 37791
rect 14691 37757 14703 37791
rect 14752 37788 14780 37819
rect 15286 37816 15292 37868
rect 15344 37816 15350 37868
rect 15930 37816 15936 37868
rect 15988 37816 15994 37868
rect 16114 37816 16120 37868
rect 16172 37816 16178 37868
rect 16206 37816 16212 37868
rect 16264 37816 16270 37868
rect 16316 37865 16344 37896
rect 16942 37884 16948 37896
rect 17000 37884 17006 37936
rect 17037 37927 17095 37933
rect 17037 37893 17049 37927
rect 17083 37924 17095 37927
rect 17405 37927 17463 37933
rect 17405 37924 17417 37927
rect 17083 37896 17417 37924
rect 17083 37893 17095 37896
rect 17037 37887 17095 37893
rect 17405 37893 17417 37896
rect 17451 37893 17463 37927
rect 17405 37887 17463 37893
rect 17512 37896 17908 37924
rect 16301 37859 16359 37865
rect 16301 37825 16313 37859
rect 16347 37825 16359 37859
rect 16301 37819 16359 37825
rect 16390 37816 16396 37868
rect 16448 37856 16454 37868
rect 16669 37859 16727 37865
rect 16669 37856 16681 37859
rect 16448 37828 16681 37856
rect 16448 37816 16454 37828
rect 16669 37825 16681 37828
rect 16715 37825 16727 37859
rect 16669 37819 16727 37825
rect 16850 37816 16856 37868
rect 16908 37816 16914 37868
rect 17221 37859 17279 37865
rect 17221 37825 17233 37859
rect 17267 37856 17279 37859
rect 17310 37856 17316 37868
rect 17267 37828 17316 37856
rect 17267 37825 17279 37828
rect 17221 37819 17279 37825
rect 17310 37816 17316 37828
rect 17368 37816 17374 37868
rect 17512 37865 17540 37896
rect 17880 37868 17908 37896
rect 17497 37859 17555 37865
rect 17497 37825 17509 37859
rect 17543 37825 17555 37859
rect 17497 37819 17555 37825
rect 17589 37859 17647 37865
rect 17589 37825 17601 37859
rect 17635 37856 17647 37859
rect 17770 37856 17776 37868
rect 17635 37828 17776 37856
rect 17635 37825 17647 37828
rect 17589 37819 17647 37825
rect 17512 37788 17540 37819
rect 17770 37816 17776 37828
rect 17828 37816 17834 37868
rect 17862 37816 17868 37868
rect 17920 37816 17926 37868
rect 14752 37760 17540 37788
rect 14645 37751 14703 37757
rect 15378 37720 15384 37732
rect 14568 37692 15384 37720
rect 13320 37680 13326 37692
rect 10652 37624 11836 37652
rect 10652 37612 10658 37624
rect 12434 37612 12440 37664
rect 12492 37652 12498 37664
rect 13541 37655 13599 37661
rect 13541 37652 13553 37655
rect 12492 37624 13553 37652
rect 12492 37612 12498 37624
rect 13541 37621 13553 37624
rect 13587 37621 13599 37655
rect 14476 37652 14504 37692
rect 15378 37680 15384 37692
rect 15436 37680 15442 37732
rect 16850 37720 16856 37732
rect 15488 37692 16856 37720
rect 15488 37652 15516 37692
rect 16850 37680 16856 37692
rect 16908 37680 16914 37732
rect 14476 37624 15516 37652
rect 13541 37615 13599 37621
rect 16482 37612 16488 37664
rect 16540 37612 16546 37664
rect 17770 37612 17776 37664
rect 17828 37612 17834 37664
rect 17972 37652 18000 37964
rect 18506 37952 18512 38004
rect 18564 37952 18570 38004
rect 19426 37952 19432 38004
rect 19484 37952 19490 38004
rect 19797 37995 19855 38001
rect 19797 37961 19809 37995
rect 19843 37992 19855 37995
rect 20990 37992 20996 38004
rect 19843 37964 20996 37992
rect 19843 37961 19855 37964
rect 19797 37955 19855 37961
rect 20990 37952 20996 37964
rect 21048 37952 21054 38004
rect 21266 37952 21272 38004
rect 21324 37992 21330 38004
rect 22005 37995 22063 38001
rect 22005 37992 22017 37995
rect 21324 37964 22017 37992
rect 21324 37952 21330 37964
rect 22005 37961 22017 37964
rect 22051 37961 22063 37995
rect 22005 37955 22063 37961
rect 22373 37995 22431 38001
rect 22373 37961 22385 37995
rect 22419 37992 22431 37995
rect 22419 37964 23520 37992
rect 22419 37961 22431 37964
rect 22373 37955 22431 37961
rect 18524 37924 18552 37952
rect 18524 37896 20484 37924
rect 20346 37816 20352 37868
rect 20404 37816 20410 37868
rect 20456 37856 20484 37896
rect 20530 37884 20536 37936
rect 20588 37924 20594 37936
rect 20588 37896 22508 37924
rect 20588 37884 20594 37896
rect 20456 37828 22094 37856
rect 19334 37748 19340 37800
rect 19392 37788 19398 37800
rect 19889 37791 19947 37797
rect 19889 37788 19901 37791
rect 19392 37760 19901 37788
rect 19392 37748 19398 37760
rect 19889 37757 19901 37760
rect 19935 37757 19947 37791
rect 19889 37751 19947 37757
rect 19904 37720 19932 37751
rect 19978 37748 19984 37800
rect 20036 37748 20042 37800
rect 20901 37791 20959 37797
rect 20901 37757 20913 37791
rect 20947 37788 20959 37791
rect 21174 37788 21180 37800
rect 20947 37760 21180 37788
rect 20947 37757 20959 37760
rect 20901 37751 20959 37757
rect 21174 37748 21180 37760
rect 21232 37748 21238 37800
rect 20530 37720 20536 37732
rect 19904 37692 20536 37720
rect 20530 37680 20536 37692
rect 20588 37680 20594 37732
rect 22066 37720 22094 37828
rect 22480 37800 22508 37896
rect 23492 37868 23520 37964
rect 25590 37952 25596 38004
rect 25648 37992 25654 38004
rect 26237 37995 26295 38001
rect 26237 37992 26249 37995
rect 25648 37964 26249 37992
rect 25648 37952 25654 37964
rect 26237 37961 26249 37964
rect 26283 37961 26295 37995
rect 26237 37955 26295 37961
rect 26789 37995 26847 38001
rect 26789 37961 26801 37995
rect 26835 37992 26847 37995
rect 27522 37992 27528 38004
rect 26835 37964 27528 37992
rect 26835 37961 26847 37964
rect 26789 37955 26847 37961
rect 27522 37952 27528 37964
rect 27580 37952 27586 38004
rect 28353 37995 28411 38001
rect 28353 37961 28365 37995
rect 28399 37992 28411 37995
rect 29454 37992 29460 38004
rect 28399 37964 29460 37992
rect 28399 37961 28411 37964
rect 28353 37955 28411 37961
rect 29454 37952 29460 37964
rect 29512 37952 29518 38004
rect 29638 37952 29644 38004
rect 29696 37952 29702 38004
rect 23569 37927 23627 37933
rect 23569 37893 23581 37927
rect 23615 37924 23627 37927
rect 24397 37927 24455 37933
rect 24397 37924 24409 37927
rect 23615 37896 24409 37924
rect 23615 37893 23627 37896
rect 23569 37887 23627 37893
rect 24397 37893 24409 37896
rect 24443 37893 24455 37927
rect 24397 37887 24455 37893
rect 25056 37896 25544 37924
rect 23014 37816 23020 37868
rect 23072 37856 23078 37868
rect 23385 37859 23443 37865
rect 23385 37856 23397 37859
rect 23072 37828 23397 37856
rect 23072 37816 23078 37828
rect 23385 37825 23397 37828
rect 23431 37825 23443 37859
rect 23385 37819 23443 37825
rect 23474 37816 23480 37868
rect 23532 37816 23538 37868
rect 23658 37816 23664 37868
rect 23716 37816 23722 37868
rect 23753 37859 23811 37865
rect 23753 37825 23765 37859
rect 23799 37856 23811 37859
rect 23934 37856 23940 37868
rect 23799 37828 23940 37856
rect 23799 37825 23811 37828
rect 23753 37819 23811 37825
rect 23934 37816 23940 37828
rect 23992 37816 23998 37868
rect 24029 37859 24087 37865
rect 24029 37825 24041 37859
rect 24075 37856 24087 37859
rect 24118 37856 24124 37868
rect 24075 37828 24124 37856
rect 24075 37825 24087 37828
rect 24029 37819 24087 37825
rect 24118 37816 24124 37828
rect 24176 37816 24182 37868
rect 25056 37865 25084 37896
rect 24213 37859 24271 37865
rect 24213 37825 24225 37859
rect 24259 37825 24271 37859
rect 24213 37819 24271 37825
rect 25041 37859 25099 37865
rect 25041 37825 25053 37859
rect 25087 37825 25099 37859
rect 25041 37819 25099 37825
rect 22462 37748 22468 37800
rect 22520 37748 22526 37800
rect 22554 37748 22560 37800
rect 22612 37748 22618 37800
rect 23492 37788 23520 37816
rect 24228 37788 24256 37819
rect 25314 37816 25320 37868
rect 25372 37816 25378 37868
rect 25516 37865 25544 37896
rect 25774 37884 25780 37936
rect 25832 37884 25838 37936
rect 29656 37924 29684 37952
rect 25976 37896 27752 37924
rect 25501 37859 25559 37865
rect 25501 37825 25513 37859
rect 25547 37856 25559 37859
rect 25866 37856 25872 37868
rect 25547 37828 25872 37856
rect 25547 37825 25559 37828
rect 25501 37819 25559 37825
rect 25866 37816 25872 37828
rect 25924 37856 25930 37868
rect 25976 37865 26004 37896
rect 25961 37859 26019 37865
rect 25961 37856 25973 37859
rect 25924 37828 25973 37856
rect 25924 37816 25930 37828
rect 25961 37825 25973 37828
rect 26007 37825 26019 37859
rect 25961 37819 26019 37825
rect 26053 37859 26111 37865
rect 26053 37825 26065 37859
rect 26099 37825 26111 37859
rect 26053 37819 26111 37825
rect 23492 37760 24256 37788
rect 25222 37748 25228 37800
rect 25280 37748 25286 37800
rect 25685 37791 25743 37797
rect 25685 37757 25697 37791
rect 25731 37788 25743 37791
rect 26068 37788 26096 37819
rect 26418 37816 26424 37868
rect 26476 37816 26482 37868
rect 26602 37816 26608 37868
rect 26660 37816 26666 37868
rect 27724 37865 27752 37896
rect 29104 37896 29684 37924
rect 27709 37859 27767 37865
rect 27709 37825 27721 37859
rect 27755 37856 27767 37859
rect 28169 37859 28227 37865
rect 28169 37856 28181 37859
rect 27755 37828 28181 37856
rect 27755 37825 27767 37828
rect 27709 37819 27767 37825
rect 28169 37825 28181 37828
rect 28215 37825 28227 37859
rect 28169 37819 28227 37825
rect 28813 37859 28871 37865
rect 28813 37825 28825 37859
rect 28859 37856 28871 37859
rect 28994 37856 29000 37868
rect 28859 37828 29000 37856
rect 28859 37825 28871 37828
rect 28813 37819 28871 37825
rect 28994 37816 29000 37828
rect 29052 37816 29058 37868
rect 29104 37865 29132 37896
rect 30374 37884 30380 37936
rect 30432 37884 30438 37936
rect 29089 37859 29147 37865
rect 29089 37825 29101 37859
rect 29135 37825 29147 37859
rect 29089 37819 29147 37825
rect 31202 37816 31208 37868
rect 31260 37816 31266 37868
rect 26142 37788 26148 37800
rect 25731 37760 26004 37788
rect 26068 37760 26148 37788
rect 25731 37757 25743 37760
rect 25685 37751 25743 37757
rect 24857 37723 24915 37729
rect 24857 37720 24869 37723
rect 22066 37692 24869 37720
rect 24857 37689 24869 37692
rect 24903 37689 24915 37723
rect 24857 37683 24915 37689
rect 25976 37664 26004 37760
rect 26142 37748 26148 37760
rect 26200 37748 26206 37800
rect 27062 37748 27068 37800
rect 27120 37788 27126 37800
rect 27525 37791 27583 37797
rect 27525 37788 27537 37791
rect 27120 37760 27537 37788
rect 27120 37748 27126 37760
rect 27525 37757 27537 37760
rect 27571 37757 27583 37791
rect 27525 37751 27583 37757
rect 27982 37748 27988 37800
rect 28040 37748 28046 37800
rect 29365 37791 29423 37797
rect 29365 37788 29377 37791
rect 29012 37760 29377 37788
rect 29012 37729 29040 37760
rect 29365 37757 29377 37760
rect 29411 37757 29423 37791
rect 29365 37751 29423 37757
rect 29454 37748 29460 37800
rect 29512 37788 29518 37800
rect 30837 37791 30895 37797
rect 30837 37788 30849 37791
rect 29512 37760 30849 37788
rect 29512 37748 29518 37760
rect 30837 37757 30849 37760
rect 30883 37757 30895 37791
rect 30837 37751 30895 37757
rect 31662 37748 31668 37800
rect 31720 37748 31726 37800
rect 28997 37723 29055 37729
rect 28997 37689 29009 37723
rect 29043 37689 29055 37723
rect 31680 37720 31708 37748
rect 28997 37683 29055 37689
rect 30392 37692 31708 37720
rect 23842 37652 23848 37664
rect 17972 37624 23848 37652
rect 23842 37612 23848 37624
rect 23900 37612 23906 37664
rect 23937 37655 23995 37661
rect 23937 37621 23949 37655
rect 23983 37652 23995 37655
rect 24578 37652 24584 37664
rect 23983 37624 24584 37652
rect 23983 37621 23995 37624
rect 23937 37615 23995 37621
rect 24578 37612 24584 37624
rect 24636 37612 24642 37664
rect 25958 37612 25964 37664
rect 26016 37612 26022 37664
rect 27893 37655 27951 37661
rect 27893 37621 27905 37655
rect 27939 37652 27951 37655
rect 30392 37652 30420 37692
rect 27939 37624 30420 37652
rect 27939 37621 27951 37624
rect 27893 37615 27951 37621
rect 30926 37612 30932 37664
rect 30984 37652 30990 37664
rect 31021 37655 31079 37661
rect 31021 37652 31033 37655
rect 30984 37624 31033 37652
rect 30984 37612 30990 37624
rect 31021 37621 31033 37624
rect 31067 37621 31079 37655
rect 31021 37615 31079 37621
rect 1104 37562 38272 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 38272 37562
rect 1104 37488 38272 37510
rect 16482 37408 16488 37460
rect 16540 37448 16546 37460
rect 17773 37451 17831 37457
rect 17773 37448 17785 37451
rect 16540 37420 17785 37448
rect 16540 37408 16546 37420
rect 17773 37417 17785 37420
rect 17819 37417 17831 37451
rect 17773 37411 17831 37417
rect 20346 37408 20352 37460
rect 20404 37408 20410 37460
rect 23845 37451 23903 37457
rect 23845 37417 23857 37451
rect 23891 37448 23903 37451
rect 24670 37448 24676 37460
rect 23891 37420 24676 37448
rect 23891 37417 23903 37420
rect 23845 37411 23903 37417
rect 24670 37408 24676 37420
rect 24728 37408 24734 37460
rect 26053 37451 26111 37457
rect 26053 37417 26065 37451
rect 26099 37448 26111 37451
rect 26418 37448 26424 37460
rect 26099 37420 26424 37448
rect 26099 37417 26111 37420
rect 26053 37411 26111 37417
rect 26418 37408 26424 37420
rect 26476 37408 26482 37460
rect 26602 37408 26608 37460
rect 26660 37448 26666 37460
rect 27341 37451 27399 37457
rect 27341 37448 27353 37451
rect 26660 37420 27353 37448
rect 26660 37408 26666 37420
rect 27341 37417 27353 37420
rect 27387 37417 27399 37451
rect 27341 37411 27399 37417
rect 20364 37380 20392 37408
rect 12406 37352 20392 37380
rect 22066 37352 26832 37380
rect 1673 37315 1731 37321
rect 1673 37281 1685 37315
rect 1719 37312 1731 37315
rect 8386 37312 8392 37324
rect 1719 37284 8392 37312
rect 1719 37281 1731 37284
rect 1673 37275 1731 37281
rect 8386 37272 8392 37284
rect 8444 37312 8450 37324
rect 12406 37312 12434 37352
rect 8444 37284 12434 37312
rect 8444 37272 8450 37284
rect 17770 37272 17776 37324
rect 17828 37312 17834 37324
rect 17865 37315 17923 37321
rect 17865 37312 17877 37315
rect 17828 37284 17877 37312
rect 17828 37272 17834 37284
rect 17865 37281 17877 37284
rect 17911 37281 17923 37315
rect 17865 37275 17923 37281
rect 17954 37272 17960 37324
rect 18012 37312 18018 37324
rect 22066 37312 22094 37352
rect 18012 37284 22094 37312
rect 22189 37315 22247 37321
rect 18012 37272 18018 37284
rect 22189 37281 22201 37315
rect 22235 37312 22247 37315
rect 22830 37312 22836 37324
rect 22235 37284 22836 37312
rect 22235 37281 22247 37284
rect 22189 37275 22247 37281
rect 22830 37272 22836 37284
rect 22888 37272 22894 37324
rect 22922 37272 22928 37324
rect 22980 37272 22986 37324
rect 23842 37272 23848 37324
rect 23900 37312 23906 37324
rect 24854 37312 24860 37324
rect 23900 37284 24860 37312
rect 23900 37272 23906 37284
rect 24854 37272 24860 37284
rect 24912 37312 24918 37324
rect 26510 37312 26516 37324
rect 24912 37284 26516 37312
rect 24912 37272 24918 37284
rect 8294 37204 8300 37256
rect 8352 37204 8358 37256
rect 8573 37247 8631 37253
rect 8573 37213 8585 37247
rect 8619 37213 8631 37247
rect 8573 37207 8631 37213
rect 8665 37247 8723 37253
rect 8665 37213 8677 37247
rect 8711 37244 8723 37247
rect 8941 37247 8999 37253
rect 8941 37244 8953 37247
rect 8711 37216 8953 37244
rect 8711 37213 8723 37216
rect 8665 37207 8723 37213
rect 8941 37213 8953 37216
rect 8987 37213 8999 37247
rect 8941 37207 8999 37213
rect 934 37136 940 37188
rect 992 37176 998 37188
rect 1489 37179 1547 37185
rect 1489 37176 1501 37179
rect 992 37148 1501 37176
rect 992 37136 998 37148
rect 1489 37145 1501 37148
rect 1535 37145 1547 37179
rect 1489 37139 1547 37145
rect 6914 37136 6920 37188
rect 6972 37176 6978 37188
rect 8588 37176 8616 37207
rect 10226 37204 10232 37256
rect 10284 37244 10290 37256
rect 18049 37247 18107 37253
rect 10284 37216 10350 37244
rect 10284 37204 10290 37216
rect 18049 37213 18061 37247
rect 18095 37244 18107 37247
rect 18325 37247 18383 37253
rect 18325 37244 18337 37247
rect 18095 37216 18337 37244
rect 18095 37213 18107 37216
rect 18049 37207 18107 37213
rect 18325 37213 18337 37216
rect 18371 37213 18383 37247
rect 18325 37207 18383 37213
rect 18509 37247 18567 37253
rect 18509 37213 18521 37247
rect 18555 37213 18567 37247
rect 18509 37207 18567 37213
rect 6972 37148 8616 37176
rect 9217 37179 9275 37185
rect 6972 37136 6978 37148
rect 9217 37145 9229 37179
rect 9263 37145 9275 37179
rect 9217 37139 9275 37145
rect 8481 37111 8539 37117
rect 8481 37077 8493 37111
rect 8527 37108 8539 37111
rect 9232 37108 9260 37139
rect 17770 37136 17776 37188
rect 17828 37136 17834 37188
rect 18524 37176 18552 37207
rect 18598 37204 18604 37256
rect 18656 37204 18662 37256
rect 20162 37204 20168 37256
rect 20220 37204 20226 37256
rect 20257 37247 20315 37253
rect 20257 37213 20269 37247
rect 20303 37244 20315 37247
rect 20441 37247 20499 37253
rect 20441 37244 20453 37247
rect 20303 37216 20453 37244
rect 20303 37213 20315 37216
rect 20257 37207 20315 37213
rect 20441 37213 20453 37216
rect 20487 37213 20499 37247
rect 20441 37207 20499 37213
rect 22462 37204 22468 37256
rect 22520 37244 22526 37256
rect 22741 37247 22799 37253
rect 22741 37244 22753 37247
rect 22520 37216 22753 37244
rect 22520 37204 22526 37216
rect 22741 37213 22753 37216
rect 22787 37213 22799 37247
rect 22741 37207 22799 37213
rect 23293 37247 23351 37253
rect 23293 37213 23305 37247
rect 23339 37244 23351 37247
rect 23382 37244 23388 37256
rect 23339 37216 23388 37244
rect 23339 37213 23351 37216
rect 23293 37207 23351 37213
rect 23382 37204 23388 37216
rect 23440 37204 23446 37256
rect 23661 37247 23719 37253
rect 23661 37213 23673 37247
rect 23707 37244 23719 37247
rect 24026 37244 24032 37256
rect 23707 37216 24032 37244
rect 23707 37213 23719 37216
rect 23661 37207 23719 37213
rect 24026 37204 24032 37216
rect 24084 37244 24090 37256
rect 24302 37244 24308 37256
rect 24084 37216 24308 37244
rect 24084 37204 24090 37216
rect 24302 37204 24308 37216
rect 24360 37204 24366 37256
rect 26436 37253 26464 37284
rect 26510 37272 26516 37284
rect 26568 37272 26574 37324
rect 26605 37315 26663 37321
rect 26605 37281 26617 37315
rect 26651 37281 26663 37315
rect 26605 37275 26663 37281
rect 26421 37247 26479 37253
rect 26421 37213 26433 37247
rect 26467 37213 26479 37247
rect 26421 37207 26479 37213
rect 19886 37176 19892 37188
rect 18156 37148 19892 37176
rect 8527 37080 9260 37108
rect 8527 37077 8539 37080
rect 8481 37071 8539 37077
rect 10686 37068 10692 37120
rect 10744 37068 10750 37120
rect 17218 37068 17224 37120
rect 17276 37108 17282 37120
rect 18156 37108 18184 37148
rect 19886 37136 19892 37148
rect 19944 37136 19950 37188
rect 20714 37136 20720 37188
rect 20772 37136 20778 37188
rect 21174 37136 21180 37188
rect 21232 37136 21238 37188
rect 23477 37179 23535 37185
rect 23477 37145 23489 37179
rect 23523 37145 23535 37179
rect 23477 37139 23535 37145
rect 23569 37179 23627 37185
rect 23569 37145 23581 37179
rect 23615 37176 23627 37179
rect 23750 37176 23756 37188
rect 23615 37148 23756 37176
rect 23615 37145 23627 37148
rect 23569 37139 23627 37145
rect 17276 37080 18184 37108
rect 18233 37111 18291 37117
rect 17276 37068 17282 37080
rect 18233 37077 18245 37111
rect 18279 37108 18291 37111
rect 18966 37108 18972 37120
rect 18279 37080 18972 37108
rect 18279 37077 18291 37080
rect 18233 37071 18291 37077
rect 18966 37068 18972 37080
rect 19024 37068 19030 37120
rect 22370 37068 22376 37120
rect 22428 37068 22434 37120
rect 23492 37108 23520 37139
rect 23750 37136 23756 37148
rect 23808 37136 23814 37188
rect 26620 37176 26648 37275
rect 26804 37244 26832 37352
rect 27985 37315 28043 37321
rect 27985 37281 27997 37315
rect 28031 37312 28043 37315
rect 28626 37312 28632 37324
rect 28031 37284 28632 37312
rect 28031 37281 28043 37284
rect 27985 37275 28043 37281
rect 28626 37272 28632 37284
rect 28684 37272 28690 37324
rect 28902 37272 28908 37324
rect 28960 37312 28966 37324
rect 29546 37312 29552 37324
rect 28960 37284 29552 37312
rect 28960 37272 28966 37284
rect 29546 37272 29552 37284
rect 29604 37312 29610 37324
rect 30193 37315 30251 37321
rect 29604 37284 29684 37312
rect 29604 37272 29610 37284
rect 27338 37244 27344 37256
rect 26804 37216 27344 37244
rect 27338 37204 27344 37216
rect 27396 37244 27402 37256
rect 27801 37247 27859 37253
rect 27801 37244 27813 37247
rect 27396 37216 27813 37244
rect 27396 37204 27402 37216
rect 27801 37213 27813 37216
rect 27847 37244 27859 37247
rect 29270 37244 29276 37256
rect 27847 37216 29276 37244
rect 27847 37213 27859 37216
rect 27801 37207 27859 37213
rect 29270 37204 29276 37216
rect 29328 37204 29334 37256
rect 29656 37253 29684 37284
rect 30193 37281 30205 37315
rect 30239 37312 30251 37315
rect 30926 37312 30932 37324
rect 30239 37284 30932 37312
rect 30239 37281 30251 37284
rect 30193 37275 30251 37281
rect 30926 37272 30932 37284
rect 30984 37272 30990 37324
rect 29641 37247 29699 37253
rect 29641 37213 29653 37247
rect 29687 37213 29699 37247
rect 29641 37207 29699 37213
rect 29733 37247 29791 37253
rect 29733 37213 29745 37247
rect 29779 37244 29791 37247
rect 29917 37247 29975 37253
rect 29917 37244 29929 37247
rect 29779 37216 29929 37244
rect 29779 37213 29791 37216
rect 29733 37207 29791 37213
rect 29917 37213 29929 37216
rect 29963 37213 29975 37247
rect 29917 37207 29975 37213
rect 32582 37204 32588 37256
rect 32640 37204 32646 37256
rect 37645 37247 37703 37253
rect 37645 37213 37657 37247
rect 37691 37213 37703 37247
rect 37645 37207 37703 37213
rect 27890 37176 27896 37188
rect 26620 37148 27896 37176
rect 27890 37136 27896 37148
rect 27948 37176 27954 37188
rect 30098 37176 30104 37188
rect 27948 37148 30104 37176
rect 27948 37136 27954 37148
rect 30098 37136 30104 37148
rect 30156 37136 30162 37188
rect 30466 37136 30472 37188
rect 30524 37176 30530 37188
rect 30524 37148 30682 37176
rect 30524 37136 30530 37148
rect 31478 37136 31484 37188
rect 31536 37176 31542 37188
rect 37660 37176 37688 37207
rect 31536 37148 37688 37176
rect 31536 37136 31542 37148
rect 24394 37108 24400 37120
rect 23492 37080 24400 37108
rect 24394 37068 24400 37080
rect 24452 37068 24458 37120
rect 26513 37111 26571 37117
rect 26513 37077 26525 37111
rect 26559 37108 26571 37111
rect 27522 37108 27528 37120
rect 26559 37080 27528 37108
rect 26559 37077 26571 37080
rect 26513 37071 26571 37077
rect 27522 37068 27528 37080
rect 27580 37108 27586 37120
rect 27709 37111 27767 37117
rect 27709 37108 27721 37111
rect 27580 37080 27721 37108
rect 27580 37068 27586 37080
rect 27709 37077 27721 37080
rect 27755 37077 27767 37111
rect 27709 37071 27767 37077
rect 30006 37068 30012 37120
rect 30064 37108 30070 37120
rect 31665 37111 31723 37117
rect 31665 37108 31677 37111
rect 30064 37080 31677 37108
rect 30064 37068 30070 37080
rect 31665 37077 31677 37080
rect 31711 37077 31723 37111
rect 31665 37071 31723 37077
rect 32490 37068 32496 37120
rect 32548 37068 32554 37120
rect 37826 37068 37832 37120
rect 37884 37068 37890 37120
rect 1104 37018 38272 37040
rect 1104 36966 4874 37018
rect 4926 36966 4938 37018
rect 4990 36966 5002 37018
rect 5054 36966 5066 37018
rect 5118 36966 5130 37018
rect 5182 36966 35594 37018
rect 35646 36966 35658 37018
rect 35710 36966 35722 37018
rect 35774 36966 35786 37018
rect 35838 36966 35850 37018
rect 35902 36966 38272 37018
rect 1104 36944 38272 36966
rect 8294 36864 8300 36916
rect 8352 36904 8358 36916
rect 9309 36907 9367 36913
rect 9309 36904 9321 36907
rect 8352 36876 9321 36904
rect 8352 36864 8358 36876
rect 9309 36873 9321 36876
rect 9355 36873 9367 36907
rect 9309 36867 9367 36873
rect 9769 36907 9827 36913
rect 9769 36873 9781 36907
rect 9815 36904 9827 36907
rect 10686 36904 10692 36916
rect 9815 36876 10692 36904
rect 9815 36873 9827 36876
rect 9769 36867 9827 36873
rect 10686 36864 10692 36876
rect 10744 36864 10750 36916
rect 20714 36864 20720 36916
rect 20772 36904 20778 36916
rect 20901 36907 20959 36913
rect 20901 36904 20913 36907
rect 20772 36876 20913 36904
rect 20772 36864 20778 36876
rect 20901 36873 20913 36876
rect 20947 36873 20959 36907
rect 22370 36904 22376 36916
rect 20901 36867 20959 36873
rect 22066 36876 22376 36904
rect 8386 36796 8392 36848
rect 8444 36836 8450 36848
rect 8757 36839 8815 36845
rect 8757 36836 8769 36839
rect 8444 36808 8769 36836
rect 8444 36796 8450 36808
rect 8757 36805 8769 36808
rect 8803 36805 8815 36839
rect 8757 36799 8815 36805
rect 7285 36771 7343 36777
rect 7285 36737 7297 36771
rect 7331 36737 7343 36771
rect 7285 36731 7343 36737
rect 9677 36771 9735 36777
rect 9677 36737 9689 36771
rect 9723 36768 9735 36771
rect 10594 36768 10600 36780
rect 9723 36740 10600 36768
rect 9723 36737 9735 36740
rect 9677 36731 9735 36737
rect 7300 36700 7328 36731
rect 10594 36728 10600 36740
rect 10652 36728 10658 36780
rect 16942 36728 16948 36780
rect 17000 36768 17006 36780
rect 18690 36768 18696 36780
rect 17000 36740 18696 36768
rect 17000 36728 17006 36740
rect 18690 36728 18696 36740
rect 18748 36728 18754 36780
rect 21085 36771 21143 36777
rect 21085 36737 21097 36771
rect 21131 36768 21143 36771
rect 22066 36768 22094 36876
rect 22370 36864 22376 36876
rect 22428 36864 22434 36916
rect 22462 36864 22468 36916
rect 22520 36904 22526 36916
rect 23382 36904 23388 36916
rect 22520 36876 23388 36904
rect 22520 36864 22526 36876
rect 23382 36864 23388 36876
rect 23440 36904 23446 36916
rect 23440 36876 24900 36904
rect 23440 36864 23446 36876
rect 24029 36839 24087 36845
rect 24029 36805 24041 36839
rect 24075 36836 24087 36839
rect 24075 36808 24808 36836
rect 24075 36805 24087 36808
rect 24029 36799 24087 36805
rect 21131 36740 22094 36768
rect 23845 36771 23903 36777
rect 21131 36737 21143 36740
rect 21085 36731 21143 36737
rect 23845 36737 23857 36771
rect 23891 36737 23903 36771
rect 23845 36731 23903 36737
rect 8021 36703 8079 36709
rect 8021 36700 8033 36703
rect 7300 36672 8033 36700
rect 8021 36669 8033 36672
rect 8067 36700 8079 36703
rect 9122 36700 9128 36712
rect 8067 36672 9128 36700
rect 8067 36669 8079 36672
rect 8021 36663 8079 36669
rect 9122 36660 9128 36672
rect 9180 36660 9186 36712
rect 9858 36660 9864 36712
rect 9916 36660 9922 36712
rect 15562 36660 15568 36712
rect 15620 36700 15626 36712
rect 17954 36700 17960 36712
rect 15620 36672 17960 36700
rect 15620 36660 15626 36672
rect 17954 36660 17960 36672
rect 18012 36660 18018 36712
rect 18708 36700 18736 36728
rect 18708 36672 20576 36700
rect 17034 36592 17040 36644
rect 17092 36632 17098 36644
rect 19702 36632 19708 36644
rect 17092 36604 19708 36632
rect 17092 36592 17098 36604
rect 19702 36592 19708 36604
rect 19760 36592 19766 36644
rect 20548 36632 20576 36672
rect 22278 36660 22284 36712
rect 22336 36700 22342 36712
rect 23661 36703 23719 36709
rect 23661 36700 23673 36703
rect 22336 36672 23673 36700
rect 22336 36660 22342 36672
rect 23661 36669 23673 36672
rect 23707 36669 23719 36703
rect 23860 36700 23888 36731
rect 24486 36728 24492 36780
rect 24544 36728 24550 36780
rect 24578 36728 24584 36780
rect 24636 36768 24642 36780
rect 24780 36777 24808 36808
rect 24673 36771 24731 36777
rect 24673 36768 24685 36771
rect 24636 36740 24685 36768
rect 24636 36728 24642 36740
rect 24673 36737 24685 36740
rect 24719 36737 24731 36771
rect 24673 36731 24731 36737
rect 24765 36771 24823 36777
rect 24765 36737 24777 36771
rect 24811 36737 24823 36771
rect 24872 36768 24900 36876
rect 27798 36864 27804 36916
rect 27856 36904 27862 36916
rect 28077 36907 28135 36913
rect 28077 36904 28089 36907
rect 27856 36876 28089 36904
rect 27856 36864 27862 36876
rect 28077 36873 28089 36876
rect 28123 36873 28135 36907
rect 28077 36867 28135 36873
rect 28994 36864 29000 36916
rect 29052 36904 29058 36916
rect 29181 36907 29239 36913
rect 29181 36904 29193 36907
rect 29052 36876 29193 36904
rect 29052 36864 29058 36876
rect 29181 36873 29193 36876
rect 29227 36873 29239 36907
rect 29181 36867 29239 36873
rect 30006 36864 30012 36916
rect 30064 36904 30070 36916
rect 30929 36907 30987 36913
rect 30929 36904 30941 36907
rect 30064 36876 30941 36904
rect 30064 36864 30070 36876
rect 30929 36873 30941 36876
rect 30975 36873 30987 36907
rect 30929 36867 30987 36873
rect 31202 36864 31208 36916
rect 31260 36904 31266 36916
rect 31297 36907 31355 36913
rect 31297 36904 31309 36907
rect 31260 36876 31309 36904
rect 31260 36864 31266 36876
rect 31297 36873 31309 36876
rect 31343 36873 31355 36907
rect 31297 36867 31355 36873
rect 31478 36864 31484 36916
rect 31536 36864 31542 36916
rect 32490 36864 32496 36916
rect 32548 36864 32554 36916
rect 25130 36796 25136 36848
rect 25188 36836 25194 36848
rect 31496 36836 31524 36864
rect 32508 36836 32536 36864
rect 25188 36808 31524 36836
rect 32324 36808 32536 36836
rect 25188 36796 25194 36808
rect 25590 36768 25596 36780
rect 24872 36740 25596 36768
rect 24765 36731 24823 36737
rect 25590 36728 25596 36740
rect 25648 36728 25654 36780
rect 27706 36728 27712 36780
rect 27764 36728 27770 36780
rect 27985 36771 28043 36777
rect 27985 36737 27997 36771
rect 28031 36768 28043 36771
rect 28166 36768 28172 36780
rect 28031 36740 28172 36768
rect 28031 36737 28043 36740
rect 27985 36731 28043 36737
rect 28166 36728 28172 36740
rect 28224 36728 28230 36780
rect 28258 36728 28264 36780
rect 28316 36728 28322 36780
rect 29362 36728 29368 36780
rect 29420 36768 29426 36780
rect 32324 36777 32352 36808
rect 29549 36771 29607 36777
rect 29549 36768 29561 36771
rect 29420 36740 29561 36768
rect 29420 36728 29426 36740
rect 29549 36737 29561 36740
rect 29595 36768 29607 36771
rect 30837 36771 30895 36777
rect 30837 36768 30849 36771
rect 29595 36740 30849 36768
rect 29595 36737 29607 36740
rect 29549 36731 29607 36737
rect 30837 36737 30849 36740
rect 30883 36737 30895 36771
rect 30837 36731 30895 36737
rect 32309 36771 32367 36777
rect 32309 36737 32321 36771
rect 32355 36737 32367 36771
rect 32309 36731 32367 36737
rect 23860 36672 23980 36700
rect 23661 36663 23719 36669
rect 23952 36632 23980 36672
rect 29638 36660 29644 36712
rect 29696 36660 29702 36712
rect 29825 36703 29883 36709
rect 29825 36669 29837 36703
rect 29871 36669 29883 36703
rect 29825 36663 29883 36669
rect 24210 36632 24216 36644
rect 20548 36604 23520 36632
rect 23952 36604 24216 36632
rect 7561 36567 7619 36573
rect 7561 36533 7573 36567
rect 7607 36564 7619 36567
rect 7650 36564 7656 36576
rect 7607 36536 7656 36564
rect 7607 36533 7619 36536
rect 7561 36527 7619 36533
rect 7650 36524 7656 36536
rect 7708 36524 7714 36576
rect 12986 36524 12992 36576
rect 13044 36564 13050 36576
rect 13722 36564 13728 36576
rect 13044 36536 13728 36564
rect 13044 36524 13050 36536
rect 13722 36524 13728 36536
rect 13780 36524 13786 36576
rect 14090 36524 14096 36576
rect 14148 36564 14154 36576
rect 14826 36564 14832 36576
rect 14148 36536 14832 36564
rect 14148 36524 14154 36536
rect 14826 36524 14832 36536
rect 14884 36524 14890 36576
rect 15746 36524 15752 36576
rect 15804 36564 15810 36576
rect 23290 36564 23296 36576
rect 15804 36536 23296 36564
rect 15804 36524 15810 36536
rect 23290 36524 23296 36536
rect 23348 36524 23354 36576
rect 23492 36564 23520 36604
rect 24210 36592 24216 36604
rect 24268 36592 24274 36644
rect 24026 36564 24032 36576
rect 23492 36536 24032 36564
rect 24026 36524 24032 36536
rect 24084 36524 24090 36576
rect 24670 36524 24676 36576
rect 24728 36524 24734 36576
rect 24946 36524 24952 36576
rect 25004 36524 25010 36576
rect 27430 36524 27436 36576
rect 27488 36564 27494 36576
rect 27617 36567 27675 36573
rect 27617 36564 27629 36567
rect 27488 36536 27629 36564
rect 27488 36524 27494 36536
rect 27617 36533 27629 36536
rect 27663 36533 27675 36567
rect 27617 36527 27675 36533
rect 28442 36524 28448 36576
rect 28500 36524 28506 36576
rect 28626 36524 28632 36576
rect 28684 36564 28690 36576
rect 29840 36564 29868 36663
rect 30098 36660 30104 36712
rect 30156 36700 30162 36712
rect 30653 36703 30711 36709
rect 30653 36700 30665 36703
rect 30156 36672 30665 36700
rect 30156 36660 30162 36672
rect 30653 36669 30665 36672
rect 30699 36669 30711 36703
rect 30653 36663 30711 36669
rect 28684 36536 29868 36564
rect 30852 36564 30880 36731
rect 33686 36728 33692 36780
rect 33744 36728 33750 36780
rect 32214 36660 32220 36712
rect 32272 36700 32278 36712
rect 32585 36703 32643 36709
rect 32585 36700 32597 36703
rect 32272 36672 32597 36700
rect 32272 36660 32278 36672
rect 32585 36669 32597 36672
rect 32631 36669 32643 36703
rect 32585 36663 32643 36669
rect 33134 36564 33140 36576
rect 30852 36536 33140 36564
rect 28684 36524 28690 36536
rect 33134 36524 33140 36536
rect 33192 36524 33198 36576
rect 34054 36524 34060 36576
rect 34112 36524 34118 36576
rect 1104 36474 38272 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 38272 36474
rect 1104 36400 38272 36422
rect 10686 36320 10692 36372
rect 10744 36320 10750 36372
rect 13814 36320 13820 36372
rect 13872 36360 13878 36372
rect 14277 36363 14335 36369
rect 14277 36360 14289 36363
rect 13872 36332 14289 36360
rect 13872 36320 13878 36332
rect 14277 36329 14289 36332
rect 14323 36329 14335 36363
rect 15930 36360 15936 36372
rect 14277 36323 14335 36329
rect 14384 36332 15936 36360
rect 9030 36184 9036 36236
rect 9088 36224 9094 36236
rect 10704 36224 10732 36320
rect 11793 36295 11851 36301
rect 11793 36261 11805 36295
rect 11839 36261 11851 36295
rect 11793 36255 11851 36261
rect 12529 36295 12587 36301
rect 12529 36261 12541 36295
rect 12575 36261 12587 36295
rect 12529 36255 12587 36261
rect 12713 36295 12771 36301
rect 12713 36261 12725 36295
rect 12759 36261 12771 36295
rect 12713 36255 12771 36261
rect 11808 36224 11836 36255
rect 12544 36224 12572 36255
rect 9088 36196 9536 36224
rect 10704 36196 11560 36224
rect 11808 36196 12572 36224
rect 12621 36227 12679 36233
rect 9088 36184 9094 36196
rect 4706 36116 4712 36168
rect 4764 36156 4770 36168
rect 9508 36165 9536 36196
rect 11532 36168 11560 36196
rect 12621 36193 12633 36227
rect 12667 36224 12679 36227
rect 12728 36224 12756 36255
rect 12667 36196 12756 36224
rect 12820 36196 13400 36224
rect 12667 36193 12679 36196
rect 12621 36187 12679 36193
rect 5721 36159 5779 36165
rect 5721 36156 5733 36159
rect 4764 36128 5733 36156
rect 4764 36116 4770 36128
rect 5721 36125 5733 36128
rect 5767 36125 5779 36159
rect 5721 36119 5779 36125
rect 5813 36159 5871 36165
rect 5813 36125 5825 36159
rect 5859 36156 5871 36159
rect 5997 36159 6055 36165
rect 5997 36156 6009 36159
rect 5859 36128 6009 36156
rect 5859 36125 5871 36128
rect 5813 36119 5871 36125
rect 5997 36125 6009 36128
rect 6043 36125 6055 36159
rect 5997 36119 6055 36125
rect 9493 36159 9551 36165
rect 9493 36125 9505 36159
rect 9539 36125 9551 36159
rect 9493 36119 9551 36125
rect 9766 36116 9772 36168
rect 9824 36116 9830 36168
rect 11238 36116 11244 36168
rect 11296 36116 11302 36168
rect 11514 36116 11520 36168
rect 11572 36116 11578 36168
rect 11609 36159 11667 36165
rect 11609 36125 11621 36159
rect 11655 36156 11667 36159
rect 11790 36156 11796 36168
rect 11655 36128 11796 36156
rect 11655 36125 11667 36128
rect 11609 36119 11667 36125
rect 11790 36116 11796 36128
rect 11848 36116 11854 36168
rect 12099 36159 12157 36165
rect 12099 36156 12111 36159
rect 12083 36125 12111 36156
rect 12145 36156 12157 36159
rect 12820 36156 12848 36196
rect 12145 36128 12848 36156
rect 12892 36159 12950 36165
rect 12145 36125 12157 36128
rect 12083 36119 12157 36125
rect 12892 36125 12904 36159
rect 12938 36125 12950 36159
rect 13262 36156 13268 36168
rect 13223 36128 13268 36156
rect 12892 36119 12950 36125
rect 6270 36048 6276 36100
rect 6328 36048 6334 36100
rect 7650 36088 7656 36100
rect 7498 36060 7656 36088
rect 6638 35980 6644 36032
rect 6696 36020 6702 36032
rect 7576 36020 7604 36060
rect 7650 36048 7656 36060
rect 7708 36088 7714 36100
rect 10226 36088 10232 36100
rect 7708 36060 10232 36088
rect 7708 36048 7714 36060
rect 10226 36048 10232 36060
rect 10284 36048 10290 36100
rect 11422 36048 11428 36100
rect 11480 36048 11486 36100
rect 11698 36048 11704 36100
rect 11756 36088 11762 36100
rect 12083 36088 12111 36119
rect 12434 36088 12440 36100
rect 11756 36060 12111 36088
rect 11756 36048 11762 36060
rect 12406 36048 12440 36088
rect 12492 36048 12498 36100
rect 12802 36048 12808 36100
rect 12860 36088 12866 36100
rect 12912 36088 12940 36119
rect 13262 36116 13268 36128
rect 13320 36116 13326 36168
rect 13372 36165 13400 36196
rect 13357 36159 13415 36165
rect 13357 36125 13369 36159
rect 13403 36125 13415 36159
rect 13357 36119 13415 36125
rect 13814 36116 13820 36168
rect 13872 36116 13878 36168
rect 14274 36116 14280 36168
rect 14332 36116 14338 36168
rect 14384 36165 14412 36332
rect 15930 36320 15936 36332
rect 15988 36320 15994 36372
rect 16408 36332 17172 36360
rect 16408 36292 16436 36332
rect 14660 36264 16436 36292
rect 16485 36295 16543 36301
rect 14660 36165 14688 36264
rect 16485 36261 16497 36295
rect 16531 36292 16543 36295
rect 17144 36292 17172 36332
rect 17770 36320 17776 36372
rect 17828 36360 17834 36372
rect 18049 36363 18107 36369
rect 18049 36360 18061 36363
rect 17828 36332 18061 36360
rect 17828 36320 17834 36332
rect 18049 36329 18061 36332
rect 18095 36329 18107 36363
rect 18049 36323 18107 36329
rect 19886 36320 19892 36372
rect 19944 36360 19950 36372
rect 24121 36363 24179 36369
rect 19944 36332 24072 36360
rect 19944 36320 19950 36332
rect 18598 36292 18604 36304
rect 16531 36264 16804 36292
rect 16531 36261 16543 36264
rect 16485 36255 16543 36261
rect 14826 36184 14832 36236
rect 14884 36224 14890 36236
rect 15562 36224 15568 36236
rect 14884 36196 15332 36224
rect 14884 36184 14890 36196
rect 14369 36159 14427 36165
rect 14369 36125 14381 36159
rect 14415 36125 14427 36159
rect 14645 36159 14703 36165
rect 14645 36156 14657 36159
rect 14369 36119 14427 36125
rect 14476 36128 14657 36156
rect 12860 36060 12940 36088
rect 12860 36048 12866 36060
rect 12986 36048 12992 36100
rect 13044 36048 13050 36100
rect 13081 36091 13139 36097
rect 13081 36057 13093 36091
rect 13127 36057 13139 36091
rect 13832 36088 13860 36116
rect 14476 36088 14504 36128
rect 14645 36125 14657 36128
rect 14691 36125 14703 36159
rect 14645 36119 14703 36125
rect 14737 36159 14795 36165
rect 14737 36125 14749 36159
rect 14783 36156 14795 36159
rect 15194 36156 15200 36168
rect 14783 36128 15200 36156
rect 14783 36125 14795 36128
rect 14737 36119 14795 36125
rect 15194 36116 15200 36128
rect 15252 36116 15258 36168
rect 15304 36165 15332 36196
rect 15396 36196 15568 36224
rect 15396 36165 15424 36196
rect 15562 36184 15568 36196
rect 15620 36184 15626 36236
rect 15672 36196 15976 36224
rect 15672 36165 15700 36196
rect 15289 36159 15347 36165
rect 15289 36125 15301 36159
rect 15335 36125 15347 36159
rect 15289 36119 15347 36125
rect 15381 36159 15439 36165
rect 15381 36125 15393 36159
rect 15427 36125 15439 36159
rect 15657 36159 15715 36165
rect 15657 36156 15669 36159
rect 15381 36119 15439 36125
rect 15488 36128 15669 36156
rect 15488 36100 15516 36128
rect 15657 36125 15669 36128
rect 15703 36125 15715 36159
rect 15657 36119 15715 36125
rect 15746 36116 15752 36168
rect 15804 36116 15810 36168
rect 15948 36165 15976 36196
rect 15933 36159 15991 36165
rect 15933 36125 15945 36159
rect 15979 36125 15991 36159
rect 15933 36119 15991 36125
rect 13832 36060 14504 36088
rect 14553 36091 14611 36097
rect 13081 36051 13139 36057
rect 14553 36057 14565 36091
rect 14599 36057 14611 36091
rect 14553 36051 14611 36057
rect 6696 35992 7604 36020
rect 6696 35980 6702 35992
rect 7742 35980 7748 36032
rect 7800 35980 7806 36032
rect 9214 35980 9220 36032
rect 9272 36020 9278 36032
rect 9401 36023 9459 36029
rect 9401 36020 9413 36023
rect 9272 35992 9413 36020
rect 9272 35980 9278 35992
rect 9401 35989 9413 35992
rect 9447 35989 9459 36023
rect 9401 35983 9459 35989
rect 9582 35980 9588 36032
rect 9640 35980 9646 36032
rect 11330 35980 11336 36032
rect 11388 36020 11394 36032
rect 11977 36023 12035 36029
rect 11977 36020 11989 36023
rect 11388 35992 11989 36020
rect 11388 35980 11394 35992
rect 11977 35989 11989 35992
rect 12023 35989 12035 36023
rect 11977 35983 12035 35989
rect 12161 36023 12219 36029
rect 12161 35989 12173 36023
rect 12207 36020 12219 36023
rect 12406 36020 12434 36048
rect 12207 35992 12434 36020
rect 12207 35989 12219 35992
rect 12161 35983 12219 35989
rect 12618 35980 12624 36032
rect 12676 36020 12682 36032
rect 13096 36020 13124 36051
rect 13814 36020 13820 36032
rect 12676 35992 13820 36020
rect 12676 35980 12682 35992
rect 13814 35980 13820 35992
rect 13872 35980 13878 36032
rect 14458 35980 14464 36032
rect 14516 36020 14522 36032
rect 14568 36020 14596 36051
rect 15470 36048 15476 36100
rect 15528 36048 15534 36100
rect 15565 36091 15623 36097
rect 15565 36057 15577 36091
rect 15611 36088 15623 36091
rect 15611 36060 15700 36088
rect 15611 36057 15623 36060
rect 15565 36051 15623 36057
rect 15672 36032 15700 36060
rect 14516 35992 14596 36020
rect 14516 35980 14522 35992
rect 15286 35980 15292 36032
rect 15344 35980 15350 36032
rect 15654 35980 15660 36032
rect 15712 35980 15718 36032
rect 15948 36020 15976 36119
rect 16206 36116 16212 36168
rect 16264 36116 16270 36168
rect 16301 36159 16359 36165
rect 16301 36125 16313 36159
rect 16347 36156 16359 36159
rect 16666 36156 16672 36168
rect 16347 36128 16672 36156
rect 16347 36125 16359 36128
rect 16301 36119 16359 36125
rect 16666 36116 16672 36128
rect 16724 36116 16730 36168
rect 16776 36165 16804 36264
rect 17144 36264 18604 36292
rect 16761 36159 16819 36165
rect 16761 36125 16773 36159
rect 16807 36125 16819 36159
rect 16761 36119 16819 36125
rect 16850 36116 16856 36168
rect 16908 36116 16914 36168
rect 17144 36165 17172 36264
rect 18598 36252 18604 36264
rect 18656 36252 18662 36304
rect 24044 36292 24072 36332
rect 24121 36329 24133 36363
rect 24167 36360 24179 36363
rect 24486 36360 24492 36372
rect 24167 36332 24492 36360
rect 24167 36329 24179 36332
rect 24121 36323 24179 36329
rect 24486 36320 24492 36332
rect 24544 36320 24550 36372
rect 27893 36363 27951 36369
rect 27893 36329 27905 36363
rect 27939 36360 27951 36363
rect 28258 36360 28264 36372
rect 27939 36332 28264 36360
rect 27939 36329 27951 36332
rect 27893 36323 27951 36329
rect 28258 36320 28264 36332
rect 28316 36320 28322 36372
rect 30098 36320 30104 36372
rect 30156 36360 30162 36372
rect 30156 36332 31754 36360
rect 30156 36320 30162 36332
rect 24210 36292 24216 36304
rect 22021 36264 23980 36292
rect 24044 36264 24216 36292
rect 17880 36196 19334 36224
rect 17310 36165 17316 36168
rect 17129 36159 17187 36165
rect 17129 36125 17141 36159
rect 17175 36125 17187 36159
rect 17129 36119 17187 36125
rect 17267 36159 17316 36165
rect 17267 36125 17279 36159
rect 17313 36125 17316 36159
rect 17267 36119 17316 36125
rect 17310 36116 17316 36119
rect 17368 36116 17374 36168
rect 17497 36159 17555 36165
rect 17497 36156 17509 36159
rect 17420 36128 17509 36156
rect 16117 36091 16175 36097
rect 16117 36057 16129 36091
rect 16163 36088 16175 36091
rect 16942 36088 16948 36100
rect 16163 36060 16948 36088
rect 16163 36057 16175 36060
rect 16117 36051 16175 36057
rect 16942 36048 16948 36060
rect 17000 36048 17006 36100
rect 17034 36048 17040 36100
rect 17092 36048 17098 36100
rect 17420 36088 17448 36128
rect 17497 36125 17509 36128
rect 17543 36125 17555 36159
rect 17497 36119 17555 36125
rect 17586 36116 17592 36168
rect 17644 36156 17650 36168
rect 17880 36165 17908 36196
rect 17865 36159 17923 36165
rect 17865 36156 17877 36159
rect 17644 36128 17877 36156
rect 17644 36116 17650 36128
rect 17865 36125 17877 36128
rect 17911 36125 17923 36159
rect 17865 36119 17923 36125
rect 18046 36116 18052 36168
rect 18104 36156 18110 36168
rect 18509 36159 18567 36165
rect 18509 36156 18521 36159
rect 18104 36128 18521 36156
rect 18104 36116 18110 36128
rect 18509 36125 18521 36128
rect 18555 36125 18567 36159
rect 18509 36119 18567 36125
rect 18690 36116 18696 36168
rect 18748 36116 18754 36168
rect 19306 36156 19334 36196
rect 19794 36184 19800 36236
rect 19852 36184 19858 36236
rect 20201 36159 20259 36165
rect 20201 36156 20213 36159
rect 19306 36128 20213 36156
rect 20201 36125 20213 36128
rect 20247 36156 20259 36159
rect 22021 36156 22049 36264
rect 20247 36128 22049 36156
rect 20247 36125 20259 36128
rect 20201 36119 20259 36125
rect 22094 36116 22100 36168
rect 22152 36156 22158 36168
rect 22830 36156 22836 36168
rect 22152 36128 22836 36156
rect 22152 36116 22158 36128
rect 22830 36116 22836 36128
rect 22888 36156 22894 36168
rect 23198 36156 23204 36168
rect 22888 36128 23204 36156
rect 22888 36116 22894 36128
rect 23198 36116 23204 36128
rect 23256 36156 23262 36168
rect 23952 36165 23980 36264
rect 24210 36252 24216 36264
rect 24268 36252 24274 36304
rect 25682 36252 25688 36304
rect 25740 36292 25746 36304
rect 26142 36292 26148 36304
rect 25740 36264 26148 36292
rect 25740 36252 25746 36264
rect 26142 36252 26148 36264
rect 26200 36252 26206 36304
rect 29822 36292 29828 36304
rect 27540 36264 29828 36292
rect 25222 36184 25228 36236
rect 25280 36224 25286 36236
rect 27540 36224 27568 36264
rect 29822 36252 29828 36264
rect 29880 36252 29886 36304
rect 25280 36196 25912 36224
rect 25280 36184 25286 36196
rect 23569 36159 23627 36165
rect 23569 36156 23581 36159
rect 23256 36128 23581 36156
rect 23256 36116 23262 36128
rect 23569 36125 23581 36128
rect 23615 36125 23627 36159
rect 23569 36119 23627 36125
rect 23937 36159 23995 36165
rect 23937 36125 23949 36159
rect 23983 36156 23995 36159
rect 24670 36156 24676 36168
rect 23983 36128 24676 36156
rect 23983 36125 23995 36128
rect 23937 36119 23995 36125
rect 24670 36116 24676 36128
rect 24728 36116 24734 36168
rect 25501 36159 25559 36165
rect 25501 36125 25513 36159
rect 25547 36156 25559 36159
rect 25590 36156 25596 36168
rect 25547 36128 25596 36156
rect 25547 36125 25559 36128
rect 25501 36119 25559 36125
rect 25590 36116 25596 36128
rect 25648 36116 25654 36168
rect 25884 36165 25912 36196
rect 27172 36196 27568 36224
rect 27172 36168 27200 36196
rect 25869 36159 25927 36165
rect 25869 36125 25881 36159
rect 25915 36156 25927 36159
rect 26326 36156 26332 36168
rect 25915 36128 26332 36156
rect 25915 36125 25927 36128
rect 25869 36119 25927 36125
rect 26326 36116 26332 36128
rect 26384 36116 26390 36168
rect 26510 36116 26516 36168
rect 26568 36156 26574 36168
rect 26568 36128 27108 36156
rect 26568 36116 26574 36128
rect 17328 36060 17448 36088
rect 17328 36020 17356 36060
rect 17678 36048 17684 36100
rect 17736 36048 17742 36100
rect 17773 36091 17831 36097
rect 17773 36057 17785 36091
rect 17819 36088 17831 36091
rect 17954 36088 17960 36100
rect 17819 36060 17960 36088
rect 17819 36057 17831 36060
rect 17773 36051 17831 36057
rect 17954 36048 17960 36060
rect 18012 36088 18018 36100
rect 18012 36060 18736 36088
rect 18012 36048 18018 36060
rect 15948 35992 17356 36020
rect 17402 35980 17408 36032
rect 17460 35980 17466 36032
rect 18598 35980 18604 36032
rect 18656 35980 18662 36032
rect 18708 36020 18736 36060
rect 18782 36048 18788 36100
rect 18840 36088 18846 36100
rect 19797 36091 19855 36097
rect 19797 36088 19809 36091
rect 18840 36060 19809 36088
rect 18840 36048 18846 36060
rect 19797 36057 19809 36060
rect 19843 36057 19855 36091
rect 19797 36051 19855 36057
rect 19886 36048 19892 36100
rect 19944 36088 19950 36100
rect 19981 36091 20039 36097
rect 19981 36088 19993 36091
rect 19944 36060 19993 36088
rect 19944 36048 19950 36060
rect 19981 36057 19993 36060
rect 20027 36057 20039 36091
rect 19981 36051 20039 36057
rect 20073 36091 20131 36097
rect 20073 36057 20085 36091
rect 20119 36088 20131 36091
rect 20530 36088 20536 36100
rect 20119 36060 20536 36088
rect 20119 36057 20131 36060
rect 20073 36051 20131 36057
rect 20530 36048 20536 36060
rect 20588 36048 20594 36100
rect 21358 36048 21364 36100
rect 21416 36088 21422 36100
rect 23753 36091 23811 36097
rect 23753 36088 23765 36091
rect 21416 36060 23765 36088
rect 21416 36048 21422 36060
rect 23753 36057 23765 36060
rect 23799 36057 23811 36091
rect 23753 36051 23811 36057
rect 23845 36091 23903 36097
rect 23845 36057 23857 36091
rect 23891 36057 23903 36091
rect 23845 36051 23903 36057
rect 22646 36020 22652 36032
rect 18708 35992 22652 36020
rect 22646 35980 22652 35992
rect 22704 35980 22710 36032
rect 23566 35980 23572 36032
rect 23624 36020 23630 36032
rect 23860 36020 23888 36051
rect 24118 36048 24124 36100
rect 24176 36088 24182 36100
rect 24486 36088 24492 36100
rect 24176 36060 24492 36088
rect 24176 36048 24182 36060
rect 24486 36048 24492 36060
rect 24544 36048 24550 36100
rect 25038 36048 25044 36100
rect 25096 36088 25102 36100
rect 25406 36088 25412 36100
rect 25096 36060 25412 36088
rect 25096 36048 25102 36060
rect 25406 36048 25412 36060
rect 25464 36088 25470 36100
rect 25685 36091 25743 36097
rect 25685 36088 25697 36091
rect 25464 36060 25697 36088
rect 25464 36048 25470 36060
rect 25685 36057 25697 36060
rect 25731 36057 25743 36091
rect 25685 36051 25743 36057
rect 25777 36091 25835 36097
rect 25777 36057 25789 36091
rect 25823 36088 25835 36091
rect 27080 36088 27108 36128
rect 27154 36116 27160 36168
rect 27212 36116 27218 36168
rect 27246 36116 27252 36168
rect 27304 36116 27310 36168
rect 27338 36116 27344 36168
rect 27396 36156 27402 36168
rect 27540 36165 27568 36196
rect 28718 36184 28724 36236
rect 28776 36184 28782 36236
rect 31726 36224 31754 36332
rect 32214 36320 32220 36372
rect 32272 36320 32278 36372
rect 34054 36320 34060 36372
rect 34112 36320 34118 36372
rect 32585 36295 32643 36301
rect 32585 36261 32597 36295
rect 32631 36261 32643 36295
rect 32585 36255 32643 36261
rect 32398 36224 32404 36236
rect 31726 36196 32404 36224
rect 32398 36184 32404 36196
rect 32456 36184 32462 36236
rect 27525 36159 27583 36165
rect 27396 36128 27441 36156
rect 27396 36116 27402 36128
rect 27525 36125 27537 36159
rect 27571 36125 27583 36159
rect 27525 36119 27583 36125
rect 27755 36159 27813 36165
rect 27755 36125 27767 36159
rect 27801 36156 27813 36159
rect 27982 36156 27988 36168
rect 27801 36128 27988 36156
rect 27801 36125 27813 36128
rect 27755 36119 27813 36125
rect 27982 36116 27988 36128
rect 28040 36116 28046 36168
rect 28534 36116 28540 36168
rect 28592 36116 28598 36168
rect 28810 36116 28816 36168
rect 28868 36156 28874 36168
rect 30006 36156 30012 36168
rect 28868 36128 30012 36156
rect 28868 36116 28874 36128
rect 30006 36116 30012 36128
rect 30064 36116 30070 36168
rect 32033 36159 32091 36165
rect 32033 36125 32045 36159
rect 32079 36156 32091 36159
rect 32600 36156 32628 36255
rect 33137 36227 33195 36233
rect 33137 36224 33149 36227
rect 32079 36128 32628 36156
rect 32692 36196 33149 36224
rect 32079 36125 32091 36128
rect 32033 36119 32091 36125
rect 27617 36091 27675 36097
rect 27617 36088 27629 36091
rect 25823 36060 27016 36088
rect 27080 36060 27629 36088
rect 25823 36057 25835 36060
rect 25777 36051 25835 36057
rect 25792 36020 25820 36051
rect 23624 35992 25820 36020
rect 23624 35980 23630 35992
rect 25866 35980 25872 36032
rect 25924 36020 25930 36032
rect 26053 36023 26111 36029
rect 26053 36020 26065 36023
rect 25924 35992 26065 36020
rect 25924 35980 25930 35992
rect 26053 35989 26065 35992
rect 26099 35989 26111 36023
rect 26988 36020 27016 36060
rect 27617 36057 27629 36060
rect 27663 36057 27675 36091
rect 27617 36051 27675 36057
rect 31846 36048 31852 36100
rect 31904 36088 31910 36100
rect 32692 36088 32720 36196
rect 33137 36193 33149 36196
rect 33183 36193 33195 36227
rect 33137 36187 33195 36193
rect 33045 36159 33103 36165
rect 33045 36156 33057 36159
rect 31904 36060 32720 36088
rect 32784 36128 33057 36156
rect 31904 36048 31910 36060
rect 30742 36020 30748 36032
rect 26988 35992 30748 36020
rect 26053 35983 26111 35989
rect 30742 35980 30748 35992
rect 30800 36020 30806 36032
rect 32784 36020 32812 36128
rect 33045 36125 33057 36128
rect 33091 36156 33103 36159
rect 34072 36156 34100 36320
rect 33091 36128 34100 36156
rect 33091 36125 33103 36128
rect 33045 36119 33103 36125
rect 30800 35992 32812 36020
rect 32953 36023 33011 36029
rect 30800 35980 30806 35992
rect 32953 35989 32965 36023
rect 32999 36020 33011 36023
rect 33134 36020 33140 36032
rect 32999 35992 33140 36020
rect 32999 35989 33011 35992
rect 32953 35983 33011 35989
rect 33134 35980 33140 35992
rect 33192 36020 33198 36032
rect 33594 36020 33600 36032
rect 33192 35992 33600 36020
rect 33192 35980 33198 35992
rect 33594 35980 33600 35992
rect 33652 35980 33658 36032
rect 1104 35930 38272 35952
rect 1104 35878 4874 35930
rect 4926 35878 4938 35930
rect 4990 35878 5002 35930
rect 5054 35878 5066 35930
rect 5118 35878 5130 35930
rect 5182 35878 35594 35930
rect 35646 35878 35658 35930
rect 35710 35878 35722 35930
rect 35774 35878 35786 35930
rect 35838 35878 35850 35930
rect 35902 35878 38272 35930
rect 1104 35856 38272 35878
rect 6270 35776 6276 35828
rect 6328 35816 6334 35828
rect 6549 35819 6607 35825
rect 6549 35816 6561 35819
rect 6328 35788 6561 35816
rect 6328 35776 6334 35788
rect 6549 35785 6561 35788
rect 6595 35785 6607 35819
rect 6549 35779 6607 35785
rect 7653 35819 7711 35825
rect 7653 35785 7665 35819
rect 7699 35816 7711 35819
rect 7742 35816 7748 35828
rect 7699 35788 7748 35816
rect 7699 35785 7711 35788
rect 7653 35779 7711 35785
rect 7742 35776 7748 35788
rect 7800 35816 7806 35828
rect 8202 35816 8208 35828
rect 7800 35788 8208 35816
rect 7800 35776 7806 35788
rect 8202 35776 8208 35788
rect 8260 35776 8266 35828
rect 9030 35776 9036 35828
rect 9088 35816 9094 35828
rect 12710 35816 12716 35828
rect 9088 35788 12716 35816
rect 9088 35776 9094 35788
rect 12710 35776 12716 35788
rect 12768 35776 12774 35828
rect 13633 35819 13691 35825
rect 13633 35816 13645 35819
rect 13188 35788 13645 35816
rect 9493 35751 9551 35757
rect 9493 35717 9505 35751
rect 9539 35748 9551 35751
rect 9582 35748 9588 35760
rect 9539 35720 9588 35748
rect 9539 35717 9551 35720
rect 9493 35711 9551 35717
rect 9582 35708 9588 35720
rect 9640 35708 9646 35760
rect 10226 35708 10232 35760
rect 10284 35708 10290 35760
rect 13188 35692 13216 35788
rect 13633 35785 13645 35788
rect 13679 35785 13691 35819
rect 13633 35779 13691 35785
rect 13909 35819 13967 35825
rect 13909 35785 13921 35819
rect 13955 35816 13967 35819
rect 14274 35816 14280 35828
rect 13955 35788 14280 35816
rect 13955 35785 13967 35788
rect 13909 35779 13967 35785
rect 14274 35776 14280 35788
rect 14332 35776 14338 35828
rect 20990 35776 20996 35828
rect 21048 35776 21054 35828
rect 22462 35776 22468 35828
rect 22520 35776 22526 35828
rect 22646 35776 22652 35828
rect 22704 35816 22710 35828
rect 27798 35816 27804 35828
rect 22704 35788 27804 35816
rect 22704 35776 22710 35788
rect 13265 35751 13323 35757
rect 13265 35717 13277 35751
rect 13311 35748 13323 35751
rect 14001 35751 14059 35757
rect 14001 35748 14013 35751
rect 13311 35720 14013 35748
rect 13311 35717 13323 35720
rect 13265 35711 13323 35717
rect 14001 35717 14013 35720
rect 14047 35717 14059 35751
rect 14001 35711 14059 35717
rect 18598 35708 18604 35760
rect 18656 35748 18662 35760
rect 19062 35751 19120 35757
rect 19062 35748 19074 35751
rect 18656 35720 19074 35748
rect 18656 35708 18662 35720
rect 19062 35717 19074 35720
rect 19108 35717 19120 35751
rect 19062 35711 19120 35717
rect 19199 35751 19257 35757
rect 19199 35717 19211 35751
rect 19245 35748 19257 35751
rect 20438 35748 20444 35760
rect 19245 35720 20444 35748
rect 19245 35717 19257 35720
rect 19199 35711 19257 35717
rect 20438 35708 20444 35720
rect 20496 35708 20502 35760
rect 20809 35751 20867 35757
rect 20809 35717 20821 35751
rect 20855 35748 20867 35751
rect 21008 35748 21036 35776
rect 22480 35748 22508 35776
rect 20855 35720 21036 35748
rect 22076 35720 22508 35748
rect 23032 35720 23612 35748
rect 20855 35717 20867 35720
rect 20809 35711 20867 35717
rect 6733 35683 6791 35689
rect 6733 35649 6745 35683
rect 6779 35680 6791 35683
rect 7745 35683 7803 35689
rect 6779 35652 7328 35680
rect 6779 35649 6791 35652
rect 6733 35643 6791 35649
rect 7300 35553 7328 35652
rect 7745 35649 7757 35683
rect 7791 35680 7803 35683
rect 7791 35652 8156 35680
rect 7791 35649 7803 35652
rect 7745 35643 7803 35649
rect 8128 35624 8156 35652
rect 9122 35640 9128 35692
rect 9180 35640 9186 35692
rect 13081 35683 13139 35689
rect 13081 35649 13093 35683
rect 13127 35680 13139 35683
rect 13170 35680 13176 35692
rect 13127 35652 13176 35680
rect 13127 35649 13139 35652
rect 13081 35643 13139 35649
rect 13170 35640 13176 35652
rect 13228 35640 13234 35692
rect 13354 35640 13360 35692
rect 13412 35680 13418 35692
rect 13541 35683 13599 35689
rect 13541 35680 13553 35683
rect 13412 35652 13553 35680
rect 13412 35640 13418 35652
rect 13541 35649 13553 35652
rect 13587 35649 13599 35683
rect 13541 35643 13599 35649
rect 13722 35640 13728 35692
rect 13780 35640 13786 35692
rect 13814 35640 13820 35692
rect 13872 35680 13878 35692
rect 14829 35683 14887 35689
rect 14829 35680 14841 35683
rect 13872 35652 14841 35680
rect 13872 35640 13878 35652
rect 14829 35649 14841 35652
rect 14875 35680 14887 35683
rect 14875 35652 18828 35680
rect 14875 35649 14887 35652
rect 14829 35643 14887 35649
rect 7834 35572 7840 35624
rect 7892 35572 7898 35624
rect 8110 35572 8116 35624
rect 8168 35572 8174 35624
rect 8294 35572 8300 35624
rect 8352 35572 8358 35624
rect 7285 35547 7343 35553
rect 7285 35513 7297 35547
rect 7331 35513 7343 35547
rect 9140 35544 9168 35640
rect 9214 35572 9220 35624
rect 9272 35572 9278 35624
rect 12897 35615 12955 35621
rect 12897 35581 12909 35615
rect 12943 35612 12955 35615
rect 13372 35612 13400 35640
rect 12943 35584 13400 35612
rect 12943 35581 12955 35584
rect 12897 35575 12955 35581
rect 16206 35572 16212 35624
rect 16264 35572 16270 35624
rect 11054 35544 11060 35556
rect 9140 35516 9260 35544
rect 7285 35507 7343 35513
rect 9232 35476 9260 35516
rect 10520 35516 11060 35544
rect 10520 35476 10548 35516
rect 11054 35504 11060 35516
rect 11112 35504 11118 35556
rect 11238 35504 11244 35556
rect 11296 35544 11302 35556
rect 13357 35547 13415 35553
rect 13357 35544 13369 35547
rect 11296 35516 13369 35544
rect 11296 35504 11302 35516
rect 13357 35513 13369 35516
rect 13403 35544 13415 35547
rect 16224 35544 16252 35572
rect 13403 35516 16252 35544
rect 13403 35513 13415 35516
rect 13357 35507 13415 35513
rect 9232 35448 10548 35476
rect 10965 35479 11023 35485
rect 10965 35445 10977 35479
rect 11011 35476 11023 35479
rect 12434 35476 12440 35488
rect 11011 35448 12440 35476
rect 11011 35445 11023 35448
rect 10965 35439 11023 35445
rect 12434 35436 12440 35448
rect 12492 35436 12498 35488
rect 18690 35436 18696 35488
rect 18748 35436 18754 35488
rect 18800 35476 18828 35652
rect 18874 35640 18880 35692
rect 18932 35640 18938 35692
rect 18969 35683 19027 35689
rect 18969 35649 18981 35683
rect 19015 35649 19027 35683
rect 18969 35643 19027 35649
rect 18984 35544 19012 35643
rect 20070 35640 20076 35692
rect 20128 35680 20134 35692
rect 20993 35683 21051 35689
rect 20993 35680 21005 35683
rect 20128 35652 21005 35680
rect 20128 35640 20134 35652
rect 20993 35649 21005 35652
rect 21039 35649 21051 35683
rect 20993 35643 21051 35649
rect 21082 35640 21088 35692
rect 21140 35640 21146 35692
rect 21174 35640 21180 35692
rect 21232 35640 21238 35692
rect 22076 35689 22104 35720
rect 21361 35683 21419 35689
rect 21361 35649 21373 35683
rect 21407 35680 21419 35683
rect 21913 35683 21971 35689
rect 21913 35680 21925 35683
rect 21407 35652 21925 35680
rect 21407 35649 21419 35652
rect 21361 35643 21419 35649
rect 21913 35649 21925 35652
rect 21959 35649 21971 35683
rect 21913 35643 21971 35649
rect 22061 35683 22119 35689
rect 22061 35649 22073 35683
rect 22107 35649 22119 35683
rect 22061 35643 22119 35649
rect 22186 35640 22192 35692
rect 22244 35640 22250 35692
rect 22278 35640 22284 35692
rect 22336 35640 22342 35692
rect 22370 35640 22376 35692
rect 22428 35689 22434 35692
rect 22428 35643 22436 35689
rect 22428 35640 22434 35643
rect 22738 35640 22744 35692
rect 22796 35680 22802 35692
rect 23032 35689 23060 35720
rect 23584 35692 23612 35720
rect 23658 35708 23664 35760
rect 23716 35748 23722 35760
rect 23716 35720 24164 35748
rect 23716 35708 23722 35720
rect 22833 35683 22891 35689
rect 22833 35680 22845 35683
rect 22796 35652 22845 35680
rect 22796 35640 22802 35652
rect 22833 35649 22845 35652
rect 22879 35649 22891 35683
rect 22833 35643 22891 35649
rect 22981 35683 23060 35689
rect 22981 35649 22993 35683
rect 23027 35652 23060 35683
rect 23027 35649 23039 35652
rect 22981 35643 23039 35649
rect 23106 35640 23112 35692
rect 23164 35640 23170 35692
rect 23198 35640 23204 35692
rect 23256 35640 23262 35692
rect 23290 35640 23296 35692
rect 23348 35689 23354 35692
rect 23348 35680 23356 35689
rect 23348 35652 23393 35680
rect 23348 35643 23356 35652
rect 23348 35640 23354 35643
rect 23566 35640 23572 35692
rect 23624 35640 23630 35692
rect 23753 35683 23811 35689
rect 23753 35680 23765 35683
rect 23676 35652 23765 35680
rect 19337 35615 19395 35621
rect 19337 35581 19349 35615
rect 19383 35612 19395 35615
rect 21542 35612 21548 35624
rect 19383 35584 21548 35612
rect 19383 35581 19395 35584
rect 19337 35575 19395 35581
rect 21542 35572 21548 35584
rect 21600 35572 21606 35624
rect 22296 35612 22324 35640
rect 23676 35612 23704 35652
rect 23753 35649 23765 35652
rect 23799 35649 23811 35683
rect 23753 35643 23811 35649
rect 23845 35683 23903 35689
rect 23845 35649 23857 35683
rect 23891 35649 23903 35683
rect 23845 35643 23903 35649
rect 21836 35584 22324 35612
rect 23032 35584 23704 35612
rect 19794 35544 19800 35556
rect 18984 35516 19800 35544
rect 19794 35504 19800 35516
rect 19852 35504 19858 35556
rect 21836 35488 21864 35584
rect 22557 35547 22615 35553
rect 22557 35513 22569 35547
rect 22603 35544 22615 35547
rect 22830 35544 22836 35556
rect 22603 35516 22836 35544
rect 22603 35513 22615 35516
rect 22557 35507 22615 35513
rect 22830 35504 22836 35516
rect 22888 35504 22894 35556
rect 23032 35488 23060 35584
rect 23382 35504 23388 35556
rect 23440 35544 23446 35556
rect 23860 35544 23888 35643
rect 23934 35640 23940 35692
rect 23992 35640 23998 35692
rect 24136 35689 24164 35720
rect 24121 35683 24179 35689
rect 24121 35649 24133 35683
rect 24167 35649 24179 35683
rect 24121 35643 24179 35649
rect 23440 35516 23888 35544
rect 24136 35544 24164 35643
rect 24854 35640 24860 35692
rect 24912 35640 24918 35692
rect 24964 35678 24992 35788
rect 27798 35776 27804 35788
rect 27856 35816 27862 35828
rect 29181 35819 29239 35825
rect 29181 35816 29193 35819
rect 27856 35788 29193 35816
rect 27856 35776 27862 35788
rect 29181 35785 29193 35788
rect 29227 35785 29239 35819
rect 29181 35779 29239 35785
rect 29564 35788 30696 35816
rect 25038 35708 25044 35760
rect 25096 35708 25102 35760
rect 25590 35748 25596 35760
rect 25424 35720 25596 35748
rect 25133 35683 25191 35689
rect 25133 35678 25145 35683
rect 24964 35650 25145 35678
rect 25133 35649 25145 35650
rect 25179 35649 25191 35683
rect 25133 35643 25191 35649
rect 25222 35640 25228 35692
rect 25280 35640 25286 35692
rect 25424 35612 25452 35720
rect 25590 35708 25596 35720
rect 25648 35748 25654 35760
rect 25648 35720 25820 35748
rect 25648 35708 25654 35720
rect 25792 35689 25820 35720
rect 28718 35708 28724 35760
rect 28776 35708 28782 35760
rect 25685 35683 25743 35689
rect 25685 35649 25697 35683
rect 25731 35649 25743 35683
rect 25685 35643 25743 35649
rect 25777 35683 25835 35689
rect 25777 35649 25789 35683
rect 25823 35649 25835 35683
rect 25777 35643 25835 35649
rect 25332 35584 25452 35612
rect 24136 35516 25084 35544
rect 23440 35504 23446 35516
rect 21450 35476 21456 35488
rect 18800 35448 21456 35476
rect 21450 35436 21456 35448
rect 21508 35436 21514 35488
rect 21818 35436 21824 35488
rect 21876 35436 21882 35488
rect 23014 35436 23020 35488
rect 23072 35436 23078 35488
rect 23474 35436 23480 35488
rect 23532 35436 23538 35488
rect 23569 35479 23627 35485
rect 23569 35445 23581 35479
rect 23615 35476 23627 35479
rect 24118 35476 24124 35488
rect 23615 35448 24124 35476
rect 23615 35445 23627 35448
rect 23569 35439 23627 35445
rect 24118 35436 24124 35448
rect 24176 35436 24182 35488
rect 25056 35476 25084 35516
rect 25332 35476 25360 35584
rect 25498 35572 25504 35624
rect 25556 35572 25562 35624
rect 25590 35572 25596 35624
rect 25648 35612 25654 35624
rect 25700 35612 25728 35643
rect 25866 35640 25872 35692
rect 25924 35680 25930 35692
rect 25961 35683 26019 35689
rect 25961 35680 25973 35683
rect 25924 35652 25973 35680
rect 25924 35640 25930 35652
rect 25961 35649 25973 35652
rect 26007 35649 26019 35683
rect 25961 35643 26019 35649
rect 26050 35640 26056 35692
rect 26108 35680 26114 35692
rect 26145 35683 26203 35689
rect 26145 35680 26157 35683
rect 26108 35652 26157 35680
rect 26108 35640 26114 35652
rect 26145 35649 26157 35652
rect 26191 35649 26203 35683
rect 26145 35643 26203 35649
rect 26234 35640 26240 35692
rect 26292 35640 26298 35692
rect 26421 35683 26479 35689
rect 26421 35649 26433 35683
rect 26467 35649 26479 35683
rect 26421 35643 26479 35649
rect 25648 35584 25728 35612
rect 26436 35612 26464 35643
rect 26510 35640 26516 35692
rect 26568 35640 26574 35692
rect 27338 35640 27344 35692
rect 27396 35640 27402 35692
rect 29564 35680 29592 35788
rect 30466 35748 30472 35760
rect 29656 35720 30472 35748
rect 29656 35689 29684 35720
rect 30466 35708 30472 35720
rect 30524 35708 30530 35760
rect 28966 35652 29592 35680
rect 29641 35683 29699 35689
rect 27356 35612 27384 35640
rect 26436 35584 27384 35612
rect 25648 35572 25654 35584
rect 27430 35572 27436 35624
rect 27488 35572 27494 35624
rect 27709 35615 27767 35621
rect 27709 35581 27721 35615
rect 27755 35612 27767 35615
rect 28166 35612 28172 35624
rect 27755 35584 28172 35612
rect 27755 35581 27767 35584
rect 27709 35575 27767 35581
rect 28166 35572 28172 35584
rect 28224 35572 28230 35624
rect 28258 35572 28264 35624
rect 28316 35612 28322 35624
rect 28966 35612 28994 35652
rect 29641 35649 29653 35683
rect 29687 35649 29699 35683
rect 29641 35643 29699 35649
rect 29734 35683 29792 35689
rect 29734 35649 29746 35683
rect 29780 35649 29792 35683
rect 29734 35643 29792 35649
rect 29748 35612 29776 35643
rect 29822 35640 29828 35692
rect 29880 35680 29886 35692
rect 29917 35683 29975 35689
rect 29917 35680 29929 35683
rect 29880 35652 29929 35680
rect 29880 35640 29886 35652
rect 29917 35649 29929 35652
rect 29963 35649 29975 35683
rect 29917 35643 29975 35649
rect 30006 35640 30012 35692
rect 30064 35640 30070 35692
rect 30190 35689 30196 35692
rect 30147 35683 30196 35689
rect 30147 35649 30159 35683
rect 30193 35649 30196 35683
rect 30147 35643 30196 35649
rect 30190 35640 30196 35643
rect 30248 35640 30254 35692
rect 30561 35683 30619 35689
rect 30561 35680 30573 35683
rect 30300 35652 30573 35680
rect 28316 35584 28994 35612
rect 29656 35584 29776 35612
rect 28316 35572 28322 35584
rect 29656 35488 29684 35584
rect 30300 35553 30328 35652
rect 30561 35649 30573 35652
rect 30607 35649 30619 35683
rect 30668 35680 30696 35788
rect 30742 35776 30748 35828
rect 30800 35776 30806 35828
rect 32582 35708 32588 35760
rect 32640 35708 32646 35760
rect 30837 35683 30895 35689
rect 30837 35680 30849 35683
rect 30668 35652 30849 35680
rect 30561 35643 30619 35649
rect 30837 35649 30849 35652
rect 30883 35649 30895 35683
rect 30837 35643 30895 35649
rect 30852 35612 30880 35643
rect 31386 35640 31392 35692
rect 31444 35640 31450 35692
rect 32600 35680 32628 35708
rect 32953 35683 33011 35689
rect 32953 35680 32965 35683
rect 32600 35652 32965 35680
rect 32953 35649 32965 35652
rect 32999 35649 33011 35683
rect 32953 35643 33011 35649
rect 33502 35640 33508 35692
rect 33560 35640 33566 35692
rect 31478 35612 31484 35624
rect 30852 35584 31484 35612
rect 31478 35572 31484 35584
rect 31536 35572 31542 35624
rect 30285 35547 30343 35553
rect 30285 35513 30297 35547
rect 30331 35513 30343 35547
rect 30285 35507 30343 35513
rect 25056 35448 25360 35476
rect 25409 35479 25467 35485
rect 25409 35445 25421 35479
rect 25455 35476 25467 35479
rect 26142 35476 26148 35488
rect 25455 35448 26148 35476
rect 25455 35445 25467 35448
rect 25409 35439 25467 35445
rect 26142 35436 26148 35448
rect 26200 35436 26206 35488
rect 26602 35436 26608 35488
rect 26660 35476 26666 35488
rect 26697 35479 26755 35485
rect 26697 35476 26709 35479
rect 26660 35448 26709 35476
rect 26660 35436 26666 35448
rect 26697 35445 26709 35448
rect 26743 35445 26755 35479
rect 26697 35439 26755 35445
rect 26878 35436 26884 35488
rect 26936 35476 26942 35488
rect 29638 35476 29644 35488
rect 26936 35448 29644 35476
rect 26936 35436 26942 35448
rect 29638 35436 29644 35448
rect 29696 35436 29702 35488
rect 30098 35436 30104 35488
rect 30156 35476 30162 35488
rect 30377 35479 30435 35485
rect 30377 35476 30389 35479
rect 30156 35448 30389 35476
rect 30156 35436 30162 35448
rect 30377 35445 30389 35448
rect 30423 35445 30435 35479
rect 30377 35439 30435 35445
rect 31018 35436 31024 35488
rect 31076 35476 31082 35488
rect 31205 35479 31263 35485
rect 31205 35476 31217 35479
rect 31076 35448 31217 35476
rect 31076 35436 31082 35448
rect 31205 35445 31217 35448
rect 31251 35445 31263 35479
rect 31205 35439 31263 35445
rect 32766 35436 32772 35488
rect 32824 35476 32830 35488
rect 32861 35479 32919 35485
rect 32861 35476 32873 35479
rect 32824 35448 32873 35476
rect 32824 35436 32830 35448
rect 32861 35445 32873 35448
rect 32907 35445 32919 35479
rect 32861 35439 32919 35445
rect 33318 35436 33324 35488
rect 33376 35436 33382 35488
rect 1104 35386 38272 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 38272 35386
rect 1104 35312 38272 35334
rect 9493 35275 9551 35281
rect 9493 35241 9505 35275
rect 9539 35272 9551 35275
rect 9766 35272 9772 35284
rect 9539 35244 9772 35272
rect 9539 35241 9551 35244
rect 9493 35235 9551 35241
rect 9766 35232 9772 35244
rect 9824 35232 9830 35284
rect 17497 35275 17555 35281
rect 17497 35241 17509 35275
rect 17543 35272 17555 35275
rect 18874 35272 18880 35284
rect 17543 35244 18880 35272
rect 17543 35241 17555 35244
rect 17497 35235 17555 35241
rect 18874 35232 18880 35244
rect 18932 35232 18938 35284
rect 27982 35232 27988 35284
rect 28040 35272 28046 35284
rect 30190 35272 30196 35284
rect 28040 35244 30196 35272
rect 28040 35232 28046 35244
rect 30190 35232 30196 35244
rect 30248 35272 30254 35284
rect 30650 35272 30656 35284
rect 30248 35244 30656 35272
rect 30248 35232 30254 35244
rect 30650 35232 30656 35244
rect 30708 35232 30714 35284
rect 30760 35244 32352 35272
rect 6914 35164 6920 35216
rect 6972 35164 6978 35216
rect 22830 35164 22836 35216
rect 22888 35204 22894 35216
rect 22888 35176 23704 35204
rect 22888 35164 22894 35176
rect 6932 35136 6960 35164
rect 6656 35108 6960 35136
rect 6656 35077 6684 35108
rect 7926 35096 7932 35148
rect 7984 35136 7990 35148
rect 7984 35108 8524 35136
rect 7984 35096 7990 35108
rect 6641 35071 6699 35077
rect 6641 35037 6653 35071
rect 6687 35037 6699 35071
rect 6641 35031 6699 35037
rect 6733 35071 6791 35077
rect 6733 35037 6745 35071
rect 6779 35068 6791 35071
rect 6917 35071 6975 35077
rect 6917 35068 6929 35071
rect 6779 35040 6929 35068
rect 6779 35037 6791 35040
rect 6733 35031 6791 35037
rect 6917 35037 6929 35040
rect 6963 35037 6975 35071
rect 6917 35031 6975 35037
rect 8294 35028 8300 35080
rect 8352 35028 8358 35080
rect 8496 35068 8524 35108
rect 9674 35096 9680 35148
rect 9732 35136 9738 35148
rect 10137 35139 10195 35145
rect 10137 35136 10149 35139
rect 9732 35108 10149 35136
rect 9732 35096 9738 35108
rect 10137 35105 10149 35108
rect 10183 35136 10195 35139
rect 10778 35136 10784 35148
rect 10183 35108 10784 35136
rect 10183 35105 10195 35108
rect 10137 35099 10195 35105
rect 10778 35096 10784 35108
rect 10836 35096 10842 35148
rect 23566 35096 23572 35148
rect 23624 35096 23630 35148
rect 23676 35145 23704 35176
rect 24118 35164 24124 35216
rect 24176 35164 24182 35216
rect 25332 35176 26740 35204
rect 23661 35139 23719 35145
rect 23661 35105 23673 35139
rect 23707 35105 23719 35139
rect 23661 35099 23719 35105
rect 9953 35071 10011 35077
rect 9953 35068 9965 35071
rect 8496 35040 9965 35068
rect 9953 35037 9965 35040
rect 9999 35037 10011 35071
rect 9953 35031 10011 35037
rect 11146 35028 11152 35080
rect 11204 35068 11210 35080
rect 11204 35040 17264 35068
rect 11204 35028 11210 35040
rect 7190 34960 7196 35012
rect 7248 34960 7254 35012
rect 9861 35003 9919 35009
rect 9861 34969 9873 35003
rect 9907 35000 9919 35003
rect 12434 35000 12440 35012
rect 9907 34972 12440 35000
rect 9907 34969 9919 34972
rect 9861 34963 9919 34969
rect 12434 34960 12440 34972
rect 12492 34960 12498 35012
rect 17236 35000 17264 35040
rect 17310 35028 17316 35080
rect 17368 35028 17374 35080
rect 23293 35071 23351 35077
rect 23293 35037 23305 35071
rect 23339 35037 23351 35071
rect 23293 35031 23351 35037
rect 23477 35071 23535 35077
rect 23477 35037 23489 35071
rect 23523 35037 23535 35071
rect 23477 35031 23535 35037
rect 23753 35071 23811 35077
rect 23753 35037 23765 35071
rect 23799 35068 23811 35071
rect 24136 35068 24164 35164
rect 25332 35080 25360 35176
rect 25608 35108 26464 35136
rect 23799 35040 24164 35068
rect 23799 35037 23811 35040
rect 23753 35031 23811 35037
rect 21818 35000 21824 35012
rect 17236 34972 21824 35000
rect 21818 34960 21824 34972
rect 21876 34960 21882 35012
rect 8478 34892 8484 34944
rect 8536 34932 8542 34944
rect 8665 34935 8723 34941
rect 8665 34932 8677 34935
rect 8536 34904 8677 34932
rect 8536 34892 8542 34904
rect 8665 34901 8677 34904
rect 8711 34901 8723 34935
rect 8665 34895 8723 34901
rect 15930 34892 15936 34944
rect 15988 34932 15994 34944
rect 19334 34932 19340 34944
rect 15988 34904 19340 34932
rect 15988 34892 15994 34904
rect 19334 34892 19340 34904
rect 19392 34892 19398 34944
rect 20714 34892 20720 34944
rect 20772 34932 20778 34944
rect 23308 34932 23336 35031
rect 23492 35000 23520 35031
rect 25314 35028 25320 35080
rect 25372 35028 25378 35080
rect 25498 35028 25504 35080
rect 25556 35028 25562 35080
rect 25608 35077 25636 35108
rect 26436 35080 26464 35108
rect 26602 35096 26608 35148
rect 26660 35096 26666 35148
rect 25593 35071 25651 35077
rect 25593 35037 25605 35071
rect 25639 35037 25651 35071
rect 25593 35031 25651 35037
rect 25685 35071 25743 35077
rect 25685 35037 25697 35071
rect 25731 35068 25743 35071
rect 25866 35068 25872 35080
rect 25731 35040 25872 35068
rect 25731 35037 25743 35040
rect 25685 35031 25743 35037
rect 25700 35000 25728 35031
rect 25866 35028 25872 35040
rect 25924 35028 25930 35080
rect 26326 35028 26332 35080
rect 26384 35028 26390 35080
rect 26418 35028 26424 35080
rect 26476 35028 26482 35080
rect 26513 35071 26571 35077
rect 26513 35037 26525 35071
rect 26559 35068 26571 35071
rect 26620 35068 26648 35096
rect 26712 35077 26740 35176
rect 28166 35164 28172 35216
rect 28224 35164 28230 35216
rect 28350 35164 28356 35216
rect 28408 35204 28414 35216
rect 30760 35204 30788 35244
rect 32324 35216 32352 35244
rect 32766 35232 32772 35284
rect 32824 35232 32830 35284
rect 28408 35176 30788 35204
rect 28408 35164 28414 35176
rect 32306 35164 32312 35216
rect 32364 35164 32370 35216
rect 27525 35139 27583 35145
rect 27525 35105 27537 35139
rect 27571 35136 27583 35139
rect 30929 35139 30987 35145
rect 27571 35108 30328 35136
rect 27571 35105 27583 35108
rect 27525 35099 27583 35105
rect 26559 35040 26648 35068
rect 26697 35071 26755 35077
rect 26559 35037 26571 35040
rect 26513 35031 26571 35037
rect 26697 35037 26709 35071
rect 26743 35037 26755 35071
rect 26697 35031 26755 35037
rect 28353 35071 28411 35077
rect 28353 35037 28365 35071
rect 28399 35037 28411 35071
rect 28353 35031 28411 35037
rect 26053 35003 26111 35009
rect 26053 35000 26065 35003
rect 23492 34972 25728 35000
rect 25884 34972 26065 35000
rect 23474 34932 23480 34944
rect 20772 34904 23480 34932
rect 20772 34892 20778 34904
rect 23474 34892 23480 34904
rect 23532 34892 23538 34944
rect 23566 34892 23572 34944
rect 23624 34932 23630 34944
rect 23937 34935 23995 34941
rect 23937 34932 23949 34935
rect 23624 34904 23949 34932
rect 23624 34892 23630 34904
rect 23937 34901 23949 34904
rect 23983 34901 23995 34935
rect 23937 34895 23995 34901
rect 25682 34892 25688 34944
rect 25740 34932 25746 34944
rect 25884 34932 25912 34972
rect 26053 34969 26065 34972
rect 26099 34969 26111 35003
rect 27522 35000 27528 35012
rect 26053 34963 26111 34969
rect 27356 34972 27528 35000
rect 27356 34944 27384 34972
rect 27522 34960 27528 34972
rect 27580 35000 27586 35012
rect 27709 35003 27767 35009
rect 27709 35000 27721 35003
rect 27580 34972 27721 35000
rect 27580 34960 27586 34972
rect 27709 34969 27721 34972
rect 27755 34969 27767 35003
rect 28368 35000 28396 35031
rect 28902 35028 28908 35080
rect 28960 35028 28966 35080
rect 27709 34963 27767 34969
rect 28092 34972 28396 35000
rect 25740 34904 25912 34932
rect 25740 34892 25746 34904
rect 25958 34892 25964 34944
rect 26016 34892 26022 34944
rect 27338 34892 27344 34944
rect 27396 34892 27402 34944
rect 27617 34935 27675 34941
rect 27617 34901 27629 34935
rect 27663 34932 27675 34935
rect 27798 34932 27804 34944
rect 27663 34904 27804 34932
rect 27663 34901 27675 34904
rect 27617 34895 27675 34901
rect 27798 34892 27804 34904
rect 27856 34892 27862 34944
rect 28092 34941 28120 34972
rect 28077 34935 28135 34941
rect 28077 34901 28089 34935
rect 28123 34901 28135 34935
rect 28077 34895 28135 34901
rect 28810 34892 28816 34944
rect 28868 34892 28874 34944
rect 30300 34932 30328 35108
rect 30929 35105 30941 35139
rect 30975 35136 30987 35139
rect 31018 35136 31024 35148
rect 30975 35108 31024 35136
rect 30975 35105 30987 35108
rect 30929 35099 30987 35105
rect 31018 35096 31024 35108
rect 31076 35096 31082 35148
rect 32677 35139 32735 35145
rect 32677 35105 32689 35139
rect 32723 35136 32735 35139
rect 32784 35136 32812 35232
rect 32723 35108 32812 35136
rect 32953 35139 33011 35145
rect 32723 35105 32735 35108
rect 32677 35099 32735 35105
rect 32953 35105 32965 35139
rect 32999 35136 33011 35139
rect 33318 35136 33324 35148
rect 32999 35108 33324 35136
rect 32999 35105 33011 35108
rect 32953 35099 33011 35105
rect 33318 35096 33324 35108
rect 33376 35096 33382 35148
rect 33410 35096 33416 35148
rect 33468 35136 33474 35148
rect 33686 35136 33692 35148
rect 33468 35108 33692 35136
rect 33468 35096 33474 35108
rect 33686 35096 33692 35108
rect 33744 35096 33750 35148
rect 30374 35028 30380 35080
rect 30432 35028 30438 35080
rect 30469 35071 30527 35077
rect 30469 35037 30481 35071
rect 30515 35068 30527 35071
rect 30653 35071 30711 35077
rect 30653 35068 30665 35071
rect 30515 35040 30665 35068
rect 30515 35037 30527 35040
rect 30469 35031 30527 35037
rect 30653 35037 30665 35040
rect 30699 35037 30711 35071
rect 30653 35031 30711 35037
rect 32490 35000 32496 35012
rect 32154 34972 32496 35000
rect 32490 34960 32496 34972
rect 32548 35000 32554 35012
rect 33410 35000 33416 35012
rect 32548 34972 33416 35000
rect 32548 34960 32554 34972
rect 33410 34960 33416 34972
rect 33468 34960 33474 35012
rect 31662 34932 31668 34944
rect 30300 34904 31668 34932
rect 31662 34892 31668 34904
rect 31720 34892 31726 34944
rect 31754 34892 31760 34944
rect 31812 34932 31818 34944
rect 32401 34935 32459 34941
rect 32401 34932 32413 34935
rect 31812 34904 32413 34932
rect 31812 34892 31818 34904
rect 32401 34901 32413 34904
rect 32447 34901 32459 34935
rect 32401 34895 32459 34901
rect 33318 34892 33324 34944
rect 33376 34932 33382 34944
rect 34425 34935 34483 34941
rect 34425 34932 34437 34935
rect 33376 34904 34437 34932
rect 33376 34892 33382 34904
rect 34425 34901 34437 34904
rect 34471 34901 34483 34935
rect 34425 34895 34483 34901
rect 1104 34842 38272 34864
rect 1104 34790 4874 34842
rect 4926 34790 4938 34842
rect 4990 34790 5002 34842
rect 5054 34790 5066 34842
rect 5118 34790 5130 34842
rect 5182 34790 35594 34842
rect 35646 34790 35658 34842
rect 35710 34790 35722 34842
rect 35774 34790 35786 34842
rect 35838 34790 35850 34842
rect 35902 34790 38272 34842
rect 1104 34768 38272 34790
rect 7190 34688 7196 34740
rect 7248 34728 7254 34740
rect 7653 34731 7711 34737
rect 7653 34728 7665 34731
rect 7248 34700 7665 34728
rect 7248 34688 7254 34700
rect 7653 34697 7665 34700
rect 7699 34697 7711 34731
rect 7653 34691 7711 34697
rect 7929 34731 7987 34737
rect 7929 34697 7941 34731
rect 7975 34697 7987 34731
rect 12158 34728 12164 34740
rect 7929 34691 7987 34697
rect 11348 34700 12164 34728
rect 5626 34552 5632 34604
rect 5684 34552 5690 34604
rect 7837 34595 7895 34601
rect 7837 34561 7849 34595
rect 7883 34592 7895 34595
rect 7944 34592 7972 34691
rect 8202 34620 8208 34672
rect 8260 34660 8266 34672
rect 8260 34632 9904 34660
rect 8260 34620 8266 34632
rect 8297 34595 8355 34601
rect 8297 34592 8309 34595
rect 7883 34564 7972 34592
rect 8220 34564 8309 34592
rect 7883 34561 7895 34564
rect 7837 34555 7895 34561
rect 8220 34536 8248 34564
rect 8297 34561 8309 34564
rect 8343 34561 8355 34595
rect 8297 34555 8355 34561
rect 8386 34552 8392 34604
rect 8444 34552 8450 34604
rect 8202 34484 8208 34536
rect 8260 34484 8266 34536
rect 8573 34527 8631 34533
rect 8573 34493 8585 34527
rect 8619 34493 8631 34527
rect 9876 34524 9904 34632
rect 11348 34592 11376 34700
rect 12158 34688 12164 34700
rect 12216 34728 12222 34740
rect 12618 34728 12624 34740
rect 12216 34700 12624 34728
rect 12216 34688 12222 34700
rect 12618 34688 12624 34700
rect 12676 34688 12682 34740
rect 16853 34731 16911 34737
rect 16853 34697 16865 34731
rect 16899 34728 16911 34731
rect 17310 34728 17316 34740
rect 16899 34700 17316 34728
rect 16899 34697 16911 34700
rect 16853 34691 16911 34697
rect 17310 34688 17316 34700
rect 17368 34688 17374 34740
rect 23750 34728 23756 34740
rect 21008 34700 23756 34728
rect 11422 34620 11428 34672
rect 11480 34660 11486 34672
rect 11882 34660 11888 34672
rect 11480 34632 11888 34660
rect 11480 34620 11486 34632
rect 11882 34620 11888 34632
rect 11940 34620 11946 34672
rect 16482 34660 16488 34672
rect 11992 34632 16488 34660
rect 11655 34595 11713 34601
rect 11655 34592 11667 34595
rect 11348 34564 11667 34592
rect 11655 34561 11667 34564
rect 11701 34561 11713 34595
rect 11655 34555 11713 34561
rect 11793 34595 11851 34601
rect 11793 34561 11805 34595
rect 11839 34592 11851 34595
rect 11992 34592 12020 34632
rect 16482 34620 16488 34632
rect 16540 34620 16546 34672
rect 16942 34620 16948 34672
rect 17000 34660 17006 34672
rect 17954 34660 17960 34672
rect 17000 34632 17960 34660
rect 17000 34620 17006 34632
rect 17954 34620 17960 34632
rect 18012 34620 18018 34672
rect 20898 34620 20904 34672
rect 20956 34660 20962 34672
rect 21008 34669 21036 34700
rect 21266 34669 21272 34672
rect 20993 34663 21051 34669
rect 20993 34660 21005 34663
rect 20956 34632 21005 34660
rect 20956 34620 20962 34632
rect 20993 34629 21005 34632
rect 21039 34629 21051 34663
rect 20993 34623 21051 34629
rect 21209 34663 21272 34669
rect 21209 34629 21221 34663
rect 21255 34629 21272 34663
rect 21209 34623 21272 34629
rect 21266 34620 21272 34623
rect 21324 34620 21330 34672
rect 21818 34620 21824 34672
rect 21876 34660 21882 34672
rect 22278 34660 22284 34672
rect 21876 34632 22284 34660
rect 21876 34620 21882 34632
rect 22278 34620 22284 34632
rect 22336 34620 22342 34672
rect 11839 34564 12020 34592
rect 12068 34595 12126 34601
rect 11839 34561 11851 34564
rect 11793 34555 11851 34561
rect 12068 34561 12080 34595
rect 12114 34561 12126 34595
rect 12068 34555 12126 34561
rect 12161 34595 12219 34601
rect 12161 34561 12173 34595
rect 12207 34592 12219 34595
rect 12250 34592 12256 34604
rect 12207 34564 12256 34592
rect 12207 34561 12219 34564
rect 12161 34555 12219 34561
rect 11808 34524 11836 34555
rect 9876 34496 11836 34524
rect 12084 34524 12112 34555
rect 12250 34552 12256 34564
rect 12308 34592 12314 34604
rect 12710 34592 12716 34604
rect 12308 34564 12716 34592
rect 12308 34552 12314 34564
rect 12710 34552 12716 34564
rect 12768 34552 12774 34604
rect 16574 34552 16580 34604
rect 16632 34592 16638 34604
rect 17129 34595 17187 34601
rect 17129 34592 17141 34595
rect 16632 34564 17141 34592
rect 16632 34552 16638 34564
rect 17129 34561 17141 34564
rect 17175 34561 17187 34595
rect 17129 34555 17187 34561
rect 12434 34524 12440 34536
rect 12084 34496 12440 34524
rect 8573 34487 8631 34493
rect 8588 34456 8616 34487
rect 12406 34484 12440 34496
rect 12492 34484 12498 34536
rect 17144 34524 17172 34555
rect 17310 34552 17316 34604
rect 17368 34592 17374 34604
rect 17678 34592 17684 34604
rect 17368 34564 17684 34592
rect 17368 34552 17374 34564
rect 17678 34552 17684 34564
rect 17736 34552 17742 34604
rect 22094 34601 22100 34604
rect 21913 34595 21971 34601
rect 21913 34592 21925 34595
rect 21376 34564 21925 34592
rect 17770 34524 17776 34536
rect 17144 34496 17776 34524
rect 17770 34484 17776 34496
rect 17828 34484 17834 34536
rect 9490 34456 9496 34468
rect 8588 34428 9496 34456
rect 9490 34416 9496 34428
rect 9548 34456 9554 34468
rect 9858 34456 9864 34468
rect 9548 34428 9864 34456
rect 9548 34416 9554 34428
rect 9858 34416 9864 34428
rect 9916 34416 9922 34468
rect 12406 34456 12434 34484
rect 13630 34456 13636 34468
rect 12406 34428 13636 34456
rect 13630 34416 13636 34428
rect 13688 34456 13694 34468
rect 21376 34465 21404 34564
rect 21913 34561 21925 34564
rect 21959 34561 21971 34595
rect 21913 34555 21971 34561
rect 22061 34595 22100 34601
rect 22061 34561 22073 34595
rect 22061 34555 22100 34561
rect 22094 34552 22100 34555
rect 22152 34552 22158 34604
rect 22189 34595 22247 34601
rect 22189 34561 22201 34595
rect 22235 34561 22247 34595
rect 22189 34555 22247 34561
rect 22378 34595 22436 34601
rect 22378 34561 22390 34595
rect 22424 34592 22436 34595
rect 22830 34592 22836 34604
rect 22424 34564 22836 34592
rect 22424 34561 22436 34564
rect 22378 34555 22436 34561
rect 22204 34524 22232 34555
rect 22830 34552 22836 34564
rect 22888 34552 22894 34604
rect 23124 34592 23152 34700
rect 23750 34688 23756 34700
rect 23808 34688 23814 34740
rect 25222 34688 25228 34740
rect 25280 34728 25286 34740
rect 25958 34728 25964 34740
rect 25280 34700 25964 34728
rect 25280 34688 25286 34700
rect 25958 34688 25964 34700
rect 26016 34688 26022 34740
rect 28810 34688 28816 34740
rect 28868 34688 28874 34740
rect 31205 34731 31263 34737
rect 31205 34697 31217 34731
rect 31251 34728 31263 34731
rect 31386 34728 31392 34740
rect 31251 34700 31392 34728
rect 31251 34697 31263 34700
rect 31205 34691 31263 34697
rect 31386 34688 31392 34700
rect 31444 34688 31450 34740
rect 33318 34688 33324 34740
rect 33376 34688 33382 34740
rect 33502 34688 33508 34740
rect 33560 34728 33566 34740
rect 33689 34731 33747 34737
rect 33689 34728 33701 34731
rect 33560 34700 33701 34728
rect 33560 34688 33566 34700
rect 33689 34697 33701 34700
rect 33735 34697 33747 34731
rect 33689 34691 33747 34697
rect 23198 34620 23204 34672
rect 23256 34660 23262 34672
rect 23661 34663 23719 34669
rect 23661 34660 23673 34663
rect 23256 34632 23673 34660
rect 23256 34620 23262 34632
rect 23661 34629 23673 34632
rect 23707 34629 23719 34663
rect 23661 34623 23719 34629
rect 28534 34620 28540 34672
rect 28592 34620 28598 34672
rect 28828 34660 28856 34688
rect 28644 34632 28856 34660
rect 31665 34663 31723 34669
rect 23385 34595 23443 34601
rect 23385 34592 23397 34595
rect 23124 34564 23397 34592
rect 23385 34561 23397 34564
rect 23431 34561 23443 34595
rect 23385 34555 23443 34561
rect 23569 34595 23627 34601
rect 23569 34561 23581 34595
rect 23615 34561 23627 34595
rect 23569 34555 23627 34561
rect 23753 34595 23811 34601
rect 23753 34561 23765 34595
rect 23799 34592 23811 34595
rect 24118 34592 24124 34604
rect 23799 34564 24124 34592
rect 23799 34561 23811 34564
rect 23753 34555 23811 34561
rect 22020 34496 22232 34524
rect 23584 34524 23612 34555
rect 24118 34552 24124 34564
rect 24176 34592 24182 34604
rect 28258 34592 28264 34604
rect 24176 34564 28264 34592
rect 24176 34552 24182 34564
rect 28258 34552 28264 34564
rect 28316 34552 28322 34604
rect 27154 34524 27160 34536
rect 23584 34496 27160 34524
rect 21361 34459 21419 34465
rect 13688 34428 18092 34456
rect 13688 34416 13694 34428
rect 18064 34400 18092 34428
rect 21361 34425 21373 34459
rect 21407 34425 21419 34459
rect 21361 34419 21419 34425
rect 22020 34400 22048 34496
rect 27154 34484 27160 34496
rect 27212 34484 27218 34536
rect 28552 34524 28580 34620
rect 28644 34601 28672 34632
rect 31665 34629 31677 34663
rect 31711 34660 31723 34663
rect 31754 34660 31760 34672
rect 31711 34632 31760 34660
rect 31711 34629 31723 34632
rect 31665 34623 31723 34629
rect 31754 34620 31760 34632
rect 31812 34620 31818 34672
rect 28629 34595 28687 34601
rect 28629 34561 28641 34595
rect 28675 34561 28687 34595
rect 28629 34555 28687 34561
rect 30024 34524 30052 34578
rect 30926 34552 30932 34604
rect 30984 34592 30990 34604
rect 31573 34595 31631 34601
rect 31573 34592 31585 34595
rect 30984 34564 31585 34592
rect 30984 34552 30990 34564
rect 31573 34561 31585 34564
rect 31619 34592 31631 34595
rect 33229 34595 33287 34601
rect 33229 34592 33241 34595
rect 31619 34564 33241 34592
rect 31619 34561 31631 34564
rect 31573 34555 31631 34561
rect 33229 34561 33241 34564
rect 33275 34592 33287 34595
rect 34146 34592 34152 34604
rect 33275 34564 34152 34592
rect 33275 34561 33287 34564
rect 33229 34555 33287 34561
rect 34146 34552 34152 34564
rect 34204 34552 34210 34604
rect 36906 34552 36912 34604
rect 36964 34592 36970 34604
rect 37553 34595 37611 34601
rect 37553 34592 37565 34595
rect 36964 34564 37565 34592
rect 36964 34552 36970 34564
rect 37553 34561 37565 34564
rect 37599 34561 37611 34595
rect 37553 34555 37611 34561
rect 28552 34496 30052 34524
rect 23474 34416 23480 34468
rect 23532 34456 23538 34468
rect 27982 34456 27988 34468
rect 23532 34428 27988 34456
rect 23532 34416 23538 34428
rect 27982 34416 27988 34428
rect 28040 34416 28046 34468
rect 30024 34456 30052 34496
rect 31846 34484 31852 34536
rect 31904 34484 31910 34536
rect 32398 34484 32404 34536
rect 32456 34524 32462 34536
rect 33137 34527 33195 34533
rect 33137 34524 33149 34527
rect 32456 34496 33149 34524
rect 32456 34484 32462 34496
rect 33137 34493 33149 34496
rect 33183 34493 33195 34527
rect 33137 34487 33195 34493
rect 37829 34527 37887 34533
rect 37829 34493 37841 34527
rect 37875 34524 37887 34527
rect 37918 34524 37924 34536
rect 37875 34496 37924 34524
rect 37875 34493 37887 34496
rect 37829 34487 37887 34493
rect 30190 34456 30196 34468
rect 30024 34428 30196 34456
rect 30190 34416 30196 34428
rect 30248 34416 30254 34468
rect 33152 34456 33180 34487
rect 37918 34484 37924 34496
rect 37976 34484 37982 34536
rect 33152 34428 33364 34456
rect 33336 34400 33364 34428
rect 5350 34348 5356 34400
rect 5408 34388 5414 34400
rect 5445 34391 5503 34397
rect 5445 34388 5457 34391
rect 5408 34360 5457 34388
rect 5408 34348 5414 34360
rect 5445 34357 5457 34360
rect 5491 34357 5503 34391
rect 5445 34351 5503 34357
rect 11514 34348 11520 34400
rect 11572 34348 11578 34400
rect 16850 34348 16856 34400
rect 16908 34348 16914 34400
rect 16942 34348 16948 34400
rect 17000 34348 17006 34400
rect 17034 34348 17040 34400
rect 17092 34348 17098 34400
rect 18046 34348 18052 34400
rect 18104 34348 18110 34400
rect 20622 34348 20628 34400
rect 20680 34388 20686 34400
rect 21177 34391 21235 34397
rect 21177 34388 21189 34391
rect 20680 34360 21189 34388
rect 20680 34348 20686 34360
rect 21177 34357 21189 34360
rect 21223 34357 21235 34391
rect 21177 34351 21235 34357
rect 22002 34348 22008 34400
rect 22060 34348 22066 34400
rect 22557 34391 22615 34397
rect 22557 34357 22569 34391
rect 22603 34388 22615 34391
rect 22646 34388 22652 34400
rect 22603 34360 22652 34388
rect 22603 34357 22615 34360
rect 22557 34351 22615 34357
rect 22646 34348 22652 34360
rect 22704 34348 22710 34400
rect 23750 34348 23756 34400
rect 23808 34388 23814 34400
rect 23937 34391 23995 34397
rect 23937 34388 23949 34391
rect 23808 34360 23949 34388
rect 23808 34348 23814 34360
rect 23937 34357 23949 34360
rect 23983 34357 23995 34391
rect 23937 34351 23995 34357
rect 24762 34348 24768 34400
rect 24820 34388 24826 34400
rect 27246 34388 27252 34400
rect 24820 34360 27252 34388
rect 24820 34348 24826 34360
rect 27246 34348 27252 34360
rect 27304 34348 27310 34400
rect 28074 34348 28080 34400
rect 28132 34388 28138 34400
rect 28886 34391 28944 34397
rect 28886 34388 28898 34391
rect 28132 34360 28898 34388
rect 28132 34348 28138 34360
rect 28886 34357 28898 34360
rect 28932 34357 28944 34391
rect 28886 34351 28944 34357
rect 30006 34348 30012 34400
rect 30064 34388 30070 34400
rect 30377 34391 30435 34397
rect 30377 34388 30389 34391
rect 30064 34360 30389 34388
rect 30064 34348 30070 34360
rect 30377 34357 30389 34360
rect 30423 34388 30435 34391
rect 30558 34388 30564 34400
rect 30423 34360 30564 34388
rect 30423 34357 30435 34360
rect 30377 34351 30435 34357
rect 30558 34348 30564 34360
rect 30616 34348 30622 34400
rect 33318 34348 33324 34400
rect 33376 34348 33382 34400
rect 1104 34298 38272 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 38272 34298
rect 1104 34224 38272 34246
rect 6730 34144 6736 34196
rect 6788 34184 6794 34196
rect 12066 34184 12072 34196
rect 6788 34156 12072 34184
rect 6788 34144 6794 34156
rect 12066 34144 12072 34156
rect 12124 34144 12130 34196
rect 14642 34144 14648 34196
rect 14700 34144 14706 34196
rect 14826 34144 14832 34196
rect 14884 34144 14890 34196
rect 16669 34187 16727 34193
rect 16669 34153 16681 34187
rect 16715 34184 16727 34187
rect 16850 34184 16856 34196
rect 16715 34156 16856 34184
rect 16715 34153 16727 34156
rect 16669 34147 16727 34153
rect 16850 34144 16856 34156
rect 16908 34144 16914 34196
rect 16942 34144 16948 34196
rect 17000 34144 17006 34196
rect 17034 34144 17040 34196
rect 17092 34144 17098 34196
rect 20530 34144 20536 34196
rect 20588 34184 20594 34196
rect 22094 34184 22100 34196
rect 20588 34156 22100 34184
rect 20588 34144 20594 34156
rect 22094 34144 22100 34156
rect 22152 34144 22158 34196
rect 22462 34144 22468 34196
rect 22520 34184 22526 34196
rect 23106 34184 23112 34196
rect 22520 34156 23112 34184
rect 22520 34144 22526 34156
rect 23106 34144 23112 34156
rect 23164 34144 23170 34196
rect 23400 34156 23612 34184
rect 11609 34119 11667 34125
rect 11609 34085 11621 34119
rect 11655 34116 11667 34119
rect 15010 34116 15016 34128
rect 11655 34088 15016 34116
rect 11655 34085 11667 34088
rect 11609 34079 11667 34085
rect 15010 34076 15016 34088
rect 15068 34076 15074 34128
rect 15933 34119 15991 34125
rect 15933 34085 15945 34119
rect 15979 34116 15991 34119
rect 16960 34116 16988 34144
rect 15979 34088 16988 34116
rect 15979 34085 15991 34088
rect 15933 34079 15991 34085
rect 5261 34051 5319 34057
rect 5261 34017 5273 34051
rect 5307 34048 5319 34051
rect 5350 34048 5356 34060
rect 5307 34020 5356 34048
rect 5307 34017 5319 34020
rect 5261 34011 5319 34017
rect 5350 34008 5356 34020
rect 5408 34008 5414 34060
rect 6914 34008 6920 34060
rect 6972 34048 6978 34060
rect 6972 34020 7328 34048
rect 6972 34008 6978 34020
rect 4706 33940 4712 33992
rect 4764 33940 4770 33992
rect 4801 33983 4859 33989
rect 4801 33949 4813 33983
rect 4847 33980 4859 33983
rect 4985 33983 5043 33989
rect 4985 33980 4997 33983
rect 4847 33952 4997 33980
rect 4847 33949 4859 33952
rect 4801 33943 4859 33949
rect 4985 33949 4997 33952
rect 5031 33949 5043 33983
rect 4985 33943 5043 33949
rect 6362 33940 6368 33992
rect 6420 33980 6426 33992
rect 6638 33980 6644 33992
rect 6420 33952 6644 33980
rect 6420 33940 6426 33952
rect 6638 33940 6644 33952
rect 6696 33940 6702 33992
rect 7300 33989 7328 34020
rect 8386 34008 8392 34060
rect 8444 34048 8450 34060
rect 8444 34020 9720 34048
rect 8444 34008 8450 34020
rect 7285 33983 7343 33989
rect 7285 33949 7297 33983
rect 7331 33980 7343 33983
rect 7558 33980 7564 33992
rect 7331 33952 7564 33980
rect 7331 33949 7343 33952
rect 7285 33943 7343 33949
rect 7558 33940 7564 33952
rect 7616 33940 7622 33992
rect 8573 33983 8631 33989
rect 8573 33949 8585 33983
rect 8619 33980 8631 33983
rect 9030 33980 9036 33992
rect 8619 33952 9036 33980
rect 8619 33949 8631 33952
rect 8573 33943 8631 33949
rect 9030 33940 9036 33952
rect 9088 33940 9094 33992
rect 9493 33983 9551 33989
rect 9493 33949 9505 33983
rect 9539 33980 9551 33983
rect 9539 33952 9628 33980
rect 9539 33949 9551 33952
rect 9493 33943 9551 33949
rect 9600 33924 9628 33952
rect 9582 33872 9588 33924
rect 9640 33872 9646 33924
rect 9692 33912 9720 34020
rect 11790 34008 11796 34060
rect 11848 34008 11854 34060
rect 13173 34051 13231 34057
rect 13173 34017 13185 34051
rect 13219 34048 13231 34051
rect 13630 34048 13636 34060
rect 13219 34020 13636 34048
rect 13219 34017 13231 34020
rect 13173 34011 13231 34017
rect 13630 34008 13636 34020
rect 13688 34008 13694 34060
rect 13725 34051 13783 34057
rect 13725 34017 13737 34051
rect 13771 34048 13783 34051
rect 14737 34051 14795 34057
rect 14737 34048 14749 34051
rect 13771 34020 14749 34048
rect 13771 34017 13783 34020
rect 13725 34011 13783 34017
rect 14737 34017 14749 34020
rect 14783 34017 14795 34051
rect 14737 34011 14795 34017
rect 15105 34051 15163 34057
rect 15105 34017 15117 34051
rect 15151 34048 15163 34051
rect 16853 34051 16911 34057
rect 15151 34020 16805 34048
rect 15151 34017 15163 34020
rect 15105 34011 15163 34017
rect 9858 33940 9864 33992
rect 9916 33940 9922 33992
rect 11514 33940 11520 33992
rect 11572 33980 11578 33992
rect 11609 33983 11667 33989
rect 11609 33980 11621 33983
rect 11572 33952 11621 33980
rect 11572 33940 11578 33952
rect 11609 33949 11621 33952
rect 11655 33949 11667 33983
rect 11808 33980 11836 34008
rect 11885 33983 11943 33989
rect 11885 33980 11897 33983
rect 11808 33952 11897 33980
rect 11609 33943 11667 33949
rect 11885 33949 11897 33952
rect 11931 33949 11943 33983
rect 11885 33943 11943 33949
rect 14369 33983 14427 33989
rect 14369 33949 14381 33983
rect 14415 33980 14427 33983
rect 14458 33980 14464 33992
rect 14415 33952 14464 33980
rect 14415 33949 14427 33952
rect 14369 33943 14427 33949
rect 14458 33940 14464 33952
rect 14516 33940 14522 33992
rect 14553 33983 14611 33989
rect 14553 33949 14565 33983
rect 14599 33980 14611 33983
rect 14599 33952 14688 33980
rect 14599 33949 14611 33952
rect 14553 33943 14611 33949
rect 13449 33915 13507 33921
rect 13449 33912 13461 33915
rect 9692 33884 11836 33912
rect 7190 33804 7196 33856
rect 7248 33804 7254 33856
rect 8662 33804 8668 33856
rect 8720 33804 8726 33856
rect 8938 33804 8944 33856
rect 8996 33804 9002 33856
rect 9398 33804 9404 33856
rect 9456 33844 9462 33856
rect 11808 33853 11836 33884
rect 13280 33884 13461 33912
rect 13280 33856 13308 33884
rect 13449 33881 13461 33884
rect 13495 33881 13507 33915
rect 13449 33875 13507 33881
rect 9677 33847 9735 33853
rect 9677 33844 9689 33847
rect 9456 33816 9689 33844
rect 9456 33804 9462 33816
rect 9677 33813 9689 33816
rect 9723 33813 9735 33847
rect 9677 33807 9735 33813
rect 11793 33847 11851 33853
rect 11793 33813 11805 33847
rect 11839 33844 11851 33847
rect 11974 33844 11980 33856
rect 11839 33816 11980 33844
rect 11839 33813 11851 33816
rect 11793 33807 11851 33813
rect 11974 33804 11980 33816
rect 12032 33804 12038 33856
rect 13262 33804 13268 33856
rect 13320 33804 13326 33856
rect 13354 33804 13360 33856
rect 13412 33804 13418 33856
rect 13541 33847 13599 33853
rect 13541 33813 13553 33847
rect 13587 33844 13599 33847
rect 13722 33844 13728 33856
rect 13587 33816 13728 33844
rect 13587 33813 13599 33816
rect 13541 33807 13599 33813
rect 13722 33804 13728 33816
rect 13780 33804 13786 33856
rect 14476 33844 14504 33940
rect 14660 33912 14688 33952
rect 15746 33940 15752 33992
rect 15804 33980 15810 33992
rect 16025 33983 16083 33989
rect 16025 33980 16037 33983
rect 15804 33952 16037 33980
rect 15804 33940 15810 33952
rect 16025 33949 16037 33952
rect 16071 33949 16083 33983
rect 16025 33943 16083 33949
rect 16206 33940 16212 33992
rect 16264 33940 16270 33992
rect 16298 33940 16304 33992
rect 16356 33940 16362 33992
rect 16393 33983 16451 33989
rect 16393 33949 16405 33983
rect 16439 33980 16451 33983
rect 16482 33980 16488 33992
rect 16439 33952 16488 33980
rect 16439 33949 16451 33952
rect 16393 33943 16451 33949
rect 16482 33940 16488 33952
rect 16540 33940 16546 33992
rect 16777 33980 16805 34020
rect 16853 34017 16865 34051
rect 16899 34048 16911 34051
rect 17052 34048 17080 34144
rect 17405 34119 17463 34125
rect 17405 34085 17417 34119
rect 17451 34116 17463 34119
rect 19429 34119 19487 34125
rect 17451 34088 19380 34116
rect 17451 34085 17463 34088
rect 17405 34079 17463 34085
rect 19245 34051 19303 34057
rect 19245 34048 19257 34051
rect 16899 34020 17080 34048
rect 17282 34020 19257 34048
rect 16899 34017 16911 34020
rect 16853 34011 16911 34017
rect 17282 33980 17310 34020
rect 19245 34017 19257 34020
rect 19291 34017 19303 34051
rect 19352 34048 19380 34088
rect 19429 34085 19441 34119
rect 19475 34116 19487 34119
rect 19889 34119 19947 34125
rect 19889 34116 19901 34119
rect 19475 34088 19901 34116
rect 19475 34085 19487 34088
rect 19429 34079 19487 34085
rect 19889 34085 19901 34088
rect 19935 34085 19947 34119
rect 23400 34116 23428 34156
rect 19889 34079 19947 34085
rect 19996 34088 23428 34116
rect 19996 34048 20024 34088
rect 20162 34048 20168 34060
rect 19352 34020 20024 34048
rect 19245 34011 19303 34017
rect 16777 33952 17310 33980
rect 17678 33940 17684 33992
rect 17736 33940 17742 33992
rect 17770 33940 17776 33992
rect 17828 33980 17834 33992
rect 17828 33952 17873 33980
rect 17828 33940 17834 33952
rect 18046 33940 18052 33992
rect 18104 33940 18110 33992
rect 18138 33940 18144 33992
rect 18196 33989 18202 33992
rect 18196 33943 18204 33989
rect 18196 33940 18202 33943
rect 18414 33940 18420 33992
rect 18472 33940 18478 33992
rect 18785 33983 18843 33989
rect 18785 33980 18797 33983
rect 18524 33952 18797 33980
rect 15381 33915 15439 33921
rect 15381 33912 15393 33915
rect 14660 33884 15393 33912
rect 15381 33881 15393 33884
rect 15427 33912 15439 33915
rect 15470 33912 15476 33924
rect 15427 33884 15476 33912
rect 15427 33881 15439 33884
rect 15381 33875 15439 33881
rect 15470 33872 15476 33884
rect 15528 33872 15534 33924
rect 15565 33915 15623 33921
rect 15565 33881 15577 33915
rect 15611 33912 15623 33915
rect 16666 33912 16672 33924
rect 15611 33884 16672 33912
rect 15611 33881 15623 33884
rect 15565 33875 15623 33881
rect 16666 33872 16672 33884
rect 16724 33912 16730 33924
rect 17221 33915 17279 33921
rect 17221 33912 17233 33915
rect 16724 33884 17233 33912
rect 16724 33872 16730 33884
rect 17221 33881 17233 33884
rect 17267 33881 17279 33915
rect 17221 33875 17279 33881
rect 17954 33872 17960 33924
rect 18012 33872 18018 33924
rect 18524 33912 18552 33952
rect 18785 33949 18797 33952
rect 18831 33949 18843 33983
rect 19521 33983 19579 33989
rect 19521 33980 19533 33983
rect 18785 33943 18843 33949
rect 18984 33952 19533 33980
rect 18248 33884 18552 33912
rect 14918 33844 14924 33856
rect 14476 33816 14924 33844
rect 14918 33804 14924 33816
rect 14976 33804 14982 33856
rect 15657 33847 15715 33853
rect 15657 33813 15669 33847
rect 15703 33844 15715 33847
rect 16942 33844 16948 33856
rect 15703 33816 16948 33844
rect 15703 33813 15715 33816
rect 15657 33807 15715 33813
rect 16942 33804 16948 33816
rect 17000 33804 17006 33856
rect 17034 33804 17040 33856
rect 17092 33804 17098 33856
rect 17126 33804 17132 33856
rect 17184 33804 17190 33856
rect 17494 33804 17500 33856
rect 17552 33844 17558 33856
rect 18248 33844 18276 33884
rect 18598 33872 18604 33924
rect 18656 33872 18662 33924
rect 18693 33915 18751 33921
rect 18693 33881 18705 33915
rect 18739 33881 18751 33915
rect 18693 33875 18751 33881
rect 17552 33816 18276 33844
rect 17552 33804 17558 33816
rect 18322 33804 18328 33856
rect 18380 33804 18386 33856
rect 18506 33804 18512 33856
rect 18564 33844 18570 33856
rect 18708 33844 18736 33875
rect 18782 33844 18788 33856
rect 18564 33816 18788 33844
rect 18564 33804 18570 33816
rect 18782 33804 18788 33816
rect 18840 33804 18846 33856
rect 18984 33853 19012 33952
rect 19521 33949 19533 33952
rect 19567 33949 19579 33983
rect 19521 33943 19579 33949
rect 19996 33912 20024 34020
rect 20088 34020 20168 34048
rect 20088 33989 20116 34020
rect 20162 34008 20168 34020
rect 20220 34008 20226 34060
rect 23584 34048 23612 34156
rect 23658 34144 23664 34196
rect 23716 34184 23722 34196
rect 24762 34184 24768 34196
rect 23716 34156 24768 34184
rect 23716 34144 23722 34156
rect 24762 34144 24768 34156
rect 24820 34144 24826 34196
rect 25406 34144 25412 34196
rect 25464 34184 25470 34196
rect 26786 34184 26792 34196
rect 25464 34156 26792 34184
rect 25464 34144 25470 34156
rect 26053 34119 26111 34125
rect 26053 34085 26065 34119
rect 26099 34085 26111 34119
rect 26053 34079 26111 34085
rect 26068 34048 26096 34079
rect 22572 34020 23244 34048
rect 23584 34020 25728 34048
rect 20073 33983 20131 33989
rect 20073 33949 20085 33983
rect 20119 33949 20131 33983
rect 20073 33943 20131 33949
rect 20254 33940 20260 33992
rect 20312 33940 20318 33992
rect 20441 33983 20499 33989
rect 20441 33949 20453 33983
rect 20487 33980 20499 33983
rect 20530 33980 20536 33992
rect 20487 33952 20536 33980
rect 20487 33949 20499 33952
rect 20441 33943 20499 33949
rect 20530 33940 20536 33952
rect 20588 33940 20594 33992
rect 20622 33940 20628 33992
rect 20680 33980 20686 33992
rect 20809 33983 20867 33989
rect 20809 33980 20821 33983
rect 20680 33952 20821 33980
rect 20680 33940 20686 33952
rect 20809 33949 20821 33952
rect 20855 33949 20867 33983
rect 20809 33943 20867 33949
rect 20898 33940 20904 33992
rect 20956 33980 20962 33992
rect 20956 33952 21036 33980
rect 20956 33940 20962 33952
rect 20165 33915 20223 33921
rect 20165 33912 20177 33915
rect 19996 33884 20177 33912
rect 20165 33881 20177 33884
rect 20211 33881 20223 33915
rect 21008 33912 21036 33952
rect 21910 33940 21916 33992
rect 21968 33940 21974 33992
rect 22462 33980 22468 33992
rect 22066 33952 22468 33980
rect 22066 33912 22094 33952
rect 22462 33940 22468 33952
rect 22520 33940 22526 33992
rect 22572 33989 22600 34020
rect 22557 33983 22615 33989
rect 22557 33949 22569 33983
rect 22603 33949 22615 33983
rect 22557 33943 22615 33949
rect 21008 33884 22094 33912
rect 20165 33875 20223 33881
rect 22278 33872 22284 33924
rect 22336 33912 22342 33924
rect 22572 33912 22600 33943
rect 22646 33940 22652 33992
rect 22704 33940 22710 33992
rect 22833 33983 22891 33989
rect 22833 33949 22845 33983
rect 22879 33949 22891 33983
rect 22833 33943 22891 33949
rect 22336 33884 22600 33912
rect 22848 33912 22876 33943
rect 22922 33940 22928 33992
rect 22980 33940 22986 33992
rect 23216 33989 23244 34020
rect 23201 33983 23259 33989
rect 23201 33949 23213 33983
rect 23247 33949 23259 33983
rect 23201 33943 23259 33949
rect 23294 33983 23352 33989
rect 23294 33949 23306 33983
rect 23340 33980 23352 33983
rect 23382 33980 23388 33992
rect 23340 33952 23388 33980
rect 23340 33949 23352 33952
rect 23294 33943 23352 33949
rect 23309 33912 23337 33943
rect 23382 33940 23388 33952
rect 23440 33940 23446 33992
rect 23569 33983 23627 33989
rect 23569 33949 23581 33983
rect 23615 33949 23627 33983
rect 23569 33943 23627 33949
rect 22848 33884 23337 33912
rect 22336 33872 22342 33884
rect 23474 33872 23480 33924
rect 23532 33872 23538 33924
rect 23584 33912 23612 33943
rect 23658 33940 23664 33992
rect 23716 33989 23722 33992
rect 23716 33980 23724 33989
rect 23716 33952 23761 33980
rect 23716 33943 23724 33952
rect 23716 33940 23722 33943
rect 23842 33940 23848 33992
rect 23900 33940 23906 33992
rect 25590 33980 25596 33992
rect 24596 33952 25596 33980
rect 23860 33912 23888 33940
rect 23584 33884 23888 33912
rect 24596 33856 24624 33952
rect 25590 33940 25596 33952
rect 25648 33940 25654 33992
rect 25700 33989 25728 34020
rect 25884 34020 26096 34048
rect 25884 33989 25912 34020
rect 25685 33983 25743 33989
rect 25685 33949 25697 33983
rect 25731 33949 25743 33983
rect 25685 33943 25743 33949
rect 25869 33983 25927 33989
rect 25869 33949 25881 33983
rect 25915 33949 25927 33983
rect 25869 33943 25927 33949
rect 18969 33847 19027 33853
rect 18969 33813 18981 33847
rect 19015 33813 19027 33847
rect 18969 33807 19027 33813
rect 19521 33847 19579 33853
rect 19521 33813 19533 33847
rect 19567 33844 19579 33847
rect 20346 33844 20352 33856
rect 19567 33816 20352 33844
rect 19567 33813 19579 33816
rect 19521 33807 19579 33813
rect 20346 33804 20352 33816
rect 20404 33804 20410 33856
rect 20806 33804 20812 33856
rect 20864 33844 20870 33856
rect 21821 33847 21879 33853
rect 21821 33844 21833 33847
rect 20864 33816 21833 33844
rect 20864 33804 20870 33816
rect 21821 33813 21833 33816
rect 21867 33844 21879 33847
rect 22922 33844 22928 33856
rect 21867 33816 22928 33844
rect 21867 33813 21879 33816
rect 21821 33807 21879 33813
rect 22922 33804 22928 33816
rect 22980 33804 22986 33856
rect 23109 33847 23167 33853
rect 23109 33813 23121 33847
rect 23155 33844 23167 33847
rect 23382 33844 23388 33856
rect 23155 33816 23388 33844
rect 23155 33813 23167 33816
rect 23109 33807 23167 33813
rect 23382 33804 23388 33816
rect 23440 33804 23446 33856
rect 23842 33804 23848 33856
rect 23900 33804 23906 33856
rect 24578 33804 24584 33856
rect 24636 33804 24642 33856
rect 25406 33804 25412 33856
rect 25464 33804 25470 33856
rect 25700 33844 25728 33943
rect 25958 33940 25964 33992
rect 26016 33940 26022 33992
rect 26234 33940 26240 33992
rect 26292 33940 26298 33992
rect 26436 33989 26464 34156
rect 26786 34144 26792 34156
rect 26844 34144 26850 34196
rect 28074 34144 28080 34196
rect 28132 34144 28138 34196
rect 28368 34156 31064 34184
rect 28368 34116 28396 34156
rect 26620 34088 28396 34116
rect 28445 34119 28503 34125
rect 26620 33989 26648 34088
rect 28445 34085 28457 34119
rect 28491 34085 28503 34119
rect 28445 34079 28503 34085
rect 26329 33983 26387 33989
rect 26329 33949 26341 33983
rect 26375 33949 26387 33983
rect 26329 33943 26387 33949
rect 26421 33983 26479 33989
rect 26421 33949 26433 33983
rect 26467 33949 26479 33983
rect 26605 33983 26663 33989
rect 26605 33980 26617 33983
rect 26421 33943 26479 33949
rect 26528 33952 26617 33980
rect 26142 33872 26148 33924
rect 26200 33912 26206 33924
rect 26344 33912 26372 33943
rect 26528 33924 26556 33952
rect 26605 33949 26617 33952
rect 26651 33949 26663 33983
rect 26605 33943 26663 33949
rect 26970 33940 26976 33992
rect 27028 33980 27034 33992
rect 27249 33983 27307 33989
rect 27249 33980 27261 33983
rect 27028 33952 27261 33980
rect 27028 33940 27034 33952
rect 27249 33949 27261 33952
rect 27295 33949 27307 33983
rect 27249 33943 27307 33949
rect 27893 33983 27951 33989
rect 27893 33949 27905 33983
rect 27939 33980 27951 33983
rect 28460 33980 28488 34079
rect 28810 34076 28816 34128
rect 28868 34116 28874 34128
rect 30926 34116 30932 34128
rect 28868 34088 30932 34116
rect 28868 34076 28874 34088
rect 30926 34076 30932 34088
rect 30984 34076 30990 34128
rect 28626 34008 28632 34060
rect 28684 34048 28690 34060
rect 28997 34051 29055 34057
rect 28997 34048 29009 34051
rect 28684 34020 29009 34048
rect 28684 34008 28690 34020
rect 28997 34017 29009 34020
rect 29043 34017 29055 34051
rect 28997 34011 29055 34017
rect 30742 34008 30748 34060
rect 30800 34048 30806 34060
rect 30800 34020 30977 34048
rect 30800 34008 30806 34020
rect 28905 33983 28963 33989
rect 28905 33980 28917 33983
rect 27939 33952 28488 33980
rect 28863 33952 28917 33980
rect 27939 33949 27951 33952
rect 27893 33943 27951 33949
rect 28905 33949 28917 33952
rect 28951 33980 28963 33983
rect 30006 33980 30012 33992
rect 28951 33952 30012 33980
rect 28951 33949 28963 33952
rect 28905 33943 28963 33949
rect 26200 33884 26372 33912
rect 26200 33872 26206 33884
rect 26510 33872 26516 33924
rect 26568 33872 26574 33924
rect 28920 33912 28948 33943
rect 30006 33940 30012 33952
rect 30064 33940 30070 33992
rect 30466 33940 30472 33992
rect 30524 33940 30530 33992
rect 30558 33940 30564 33992
rect 30616 33989 30622 33992
rect 30949 33989 30977 34020
rect 30616 33983 30647 33989
rect 30635 33949 30647 33983
rect 30616 33943 30647 33949
rect 30934 33983 30992 33989
rect 30934 33949 30946 33983
rect 30980 33949 30992 33983
rect 30934 33943 30992 33949
rect 30616 33940 30622 33943
rect 26620 33884 28948 33912
rect 26620 33844 26648 33884
rect 29822 33872 29828 33924
rect 29880 33872 29886 33924
rect 30745 33915 30803 33921
rect 30745 33881 30757 33915
rect 30791 33881 30803 33915
rect 30745 33875 30803 33881
rect 30837 33915 30895 33921
rect 30837 33881 30849 33915
rect 30883 33912 30895 33915
rect 31036 33912 31064 34156
rect 31113 34119 31171 34125
rect 31113 34085 31125 34119
rect 31159 34116 31171 34119
rect 34057 34119 34115 34125
rect 31159 34088 31754 34116
rect 31159 34085 31171 34088
rect 31113 34079 31171 34085
rect 31726 34048 31754 34088
rect 34057 34085 34069 34119
rect 34103 34085 34115 34119
rect 34057 34079 34115 34085
rect 34072 34048 34100 34079
rect 34977 34051 35035 34057
rect 34977 34048 34989 34051
rect 31726 34020 31800 34048
rect 34072 34020 34989 34048
rect 31478 33940 31484 33992
rect 31536 33940 31542 33992
rect 31772 33989 31800 34020
rect 34977 34017 34989 34020
rect 35023 34017 35035 34051
rect 34977 34011 35035 34017
rect 31757 33983 31815 33989
rect 31757 33949 31769 33983
rect 31803 33949 31815 33983
rect 31757 33943 31815 33949
rect 33410 33940 33416 33992
rect 33468 33940 33474 33992
rect 33870 33940 33876 33992
rect 33928 33940 33934 33992
rect 34333 33983 34391 33989
rect 34333 33949 34345 33983
rect 34379 33949 34391 33983
rect 34333 33943 34391 33949
rect 34425 33983 34483 33989
rect 34425 33949 34437 33983
rect 34471 33980 34483 33983
rect 34701 33983 34759 33989
rect 34701 33980 34713 33983
rect 34471 33952 34713 33980
rect 34471 33949 34483 33952
rect 34425 33943 34483 33949
rect 34701 33949 34713 33952
rect 34747 33949 34759 33983
rect 34701 33943 34759 33949
rect 33428 33912 33456 33940
rect 30883 33884 33456 33912
rect 30883 33881 30895 33884
rect 30837 33875 30895 33881
rect 25700 33816 26648 33844
rect 27154 33804 27160 33856
rect 27212 33804 27218 33856
rect 28810 33804 28816 33856
rect 28868 33804 28874 33856
rect 29840 33844 29868 33872
rect 30760 33844 30788 33875
rect 34348 33856 34376 33943
rect 35986 33872 35992 33924
rect 36044 33872 36050 33924
rect 36630 33872 36636 33924
rect 36688 33912 36694 33924
rect 36725 33915 36783 33921
rect 36725 33912 36737 33915
rect 36688 33884 36737 33912
rect 36688 33872 36694 33884
rect 36725 33881 36737 33884
rect 36771 33881 36783 33915
rect 36725 33875 36783 33881
rect 29840 33816 30788 33844
rect 31570 33804 31576 33856
rect 31628 33804 31634 33856
rect 31941 33847 31999 33853
rect 31941 33813 31953 33847
rect 31987 33844 31999 33847
rect 32214 33844 32220 33856
rect 31987 33816 32220 33844
rect 31987 33813 31999 33816
rect 31941 33807 31999 33813
rect 32214 33804 32220 33816
rect 32272 33804 32278 33856
rect 34330 33804 34336 33856
rect 34388 33804 34394 33856
rect 1104 33754 38272 33776
rect 1104 33702 4874 33754
rect 4926 33702 4938 33754
rect 4990 33702 5002 33754
rect 5054 33702 5066 33754
rect 5118 33702 5130 33754
rect 5182 33702 35594 33754
rect 35646 33702 35658 33754
rect 35710 33702 35722 33754
rect 35774 33702 35786 33754
rect 35838 33702 35850 33754
rect 35902 33702 38272 33754
rect 1104 33680 38272 33702
rect 5445 33643 5503 33649
rect 5445 33609 5457 33643
rect 5491 33640 5503 33643
rect 5626 33640 5632 33652
rect 5491 33612 5632 33640
rect 5491 33609 5503 33612
rect 5445 33603 5503 33609
rect 5626 33600 5632 33612
rect 5684 33600 5690 33652
rect 5813 33643 5871 33649
rect 5813 33609 5825 33643
rect 5859 33640 5871 33643
rect 6730 33640 6736 33652
rect 5859 33612 6736 33640
rect 5859 33609 5871 33612
rect 5813 33603 5871 33609
rect 6730 33600 6736 33612
rect 6788 33600 6794 33652
rect 7190 33600 7196 33652
rect 7248 33600 7254 33652
rect 8662 33600 8668 33652
rect 8720 33600 8726 33652
rect 9398 33640 9404 33652
rect 9232 33612 9404 33640
rect 7208 33572 7236 33600
rect 7024 33544 7236 33572
rect 7024 33513 7052 33544
rect 8294 33532 8300 33584
rect 8352 33532 8358 33584
rect 7009 33507 7067 33513
rect 7009 33473 7021 33507
rect 7055 33473 7067 33507
rect 8680 33504 8708 33600
rect 9232 33581 9260 33612
rect 9398 33600 9404 33612
rect 9456 33600 9462 33652
rect 13170 33600 13176 33652
rect 13228 33640 13234 33652
rect 14277 33643 14335 33649
rect 14277 33640 14289 33643
rect 13228 33612 14289 33640
rect 13228 33600 13234 33612
rect 14277 33609 14289 33612
rect 14323 33609 14335 33643
rect 14277 33603 14335 33609
rect 14553 33643 14611 33649
rect 14553 33609 14565 33643
rect 14599 33640 14611 33643
rect 14642 33640 14648 33652
rect 14599 33612 14648 33640
rect 14599 33609 14611 33612
rect 14553 33603 14611 33609
rect 14642 33600 14648 33612
rect 14700 33600 14706 33652
rect 16482 33600 16488 33652
rect 16540 33640 16546 33652
rect 16540 33612 16712 33640
rect 16540 33600 16546 33612
rect 9217 33575 9275 33581
rect 9217 33541 9229 33575
rect 9263 33541 9275 33575
rect 9217 33535 9275 33541
rect 10226 33532 10232 33584
rect 10284 33532 10290 33584
rect 13354 33532 13360 33584
rect 13412 33572 13418 33584
rect 14185 33575 14243 33581
rect 14185 33572 14197 33575
rect 13412 33544 14197 33572
rect 13412 33532 13418 33544
rect 14185 33541 14197 33544
rect 14231 33541 14243 33575
rect 16574 33572 16580 33584
rect 14185 33535 14243 33541
rect 14292 33544 16580 33572
rect 8941 33507 8999 33513
rect 8941 33504 8953 33507
rect 8680 33476 8953 33504
rect 7009 33467 7067 33473
rect 8941 33473 8953 33476
rect 8987 33473 8999 33507
rect 8941 33467 8999 33473
rect 11974 33464 11980 33516
rect 12032 33504 12038 33516
rect 14001 33507 14059 33513
rect 14001 33504 14013 33507
rect 12032 33476 14013 33504
rect 12032 33464 12038 33476
rect 14001 33473 14013 33476
rect 14047 33504 14059 33507
rect 14292 33504 14320 33544
rect 16574 33532 16580 33544
rect 16632 33532 16638 33584
rect 16684 33572 16712 33612
rect 16850 33600 16856 33652
rect 16908 33640 16914 33652
rect 17034 33640 17040 33652
rect 16908 33612 17040 33640
rect 16908 33600 16914 33612
rect 17034 33600 17040 33612
rect 17092 33640 17098 33652
rect 17421 33643 17479 33649
rect 17421 33640 17433 33643
rect 17092 33612 17433 33640
rect 17092 33600 17098 33612
rect 17421 33609 17433 33612
rect 17467 33609 17479 33643
rect 17421 33603 17479 33609
rect 17589 33643 17647 33649
rect 17589 33609 17601 33643
rect 17635 33640 17647 33643
rect 17678 33640 17684 33652
rect 17635 33612 17684 33640
rect 17635 33609 17647 33612
rect 17589 33603 17647 33609
rect 17678 33600 17684 33612
rect 17736 33600 17742 33652
rect 19334 33600 19340 33652
rect 19392 33640 19398 33652
rect 19392 33612 19932 33640
rect 19392 33600 19398 33612
rect 17221 33575 17279 33581
rect 17221 33572 17233 33575
rect 16684 33544 17233 33572
rect 17221 33541 17233 33544
rect 17267 33572 17279 33575
rect 18414 33572 18420 33584
rect 17267 33544 18420 33572
rect 17267 33541 17279 33544
rect 17221 33535 17279 33541
rect 18414 33532 18420 33544
rect 18472 33532 18478 33584
rect 14047 33476 14320 33504
rect 14047 33473 14059 33476
rect 14001 33467 14059 33473
rect 14366 33464 14372 33516
rect 14424 33464 14430 33516
rect 14734 33464 14740 33516
rect 14792 33504 14798 33516
rect 18598 33504 18604 33516
rect 14792 33476 18604 33504
rect 14792 33464 14798 33476
rect 18598 33464 18604 33476
rect 18656 33464 18662 33516
rect 19702 33513 19708 33516
rect 19696 33467 19708 33513
rect 19702 33464 19708 33467
rect 19760 33464 19766 33516
rect 19904 33513 19932 33612
rect 20254 33600 20260 33652
rect 20312 33640 20318 33652
rect 21085 33643 21143 33649
rect 21085 33640 21097 33643
rect 20312 33612 21097 33640
rect 20312 33600 20318 33612
rect 21085 33609 21097 33612
rect 21131 33609 21143 33643
rect 21085 33603 21143 33609
rect 20809 33575 20867 33581
rect 20809 33572 20821 33575
rect 20272 33544 20821 33572
rect 20272 33513 20300 33544
rect 20809 33541 20821 33544
rect 20855 33541 20867 33575
rect 21100 33572 21128 33603
rect 21266 33600 21272 33652
rect 21324 33640 21330 33652
rect 21910 33640 21916 33652
rect 21324 33612 21916 33640
rect 21324 33600 21330 33612
rect 21910 33600 21916 33612
rect 21968 33600 21974 33652
rect 22094 33600 22100 33652
rect 22152 33640 22158 33652
rect 26142 33640 26148 33652
rect 22152 33612 26148 33640
rect 22152 33600 22158 33612
rect 26142 33600 26148 33612
rect 26200 33640 26206 33652
rect 31570 33640 31576 33652
rect 26200 33612 31576 33640
rect 26200 33600 26206 33612
rect 31570 33600 31576 33612
rect 31628 33600 31634 33652
rect 33226 33640 33232 33652
rect 31726 33612 33232 33640
rect 21358 33572 21364 33584
rect 21100 33544 21364 33572
rect 20809 33535 20867 33541
rect 21358 33532 21364 33544
rect 21416 33532 21422 33584
rect 21453 33575 21511 33581
rect 21453 33541 21465 33575
rect 21499 33572 21511 33575
rect 21542 33572 21548 33584
rect 21499 33544 21548 33572
rect 21499 33541 21511 33544
rect 21453 33535 21511 33541
rect 21542 33532 21548 33544
rect 21600 33532 21606 33584
rect 23198 33532 23204 33584
rect 23256 33572 23262 33584
rect 25225 33575 25283 33581
rect 23256 33544 25176 33572
rect 23256 33532 23262 33544
rect 19889 33507 19947 33513
rect 19889 33473 19901 33507
rect 19935 33473 19947 33507
rect 19889 33467 19947 33473
rect 20257 33507 20315 33513
rect 20257 33473 20269 33507
rect 20303 33473 20315 33507
rect 20257 33467 20315 33473
rect 20346 33464 20352 33516
rect 20404 33464 20410 33516
rect 20625 33507 20683 33513
rect 20625 33473 20637 33507
rect 20671 33473 20683 33507
rect 20625 33467 20683 33473
rect 5902 33396 5908 33448
rect 5960 33396 5966 33448
rect 6089 33439 6147 33445
rect 6089 33405 6101 33439
rect 6135 33436 6147 33439
rect 6135 33408 6960 33436
rect 6135 33405 6147 33408
rect 6089 33399 6147 33405
rect 6932 33300 6960 33408
rect 7282 33396 7288 33448
rect 7340 33396 7346 33448
rect 8757 33439 8815 33445
rect 8757 33405 8769 33439
rect 8803 33436 8815 33439
rect 9582 33436 9588 33448
rect 8803 33408 9588 33436
rect 8803 33405 8815 33408
rect 8757 33399 8815 33405
rect 9582 33396 9588 33408
rect 9640 33436 9646 33448
rect 18414 33436 18420 33448
rect 9640 33408 18420 33436
rect 9640 33396 9646 33408
rect 18414 33396 18420 33408
rect 18472 33396 18478 33448
rect 19058 33396 19064 33448
rect 19116 33396 19122 33448
rect 19334 33396 19340 33448
rect 19392 33436 19398 33448
rect 19610 33436 19616 33448
rect 19392 33408 19616 33436
rect 19392 33396 19398 33408
rect 19610 33396 19616 33408
rect 19668 33436 19674 33448
rect 20640 33436 20668 33467
rect 20714 33464 20720 33516
rect 20772 33464 20778 33516
rect 20901 33507 20959 33513
rect 20901 33473 20913 33507
rect 20947 33473 20959 33507
rect 20901 33467 20959 33473
rect 20916 33436 20944 33467
rect 21818 33464 21824 33516
rect 21876 33464 21882 33516
rect 22005 33507 22063 33513
rect 22005 33504 22017 33507
rect 21963 33476 22017 33504
rect 22005 33473 22017 33476
rect 22051 33504 22063 33507
rect 22051 33476 23704 33504
rect 22051 33473 22063 33476
rect 22005 33467 22063 33473
rect 22020 33436 22048 33467
rect 19668 33408 20760 33436
rect 20916 33408 22048 33436
rect 19668 33396 19674 33408
rect 17034 33328 17040 33380
rect 17092 33368 17098 33380
rect 17954 33368 17960 33380
rect 17092 33340 17960 33368
rect 17092 33328 17098 33340
rect 17954 33328 17960 33340
rect 18012 33368 18018 33380
rect 19518 33368 19524 33380
rect 18012 33340 19524 33368
rect 18012 33328 18018 33340
rect 19518 33328 19524 33340
rect 19576 33328 19582 33380
rect 19886 33328 19892 33380
rect 19944 33368 19950 33380
rect 20622 33368 20628 33380
rect 19944 33340 20628 33368
rect 19944 33328 19950 33340
rect 20622 33328 20628 33340
rect 20680 33328 20686 33380
rect 20732 33368 20760 33408
rect 23474 33396 23480 33448
rect 23532 33396 23538 33448
rect 23566 33396 23572 33448
rect 23624 33396 23630 33448
rect 23676 33436 23704 33476
rect 23750 33464 23756 33516
rect 23808 33464 23814 33516
rect 23842 33464 23848 33516
rect 23900 33464 23906 33516
rect 25148 33504 25176 33544
rect 25225 33541 25237 33575
rect 25271 33572 25283 33575
rect 25314 33572 25320 33584
rect 25271 33544 25320 33572
rect 25271 33541 25283 33544
rect 25225 33535 25283 33541
rect 25314 33532 25320 33544
rect 25372 33572 25378 33584
rect 25498 33572 25504 33584
rect 25372 33544 25504 33572
rect 25372 33532 25378 33544
rect 25498 33532 25504 33544
rect 25556 33532 25562 33584
rect 27154 33572 27160 33584
rect 26988 33544 27160 33572
rect 26510 33504 26516 33516
rect 25148 33476 26516 33504
rect 26510 33464 26516 33476
rect 26568 33464 26574 33516
rect 26602 33464 26608 33516
rect 26660 33464 26666 33516
rect 26988 33513 27016 33544
rect 27154 33532 27160 33544
rect 27212 33532 27218 33584
rect 28534 33572 28540 33584
rect 28474 33544 28540 33572
rect 28534 33532 28540 33544
rect 28592 33572 28598 33584
rect 28994 33572 29000 33584
rect 28592 33544 29000 33572
rect 28592 33532 28598 33544
rect 28994 33532 29000 33544
rect 29052 33532 29058 33584
rect 26973 33507 27031 33513
rect 26973 33473 26985 33507
rect 27019 33473 27031 33507
rect 26973 33467 27031 33473
rect 27249 33439 27307 33445
rect 27249 33436 27261 33439
rect 23676 33408 25544 33436
rect 20898 33368 20904 33380
rect 20732 33340 20904 33368
rect 20898 33328 20904 33340
rect 20956 33328 20962 33380
rect 21821 33371 21879 33377
rect 21821 33368 21833 33371
rect 21192 33340 21833 33368
rect 7006 33300 7012 33312
rect 6932 33272 7012 33300
rect 7006 33260 7012 33272
rect 7064 33300 7070 33312
rect 7834 33300 7840 33312
rect 7064 33272 7840 33300
rect 7064 33260 7070 33272
rect 7834 33260 7840 33272
rect 7892 33260 7898 33312
rect 10689 33303 10747 33309
rect 10689 33269 10701 33303
rect 10735 33300 10747 33303
rect 11606 33300 11612 33312
rect 10735 33272 11612 33300
rect 10735 33269 10747 33272
rect 10689 33263 10747 33269
rect 11606 33260 11612 33272
rect 11664 33260 11670 33312
rect 16206 33260 16212 33312
rect 16264 33300 16270 33312
rect 17405 33303 17463 33309
rect 17405 33300 17417 33303
rect 16264 33272 17417 33300
rect 16264 33260 16270 33272
rect 17405 33269 17417 33272
rect 17451 33269 17463 33303
rect 17405 33263 17463 33269
rect 18138 33260 18144 33312
rect 18196 33300 18202 33312
rect 20346 33300 20352 33312
rect 18196 33272 20352 33300
rect 18196 33260 18202 33272
rect 20346 33260 20352 33272
rect 20404 33260 20410 33312
rect 20438 33260 20444 33312
rect 20496 33300 20502 33312
rect 21192 33300 21220 33340
rect 21821 33337 21833 33340
rect 21867 33368 21879 33371
rect 24857 33371 24915 33377
rect 24857 33368 24869 33371
rect 21867 33340 24869 33368
rect 21867 33337 21879 33340
rect 21821 33331 21879 33337
rect 24857 33337 24869 33340
rect 24903 33337 24915 33371
rect 25314 33368 25320 33380
rect 24857 33331 24915 33337
rect 25240 33340 25320 33368
rect 20496 33272 21220 33300
rect 21269 33303 21327 33309
rect 20496 33260 20502 33272
rect 21269 33269 21281 33303
rect 21315 33300 21327 33303
rect 21450 33300 21456 33312
rect 21315 33272 21456 33300
rect 21315 33269 21327 33272
rect 21269 33263 21327 33269
rect 21450 33260 21456 33272
rect 21508 33260 21514 33312
rect 22922 33260 22928 33312
rect 22980 33300 22986 33312
rect 23750 33300 23756 33312
rect 22980 33272 23756 33300
rect 22980 33260 22986 33272
rect 23750 33260 23756 33272
rect 23808 33260 23814 33312
rect 24026 33260 24032 33312
rect 24084 33260 24090 33312
rect 25240 33309 25268 33340
rect 25314 33328 25320 33340
rect 25372 33328 25378 33380
rect 25225 33303 25283 33309
rect 25225 33269 25237 33303
rect 25271 33269 25283 33303
rect 25225 33263 25283 33269
rect 25406 33260 25412 33312
rect 25464 33260 25470 33312
rect 25516 33300 25544 33408
rect 26804 33408 27261 33436
rect 26804 33377 26832 33408
rect 27249 33405 27261 33408
rect 27295 33405 27307 33439
rect 27249 33399 27307 33405
rect 27798 33396 27804 33448
rect 27856 33436 27862 33448
rect 28997 33439 29055 33445
rect 28997 33436 29009 33439
rect 27856 33408 29009 33436
rect 27856 33396 27862 33408
rect 28997 33405 29009 33408
rect 29043 33405 29055 33439
rect 28997 33399 29055 33405
rect 26789 33371 26847 33377
rect 26789 33337 26801 33371
rect 26835 33337 26847 33371
rect 31726 33368 31754 33612
rect 33226 33600 33232 33612
rect 33284 33600 33290 33652
rect 33321 33643 33379 33649
rect 33321 33609 33333 33643
rect 33367 33640 33379 33643
rect 33594 33640 33600 33652
rect 33367 33612 33600 33640
rect 33367 33609 33379 33612
rect 33321 33603 33379 33609
rect 33594 33600 33600 33612
rect 33652 33600 33658 33652
rect 33781 33643 33839 33649
rect 33781 33609 33793 33643
rect 33827 33640 33839 33643
rect 33870 33640 33876 33652
rect 33827 33612 33876 33640
rect 33827 33609 33839 33612
rect 33781 33603 33839 33609
rect 33870 33600 33876 33612
rect 33928 33600 33934 33652
rect 34146 33600 34152 33652
rect 34204 33600 34210 33652
rect 34609 33643 34667 33649
rect 34609 33609 34621 33643
rect 34655 33609 34667 33643
rect 34609 33603 34667 33609
rect 33244 33572 33272 33600
rect 34241 33575 34299 33581
rect 34241 33572 34253 33575
rect 33244 33544 34253 33572
rect 34241 33541 34253 33544
rect 34287 33541 34299 33575
rect 34241 33535 34299 33541
rect 32306 33464 32312 33516
rect 32364 33504 32370 33516
rect 33413 33507 33471 33513
rect 33413 33504 33425 33507
rect 32364 33476 33425 33504
rect 32364 33464 32370 33476
rect 33413 33473 33425 33476
rect 33459 33504 33471 33507
rect 34624 33504 34652 33603
rect 36906 33600 36912 33652
rect 36964 33600 36970 33652
rect 34701 33507 34759 33513
rect 34701 33504 34713 33507
rect 33459 33476 34192 33504
rect 34624 33476 34713 33504
rect 33459 33473 33471 33476
rect 33413 33467 33471 33473
rect 33229 33439 33287 33445
rect 33229 33405 33241 33439
rect 33275 33405 33287 33439
rect 33229 33399 33287 33405
rect 26789 33331 26847 33337
rect 28276 33340 31754 33368
rect 33244 33368 33272 33399
rect 34054 33396 34060 33448
rect 34112 33396 34118 33448
rect 34164 33436 34192 33476
rect 34701 33473 34713 33476
rect 34747 33473 34759 33507
rect 34701 33467 34759 33473
rect 36630 33464 36636 33516
rect 36688 33464 36694 33516
rect 36722 33464 36728 33516
rect 36780 33464 36786 33516
rect 36648 33436 36676 33464
rect 34164 33408 36676 33436
rect 34072 33368 34100 33396
rect 35986 33368 35992 33380
rect 33244 33340 34100 33368
rect 34164 33340 35992 33368
rect 28276 33300 28304 33340
rect 25516 33272 28304 33300
rect 28534 33260 28540 33312
rect 28592 33300 28598 33312
rect 28718 33300 28724 33312
rect 28592 33272 28724 33300
rect 28592 33260 28598 33272
rect 28718 33260 28724 33272
rect 28776 33260 28782 33312
rect 30190 33260 30196 33312
rect 30248 33300 30254 33312
rect 34164 33300 34192 33340
rect 35986 33328 35992 33340
rect 36044 33328 36050 33380
rect 30248 33272 34192 33300
rect 30248 33260 30254 33272
rect 34790 33260 34796 33312
rect 34848 33300 34854 33312
rect 34885 33303 34943 33309
rect 34885 33300 34897 33303
rect 34848 33272 34897 33300
rect 34848 33260 34854 33272
rect 34885 33269 34897 33272
rect 34931 33269 34943 33303
rect 34885 33263 34943 33269
rect 1104 33210 38272 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 38272 33210
rect 1104 33136 38272 33158
rect 7282 33056 7288 33108
rect 7340 33096 7346 33108
rect 7653 33099 7711 33105
rect 7653 33096 7665 33099
rect 7340 33068 7665 33096
rect 7340 33056 7346 33068
rect 7653 33065 7665 33068
rect 7699 33065 7711 33099
rect 8938 33096 8944 33108
rect 7653 33059 7711 33065
rect 7944 33068 8944 33096
rect 4614 32960 4620 32972
rect 4080 32932 4620 32960
rect 4080 32901 4108 32932
rect 4614 32920 4620 32932
rect 4672 32920 4678 32972
rect 6089 32963 6147 32969
rect 6089 32929 6101 32963
rect 6135 32960 6147 32963
rect 6730 32960 6736 32972
rect 6135 32932 6736 32960
rect 6135 32929 6147 32932
rect 6089 32923 6147 32929
rect 6730 32920 6736 32932
rect 6788 32920 6794 32972
rect 6822 32920 6828 32972
rect 6880 32920 6886 32972
rect 4065 32895 4123 32901
rect 4065 32861 4077 32895
rect 4111 32861 4123 32895
rect 4065 32855 4123 32861
rect 4157 32895 4215 32901
rect 4157 32861 4169 32895
rect 4203 32892 4215 32895
rect 4341 32895 4399 32901
rect 4341 32892 4353 32895
rect 4203 32864 4353 32892
rect 4203 32861 4215 32864
rect 4157 32855 4215 32861
rect 4341 32861 4353 32864
rect 4387 32861 4399 32895
rect 4341 32855 4399 32861
rect 5902 32852 5908 32904
rect 5960 32892 5966 32904
rect 6638 32892 6644 32904
rect 5960 32864 6644 32892
rect 5960 32852 5966 32864
rect 6638 32852 6644 32864
rect 6696 32852 6702 32904
rect 7944 32901 7972 33068
rect 8938 33056 8944 33068
rect 8996 33056 9002 33108
rect 9858 33056 9864 33108
rect 9916 33096 9922 33108
rect 10137 33099 10195 33105
rect 10137 33096 10149 33099
rect 9916 33068 10149 33096
rect 9916 33056 9922 33068
rect 10137 33065 10149 33068
rect 10183 33065 10195 33099
rect 10137 33059 10195 33065
rect 11606 33056 11612 33108
rect 11664 33096 11670 33108
rect 11664 33068 14228 33096
rect 11664 33056 11670 33068
rect 8113 32963 8171 32969
rect 8113 32929 8125 32963
rect 8159 32960 8171 32963
rect 8389 32963 8447 32969
rect 8389 32960 8401 32963
rect 8159 32932 8401 32960
rect 8159 32929 8171 32932
rect 8113 32923 8171 32929
rect 8389 32929 8401 32932
rect 8435 32929 8447 32963
rect 8389 32923 8447 32929
rect 9585 32963 9643 32969
rect 9585 32929 9597 32963
rect 9631 32960 9643 32963
rect 9674 32960 9680 32972
rect 9631 32932 9680 32960
rect 9631 32929 9643 32932
rect 9585 32923 9643 32929
rect 9674 32920 9680 32932
rect 9732 32920 9738 32972
rect 11624 32960 11652 33056
rect 11698 32988 11704 33040
rect 11756 33028 11762 33040
rect 12158 33028 12164 33040
rect 11756 33000 12164 33028
rect 11756 32988 11762 33000
rect 12158 32988 12164 33000
rect 12216 32988 12222 33040
rect 9784 32932 11837 32960
rect 7837 32895 7895 32901
rect 7837 32861 7849 32895
rect 7883 32861 7895 32895
rect 7837 32855 7895 32861
rect 7929 32895 7987 32901
rect 7929 32861 7941 32895
rect 7975 32861 7987 32895
rect 7929 32855 7987 32861
rect 4617 32827 4675 32833
rect 4617 32793 4629 32827
rect 4663 32824 4675 32827
rect 4706 32824 4712 32836
rect 4663 32796 4712 32824
rect 4663 32793 4675 32796
rect 4617 32787 4675 32793
rect 4706 32784 4712 32796
rect 4764 32784 4770 32836
rect 6362 32824 6368 32836
rect 5842 32796 6368 32824
rect 6362 32784 6368 32796
rect 6420 32784 6426 32836
rect 7852 32824 7880 32855
rect 8202 32852 8208 32904
rect 8260 32852 8266 32904
rect 8478 32852 8484 32904
rect 8536 32852 8542 32904
rect 9784 32901 9812 32932
rect 9769 32895 9827 32901
rect 9769 32861 9781 32895
rect 9815 32861 9827 32895
rect 9769 32855 9827 32861
rect 11422 32852 11428 32904
rect 11480 32892 11486 32904
rect 11809 32901 11837 32932
rect 11701 32895 11759 32901
rect 11701 32892 11713 32895
rect 11480 32864 11713 32892
rect 11480 32852 11486 32864
rect 11701 32861 11713 32864
rect 11747 32861 11759 32895
rect 11701 32855 11759 32861
rect 11794 32895 11852 32901
rect 11794 32861 11806 32895
rect 11840 32861 11852 32895
rect 11794 32855 11852 32861
rect 11882 32852 11888 32904
rect 11940 32892 11946 32904
rect 12176 32901 12204 32988
rect 11977 32895 12035 32901
rect 11977 32892 11989 32895
rect 11940 32864 11989 32892
rect 11940 32852 11946 32864
rect 11977 32861 11989 32864
rect 12023 32861 12035 32895
rect 11977 32855 12035 32861
rect 12166 32895 12224 32901
rect 12166 32861 12178 32895
rect 12212 32861 12224 32895
rect 12166 32855 12224 32861
rect 8386 32824 8392 32836
rect 7852 32796 8392 32824
rect 8386 32784 8392 32796
rect 8444 32784 8450 32836
rect 8570 32784 8576 32836
rect 8628 32824 8634 32836
rect 10962 32824 10968 32836
rect 8628 32796 10968 32824
rect 8628 32784 8634 32796
rect 10962 32784 10968 32796
rect 11020 32784 11026 32836
rect 12066 32784 12072 32836
rect 12124 32784 12130 32836
rect 6270 32716 6276 32768
rect 6328 32716 6334 32768
rect 8846 32716 8852 32768
rect 8904 32756 8910 32768
rect 9677 32759 9735 32765
rect 9677 32756 9689 32759
rect 8904 32728 9689 32756
rect 8904 32716 8910 32728
rect 9677 32725 9689 32728
rect 9723 32725 9735 32759
rect 9677 32719 9735 32725
rect 11606 32716 11612 32768
rect 11664 32756 11670 32768
rect 12250 32756 12256 32768
rect 11664 32728 12256 32756
rect 11664 32716 11670 32728
rect 12250 32716 12256 32728
rect 12308 32716 12314 32768
rect 12342 32716 12348 32768
rect 12400 32716 12406 32768
rect 14200 32756 14228 33068
rect 17402 33056 17408 33108
rect 17460 33096 17466 33108
rect 17460 33068 18276 33096
rect 17460 33056 17466 33068
rect 16758 32988 16764 33040
rect 16816 33028 16822 33040
rect 17678 33028 17684 33040
rect 16816 33000 17684 33028
rect 16816 32988 16822 33000
rect 16960 32969 16988 33000
rect 17678 32988 17684 33000
rect 17736 33028 17742 33040
rect 18138 33028 18144 33040
rect 17736 33000 18144 33028
rect 17736 32988 17742 33000
rect 18138 32988 18144 33000
rect 18196 32988 18202 33040
rect 16945 32963 17003 32969
rect 16945 32929 16957 32963
rect 16991 32929 17003 32963
rect 18248 32960 18276 33068
rect 18322 33056 18328 33108
rect 18380 33096 18386 33108
rect 18601 33099 18659 33105
rect 18601 33096 18613 33099
rect 18380 33068 18613 33096
rect 18380 33056 18386 33068
rect 18601 33065 18613 33068
rect 18647 33065 18659 33099
rect 18601 33059 18659 33065
rect 20346 33056 20352 33108
rect 20404 33096 20410 33108
rect 20404 33068 20668 33096
rect 20404 33056 20410 33068
rect 18432 33000 19472 33028
rect 18248 32932 18368 32960
rect 16945 32923 17003 32929
rect 15838 32852 15844 32904
rect 15896 32892 15902 32904
rect 16206 32892 16212 32904
rect 15896 32864 16212 32892
rect 15896 32852 15902 32864
rect 16206 32852 16212 32864
rect 16264 32852 16270 32904
rect 17313 32895 17371 32901
rect 17313 32861 17325 32895
rect 17359 32892 17371 32895
rect 17954 32892 17960 32904
rect 17359 32864 17960 32892
rect 17359 32861 17371 32864
rect 17313 32855 17371 32861
rect 17954 32852 17960 32864
rect 18012 32852 18018 32904
rect 18340 32901 18368 32932
rect 18432 32904 18460 33000
rect 18598 32920 18604 32972
rect 18656 32960 18662 32972
rect 19334 32960 19340 32972
rect 18656 32932 19340 32960
rect 18656 32920 18662 32932
rect 19334 32920 19340 32932
rect 19392 32920 19398 32972
rect 18325 32895 18383 32901
rect 18325 32861 18337 32895
rect 18371 32861 18383 32895
rect 18325 32855 18383 32861
rect 18414 32852 18420 32904
rect 18472 32852 18478 32904
rect 18693 32895 18751 32901
rect 18693 32861 18705 32895
rect 18739 32892 18751 32895
rect 18874 32892 18880 32904
rect 18739 32864 18880 32892
rect 18739 32861 18751 32864
rect 18693 32855 18751 32861
rect 18874 32852 18880 32864
rect 18932 32852 18938 32904
rect 19444 32902 19472 33000
rect 19702 32988 19708 33040
rect 19760 32988 19766 33040
rect 19797 33031 19855 33037
rect 19797 32997 19809 33031
rect 19843 33028 19855 33031
rect 20530 33028 20536 33040
rect 19843 33000 20536 33028
rect 19843 32997 19855 33000
rect 19797 32991 19855 32997
rect 20530 32988 20536 33000
rect 20588 32988 20594 33040
rect 19610 32920 19616 32972
rect 19668 32920 19674 32972
rect 20640 32960 20668 33068
rect 20898 33056 20904 33108
rect 20956 33096 20962 33108
rect 23474 33096 23480 33108
rect 20956 33068 23480 33096
rect 20956 33056 20962 33068
rect 23474 33056 23480 33068
rect 23532 33056 23538 33108
rect 26602 33056 26608 33108
rect 26660 33056 26666 33108
rect 30006 33056 30012 33108
rect 30064 33096 30070 33108
rect 30466 33096 30472 33108
rect 30064 33068 30472 33096
rect 30064 33056 30070 33068
rect 30466 33056 30472 33068
rect 30524 33056 30530 33108
rect 31846 33096 31852 33108
rect 30668 33068 31852 33096
rect 30668 33040 30696 33068
rect 31846 33056 31852 33068
rect 31904 33056 31910 33108
rect 34790 33056 34796 33108
rect 34848 33056 34854 33108
rect 20714 32988 20720 33040
rect 20772 32988 20778 33040
rect 30650 32988 30656 33040
rect 30708 32988 30714 33040
rect 24578 32960 24584 32972
rect 19996 32932 20484 32960
rect 19996 32904 20024 32932
rect 19444 32892 19564 32902
rect 19889 32895 19947 32901
rect 19889 32892 19901 32895
rect 19444 32874 19901 32892
rect 19536 32864 19901 32874
rect 19889 32861 19901 32864
rect 19935 32861 19947 32895
rect 19889 32855 19947 32861
rect 19978 32852 19984 32904
rect 20036 32852 20042 32904
rect 20162 32852 20168 32904
rect 20220 32852 20226 32904
rect 20456 32901 20484 32932
rect 20640 32932 24584 32960
rect 20441 32895 20499 32901
rect 20441 32861 20453 32895
rect 20487 32861 20499 32895
rect 20441 32855 20499 32861
rect 20533 32895 20591 32901
rect 20533 32861 20545 32895
rect 20579 32892 20591 32895
rect 20640 32892 20668 32932
rect 24578 32920 24584 32932
rect 24636 32960 24642 32972
rect 26050 32960 26056 32972
rect 24636 32932 26056 32960
rect 24636 32920 24642 32932
rect 26050 32920 26056 32932
rect 26108 32920 26114 32972
rect 27246 32920 27252 32972
rect 27304 32920 27310 32972
rect 27798 32960 27804 32972
rect 27448 32932 27804 32960
rect 20579 32864 20668 32892
rect 20579 32861 20591 32864
rect 20533 32855 20591 32861
rect 21450 32852 21456 32904
rect 21508 32852 21514 32904
rect 21910 32852 21916 32904
rect 21968 32892 21974 32904
rect 22097 32895 22155 32901
rect 22097 32892 22109 32895
rect 21968 32864 22109 32892
rect 21968 32852 21974 32864
rect 22097 32861 22109 32864
rect 22143 32892 22155 32895
rect 22186 32892 22192 32904
rect 22143 32864 22192 32892
rect 22143 32861 22155 32864
rect 22097 32855 22155 32861
rect 22186 32852 22192 32864
rect 22244 32852 22250 32904
rect 23382 32852 23388 32904
rect 23440 32852 23446 32904
rect 24486 32852 24492 32904
rect 24544 32852 24550 32904
rect 27448 32892 27476 32932
rect 27798 32920 27804 32932
rect 27856 32920 27862 32972
rect 34808 32960 34836 33056
rect 34977 32963 35035 32969
rect 34977 32960 34989 32963
rect 30392 32932 33548 32960
rect 34808 32932 34989 32960
rect 26988 32864 27476 32892
rect 16850 32784 16856 32836
rect 16908 32824 16914 32836
rect 17586 32824 17592 32836
rect 16908 32796 17592 32824
rect 16908 32784 16914 32796
rect 17586 32784 17592 32796
rect 17644 32784 17650 32836
rect 18782 32784 18788 32836
rect 18840 32784 18846 32836
rect 19334 32824 19340 32836
rect 19306 32784 19340 32824
rect 19392 32784 19398 32836
rect 19518 32784 19524 32836
rect 19576 32824 19582 32836
rect 20349 32827 20407 32833
rect 20349 32824 20361 32827
rect 19576 32796 20361 32824
rect 19576 32784 19582 32796
rect 20349 32793 20361 32796
rect 20395 32793 20407 32827
rect 20349 32787 20407 32793
rect 19306 32756 19334 32784
rect 19978 32756 19984 32768
rect 14200 32728 19984 32756
rect 19978 32716 19984 32728
rect 20036 32716 20042 32768
rect 20364 32756 20392 32787
rect 21542 32784 21548 32836
rect 21600 32824 21606 32836
rect 23201 32827 23259 32833
rect 23201 32824 23213 32827
rect 21600 32796 23213 32824
rect 21600 32784 21606 32796
rect 23201 32793 23213 32796
rect 23247 32824 23259 32827
rect 24504 32824 24532 32852
rect 23247 32796 24532 32824
rect 23247 32793 23259 32796
rect 23201 32787 23259 32793
rect 20993 32759 21051 32765
rect 20993 32756 21005 32759
rect 20364 32728 21005 32756
rect 20993 32725 21005 32728
rect 21039 32756 21051 32759
rect 22002 32756 22008 32768
rect 21039 32728 22008 32756
rect 21039 32725 21051 32728
rect 20993 32719 21051 32725
rect 22002 32716 22008 32728
rect 22060 32716 22066 32768
rect 23566 32716 23572 32768
rect 23624 32716 23630 32768
rect 23750 32716 23756 32768
rect 23808 32756 23814 32768
rect 25038 32756 25044 32768
rect 23808 32728 25044 32756
rect 23808 32716 23814 32728
rect 25038 32716 25044 32728
rect 25096 32756 25102 32768
rect 25958 32756 25964 32768
rect 25096 32728 25964 32756
rect 25096 32716 25102 32728
rect 25958 32716 25964 32728
rect 26016 32716 26022 32768
rect 26326 32716 26332 32768
rect 26384 32756 26390 32768
rect 26694 32756 26700 32768
rect 26384 32728 26700 32756
rect 26384 32716 26390 32728
rect 26694 32716 26700 32728
rect 26752 32756 26758 32768
rect 26988 32765 27016 32864
rect 27522 32852 27528 32904
rect 27580 32852 27586 32904
rect 30392 32901 30420 32932
rect 30377 32895 30435 32901
rect 30377 32892 30389 32895
rect 30300 32864 30389 32892
rect 27801 32827 27859 32833
rect 27801 32793 27813 32827
rect 27847 32824 27859 32827
rect 28074 32824 28080 32836
rect 27847 32796 28080 32824
rect 27847 32793 27859 32796
rect 27801 32787 27859 32793
rect 28074 32784 28080 32796
rect 28132 32784 28138 32836
rect 28534 32784 28540 32836
rect 28592 32784 28598 32836
rect 30300 32768 30328 32864
rect 30377 32861 30389 32864
rect 30423 32861 30435 32895
rect 30377 32855 30435 32861
rect 30926 32852 30932 32904
rect 30984 32852 30990 32904
rect 31202 32852 31208 32904
rect 31260 32852 31266 32904
rect 32490 32852 32496 32904
rect 32548 32892 32554 32904
rect 32950 32892 32956 32904
rect 32548 32864 32956 32892
rect 32548 32852 32554 32864
rect 32950 32852 32956 32864
rect 33008 32852 33014 32904
rect 33520 32892 33548 32932
rect 34977 32929 34989 32932
rect 35023 32929 35035 32963
rect 34977 32923 35035 32929
rect 34330 32892 34336 32904
rect 33520 32864 34336 32892
rect 34330 32852 34336 32864
rect 34388 32852 34394 32904
rect 34425 32895 34483 32901
rect 34425 32861 34437 32895
rect 34471 32892 34483 32895
rect 34701 32895 34759 32901
rect 34701 32892 34713 32895
rect 34471 32864 34713 32892
rect 34471 32861 34483 32864
rect 34425 32855 34483 32861
rect 34701 32861 34713 32864
rect 34747 32861 34759 32895
rect 34701 32855 34759 32861
rect 35986 32852 35992 32904
rect 36044 32892 36050 32904
rect 36044 32864 36110 32892
rect 36044 32852 36050 32864
rect 31481 32827 31539 32833
rect 31481 32793 31493 32827
rect 31527 32793 31539 32827
rect 36725 32827 36783 32833
rect 36725 32824 36737 32827
rect 31481 32787 31539 32793
rect 36280 32796 36737 32824
rect 26973 32759 27031 32765
rect 26973 32756 26985 32759
rect 26752 32728 26985 32756
rect 26752 32716 26758 32728
rect 26973 32725 26985 32728
rect 27019 32725 27031 32759
rect 26973 32719 27031 32725
rect 27065 32759 27123 32765
rect 27065 32725 27077 32759
rect 27111 32756 27123 32759
rect 27338 32756 27344 32768
rect 27111 32728 27344 32756
rect 27111 32725 27123 32728
rect 27065 32719 27123 32725
rect 27338 32716 27344 32728
rect 27396 32716 27402 32768
rect 28718 32716 28724 32768
rect 28776 32756 28782 32768
rect 29273 32759 29331 32765
rect 29273 32756 29285 32759
rect 28776 32728 29285 32756
rect 28776 32716 28782 32728
rect 29273 32725 29285 32728
rect 29319 32725 29331 32759
rect 29273 32719 29331 32725
rect 30190 32716 30196 32768
rect 30248 32716 30254 32768
rect 30282 32716 30288 32768
rect 30340 32716 30346 32768
rect 31113 32759 31171 32765
rect 31113 32725 31125 32759
rect 31159 32756 31171 32759
rect 31496 32756 31524 32787
rect 36280 32768 36308 32796
rect 36725 32793 36737 32796
rect 36771 32793 36783 32827
rect 36725 32787 36783 32793
rect 31159 32728 31524 32756
rect 31159 32725 31171 32728
rect 31113 32719 31171 32725
rect 31846 32716 31852 32768
rect 31904 32756 31910 32768
rect 32953 32759 33011 32765
rect 32953 32756 32965 32759
rect 31904 32728 32965 32756
rect 31904 32716 31910 32728
rect 32953 32725 32965 32728
rect 32999 32725 33011 32759
rect 32953 32719 33011 32725
rect 36262 32716 36268 32768
rect 36320 32716 36326 32768
rect 1104 32666 38272 32688
rect 1104 32614 4874 32666
rect 4926 32614 4938 32666
rect 4990 32614 5002 32666
rect 5054 32614 5066 32666
rect 5118 32614 5130 32666
rect 5182 32614 35594 32666
rect 35646 32614 35658 32666
rect 35710 32614 35722 32666
rect 35774 32614 35786 32666
rect 35838 32614 35850 32666
rect 35902 32614 38272 32666
rect 1104 32592 38272 32614
rect 4706 32512 4712 32564
rect 4764 32552 4770 32564
rect 4985 32555 5043 32561
rect 4985 32552 4997 32555
rect 4764 32524 4997 32552
rect 4764 32512 4770 32524
rect 4985 32521 4997 32524
rect 5031 32521 5043 32555
rect 4985 32515 5043 32521
rect 6270 32512 6276 32564
rect 6328 32512 6334 32564
rect 6730 32512 6736 32564
rect 6788 32512 6794 32564
rect 11606 32512 11612 32564
rect 11664 32512 11670 32564
rect 11790 32512 11796 32564
rect 11848 32512 11854 32564
rect 12069 32555 12127 32561
rect 12069 32521 12081 32555
rect 12115 32552 12127 32555
rect 12115 32524 12296 32552
rect 12115 32521 12127 32524
rect 12069 32515 12127 32521
rect 5169 32419 5227 32425
rect 5169 32385 5181 32419
rect 5215 32416 5227 32419
rect 6288 32416 6316 32512
rect 5215 32388 6316 32416
rect 5215 32385 5227 32388
rect 5169 32379 5227 32385
rect 6748 32348 6776 32512
rect 11624 32484 11652 32512
rect 11701 32487 11759 32493
rect 11701 32484 11713 32487
rect 11624 32456 11713 32484
rect 11701 32453 11713 32456
rect 11747 32453 11759 32487
rect 11808 32484 11836 32512
rect 12268 32493 12296 32524
rect 12342 32512 12348 32564
rect 12400 32552 12406 32564
rect 17681 32555 17739 32561
rect 12400 32524 12480 32552
rect 12400 32512 12406 32524
rect 12452 32493 12480 32524
rect 16776 32524 17356 32552
rect 16776 32496 16804 32524
rect 12253 32487 12311 32493
rect 11808 32456 11928 32484
rect 11701 32447 11759 32453
rect 11517 32419 11575 32425
rect 11517 32385 11529 32419
rect 11563 32416 11575 32419
rect 11606 32416 11612 32428
rect 11563 32388 11612 32416
rect 11563 32385 11575 32388
rect 11517 32379 11575 32385
rect 11606 32376 11612 32388
rect 11664 32376 11670 32428
rect 11900 32425 11928 32456
rect 12253 32453 12265 32487
rect 12299 32453 12311 32487
rect 12253 32447 12311 32453
rect 12437 32487 12495 32493
rect 12437 32453 12449 32487
rect 12483 32453 12495 32487
rect 12437 32447 12495 32453
rect 16669 32487 16727 32493
rect 16669 32453 16681 32487
rect 16715 32484 16727 32487
rect 16758 32484 16764 32496
rect 16715 32456 16764 32484
rect 16715 32453 16727 32456
rect 16669 32447 16727 32453
rect 16758 32444 16764 32456
rect 16816 32444 16822 32496
rect 17328 32493 17356 32524
rect 17681 32521 17693 32555
rect 17727 32552 17739 32555
rect 17862 32552 17868 32564
rect 17727 32524 17868 32552
rect 17727 32521 17739 32524
rect 17681 32515 17739 32521
rect 17862 32512 17868 32524
rect 17920 32512 17926 32564
rect 18690 32512 18696 32564
rect 18748 32512 18754 32564
rect 18874 32512 18880 32564
rect 18932 32512 18938 32564
rect 19978 32512 19984 32564
rect 20036 32512 20042 32564
rect 22278 32552 22284 32564
rect 21100 32524 22284 32552
rect 16853 32487 16911 32493
rect 16853 32453 16865 32487
rect 16899 32453 16911 32487
rect 16853 32447 16911 32453
rect 17313 32487 17371 32493
rect 17313 32453 17325 32487
rect 17359 32453 17371 32487
rect 17313 32447 17371 32453
rect 17497 32487 17555 32493
rect 17497 32453 17509 32487
rect 17543 32484 17555 32487
rect 17586 32484 17592 32496
rect 17543 32456 17592 32484
rect 17543 32453 17555 32456
rect 17497 32447 17555 32453
rect 11793 32419 11851 32425
rect 11793 32385 11805 32419
rect 11839 32385 11851 32419
rect 11793 32379 11851 32385
rect 11885 32419 11943 32425
rect 11885 32385 11897 32419
rect 11931 32385 11943 32419
rect 11885 32379 11943 32385
rect 11808 32348 11836 32379
rect 15470 32376 15476 32428
rect 15528 32416 15534 32428
rect 15746 32416 15752 32428
rect 15528 32388 15752 32416
rect 15528 32376 15534 32388
rect 15746 32376 15752 32388
rect 15804 32416 15810 32428
rect 16868 32416 16896 32447
rect 17586 32444 17592 32456
rect 17644 32444 17650 32496
rect 17954 32444 17960 32496
rect 18012 32444 18018 32496
rect 18708 32484 18736 32512
rect 18892 32484 18920 32512
rect 21100 32496 21128 32524
rect 22278 32512 22284 32524
rect 22336 32512 22342 32564
rect 23382 32552 23388 32564
rect 23124 32524 23388 32552
rect 21082 32484 21088 32496
rect 18616 32456 18736 32484
rect 18800 32456 21088 32484
rect 17972 32416 18000 32444
rect 15804 32388 18000 32416
rect 15804 32376 15810 32388
rect 18414 32376 18420 32428
rect 18472 32376 18478 32428
rect 18616 32425 18644 32456
rect 18601 32419 18659 32425
rect 18601 32385 18613 32419
rect 18647 32385 18659 32419
rect 18601 32379 18659 32385
rect 18693 32419 18751 32425
rect 18693 32385 18705 32419
rect 18739 32416 18751 32419
rect 18800 32416 18828 32456
rect 21082 32444 21088 32456
rect 21140 32444 21146 32496
rect 21634 32484 21640 32496
rect 21284 32456 21640 32484
rect 18739 32388 18828 32416
rect 18739 32385 18751 32388
rect 18693 32379 18751 32385
rect 18874 32376 18880 32428
rect 18932 32376 18938 32428
rect 18969 32419 19027 32425
rect 18969 32385 18981 32419
rect 19015 32385 19027 32419
rect 18969 32379 19027 32385
rect 6748 32320 17908 32348
rect 5718 32240 5724 32292
rect 5776 32280 5782 32292
rect 8294 32280 8300 32292
rect 5776 32252 8300 32280
rect 5776 32240 5782 32252
rect 8294 32240 8300 32252
rect 8352 32240 8358 32292
rect 12618 32240 12624 32292
rect 12676 32240 12682 32292
rect 16114 32240 16120 32292
rect 16172 32280 16178 32292
rect 17037 32283 17095 32289
rect 17037 32280 17049 32283
rect 16172 32252 17049 32280
rect 16172 32240 16178 32252
rect 17037 32249 17049 32252
rect 17083 32280 17095 32283
rect 17126 32280 17132 32292
rect 17083 32252 17132 32280
rect 17083 32249 17095 32252
rect 17037 32243 17095 32249
rect 17126 32240 17132 32252
rect 17184 32240 17190 32292
rect 17880 32280 17908 32320
rect 18230 32308 18236 32360
rect 18288 32348 18294 32360
rect 18984 32348 19012 32379
rect 20438 32376 20444 32428
rect 20496 32376 20502 32428
rect 21284 32425 21312 32456
rect 21634 32444 21640 32456
rect 21692 32444 21698 32496
rect 23124 32493 23152 32524
rect 23382 32512 23388 32524
rect 23440 32512 23446 32564
rect 23566 32512 23572 32564
rect 23624 32552 23630 32564
rect 23624 32524 23796 32552
rect 23624 32512 23630 32524
rect 23109 32487 23167 32493
rect 23109 32484 23121 32487
rect 22020 32456 23121 32484
rect 21269 32419 21327 32425
rect 21269 32385 21281 32419
rect 21315 32385 21327 32419
rect 21269 32379 21327 32385
rect 21358 32376 21364 32428
rect 21416 32416 21422 32428
rect 21913 32419 21971 32425
rect 21913 32416 21925 32419
rect 21416 32388 21925 32416
rect 21416 32376 21422 32388
rect 21913 32385 21925 32388
rect 21959 32385 21971 32419
rect 21913 32379 21971 32385
rect 18288 32320 19012 32348
rect 20456 32348 20484 32376
rect 22020 32348 22048 32456
rect 23109 32453 23121 32456
rect 23155 32453 23167 32487
rect 23109 32447 23167 32453
rect 23198 32444 23204 32496
rect 23256 32444 23262 32496
rect 23768 32484 23796 32524
rect 27522 32512 27528 32564
rect 27580 32552 27586 32564
rect 27801 32555 27859 32561
rect 27801 32552 27813 32555
rect 27580 32524 27813 32552
rect 27580 32512 27586 32524
rect 27801 32521 27813 32524
rect 27847 32521 27859 32555
rect 27801 32515 27859 32521
rect 28074 32512 28080 32564
rect 28132 32552 28138 32564
rect 28997 32555 29055 32561
rect 28997 32552 29009 32555
rect 28132 32524 29009 32552
rect 28132 32512 28138 32524
rect 28997 32521 29009 32524
rect 29043 32521 29055 32555
rect 28997 32515 29055 32521
rect 31202 32512 31208 32564
rect 31260 32552 31266 32564
rect 31389 32555 31447 32561
rect 31389 32552 31401 32555
rect 31260 32524 31401 32552
rect 31260 32512 31266 32524
rect 31389 32521 31401 32524
rect 31435 32521 31447 32555
rect 31389 32515 31447 32521
rect 35989 32555 36047 32561
rect 35989 32521 36001 32555
rect 36035 32552 36047 32555
rect 36722 32552 36728 32564
rect 36035 32524 36728 32552
rect 36035 32521 36047 32524
rect 35989 32515 36047 32521
rect 36722 32512 36728 32524
rect 36780 32512 36786 32564
rect 23308 32456 23612 32484
rect 23768 32456 23934 32484
rect 22738 32376 22744 32428
rect 22796 32416 22802 32428
rect 22922 32416 22928 32428
rect 22796 32388 22928 32416
rect 22796 32376 22802 32388
rect 22922 32376 22928 32388
rect 22980 32376 22986 32428
rect 23014 32376 23020 32428
rect 23072 32376 23078 32428
rect 20456 32320 22048 32348
rect 18288 32308 18294 32320
rect 22278 32308 22284 32360
rect 22336 32348 22342 32360
rect 23308 32348 23336 32456
rect 23385 32419 23443 32425
rect 23385 32385 23397 32419
rect 23431 32416 23443 32419
rect 23431 32388 23521 32416
rect 23431 32385 23443 32388
rect 23385 32379 23443 32385
rect 22336 32320 23336 32348
rect 22336 32308 22342 32320
rect 17880 32252 19012 32280
rect 6546 32172 6552 32224
rect 6604 32212 6610 32224
rect 11606 32212 11612 32224
rect 6604 32184 11612 32212
rect 6604 32172 6610 32184
rect 11606 32172 11612 32184
rect 11664 32172 11670 32224
rect 16666 32172 16672 32224
rect 16724 32212 16730 32224
rect 16853 32215 16911 32221
rect 16853 32212 16865 32215
rect 16724 32184 16865 32212
rect 16724 32172 16730 32184
rect 16853 32181 16865 32184
rect 16899 32212 16911 32215
rect 16942 32212 16948 32224
rect 16899 32184 16948 32212
rect 16899 32181 16911 32184
rect 16853 32175 16911 32181
rect 16942 32172 16948 32184
rect 17000 32212 17006 32224
rect 17463 32215 17521 32221
rect 17463 32212 17475 32215
rect 17000 32184 17475 32212
rect 17000 32172 17006 32184
rect 17463 32181 17475 32184
rect 17509 32181 17521 32215
rect 18984 32212 19012 32252
rect 19058 32240 19064 32292
rect 19116 32280 19122 32292
rect 23198 32280 23204 32292
rect 19116 32252 23204 32280
rect 19116 32240 19122 32252
rect 23198 32240 23204 32252
rect 23256 32240 23262 32292
rect 23493 32280 23521 32388
rect 23584 32348 23612 32456
rect 23750 32376 23756 32428
rect 23808 32376 23814 32428
rect 23906 32425 23934 32456
rect 27706 32444 27712 32496
rect 27764 32484 27770 32496
rect 32582 32484 32588 32496
rect 27764 32456 32588 32484
rect 27764 32444 27770 32456
rect 23891 32419 23949 32425
rect 23891 32385 23903 32419
rect 23937 32385 23949 32419
rect 23891 32379 23949 32385
rect 24029 32419 24087 32425
rect 24029 32385 24041 32419
rect 24075 32385 24087 32419
rect 24029 32379 24087 32385
rect 24044 32348 24072 32379
rect 24118 32376 24124 32428
rect 24176 32376 24182 32428
rect 27724 32416 27752 32444
rect 27893 32419 27951 32425
rect 27893 32416 27905 32419
rect 27724 32388 27905 32416
rect 27893 32385 27905 32388
rect 27939 32385 27951 32419
rect 28537 32419 28595 32425
rect 28537 32416 28549 32419
rect 27893 32379 27951 32385
rect 28000 32388 28549 32416
rect 23584 32320 24072 32348
rect 24394 32308 24400 32360
rect 24452 32348 24458 32360
rect 26510 32348 26516 32360
rect 24452 32320 26516 32348
rect 24452 32308 24458 32320
rect 26510 32308 26516 32320
rect 26568 32348 26574 32360
rect 28000 32348 28028 32388
rect 28537 32385 28549 32388
rect 28583 32416 28595 32419
rect 28718 32416 28724 32428
rect 28583 32388 28724 32416
rect 28583 32385 28595 32388
rect 28537 32379 28595 32385
rect 28718 32376 28724 32388
rect 28776 32376 28782 32428
rect 29181 32419 29239 32425
rect 29181 32416 29193 32419
rect 28920 32388 29193 32416
rect 26568 32320 28028 32348
rect 28261 32351 28319 32357
rect 26568 32308 26574 32320
rect 28261 32317 28273 32351
rect 28307 32317 28319 32351
rect 28261 32311 28319 32317
rect 23493 32252 24992 32280
rect 24964 32224 24992 32252
rect 27890 32240 27896 32292
rect 27948 32280 27954 32292
rect 28276 32280 28304 32311
rect 28442 32308 28448 32360
rect 28500 32308 28506 32360
rect 28920 32289 28948 32388
rect 29181 32385 29193 32388
rect 29227 32385 29239 32419
rect 29181 32379 29239 32385
rect 30834 32376 30840 32428
rect 30892 32376 30898 32428
rect 30926 32376 30932 32428
rect 30984 32376 30990 32428
rect 31496 32425 31524 32456
rect 32582 32444 32588 32456
rect 32640 32484 32646 32496
rect 34606 32484 34612 32496
rect 32640 32456 34612 32484
rect 32640 32444 32646 32456
rect 34606 32444 34612 32456
rect 34664 32444 34670 32496
rect 36262 32484 36268 32496
rect 35636 32456 36268 32484
rect 31481 32419 31539 32425
rect 31481 32385 31493 32419
rect 31527 32385 31539 32419
rect 31481 32379 31539 32385
rect 32122 32376 32128 32428
rect 32180 32376 32186 32428
rect 32214 32376 32220 32428
rect 32272 32416 32278 32428
rect 32401 32419 32459 32425
rect 32401 32416 32413 32419
rect 32272 32388 32413 32416
rect 32272 32376 32278 32388
rect 32401 32385 32413 32388
rect 32447 32385 32459 32419
rect 32401 32379 32459 32385
rect 33134 32376 33140 32428
rect 33192 32376 33198 32428
rect 33226 32376 33232 32428
rect 33284 32416 33290 32428
rect 35636 32425 35664 32456
rect 36262 32444 36268 32456
rect 36320 32444 36326 32496
rect 33413 32419 33471 32425
rect 33413 32416 33425 32419
rect 33284 32388 33425 32416
rect 33284 32376 33290 32388
rect 33413 32385 33425 32388
rect 33459 32416 33471 32419
rect 35621 32419 35679 32425
rect 35621 32416 35633 32419
rect 33459 32388 35633 32416
rect 33459 32385 33471 32388
rect 33413 32379 33471 32385
rect 35621 32385 35633 32388
rect 35667 32385 35679 32419
rect 35621 32379 35679 32385
rect 35805 32419 35863 32425
rect 35805 32385 35817 32419
rect 35851 32385 35863 32419
rect 35805 32379 35863 32385
rect 30650 32308 30656 32360
rect 30708 32308 30714 32360
rect 30745 32351 30803 32357
rect 30745 32317 30757 32351
rect 30791 32317 30803 32351
rect 30745 32311 30803 32317
rect 27948 32252 28304 32280
rect 28905 32283 28963 32289
rect 27948 32240 27954 32252
rect 28905 32249 28917 32283
rect 28951 32249 28963 32283
rect 28905 32243 28963 32249
rect 20162 32212 20168 32224
rect 18984 32184 20168 32212
rect 17463 32175 17521 32181
rect 20162 32172 20168 32184
rect 20220 32212 20226 32224
rect 20898 32212 20904 32224
rect 20220 32184 20904 32212
rect 20220 32172 20226 32184
rect 20898 32172 20904 32184
rect 20956 32172 20962 32224
rect 22186 32172 22192 32224
rect 22244 32172 22250 32224
rect 22830 32172 22836 32224
rect 22888 32172 22894 32224
rect 24302 32172 24308 32224
rect 24360 32172 24366 32224
rect 24946 32172 24952 32224
rect 25004 32212 25010 32224
rect 26234 32212 26240 32224
rect 25004 32184 26240 32212
rect 25004 32172 25010 32184
rect 26234 32172 26240 32184
rect 26292 32212 26298 32224
rect 30760 32212 30788 32311
rect 30944 32280 30972 32376
rect 32140 32348 32168 32376
rect 32140 32320 32260 32348
rect 31205 32283 31263 32289
rect 31205 32280 31217 32283
rect 30944 32252 31217 32280
rect 31205 32249 31217 32252
rect 31251 32249 31263 32283
rect 31846 32280 31852 32292
rect 31205 32243 31263 32249
rect 31726 32252 31852 32280
rect 31726 32212 31754 32252
rect 31846 32240 31852 32252
rect 31904 32240 31910 32292
rect 32122 32240 32128 32292
rect 32180 32240 32186 32292
rect 32232 32280 32260 32320
rect 32306 32308 32312 32360
rect 32364 32348 32370 32360
rect 32677 32351 32735 32357
rect 32677 32348 32689 32351
rect 32364 32320 32689 32348
rect 32364 32308 32370 32320
rect 32677 32317 32689 32320
rect 32723 32317 32735 32351
rect 32677 32311 32735 32317
rect 35820 32280 35848 32379
rect 32232 32252 35848 32280
rect 26292 32184 31754 32212
rect 26292 32172 26298 32184
rect 1104 32122 38272 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 38272 32122
rect 1104 32048 38272 32070
rect 4614 32008 4620 32020
rect 4080 31980 4620 32008
rect 4080 31872 4108 31980
rect 4614 31968 4620 31980
rect 4672 32008 4678 32020
rect 7190 32008 7196 32020
rect 4672 31980 7196 32008
rect 4672 31968 4678 31980
rect 7190 31968 7196 31980
rect 7248 31968 7254 32020
rect 17402 31968 17408 32020
rect 17460 32008 17466 32020
rect 17460 31980 19012 32008
rect 17460 31968 17466 31980
rect 7466 31900 7472 31952
rect 7524 31940 7530 31952
rect 8478 31940 8484 31952
rect 7524 31912 8484 31940
rect 7524 31900 7530 31912
rect 8478 31900 8484 31912
rect 8536 31900 8542 31952
rect 18690 31900 18696 31952
rect 18748 31900 18754 31952
rect 18984 31940 19012 31980
rect 19058 31968 19064 32020
rect 19116 31968 19122 32020
rect 20806 32008 20812 32020
rect 19168 31980 20812 32008
rect 19168 31940 19196 31980
rect 20806 31968 20812 31980
rect 20864 31968 20870 32020
rect 22002 31968 22008 32020
rect 22060 32008 22066 32020
rect 22060 31980 24256 32008
rect 22060 31968 22066 31980
rect 18984 31912 19196 31940
rect 19981 31943 20039 31949
rect 19981 31909 19993 31943
rect 20027 31940 20039 31943
rect 20254 31940 20260 31952
rect 20027 31912 20260 31940
rect 20027 31909 20039 31912
rect 19981 31903 20039 31909
rect 20254 31900 20260 31912
rect 20312 31900 20318 31952
rect 20622 31900 20628 31952
rect 20680 31940 20686 31952
rect 22278 31940 22284 31952
rect 20680 31912 22284 31940
rect 20680 31900 20686 31912
rect 22278 31900 22284 31912
rect 22336 31900 22342 31952
rect 22738 31900 22744 31952
rect 22796 31940 22802 31952
rect 23014 31940 23020 31952
rect 22796 31912 23020 31940
rect 22796 31900 22802 31912
rect 23014 31900 23020 31912
rect 23072 31900 23078 31952
rect 23934 31900 23940 31952
rect 23992 31900 23998 31952
rect 24228 31940 24256 31980
rect 24302 31968 24308 32020
rect 24360 32008 24366 32020
rect 24360 31980 25360 32008
rect 24360 31968 24366 31980
rect 24394 31940 24400 31952
rect 24228 31912 24400 31940
rect 24394 31900 24400 31912
rect 24452 31900 24458 31952
rect 25332 31949 25360 31980
rect 26970 31968 26976 32020
rect 27028 32008 27034 32020
rect 30282 32008 30288 32020
rect 27028 31980 30288 32008
rect 27028 31968 27034 31980
rect 30282 31968 30288 31980
rect 30340 31968 30346 32020
rect 31846 31968 31852 32020
rect 31904 31968 31910 32020
rect 24949 31943 25007 31949
rect 24949 31909 24961 31943
rect 24995 31909 25007 31943
rect 24949 31903 25007 31909
rect 25317 31943 25375 31949
rect 25317 31909 25329 31943
rect 25363 31909 25375 31943
rect 25317 31903 25375 31909
rect 3988 31844 4108 31872
rect 7193 31875 7251 31881
rect 3988 31813 4016 31844
rect 7193 31841 7205 31875
rect 7239 31872 7251 31875
rect 7239 31844 7880 31872
rect 7239 31841 7251 31844
rect 7193 31835 7251 31841
rect 3973 31807 4031 31813
rect 3973 31773 3985 31807
rect 4019 31773 4031 31807
rect 3973 31767 4031 31773
rect 4065 31807 4123 31813
rect 4065 31773 4077 31807
rect 4111 31804 4123 31807
rect 4249 31807 4307 31813
rect 4249 31804 4261 31807
rect 4111 31776 4261 31804
rect 4111 31773 4123 31776
rect 4065 31767 4123 31773
rect 4249 31773 4261 31776
rect 4295 31773 4307 31807
rect 5810 31804 5816 31816
rect 5658 31776 5816 31804
rect 4249 31767 4307 31773
rect 5810 31764 5816 31776
rect 5868 31764 5874 31816
rect 6273 31807 6331 31813
rect 6273 31773 6285 31807
rect 6319 31804 6331 31807
rect 6546 31804 6552 31816
rect 6319 31776 6552 31804
rect 6319 31773 6331 31776
rect 6273 31767 6331 31773
rect 6546 31764 6552 31776
rect 6604 31764 6610 31816
rect 6638 31764 6644 31816
rect 6696 31804 6702 31816
rect 6696 31776 7052 31804
rect 6696 31764 6702 31776
rect 4525 31739 4583 31745
rect 4525 31705 4537 31739
rect 4571 31705 4583 31739
rect 7024 31736 7052 31776
rect 7466 31764 7472 31816
rect 7524 31764 7530 31816
rect 7561 31807 7619 31813
rect 7561 31773 7573 31807
rect 7607 31773 7619 31807
rect 7561 31767 7619 31773
rect 7576 31736 7604 31767
rect 7650 31764 7656 31816
rect 7708 31764 7714 31816
rect 7852 31813 7880 31844
rect 7944 31844 8892 31872
rect 7837 31807 7895 31813
rect 7837 31773 7849 31807
rect 7883 31773 7895 31807
rect 7837 31767 7895 31773
rect 7944 31736 7972 31844
rect 8864 31816 8892 31844
rect 11606 31832 11612 31884
rect 11664 31872 11670 31884
rect 20640 31872 20668 31900
rect 22756 31872 22784 31900
rect 23566 31872 23572 31884
rect 11664 31844 20668 31872
rect 22572 31844 22784 31872
rect 22812 31844 23572 31872
rect 11664 31832 11670 31844
rect 8110 31764 8116 31816
rect 8168 31764 8174 31816
rect 8478 31764 8484 31816
rect 8536 31764 8542 31816
rect 8846 31764 8852 31816
rect 8904 31764 8910 31816
rect 9030 31764 9036 31816
rect 9088 31804 9094 31816
rect 9217 31807 9275 31813
rect 9217 31804 9229 31807
rect 9088 31776 9229 31804
rect 9088 31764 9094 31776
rect 9217 31773 9229 31776
rect 9263 31773 9275 31807
rect 9217 31767 9275 31773
rect 9309 31807 9367 31813
rect 9309 31773 9321 31807
rect 9355 31804 9367 31807
rect 9493 31807 9551 31813
rect 9493 31804 9505 31807
rect 9355 31776 9505 31804
rect 9355 31773 9367 31776
rect 9309 31767 9367 31773
rect 9493 31773 9505 31776
rect 9539 31773 9551 31807
rect 9493 31767 9551 31773
rect 13096 31776 13584 31804
rect 7024 31708 7972 31736
rect 4525 31699 4583 31705
rect 4540 31668 4568 31699
rect 9766 31696 9772 31748
rect 9824 31696 9830 31748
rect 10226 31696 10232 31748
rect 10284 31696 10290 31748
rect 11790 31696 11796 31748
rect 11848 31736 11854 31748
rect 13096 31745 13124 31776
rect 13081 31739 13139 31745
rect 13081 31736 13093 31739
rect 11848 31708 13093 31736
rect 11848 31696 11854 31708
rect 13081 31705 13093 31708
rect 13127 31705 13139 31739
rect 13081 31699 13139 31705
rect 13170 31696 13176 31748
rect 13228 31736 13234 31748
rect 13357 31739 13415 31745
rect 13357 31736 13369 31739
rect 13228 31708 13369 31736
rect 13228 31696 13234 31708
rect 13357 31705 13369 31708
rect 13403 31705 13415 31739
rect 13556 31736 13584 31776
rect 13630 31764 13636 31816
rect 13688 31764 13694 31816
rect 17586 31764 17592 31816
rect 17644 31804 17650 31816
rect 18782 31804 18788 31816
rect 17644 31776 18788 31804
rect 17644 31764 17650 31776
rect 18782 31764 18788 31776
rect 18840 31764 18846 31816
rect 18874 31764 18880 31816
rect 18932 31764 18938 31816
rect 19061 31807 19119 31813
rect 19061 31773 19073 31807
rect 19107 31804 19119 31807
rect 21269 31807 21327 31813
rect 19107 31776 19196 31804
rect 19107 31773 19119 31776
rect 19061 31767 19119 31773
rect 19168 31748 19196 31776
rect 21269 31773 21281 31807
rect 21315 31804 21327 31807
rect 21726 31804 21732 31816
rect 21315 31776 21732 31804
rect 21315 31773 21327 31776
rect 21269 31767 21327 31773
rect 21726 31764 21732 31776
rect 21784 31764 21790 31816
rect 21910 31764 21916 31816
rect 21968 31764 21974 31816
rect 22002 31764 22008 31816
rect 22060 31764 22066 31816
rect 22094 31764 22100 31816
rect 22152 31804 22158 31816
rect 22189 31807 22247 31813
rect 22189 31804 22201 31807
rect 22152 31776 22201 31804
rect 22152 31764 22158 31776
rect 22189 31773 22201 31776
rect 22235 31773 22247 31807
rect 22189 31767 22247 31773
rect 22278 31764 22284 31816
rect 22336 31764 22342 31816
rect 22370 31764 22376 31816
rect 22428 31813 22434 31816
rect 22428 31804 22436 31813
rect 22428 31776 22473 31804
rect 22428 31767 22436 31776
rect 22428 31764 22434 31767
rect 14550 31736 14556 31748
rect 13556 31708 14556 31736
rect 13357 31699 13415 31705
rect 14550 31696 14556 31708
rect 14608 31696 14614 31748
rect 16482 31696 16488 31748
rect 16540 31736 16546 31748
rect 18138 31736 18144 31748
rect 16540 31708 18144 31736
rect 16540 31696 16546 31708
rect 18138 31696 18144 31708
rect 18196 31696 18202 31748
rect 19150 31696 19156 31748
rect 19208 31736 19214 31748
rect 21818 31736 21824 31748
rect 19208 31708 21824 31736
rect 19208 31696 19214 31708
rect 21818 31696 21824 31708
rect 21876 31696 21882 31748
rect 22572 31736 22600 31844
rect 22646 31764 22652 31816
rect 22704 31764 22710 31816
rect 22812 31813 22840 31844
rect 23198 31813 23204 31816
rect 22797 31807 22855 31813
rect 22797 31773 22809 31807
rect 22843 31773 22855 31807
rect 22797 31767 22855 31773
rect 23155 31807 23204 31813
rect 23155 31773 23167 31807
rect 23201 31773 23204 31807
rect 23155 31767 23204 31773
rect 23198 31764 23204 31767
rect 23256 31764 23262 31816
rect 23382 31764 23388 31816
rect 23440 31764 23446 31816
rect 23493 31813 23521 31844
rect 23566 31832 23572 31844
rect 23624 31832 23630 31884
rect 23952 31872 23980 31900
rect 23676 31844 23980 31872
rect 23478 31807 23536 31813
rect 23478 31773 23490 31807
rect 23524 31804 23536 31807
rect 23524 31776 23558 31804
rect 23524 31773 23536 31776
rect 23478 31767 23536 31773
rect 23676 31748 23704 31844
rect 23891 31807 23949 31813
rect 23891 31773 23903 31807
rect 23937 31804 23949 31807
rect 24210 31804 24216 31816
rect 23937 31776 24216 31804
rect 23937 31773 23949 31776
rect 23891 31767 23949 31773
rect 24210 31764 24216 31776
rect 24268 31764 24274 31816
rect 24412 31813 24440 31900
rect 24964 31872 24992 31903
rect 25406 31900 25412 31952
rect 25464 31940 25470 31952
rect 26789 31943 26847 31949
rect 26789 31940 26801 31943
rect 25464 31912 26801 31940
rect 25464 31900 25470 31912
rect 26789 31909 26801 31912
rect 26835 31909 26847 31943
rect 26789 31903 26847 31909
rect 28718 31900 28724 31952
rect 28776 31940 28782 31952
rect 28776 31912 29960 31940
rect 28776 31900 28782 31912
rect 28902 31872 28908 31884
rect 24964 31844 25452 31872
rect 24397 31807 24455 31813
rect 24397 31773 24409 31807
rect 24443 31773 24455 31807
rect 24397 31767 24455 31773
rect 24486 31764 24492 31816
rect 24544 31804 24550 31816
rect 24544 31776 24624 31804
rect 24544 31764 24550 31776
rect 22925 31739 22983 31745
rect 22925 31736 22937 31739
rect 22572 31708 22937 31736
rect 22925 31705 22937 31708
rect 22971 31705 22983 31739
rect 22925 31699 22983 31705
rect 23017 31739 23075 31745
rect 23017 31705 23029 31739
rect 23063 31705 23075 31739
rect 23017 31699 23075 31705
rect 7285 31671 7343 31677
rect 7285 31668 7297 31671
rect 4540 31640 7297 31668
rect 7285 31637 7297 31640
rect 7331 31637 7343 31671
rect 7285 31631 7343 31637
rect 7834 31628 7840 31680
rect 7892 31668 7898 31680
rect 8021 31671 8079 31677
rect 8021 31668 8033 31671
rect 7892 31640 8033 31668
rect 7892 31628 7898 31640
rect 8021 31637 8033 31640
rect 8067 31637 8079 31671
rect 8021 31631 8079 31637
rect 8294 31628 8300 31680
rect 8352 31628 8358 31680
rect 11241 31671 11299 31677
rect 11241 31637 11253 31671
rect 11287 31668 11299 31671
rect 11514 31668 11520 31680
rect 11287 31640 11520 31668
rect 11287 31637 11299 31640
rect 11241 31631 11299 31637
rect 11514 31628 11520 31640
rect 11572 31628 11578 31680
rect 12986 31628 12992 31680
rect 13044 31668 13050 31680
rect 13265 31671 13323 31677
rect 13265 31668 13277 31671
rect 13044 31640 13277 31668
rect 13044 31628 13050 31640
rect 13265 31637 13277 31640
rect 13311 31637 13323 31671
rect 13265 31631 13323 31637
rect 13449 31671 13507 31677
rect 13449 31637 13461 31671
rect 13495 31668 13507 31671
rect 13906 31668 13912 31680
rect 13495 31640 13912 31668
rect 13495 31637 13507 31640
rect 13449 31631 13507 31637
rect 13906 31628 13912 31640
rect 13964 31668 13970 31680
rect 14366 31668 14372 31680
rect 13964 31640 14372 31668
rect 13964 31628 13970 31640
rect 14366 31628 14372 31640
rect 14424 31628 14430 31680
rect 16942 31628 16948 31680
rect 17000 31668 17006 31680
rect 19610 31668 19616 31680
rect 17000 31640 19616 31668
rect 17000 31628 17006 31640
rect 19610 31628 19616 31640
rect 19668 31668 19674 31680
rect 19886 31668 19892 31680
rect 19668 31640 19892 31668
rect 19668 31628 19674 31640
rect 19886 31628 19892 31640
rect 19944 31628 19950 31680
rect 20438 31628 20444 31680
rect 20496 31668 20502 31680
rect 21358 31668 21364 31680
rect 20496 31640 21364 31668
rect 20496 31628 20502 31640
rect 21358 31628 21364 31640
rect 21416 31628 21422 31680
rect 21836 31668 21864 31696
rect 22002 31668 22008 31680
rect 21836 31640 22008 31668
rect 22002 31628 22008 31640
rect 22060 31628 22066 31680
rect 22554 31628 22560 31680
rect 22612 31628 22618 31680
rect 22646 31628 22652 31680
rect 22704 31668 22710 31680
rect 23032 31668 23060 31699
rect 23658 31696 23664 31748
rect 23716 31696 23722 31748
rect 23750 31696 23756 31748
rect 23808 31696 23814 31748
rect 24596 31745 24624 31776
rect 24762 31764 24768 31816
rect 24820 31764 24826 31816
rect 24946 31764 24952 31816
rect 25004 31764 25010 31816
rect 25130 31764 25136 31816
rect 25188 31764 25194 31816
rect 25225 31807 25283 31813
rect 25225 31773 25237 31807
rect 25271 31773 25283 31807
rect 25225 31767 25283 31773
rect 24581 31739 24639 31745
rect 24581 31705 24593 31739
rect 24627 31705 24639 31739
rect 24581 31699 24639 31705
rect 24673 31739 24731 31745
rect 24673 31705 24685 31739
rect 24719 31736 24731 31739
rect 24964 31736 24992 31764
rect 24719 31708 24992 31736
rect 24719 31705 24731 31708
rect 24673 31699 24731 31705
rect 22704 31640 23060 31668
rect 22704 31628 22710 31640
rect 23198 31628 23204 31680
rect 23256 31668 23262 31680
rect 23293 31671 23351 31677
rect 23293 31668 23305 31671
rect 23256 31640 23305 31668
rect 23256 31628 23262 31640
rect 23293 31637 23305 31640
rect 23339 31637 23351 31671
rect 23293 31631 23351 31637
rect 24029 31671 24087 31677
rect 24029 31637 24041 31671
rect 24075 31668 24087 31671
rect 25240 31668 25268 31767
rect 25314 31764 25320 31816
rect 25372 31764 25378 31816
rect 25424 31813 25452 31844
rect 28000 31844 28908 31872
rect 25409 31807 25467 31813
rect 25409 31773 25421 31807
rect 25455 31773 25467 31807
rect 25409 31767 25467 31773
rect 26142 31764 26148 31816
rect 26200 31764 26206 31816
rect 26234 31764 26240 31816
rect 26292 31764 26298 31816
rect 26510 31764 26516 31816
rect 26568 31764 26574 31816
rect 26970 31764 26976 31816
rect 27028 31764 27034 31816
rect 28000 31813 28028 31844
rect 28902 31832 28908 31844
rect 28960 31832 28966 31884
rect 29472 31844 29712 31872
rect 29472 31816 29500 31844
rect 27985 31807 28043 31813
rect 27985 31773 27997 31807
rect 28031 31773 28043 31807
rect 27985 31767 28043 31773
rect 28258 31764 28264 31816
rect 28316 31764 28322 31816
rect 29454 31764 29460 31816
rect 29512 31764 29518 31816
rect 29684 31813 29712 31844
rect 29549 31807 29607 31813
rect 29549 31773 29561 31807
rect 29595 31804 29607 31807
rect 29684 31807 29745 31813
rect 29595 31776 29629 31804
rect 29684 31776 29699 31807
rect 29595 31773 29607 31776
rect 29549 31767 29607 31773
rect 29687 31773 29699 31776
rect 29733 31773 29745 31807
rect 29687 31767 29745 31773
rect 25332 31736 25360 31764
rect 26160 31736 26188 31764
rect 25332 31708 26188 31736
rect 26329 31739 26387 31745
rect 26329 31705 26341 31739
rect 26375 31736 26387 31739
rect 26786 31736 26792 31748
rect 26375 31708 26792 31736
rect 26375 31705 26387 31708
rect 26329 31699 26387 31705
rect 24075 31640 25268 31668
rect 24075 31637 24087 31640
rect 24029 31631 24087 31637
rect 25590 31628 25596 31680
rect 25648 31628 25654 31680
rect 25961 31671 26019 31677
rect 25961 31637 25973 31671
rect 26007 31668 26019 31671
rect 26142 31668 26148 31680
rect 26007 31640 26148 31668
rect 26007 31637 26019 31640
rect 25961 31631 26019 31637
rect 26142 31628 26148 31640
rect 26200 31628 26206 31680
rect 26234 31628 26240 31680
rect 26292 31668 26298 31680
rect 26344 31668 26372 31699
rect 26786 31696 26792 31708
rect 26844 31696 26850 31748
rect 26292 31640 26372 31668
rect 26292 31628 26298 31640
rect 27706 31628 27712 31680
rect 27764 31668 27770 31680
rect 27893 31671 27951 31677
rect 27893 31668 27905 31671
rect 27764 31640 27905 31668
rect 27764 31628 27770 31640
rect 27893 31637 27905 31640
rect 27939 31637 27951 31671
rect 27893 31631 27951 31637
rect 27982 31628 27988 31680
rect 28040 31668 28046 31680
rect 28077 31671 28135 31677
rect 28077 31668 28089 31671
rect 28040 31640 28089 31668
rect 28040 31628 28046 31640
rect 28077 31637 28089 31640
rect 28123 31637 28135 31671
rect 28077 31631 28135 31637
rect 29086 31628 29092 31680
rect 29144 31668 29150 31680
rect 29564 31668 29592 31767
rect 29822 31764 29828 31816
rect 29880 31764 29886 31816
rect 29932 31813 29960 31912
rect 30208 31912 30788 31940
rect 29917 31807 29975 31813
rect 29917 31773 29929 31807
rect 29963 31773 29975 31807
rect 29917 31767 29975 31773
rect 30055 31807 30113 31813
rect 30055 31773 30067 31807
rect 30101 31804 30113 31807
rect 30208 31804 30236 31912
rect 30282 31832 30288 31884
rect 30340 31872 30346 31884
rect 30340 31844 30512 31872
rect 30340 31832 30346 31844
rect 30484 31813 30512 31844
rect 30760 31816 30788 31912
rect 31128 31844 31800 31872
rect 30101 31776 30236 31804
rect 30469 31807 30527 31813
rect 30101 31773 30113 31776
rect 30055 31767 30113 31773
rect 30469 31773 30481 31807
rect 30515 31773 30527 31807
rect 30469 31767 30527 31773
rect 30742 31764 30748 31816
rect 30800 31764 30806 31816
rect 31128 31736 31156 31844
rect 31478 31764 31484 31816
rect 31536 31764 31542 31816
rect 31772 31813 31800 31844
rect 31757 31807 31815 31813
rect 31757 31773 31769 31807
rect 31803 31773 31815 31807
rect 31757 31767 31815 31773
rect 30208 31708 31156 31736
rect 31573 31739 31631 31745
rect 30006 31668 30012 31680
rect 29144 31640 30012 31668
rect 29144 31628 29150 31640
rect 30006 31628 30012 31640
rect 30064 31628 30070 31680
rect 30208 31677 30236 31708
rect 31573 31705 31585 31739
rect 31619 31736 31631 31739
rect 31864 31736 31892 31968
rect 31938 31764 31944 31816
rect 31996 31764 32002 31816
rect 34606 31764 34612 31816
rect 34664 31804 34670 31816
rect 34885 31807 34943 31813
rect 34885 31804 34897 31807
rect 34664 31776 34897 31804
rect 34664 31764 34670 31776
rect 34885 31773 34897 31776
rect 34931 31804 34943 31807
rect 34977 31807 35035 31813
rect 34977 31804 34989 31807
rect 34931 31776 34989 31804
rect 34931 31773 34943 31776
rect 34885 31767 34943 31773
rect 34977 31773 34989 31776
rect 35023 31773 35035 31807
rect 34977 31767 35035 31773
rect 35434 31764 35440 31816
rect 35492 31764 35498 31816
rect 31619 31708 31892 31736
rect 31619 31705 31631 31708
rect 31573 31699 31631 31705
rect 34514 31696 34520 31748
rect 34572 31736 34578 31748
rect 35069 31739 35127 31745
rect 35069 31736 35081 31739
rect 34572 31708 35081 31736
rect 34572 31696 34578 31708
rect 35069 31705 35081 31708
rect 35115 31705 35127 31739
rect 35069 31699 35127 31705
rect 30193 31671 30251 31677
rect 30193 31637 30205 31671
rect 30239 31637 30251 31671
rect 30193 31631 30251 31637
rect 30374 31628 30380 31680
rect 30432 31628 30438 31680
rect 34790 31628 34796 31680
rect 34848 31628 34854 31680
rect 35250 31628 35256 31680
rect 35308 31628 35314 31680
rect 1104 31578 38272 31600
rect 1104 31526 4874 31578
rect 4926 31526 4938 31578
rect 4990 31526 5002 31578
rect 5054 31526 5066 31578
rect 5118 31526 5130 31578
rect 5182 31526 35594 31578
rect 35646 31526 35658 31578
rect 35710 31526 35722 31578
rect 35774 31526 35786 31578
rect 35838 31526 35850 31578
rect 35902 31526 38272 31578
rect 1104 31504 38272 31526
rect 8294 31464 8300 31476
rect 8128 31436 8300 31464
rect 8128 31405 8156 31436
rect 8294 31424 8300 31436
rect 8352 31424 8358 31476
rect 9766 31424 9772 31476
rect 9824 31464 9830 31476
rect 9861 31467 9919 31473
rect 9861 31464 9873 31467
rect 9824 31436 9873 31464
rect 9824 31424 9830 31436
rect 9861 31433 9873 31436
rect 9907 31433 9919 31467
rect 9861 31427 9919 31433
rect 10137 31467 10195 31473
rect 10137 31433 10149 31467
rect 10183 31433 10195 31467
rect 10137 31427 10195 31433
rect 10597 31467 10655 31473
rect 10597 31433 10609 31467
rect 10643 31464 10655 31467
rect 10870 31464 10876 31476
rect 10643 31436 10876 31464
rect 10643 31433 10655 31436
rect 10597 31427 10655 31433
rect 8113 31399 8171 31405
rect 8113 31365 8125 31399
rect 8159 31365 8171 31399
rect 8113 31359 8171 31365
rect 8570 31356 8576 31408
rect 8628 31356 8634 31408
rect 10045 31331 10103 31337
rect 10045 31297 10057 31331
rect 10091 31328 10103 31331
rect 10152 31328 10180 31427
rect 10870 31424 10876 31436
rect 10928 31424 10934 31476
rect 11606 31424 11612 31476
rect 11664 31464 11670 31476
rect 11974 31464 11980 31476
rect 11664 31436 11980 31464
rect 11664 31424 11670 31436
rect 11974 31424 11980 31436
rect 12032 31424 12038 31476
rect 12986 31424 12992 31476
rect 13044 31464 13050 31476
rect 13354 31464 13360 31476
rect 13044 31436 13360 31464
rect 13044 31424 13050 31436
rect 13354 31424 13360 31436
rect 13412 31424 13418 31476
rect 13446 31424 13452 31476
rect 13504 31424 13510 31476
rect 16206 31464 16212 31476
rect 14660 31436 16212 31464
rect 11790 31396 11796 31408
rect 10091 31300 10180 31328
rect 10428 31368 11796 31396
rect 10091 31297 10103 31300
rect 10045 31291 10103 31297
rect 7834 31220 7840 31272
rect 7892 31220 7898 31272
rect 9398 31220 9404 31272
rect 9456 31260 9462 31272
rect 9585 31263 9643 31269
rect 9585 31260 9597 31263
rect 9456 31232 9597 31260
rect 9456 31220 9462 31232
rect 9585 31229 9597 31232
rect 9631 31260 9643 31263
rect 10428 31260 10456 31368
rect 11790 31356 11796 31368
rect 11848 31356 11854 31408
rect 10505 31331 10563 31337
rect 10505 31297 10517 31331
rect 10551 31328 10563 31331
rect 11514 31328 11520 31340
rect 10551 31300 11520 31328
rect 10551 31297 10563 31300
rect 10505 31291 10563 31297
rect 11514 31288 11520 31300
rect 11572 31288 11578 31340
rect 11606 31288 11612 31340
rect 11664 31328 11670 31340
rect 11701 31331 11759 31337
rect 11701 31328 11713 31331
rect 11664 31300 11713 31328
rect 11664 31288 11670 31300
rect 11701 31297 11713 31300
rect 11747 31297 11759 31331
rect 11701 31291 11759 31297
rect 11882 31288 11888 31340
rect 11940 31328 11946 31340
rect 12342 31328 12348 31340
rect 11940 31300 12348 31328
rect 11940 31288 11946 31300
rect 12342 31288 12348 31300
rect 12400 31288 12406 31340
rect 14660 31328 14688 31436
rect 16206 31424 16212 31436
rect 16264 31464 16270 31476
rect 17678 31464 17684 31476
rect 16264 31436 17080 31464
rect 16264 31424 16270 31436
rect 14737 31399 14795 31405
rect 14737 31365 14749 31399
rect 14783 31396 14795 31399
rect 14783 31368 16897 31396
rect 14783 31365 14795 31368
rect 14737 31359 14795 31365
rect 13372 31300 14688 31328
rect 9631 31232 10456 31260
rect 9631 31229 9643 31232
rect 9585 31223 9643 31229
rect 10778 31220 10784 31272
rect 10836 31220 10842 31272
rect 11532 31260 11560 31288
rect 13372 31272 13400 31300
rect 15470 31288 15476 31340
rect 15528 31288 15534 31340
rect 15657 31331 15715 31337
rect 15657 31297 15669 31331
rect 15703 31328 15715 31331
rect 15746 31328 15752 31340
rect 15703 31300 15752 31328
rect 15703 31297 15715 31300
rect 15657 31291 15715 31297
rect 15746 31288 15752 31300
rect 15804 31288 15810 31340
rect 15933 31331 15991 31337
rect 15933 31297 15945 31331
rect 15979 31328 15991 31331
rect 16022 31328 16028 31340
rect 15979 31300 16028 31328
rect 15979 31297 15991 31300
rect 15933 31291 15991 31297
rect 16022 31288 16028 31300
rect 16080 31288 16086 31340
rect 16114 31288 16120 31340
rect 16172 31288 16178 31340
rect 16206 31288 16212 31340
rect 16264 31288 16270 31340
rect 16301 31331 16359 31337
rect 16301 31297 16313 31331
rect 16347 31328 16359 31331
rect 16482 31328 16488 31340
rect 16347 31300 16488 31328
rect 16347 31297 16359 31300
rect 16301 31291 16359 31297
rect 16482 31288 16488 31300
rect 16540 31288 16546 31340
rect 16669 31331 16727 31337
rect 16669 31297 16681 31331
rect 16715 31297 16727 31331
rect 16669 31291 16727 31297
rect 16762 31331 16820 31337
rect 16762 31297 16774 31331
rect 16808 31297 16820 31331
rect 16762 31291 16820 31297
rect 13354 31260 13360 31272
rect 11532 31232 13360 31260
rect 13354 31220 13360 31232
rect 13412 31220 13418 31272
rect 15381 31263 15439 31269
rect 15381 31260 15393 31263
rect 14660 31232 15393 31260
rect 9674 31152 9680 31204
rect 9732 31192 9738 31204
rect 10796 31192 10824 31220
rect 9732 31164 10824 31192
rect 9732 31152 9738 31164
rect 14660 31136 14688 31232
rect 15381 31229 15393 31232
rect 15427 31229 15439 31263
rect 15381 31223 15439 31229
rect 15841 31263 15899 31269
rect 15841 31229 15853 31263
rect 15887 31260 15899 31263
rect 16684 31260 16712 31291
rect 15887 31232 16712 31260
rect 15887 31229 15899 31232
rect 15841 31223 15899 31229
rect 16777 31136 16805 31291
rect 16869 31260 16897 31368
rect 16942 31356 16948 31408
rect 17000 31356 17006 31408
rect 17052 31337 17080 31436
rect 17190 31436 17684 31464
rect 17190 31337 17218 31436
rect 17678 31424 17684 31436
rect 17736 31424 17742 31476
rect 18690 31424 18696 31476
rect 18748 31424 18754 31476
rect 18782 31424 18788 31476
rect 18840 31464 18846 31476
rect 19426 31464 19432 31476
rect 18840 31436 19432 31464
rect 18840 31424 18846 31436
rect 19426 31424 19432 31436
rect 19484 31424 19490 31476
rect 19794 31424 19800 31476
rect 19852 31464 19858 31476
rect 19889 31467 19947 31473
rect 19889 31464 19901 31467
rect 19852 31436 19901 31464
rect 19852 31424 19858 31436
rect 19889 31433 19901 31436
rect 19935 31464 19947 31467
rect 20346 31464 20352 31476
rect 19935 31436 20352 31464
rect 19935 31433 19947 31436
rect 19889 31427 19947 31433
rect 20346 31424 20352 31436
rect 20404 31424 20410 31476
rect 20806 31424 20812 31476
rect 20864 31424 20870 31476
rect 20993 31467 21051 31473
rect 20993 31433 21005 31467
rect 21039 31464 21051 31467
rect 21450 31464 21456 31476
rect 21039 31436 21128 31464
rect 21039 31433 21051 31436
rect 20993 31427 21051 31433
rect 19978 31396 19984 31408
rect 17282 31368 19984 31396
rect 17037 31331 17095 31337
rect 17037 31297 17049 31331
rect 17083 31297 17095 31331
rect 17037 31291 17095 31297
rect 17175 31331 17233 31337
rect 17175 31297 17187 31331
rect 17221 31297 17233 31331
rect 17175 31291 17233 31297
rect 17282 31260 17310 31368
rect 19978 31356 19984 31368
rect 20036 31356 20042 31408
rect 20824 31396 20852 31424
rect 20548 31368 20852 31396
rect 17402 31288 17408 31340
rect 17460 31288 17466 31340
rect 17586 31288 17592 31340
rect 17644 31288 17650 31340
rect 17681 31331 17739 31337
rect 17681 31297 17693 31331
rect 17727 31297 17739 31331
rect 17681 31291 17739 31297
rect 17773 31331 17831 31337
rect 17773 31297 17785 31331
rect 17819 31328 17831 31331
rect 17862 31328 17868 31340
rect 17819 31300 17868 31328
rect 17819 31297 17831 31300
rect 17773 31291 17831 31297
rect 16869 31232 17310 31260
rect 17696 31260 17724 31291
rect 17862 31288 17868 31300
rect 17920 31288 17926 31340
rect 18414 31288 18420 31340
rect 18472 31288 18478 31340
rect 18509 31331 18567 31337
rect 18509 31297 18521 31331
rect 18555 31297 18567 31331
rect 18509 31291 18567 31297
rect 18432 31260 18460 31288
rect 17696 31232 18460 31260
rect 17313 31195 17371 31201
rect 17313 31161 17325 31195
rect 17359 31192 17371 31195
rect 18138 31192 18144 31204
rect 17359 31164 18144 31192
rect 17359 31161 17371 31164
rect 17313 31155 17371 31161
rect 18138 31152 18144 31164
rect 18196 31152 18202 31204
rect 18524 31192 18552 31291
rect 18782 31288 18788 31340
rect 18840 31288 18846 31340
rect 19242 31288 19248 31340
rect 19300 31328 19306 31340
rect 19429 31331 19487 31337
rect 19429 31328 19441 31331
rect 19300 31300 19441 31328
rect 19300 31288 19306 31300
rect 19429 31297 19441 31300
rect 19475 31297 19487 31331
rect 19429 31291 19487 31297
rect 19610 31288 19616 31340
rect 19668 31328 19674 31340
rect 20548 31337 20576 31368
rect 19705 31331 19763 31337
rect 19705 31328 19717 31331
rect 19668 31300 19717 31328
rect 19668 31288 19674 31300
rect 19705 31297 19717 31300
rect 19751 31297 19763 31331
rect 19705 31291 19763 31297
rect 20533 31331 20591 31337
rect 20533 31297 20545 31331
rect 20579 31297 20591 31331
rect 20533 31291 20591 31297
rect 20622 31288 20628 31340
rect 20680 31288 20686 31340
rect 20714 31288 20720 31340
rect 20772 31328 20778 31340
rect 20809 31331 20867 31337
rect 20809 31328 20821 31331
rect 20772 31300 20821 31328
rect 20772 31288 20778 31300
rect 20809 31297 20821 31300
rect 20855 31297 20867 31331
rect 20809 31291 20867 31297
rect 20901 31331 20959 31337
rect 20901 31297 20913 31331
rect 20947 31328 20959 31331
rect 21100 31328 21128 31436
rect 21376 31436 21456 31464
rect 21376 31396 21404 31436
rect 21450 31424 21456 31436
rect 21508 31464 21514 31476
rect 22097 31467 22155 31473
rect 22097 31464 22109 31467
rect 21508 31436 22109 31464
rect 21508 31424 21514 31436
rect 22097 31433 22109 31436
rect 22143 31433 22155 31467
rect 22097 31427 22155 31433
rect 22186 31424 22192 31476
rect 22244 31424 22250 31476
rect 22373 31467 22431 31473
rect 22373 31433 22385 31467
rect 22419 31464 22431 31467
rect 23290 31464 23296 31476
rect 22419 31436 23296 31464
rect 22419 31433 22431 31436
rect 22373 31427 22431 31433
rect 23290 31424 23296 31436
rect 23348 31424 23354 31476
rect 28994 31464 29000 31476
rect 27724 31436 29000 31464
rect 21284 31368 21404 31396
rect 21821 31399 21879 31405
rect 20947 31300 21128 31328
rect 20947 31297 20959 31300
rect 20901 31291 20959 31297
rect 21174 31288 21180 31340
rect 21232 31288 21238 31340
rect 21284 31337 21312 31368
rect 21821 31365 21833 31399
rect 21867 31396 21879 31399
rect 21867 31368 22140 31396
rect 21867 31365 21879 31368
rect 21821 31359 21879 31365
rect 21269 31331 21327 31337
rect 21269 31297 21281 31331
rect 21315 31297 21327 31331
rect 21269 31291 21327 31297
rect 20346 31220 20352 31272
rect 20404 31260 20410 31272
rect 21284 31260 21312 31291
rect 21542 31288 21548 31340
rect 21600 31328 21606 31340
rect 22005 31331 22063 31337
rect 22005 31328 22017 31331
rect 21600 31300 22017 31328
rect 21600 31288 21606 31300
rect 22005 31297 22017 31300
rect 22051 31297 22063 31331
rect 22005 31291 22063 31297
rect 22112 31328 22140 31368
rect 22278 31356 22284 31408
rect 22336 31396 22342 31408
rect 23385 31399 23443 31405
rect 23385 31396 23397 31399
rect 22336 31368 23397 31396
rect 22336 31356 22342 31368
rect 23385 31365 23397 31368
rect 23431 31365 23443 31399
rect 23385 31359 23443 31365
rect 25133 31399 25191 31405
rect 25133 31365 25145 31399
rect 25179 31396 25191 31399
rect 25498 31396 25504 31408
rect 25179 31368 25504 31396
rect 25179 31365 25191 31368
rect 25133 31359 25191 31365
rect 25498 31356 25504 31368
rect 25556 31396 25562 31408
rect 27614 31396 27620 31408
rect 25556 31368 27620 31396
rect 25556 31356 25562 31368
rect 27614 31356 27620 31368
rect 27672 31356 27678 31408
rect 22646 31328 22652 31340
rect 22112 31300 22652 31328
rect 20404 31232 21312 31260
rect 20404 31220 20410 31232
rect 21358 31220 21364 31272
rect 21416 31220 21422 31272
rect 21453 31263 21511 31269
rect 21453 31229 21465 31263
rect 21499 31260 21511 31263
rect 21726 31260 21732 31272
rect 21499 31232 21732 31260
rect 21499 31229 21511 31232
rect 21453 31223 21511 31229
rect 21726 31220 21732 31232
rect 21784 31220 21790 31272
rect 22112 31260 22140 31300
rect 22646 31288 22652 31300
rect 22704 31288 22710 31340
rect 22830 31288 22836 31340
rect 22888 31288 22894 31340
rect 23017 31331 23075 31337
rect 23017 31297 23029 31331
rect 23063 31328 23075 31331
rect 23198 31328 23204 31340
rect 23063 31300 23204 31328
rect 23063 31297 23075 31300
rect 23017 31291 23075 31297
rect 23198 31288 23204 31300
rect 23256 31288 23262 31340
rect 23290 31288 23296 31340
rect 23348 31288 23354 31340
rect 25406 31288 25412 31340
rect 25464 31288 25470 31340
rect 25590 31288 25596 31340
rect 25648 31288 25654 31340
rect 25961 31331 26019 31337
rect 25961 31328 25973 31331
rect 25700 31300 25973 31328
rect 21836 31232 22140 31260
rect 18524 31164 18828 31192
rect 18800 31136 18828 31164
rect 20898 31152 20904 31204
rect 20956 31192 20962 31204
rect 21836 31192 21864 31232
rect 22554 31220 22560 31272
rect 22612 31260 22618 31272
rect 22925 31263 22983 31269
rect 22925 31260 22937 31263
rect 22612 31232 22937 31260
rect 22612 31220 22618 31232
rect 22925 31229 22937 31232
rect 22971 31229 22983 31263
rect 22925 31223 22983 31229
rect 23109 31263 23167 31269
rect 23109 31229 23121 31263
rect 23155 31260 23167 31263
rect 23382 31260 23388 31272
rect 23155 31232 23388 31260
rect 23155 31229 23167 31232
rect 23109 31223 23167 31229
rect 23382 31220 23388 31232
rect 23440 31260 23446 31272
rect 24578 31260 24584 31272
rect 23440 31232 24584 31260
rect 23440 31220 23446 31232
rect 24578 31220 24584 31232
rect 24636 31220 24642 31272
rect 25700 31192 25728 31300
rect 25961 31297 25973 31300
rect 26007 31297 26019 31331
rect 25961 31291 26019 31297
rect 26326 31288 26332 31340
rect 26384 31288 26390 31340
rect 26973 31331 27031 31337
rect 26973 31328 26985 31331
rect 26436 31300 26985 31328
rect 26436 31260 26464 31300
rect 26973 31297 26985 31300
rect 27019 31297 27031 31331
rect 26973 31291 27031 31297
rect 27154 31288 27160 31340
rect 27212 31288 27218 31340
rect 27249 31331 27307 31337
rect 27249 31297 27261 31331
rect 27295 31297 27307 31331
rect 27249 31291 27307 31297
rect 27341 31331 27399 31337
rect 27341 31297 27353 31331
rect 27387 31297 27399 31331
rect 27341 31291 27399 31297
rect 20956 31164 21864 31192
rect 22066 31164 25728 31192
rect 26260 31232 26464 31260
rect 20956 31152 20962 31164
rect 12069 31127 12127 31133
rect 12069 31093 12081 31127
rect 12115 31124 12127 31127
rect 13538 31124 13544 31136
rect 12115 31096 13544 31124
rect 12115 31093 12127 31096
rect 12069 31087 12127 31093
rect 13538 31084 13544 31096
rect 13596 31084 13602 31136
rect 14642 31084 14648 31136
rect 14700 31084 14706 31136
rect 16482 31084 16488 31136
rect 16540 31084 16546 31136
rect 16758 31084 16764 31136
rect 16816 31084 16822 31136
rect 17957 31127 18015 31133
rect 17957 31093 17969 31127
rect 18003 31124 18015 31127
rect 18046 31124 18052 31136
rect 18003 31096 18052 31124
rect 18003 31093 18015 31096
rect 17957 31087 18015 31093
rect 18046 31084 18052 31096
rect 18104 31084 18110 31136
rect 18322 31084 18328 31136
rect 18380 31084 18386 31136
rect 18782 31084 18788 31136
rect 18840 31084 18846 31136
rect 20349 31127 20407 31133
rect 20349 31093 20361 31127
rect 20395 31124 20407 31127
rect 22066 31124 22094 31164
rect 20395 31096 22094 31124
rect 20395 31093 20407 31096
rect 20349 31087 20407 31093
rect 22646 31084 22652 31136
rect 22704 31084 22710 31136
rect 25406 31084 25412 31136
rect 25464 31124 25470 31136
rect 25958 31124 25964 31136
rect 25464 31096 25964 31124
rect 25464 31084 25470 31096
rect 25958 31084 25964 31096
rect 26016 31124 26022 31136
rect 26260 31124 26288 31232
rect 26510 31220 26516 31272
rect 26568 31260 26574 31272
rect 27264 31260 27292 31291
rect 26568 31232 27292 31260
rect 26568 31220 26574 31232
rect 26694 31152 26700 31204
rect 26752 31152 26758 31204
rect 27356 31192 27384 31291
rect 27522 31288 27528 31340
rect 27580 31328 27586 31340
rect 27724 31328 27752 31436
rect 27982 31356 27988 31408
rect 28040 31356 28046 31408
rect 28368 31396 28396 31436
rect 28994 31424 29000 31436
rect 29052 31464 29058 31476
rect 29052 31436 29316 31464
rect 29052 31424 29058 31436
rect 29288 31396 29316 31436
rect 34790 31424 34796 31476
rect 34848 31424 34854 31476
rect 34808 31396 34836 31424
rect 28368 31368 28474 31396
rect 29288 31368 30682 31396
rect 32876 31368 32982 31396
rect 34440 31368 34836 31396
rect 32876 31340 32904 31368
rect 27580 31300 27752 31328
rect 27580 31288 27586 31300
rect 29638 31288 29644 31340
rect 29696 31288 29702 31340
rect 29917 31331 29975 31337
rect 29917 31328 29929 31331
rect 29748 31300 29929 31328
rect 27706 31220 27712 31272
rect 27764 31220 27770 31272
rect 26804 31164 27384 31192
rect 26804 31136 26832 31164
rect 26016 31096 26288 31124
rect 26016 31084 26022 31096
rect 26326 31084 26332 31136
rect 26384 31124 26390 31136
rect 26602 31124 26608 31136
rect 26384 31096 26608 31124
rect 26384 31084 26390 31096
rect 26602 31084 26608 31096
rect 26660 31084 26666 31136
rect 26786 31084 26792 31136
rect 26844 31084 26850 31136
rect 27617 31127 27675 31133
rect 27617 31093 27629 31127
rect 27663 31124 27675 31127
rect 27706 31124 27712 31136
rect 27663 31096 27712 31124
rect 27663 31093 27675 31096
rect 27617 31087 27675 31093
rect 27706 31084 27712 31096
rect 27764 31084 27770 31136
rect 29454 31084 29460 31136
rect 29512 31084 29518 31136
rect 29748 31124 29776 31300
rect 29917 31297 29929 31300
rect 29963 31297 29975 31331
rect 29917 31291 29975 31297
rect 31662 31288 31668 31340
rect 31720 31328 31726 31340
rect 32401 31331 32459 31337
rect 32401 31328 32413 31331
rect 31720 31300 32413 31328
rect 31720 31288 31726 31300
rect 32401 31297 32413 31300
rect 32447 31297 32459 31331
rect 32401 31291 32459 31297
rect 32858 31288 32864 31340
rect 32916 31288 32922 31340
rect 34440 31337 34468 31368
rect 34425 31331 34483 31337
rect 34425 31297 34437 31331
rect 34471 31297 34483 31331
rect 34425 31291 34483 31297
rect 34514 31288 34520 31340
rect 34572 31288 34578 31340
rect 35926 31300 36032 31328
rect 30193 31263 30251 31269
rect 30193 31260 30205 31263
rect 29840 31232 30205 31260
rect 29840 31201 29868 31232
rect 30193 31229 30205 31232
rect 30239 31229 30251 31263
rect 30193 31223 30251 31229
rect 31941 31263 31999 31269
rect 31941 31229 31953 31263
rect 31987 31260 31999 31263
rect 32490 31260 32496 31272
rect 31987 31232 32496 31260
rect 31987 31229 31999 31232
rect 31941 31223 31999 31229
rect 32490 31220 32496 31232
rect 32548 31220 32554 31272
rect 34146 31220 34152 31272
rect 34204 31220 34210 31272
rect 34793 31263 34851 31269
rect 34793 31229 34805 31263
rect 34839 31260 34851 31263
rect 35250 31260 35256 31272
rect 34839 31232 35256 31260
rect 34839 31229 34851 31232
rect 34793 31223 34851 31229
rect 35250 31220 35256 31232
rect 35308 31220 35314 31272
rect 29825 31195 29883 31201
rect 29825 31161 29837 31195
rect 29871 31161 29883 31195
rect 29825 31155 29883 31161
rect 36004 31136 36032 31300
rect 36541 31263 36599 31269
rect 36541 31229 36553 31263
rect 36587 31229 36599 31263
rect 36541 31223 36599 31229
rect 36556 31136 36584 31223
rect 30374 31124 30380 31136
rect 29748 31096 30380 31124
rect 30374 31084 30380 31096
rect 30432 31084 30438 31136
rect 31754 31084 31760 31136
rect 31812 31124 31818 31136
rect 32030 31124 32036 31136
rect 31812 31096 32036 31124
rect 31812 31084 31818 31096
rect 32030 31084 32036 31096
rect 32088 31084 32094 31136
rect 35986 31084 35992 31136
rect 36044 31084 36050 31136
rect 36538 31084 36544 31136
rect 36596 31084 36602 31136
rect 1104 31034 38272 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 38272 31034
rect 1104 30960 38272 30982
rect 7834 30880 7840 30932
rect 7892 30880 7898 30932
rect 8478 30880 8484 30932
rect 8536 30920 8542 30932
rect 8941 30923 8999 30929
rect 8941 30920 8953 30923
rect 8536 30892 8953 30920
rect 8536 30880 8542 30892
rect 8941 30889 8953 30892
rect 8987 30889 8999 30923
rect 8941 30883 8999 30889
rect 13354 30880 13360 30932
rect 13412 30880 13418 30932
rect 13630 30880 13636 30932
rect 13688 30920 13694 30932
rect 14461 30923 14519 30929
rect 14461 30920 14473 30923
rect 13688 30892 14473 30920
rect 13688 30880 13694 30892
rect 14461 30889 14473 30892
rect 14507 30889 14519 30923
rect 14461 30883 14519 30889
rect 14550 30880 14556 30932
rect 14608 30880 14614 30932
rect 16485 30923 16543 30929
rect 16485 30889 16497 30923
rect 16531 30920 16543 30923
rect 17586 30920 17592 30932
rect 16531 30892 17592 30920
rect 16531 30889 16543 30892
rect 16485 30883 16543 30889
rect 17586 30880 17592 30892
rect 17644 30880 17650 30932
rect 18506 30880 18512 30932
rect 18564 30920 18570 30932
rect 19150 30920 19156 30932
rect 18564 30892 19156 30920
rect 18564 30880 18570 30892
rect 19150 30880 19156 30892
rect 19208 30920 19214 30932
rect 19337 30923 19395 30929
rect 19337 30920 19349 30923
rect 19208 30892 19349 30920
rect 19208 30880 19214 30892
rect 19337 30889 19349 30892
rect 19383 30889 19395 30923
rect 21269 30923 21327 30929
rect 19337 30883 19395 30889
rect 20548 30892 21036 30920
rect 7374 30744 7380 30796
rect 7432 30784 7438 30796
rect 8389 30787 8447 30793
rect 8389 30784 8401 30787
rect 7432 30756 8401 30784
rect 7432 30744 7438 30756
rect 8389 30753 8401 30756
rect 8435 30753 8447 30787
rect 8389 30747 8447 30753
rect 8570 30744 8576 30796
rect 8628 30744 8634 30796
rect 9398 30744 9404 30796
rect 9456 30744 9462 30796
rect 9490 30744 9496 30796
rect 9548 30744 9554 30796
rect 13372 30793 13400 30880
rect 14568 30852 14596 30880
rect 16758 30852 16764 30864
rect 14568 30824 16764 30852
rect 13357 30787 13415 30793
rect 13357 30753 13369 30787
rect 13403 30753 13415 30787
rect 13357 30747 13415 30753
rect 13909 30787 13967 30793
rect 13909 30753 13921 30787
rect 13955 30784 13967 30787
rect 14553 30787 14611 30793
rect 14553 30784 14565 30787
rect 13955 30756 14565 30784
rect 13955 30753 13967 30756
rect 13909 30747 13967 30753
rect 14553 30753 14565 30756
rect 14599 30753 14611 30787
rect 14553 30747 14611 30753
rect 4525 30719 4583 30725
rect 4525 30685 4537 30719
rect 4571 30716 4583 30719
rect 4571 30688 4660 30716
rect 4571 30685 4583 30688
rect 4525 30679 4583 30685
rect 4632 30592 4660 30688
rect 4798 30676 4804 30728
rect 4856 30716 4862 30728
rect 5626 30716 5632 30728
rect 4856 30688 5632 30716
rect 4856 30676 4862 30688
rect 5626 30676 5632 30688
rect 5684 30676 5690 30728
rect 5721 30719 5779 30725
rect 5721 30685 5733 30719
rect 5767 30716 5779 30719
rect 5905 30719 5963 30725
rect 5905 30716 5917 30719
rect 5767 30688 5917 30716
rect 5767 30685 5779 30688
rect 5721 30679 5779 30685
rect 5905 30685 5917 30688
rect 5951 30685 5963 30719
rect 8588 30716 8616 30744
rect 14369 30719 14427 30725
rect 7314 30702 8616 30716
rect 5905 30679 5963 30685
rect 7300 30688 8616 30702
rect 12406 30688 14320 30716
rect 6178 30608 6184 30660
rect 6236 30608 6242 30660
rect 4246 30540 4252 30592
rect 4304 30580 4310 30592
rect 4433 30583 4491 30589
rect 4433 30580 4445 30583
rect 4304 30552 4445 30580
rect 4304 30540 4310 30552
rect 4433 30549 4445 30552
rect 4479 30549 4491 30583
rect 4433 30543 4491 30549
rect 4614 30540 4620 30592
rect 4672 30540 4678 30592
rect 6362 30540 6368 30592
rect 6420 30580 6426 30592
rect 7300 30580 7328 30688
rect 8205 30651 8263 30657
rect 8205 30648 8217 30651
rect 7668 30620 8217 30648
rect 7668 30589 7696 30620
rect 8205 30617 8217 30620
rect 8251 30648 8263 30651
rect 11698 30648 11704 30660
rect 8251 30620 11704 30648
rect 8251 30617 8263 30620
rect 8205 30611 8263 30617
rect 11698 30608 11704 30620
rect 11756 30648 11762 30660
rect 12406 30648 12434 30688
rect 11756 30620 12434 30648
rect 11756 30608 11762 30620
rect 12986 30608 12992 30660
rect 13044 30608 13050 30660
rect 13170 30608 13176 30660
rect 13228 30648 13234 30660
rect 13228 30620 13676 30648
rect 13228 30608 13234 30620
rect 6420 30552 7328 30580
rect 7653 30583 7711 30589
rect 6420 30540 6426 30552
rect 7653 30549 7665 30583
rect 7699 30549 7711 30583
rect 7653 30543 7711 30549
rect 7742 30540 7748 30592
rect 7800 30580 7806 30592
rect 8297 30583 8355 30589
rect 8297 30580 8309 30583
rect 7800 30552 8309 30580
rect 7800 30540 7806 30552
rect 8297 30549 8309 30552
rect 8343 30580 8355 30583
rect 9309 30583 9367 30589
rect 9309 30580 9321 30583
rect 8343 30552 9321 30580
rect 8343 30549 8355 30552
rect 8297 30543 8355 30549
rect 9309 30549 9321 30552
rect 9355 30580 9367 30583
rect 10870 30580 10876 30592
rect 9355 30552 10876 30580
rect 9355 30549 9367 30552
rect 9309 30543 9367 30549
rect 10870 30540 10876 30552
rect 10928 30540 10934 30592
rect 13004 30580 13032 30608
rect 13648 30592 13676 30620
rect 13722 30608 13728 30660
rect 13780 30648 13786 30660
rect 14292 30648 14320 30688
rect 14369 30685 14381 30719
rect 14415 30716 14427 30719
rect 14458 30716 14464 30728
rect 14415 30688 14464 30716
rect 14415 30685 14427 30688
rect 14369 30679 14427 30685
rect 14458 30676 14464 30688
rect 14516 30676 14522 30728
rect 14642 30676 14648 30728
rect 14700 30676 14706 30728
rect 14734 30676 14740 30728
rect 14792 30716 14798 30728
rect 14829 30719 14887 30725
rect 14829 30716 14841 30719
rect 14792 30688 14841 30716
rect 14792 30676 14798 30688
rect 14829 30685 14841 30688
rect 14875 30685 14887 30719
rect 16301 30719 16359 30725
rect 16301 30716 16313 30719
rect 14829 30679 14887 30685
rect 14936 30688 16313 30716
rect 14660 30648 14688 30676
rect 14936 30648 14964 30688
rect 16301 30685 16313 30688
rect 16347 30685 16359 30719
rect 16301 30679 16359 30685
rect 16574 30676 16580 30728
rect 16632 30676 16638 30728
rect 16685 30725 16713 30824
rect 16758 30812 16764 30824
rect 16816 30812 16822 30864
rect 17310 30852 17316 30864
rect 16869 30824 17316 30852
rect 16869 30725 16897 30824
rect 17310 30812 17316 30824
rect 17368 30812 17374 30864
rect 18874 30812 18880 30864
rect 18932 30852 18938 30864
rect 20548 30852 20576 30892
rect 18932 30824 20576 30852
rect 18932 30812 18938 30824
rect 20714 30812 20720 30864
rect 20772 30812 20778 30864
rect 21008 30852 21036 30892
rect 21269 30889 21281 30923
rect 21315 30920 21327 30923
rect 21910 30920 21916 30932
rect 21315 30892 21916 30920
rect 21315 30889 21327 30892
rect 21269 30883 21327 30889
rect 21910 30880 21916 30892
rect 21968 30880 21974 30932
rect 22002 30880 22008 30932
rect 22060 30920 22066 30932
rect 22060 30892 24348 30920
rect 22060 30880 22066 30892
rect 21008 30824 21772 30852
rect 16942 30744 16948 30796
rect 17000 30784 17006 30796
rect 21744 30793 21772 30824
rect 21729 30787 21787 30793
rect 17000 30756 21680 30784
rect 17000 30744 17006 30756
rect 17126 30725 17132 30728
rect 16670 30719 16728 30725
rect 16670 30685 16682 30719
rect 16716 30685 16728 30719
rect 16670 30679 16728 30685
rect 16853 30719 16911 30725
rect 16853 30685 16865 30719
rect 16899 30685 16911 30719
rect 16853 30679 16911 30685
rect 17083 30719 17132 30725
rect 17083 30685 17095 30719
rect 17129 30685 17132 30719
rect 17083 30679 17132 30685
rect 17126 30676 17132 30679
rect 17184 30676 17190 30728
rect 17954 30676 17960 30728
rect 18012 30716 18018 30728
rect 19242 30716 19248 30728
rect 18012 30688 19248 30716
rect 18012 30676 18018 30688
rect 19242 30676 19248 30688
rect 19300 30716 19306 30728
rect 19337 30719 19395 30725
rect 19337 30716 19349 30719
rect 19300 30688 19349 30716
rect 19300 30676 19306 30688
rect 19337 30685 19349 30688
rect 19383 30685 19395 30719
rect 19337 30679 19395 30685
rect 20070 30676 20076 30728
rect 20128 30676 20134 30728
rect 20346 30676 20352 30728
rect 20404 30676 20410 30728
rect 20530 30676 20536 30728
rect 20588 30716 20594 30728
rect 21358 30716 21364 30728
rect 20588 30688 21364 30716
rect 20588 30676 20594 30688
rect 21358 30676 21364 30688
rect 21416 30676 21422 30728
rect 21652 30716 21680 30756
rect 21729 30753 21741 30787
rect 21775 30784 21787 30787
rect 22554 30784 22560 30796
rect 21775 30756 22560 30784
rect 21775 30753 21787 30756
rect 21729 30747 21787 30753
rect 22554 30744 22560 30756
rect 22612 30784 22618 30796
rect 23290 30784 23296 30796
rect 22612 30756 23296 30784
rect 22612 30744 22618 30756
rect 23290 30744 23296 30756
rect 23348 30744 23354 30796
rect 23382 30716 23388 30728
rect 21652 30688 23388 30716
rect 23382 30676 23388 30688
rect 23440 30676 23446 30728
rect 24320 30716 24348 30892
rect 24486 30880 24492 30932
rect 24544 30880 24550 30932
rect 24857 30923 24915 30929
rect 24857 30889 24869 30923
rect 24903 30920 24915 30923
rect 25130 30920 25136 30932
rect 24903 30892 25136 30920
rect 24903 30889 24915 30892
rect 24857 30883 24915 30889
rect 25130 30880 25136 30892
rect 25188 30880 25194 30932
rect 26605 30923 26663 30929
rect 25976 30892 26556 30920
rect 25976 30852 26004 30892
rect 24596 30824 26004 30852
rect 24596 30796 24624 30824
rect 26050 30812 26056 30864
rect 26108 30812 26114 30864
rect 26528 30852 26556 30892
rect 26605 30889 26617 30923
rect 26651 30920 26663 30923
rect 27154 30920 27160 30932
rect 26651 30892 27160 30920
rect 26651 30889 26663 30892
rect 26605 30883 26663 30889
rect 27154 30880 27160 30892
rect 27212 30880 27218 30932
rect 28077 30923 28135 30929
rect 28077 30889 28089 30923
rect 28123 30920 28135 30923
rect 28258 30920 28264 30932
rect 28123 30892 28264 30920
rect 28123 30889 28135 30892
rect 28077 30883 28135 30889
rect 28258 30880 28264 30892
rect 28316 30880 28322 30932
rect 29638 30880 29644 30932
rect 29696 30920 29702 30932
rect 30101 30923 30159 30929
rect 30101 30920 30113 30923
rect 29696 30892 30113 30920
rect 29696 30880 29702 30892
rect 30101 30889 30113 30892
rect 30147 30889 30159 30923
rect 30101 30883 30159 30889
rect 30650 30880 30656 30932
rect 30708 30920 30714 30932
rect 34057 30923 34115 30929
rect 30708 30892 34008 30920
rect 30708 30880 30714 30892
rect 26786 30852 26792 30864
rect 26528 30824 26792 30852
rect 26786 30812 26792 30824
rect 26844 30852 26850 30864
rect 32490 30852 32496 30864
rect 26844 30824 32496 30852
rect 26844 30812 26850 30824
rect 24578 30744 24584 30796
rect 24636 30744 24642 30796
rect 26068 30784 26096 30812
rect 26068 30756 26464 30784
rect 26436 30728 26464 30756
rect 27798 30744 27804 30796
rect 27856 30784 27862 30796
rect 28626 30784 28632 30796
rect 27856 30756 28632 30784
rect 27856 30744 27862 30756
rect 28626 30744 28632 30756
rect 28684 30744 28690 30796
rect 24394 30716 24400 30728
rect 24320 30688 24400 30716
rect 24394 30676 24400 30688
rect 24452 30716 24458 30728
rect 24489 30719 24547 30725
rect 24489 30716 24501 30719
rect 24452 30688 24501 30716
rect 24452 30676 24458 30688
rect 24489 30685 24501 30688
rect 24535 30685 24547 30719
rect 24489 30679 24547 30685
rect 26053 30719 26111 30725
rect 26053 30685 26065 30719
rect 26099 30685 26111 30719
rect 26053 30679 26111 30685
rect 13780 30620 14228 30648
rect 14292 30620 14964 30648
rect 16117 30651 16175 30657
rect 13780 30608 13786 30620
rect 13354 30580 13360 30592
rect 13004 30552 13360 30580
rect 13354 30540 13360 30552
rect 13412 30580 13418 30592
rect 13541 30583 13599 30589
rect 13541 30580 13553 30583
rect 13412 30552 13553 30580
rect 13412 30540 13418 30552
rect 13541 30549 13553 30552
rect 13587 30549 13599 30583
rect 13541 30543 13599 30549
rect 13630 30540 13636 30592
rect 13688 30540 13694 30592
rect 14090 30540 14096 30592
rect 14148 30540 14154 30592
rect 14200 30580 14228 30620
rect 16117 30617 16129 30651
rect 16163 30648 16175 30651
rect 16945 30651 17003 30657
rect 16163 30620 16344 30648
rect 16163 30617 16175 30620
rect 16117 30611 16175 30617
rect 16316 30592 16344 30620
rect 16945 30617 16957 30651
rect 16991 30617 17003 30651
rect 16945 30611 17003 30617
rect 14366 30580 14372 30592
rect 14200 30552 14372 30580
rect 14366 30540 14372 30552
rect 14424 30540 14430 30592
rect 14458 30540 14464 30592
rect 14516 30580 14522 30592
rect 14826 30580 14832 30592
rect 14516 30552 14832 30580
rect 14516 30540 14522 30552
rect 14826 30540 14832 30552
rect 14884 30540 14890 30592
rect 16298 30540 16304 30592
rect 16356 30540 16362 30592
rect 16666 30540 16672 30592
rect 16724 30580 16730 30592
rect 16960 30580 16988 30611
rect 18138 30608 18144 30660
rect 18196 30648 18202 30660
rect 18598 30648 18604 30660
rect 18196 30620 18604 30648
rect 18196 30608 18202 30620
rect 18598 30608 18604 30620
rect 18656 30608 18662 30660
rect 19058 30608 19064 30660
rect 19116 30608 19122 30660
rect 19886 30608 19892 30660
rect 19944 30648 19950 30660
rect 20088 30648 20116 30676
rect 19944 30620 20392 30648
rect 19944 30608 19950 30620
rect 16724 30552 16988 30580
rect 16724 30540 16730 30552
rect 17218 30540 17224 30592
rect 17276 30540 17282 30592
rect 17773 30583 17831 30589
rect 17773 30549 17785 30583
rect 17819 30580 17831 30583
rect 17954 30580 17960 30592
rect 17819 30552 17960 30580
rect 17819 30549 17831 30552
rect 17773 30543 17831 30549
rect 17954 30540 17960 30552
rect 18012 30580 18018 30592
rect 20162 30580 20168 30592
rect 18012 30552 20168 30580
rect 18012 30540 18018 30552
rect 20162 30540 20168 30552
rect 20220 30540 20226 30592
rect 20364 30580 20392 30620
rect 20622 30608 20628 30660
rect 20680 30648 20686 30660
rect 21174 30648 21180 30660
rect 20680 30620 21180 30648
rect 20680 30608 20686 30620
rect 21174 30608 21180 30620
rect 21232 30608 21238 30660
rect 21545 30651 21603 30657
rect 21545 30648 21557 30651
rect 21284 30620 21557 30648
rect 20714 30580 20720 30592
rect 20364 30552 20720 30580
rect 20714 30540 20720 30552
rect 20772 30580 20778 30592
rect 20901 30583 20959 30589
rect 20901 30580 20913 30583
rect 20772 30552 20913 30580
rect 20772 30540 20778 30552
rect 20901 30549 20913 30552
rect 20947 30549 20959 30583
rect 20901 30543 20959 30549
rect 20990 30540 20996 30592
rect 21048 30540 21054 30592
rect 21082 30540 21088 30592
rect 21140 30580 21146 30592
rect 21284 30580 21312 30620
rect 21545 30617 21557 30620
rect 21591 30617 21603 30651
rect 21545 30611 21603 30617
rect 23566 30608 23572 30660
rect 23624 30648 23630 30660
rect 23624 30620 24164 30648
rect 23624 30608 23630 30620
rect 21140 30552 21312 30580
rect 21140 30540 21146 30552
rect 21634 30540 21640 30592
rect 21692 30580 21698 30592
rect 24026 30580 24032 30592
rect 21692 30552 24032 30580
rect 21692 30540 21698 30552
rect 24026 30540 24032 30552
rect 24084 30540 24090 30592
rect 24136 30580 24164 30620
rect 25038 30608 25044 30660
rect 25096 30648 25102 30660
rect 26068 30648 26096 30679
rect 26142 30676 26148 30728
rect 26200 30676 26206 30728
rect 26329 30719 26387 30725
rect 26329 30685 26341 30719
rect 26375 30685 26387 30719
rect 26329 30679 26387 30685
rect 25096 30620 26096 30648
rect 26344 30648 26372 30679
rect 26418 30676 26424 30728
rect 26476 30676 26482 30728
rect 27246 30676 27252 30728
rect 27304 30716 27310 30728
rect 27430 30716 27436 30728
rect 27304 30688 27436 30716
rect 27304 30676 27310 30688
rect 27430 30676 27436 30688
rect 27488 30676 27494 30728
rect 30469 30719 30527 30725
rect 30469 30685 30481 30719
rect 30515 30716 30527 30719
rect 30576 30716 30604 30824
rect 32490 30812 32496 30824
rect 32548 30812 32554 30864
rect 33781 30855 33839 30861
rect 33060 30824 33548 30852
rect 30745 30787 30803 30793
rect 30745 30753 30757 30787
rect 30791 30784 30803 30787
rect 33060 30784 33088 30824
rect 33520 30796 33548 30824
rect 33781 30821 33793 30855
rect 33827 30821 33839 30855
rect 33781 30815 33839 30821
rect 30791 30756 33088 30784
rect 30791 30753 30803 30756
rect 30745 30747 30803 30753
rect 33134 30744 33140 30796
rect 33192 30744 33198 30796
rect 33502 30744 33508 30796
rect 33560 30744 33566 30796
rect 30515 30688 30604 30716
rect 30852 30688 31064 30716
rect 30515 30685 30527 30688
rect 30469 30679 30527 30685
rect 28537 30651 28595 30657
rect 28537 30648 28549 30651
rect 26344 30620 28549 30648
rect 25096 30608 25102 30620
rect 26344 30580 26372 30620
rect 28537 30617 28549 30620
rect 28583 30648 28595 30651
rect 29454 30648 29460 30660
rect 28583 30620 29460 30648
rect 28583 30617 28595 30620
rect 28537 30611 28595 30617
rect 29454 30608 29460 30620
rect 29512 30608 29518 30660
rect 30374 30608 30380 30660
rect 30432 30648 30438 30660
rect 30852 30648 30880 30688
rect 30432 30620 30880 30648
rect 30432 30608 30438 30620
rect 30926 30608 30932 30660
rect 30984 30608 30990 30660
rect 31036 30648 31064 30688
rect 31110 30676 31116 30728
rect 31168 30716 31174 30728
rect 31662 30716 31668 30728
rect 31168 30688 31668 30716
rect 31168 30676 31174 30688
rect 31662 30676 31668 30688
rect 31720 30716 31726 30728
rect 33413 30719 33471 30725
rect 33413 30716 33425 30719
rect 31720 30688 33425 30716
rect 31720 30676 31726 30688
rect 33413 30685 33425 30688
rect 33459 30685 33471 30719
rect 33796 30716 33824 30815
rect 33980 30796 34008 30892
rect 34057 30889 34069 30923
rect 34103 30920 34115 30923
rect 34146 30920 34152 30932
rect 34103 30892 34152 30920
rect 34103 30889 34115 30892
rect 34057 30883 34115 30889
rect 34146 30880 34152 30892
rect 34204 30880 34210 30932
rect 35434 30880 35440 30932
rect 35492 30880 35498 30932
rect 33962 30744 33968 30796
rect 34020 30784 34026 30796
rect 34793 30787 34851 30793
rect 34793 30784 34805 30787
rect 34020 30756 34805 30784
rect 34020 30744 34026 30756
rect 34793 30753 34805 30756
rect 34839 30753 34851 30787
rect 34793 30747 34851 30753
rect 33873 30719 33931 30725
rect 33873 30716 33885 30719
rect 33796 30688 33885 30716
rect 33413 30679 33471 30685
rect 33873 30685 33885 30688
rect 33919 30685 33931 30719
rect 33873 30679 33931 30685
rect 31570 30648 31576 30660
rect 31036 30620 31576 30648
rect 31570 30608 31576 30620
rect 31628 30648 31634 30660
rect 34977 30651 35035 30657
rect 34977 30648 34989 30651
rect 31628 30620 34989 30648
rect 31628 30608 31634 30620
rect 34977 30617 34989 30620
rect 35023 30648 35035 30651
rect 36538 30648 36544 30660
rect 35023 30620 36544 30648
rect 35023 30617 35035 30620
rect 34977 30611 35035 30617
rect 36538 30608 36544 30620
rect 36596 30608 36602 30660
rect 24136 30552 26372 30580
rect 28442 30540 28448 30592
rect 28500 30580 28506 30592
rect 30561 30583 30619 30589
rect 30561 30580 30573 30583
rect 28500 30552 30573 30580
rect 28500 30540 28506 30552
rect 30561 30549 30573 30552
rect 30607 30580 30619 30583
rect 31018 30580 31024 30592
rect 30607 30552 31024 30580
rect 30607 30549 30619 30552
rect 30561 30543 30619 30549
rect 31018 30540 31024 30552
rect 31076 30540 31082 30592
rect 31294 30540 31300 30592
rect 31352 30580 31358 30592
rect 32217 30583 32275 30589
rect 32217 30580 32229 30583
rect 31352 30552 32229 30580
rect 31352 30540 31358 30552
rect 32217 30549 32229 30552
rect 32263 30549 32275 30583
rect 32217 30543 32275 30549
rect 33318 30540 33324 30592
rect 33376 30580 33382 30592
rect 35069 30583 35127 30589
rect 35069 30580 35081 30583
rect 33376 30552 35081 30580
rect 33376 30540 33382 30552
rect 35069 30549 35081 30552
rect 35115 30549 35127 30583
rect 35069 30543 35127 30549
rect 1104 30490 38272 30512
rect 1104 30438 4874 30490
rect 4926 30438 4938 30490
rect 4990 30438 5002 30490
rect 5054 30438 5066 30490
rect 5118 30438 5130 30490
rect 5182 30438 35594 30490
rect 35646 30438 35658 30490
rect 35710 30438 35722 30490
rect 35774 30438 35786 30490
rect 35838 30438 35850 30490
rect 35902 30438 38272 30490
rect 1104 30416 38272 30438
rect 5997 30379 6055 30385
rect 5997 30345 6009 30379
rect 6043 30345 6055 30379
rect 5997 30339 6055 30345
rect 5258 30268 5264 30320
rect 5316 30268 5322 30320
rect 6012 30240 6040 30339
rect 6178 30336 6184 30388
rect 6236 30376 6242 30388
rect 6457 30379 6515 30385
rect 6457 30376 6469 30379
rect 6236 30348 6469 30376
rect 6236 30336 6242 30348
rect 6457 30345 6469 30348
rect 6503 30345 6515 30379
rect 7834 30376 7840 30388
rect 6457 30339 6515 30345
rect 7208 30348 7840 30376
rect 6641 30243 6699 30249
rect 6012 30212 6592 30240
rect 4246 30132 4252 30184
rect 4304 30132 4310 30184
rect 4525 30175 4583 30181
rect 4525 30141 4537 30175
rect 4571 30172 4583 30175
rect 6564 30172 6592 30212
rect 6641 30209 6653 30243
rect 6687 30240 6699 30243
rect 7208 30240 7236 30348
rect 7834 30336 7840 30348
rect 7892 30336 7898 30388
rect 9582 30336 9588 30388
rect 9640 30376 9646 30388
rect 13446 30376 13452 30388
rect 9640 30348 13452 30376
rect 9640 30336 9646 30348
rect 13446 30336 13452 30348
rect 13504 30336 13510 30388
rect 13630 30336 13636 30388
rect 13688 30376 13694 30388
rect 14550 30376 14556 30388
rect 13688 30348 14556 30376
rect 13688 30336 13694 30348
rect 14550 30336 14556 30348
rect 14608 30336 14614 30388
rect 14918 30336 14924 30388
rect 14976 30376 14982 30388
rect 18874 30376 18880 30388
rect 14976 30348 18880 30376
rect 14976 30336 14982 30348
rect 18874 30336 18880 30348
rect 18932 30336 18938 30388
rect 23842 30376 23848 30388
rect 19306 30348 23848 30376
rect 7377 30311 7435 30317
rect 7377 30277 7389 30311
rect 7423 30308 7435 30311
rect 7423 30280 8064 30308
rect 7423 30277 7435 30280
rect 7377 30271 7435 30277
rect 6687 30212 7236 30240
rect 6687 30209 6699 30212
rect 6641 30203 6699 30209
rect 7466 30200 7472 30252
rect 7524 30240 7530 30252
rect 7653 30243 7711 30249
rect 7653 30240 7665 30243
rect 7524 30212 7665 30240
rect 7524 30200 7530 30212
rect 7653 30209 7665 30212
rect 7699 30209 7711 30243
rect 7653 30203 7711 30209
rect 7742 30200 7748 30252
rect 7800 30200 7806 30252
rect 7837 30243 7895 30249
rect 7837 30209 7849 30243
rect 7883 30240 7895 30243
rect 7926 30240 7932 30252
rect 7883 30212 7932 30240
rect 7883 30209 7895 30212
rect 7837 30203 7895 30209
rect 7926 30200 7932 30212
rect 7984 30200 7990 30252
rect 8036 30249 8064 30280
rect 8386 30268 8392 30320
rect 8444 30308 8450 30320
rect 8444 30280 8616 30308
rect 8444 30268 8450 30280
rect 8588 30252 8616 30280
rect 9950 30268 9956 30320
rect 10008 30308 10014 30320
rect 12989 30311 13047 30317
rect 12989 30308 13001 30311
rect 10008 30280 13001 30308
rect 10008 30268 10014 30280
rect 12989 30277 13001 30280
rect 13035 30277 13047 30311
rect 12989 30271 13047 30277
rect 14752 30280 19104 30308
rect 8021 30243 8079 30249
rect 8021 30209 8033 30243
rect 8067 30209 8079 30243
rect 8021 30203 8079 30209
rect 8570 30200 8576 30252
rect 8628 30200 8634 30252
rect 9490 30200 9496 30252
rect 9548 30240 9554 30252
rect 10042 30240 10048 30252
rect 9548 30212 10048 30240
rect 9548 30200 9554 30212
rect 10042 30200 10048 30212
rect 10100 30200 10106 30252
rect 11422 30200 11428 30252
rect 11480 30240 11486 30252
rect 11609 30243 11667 30249
rect 11609 30240 11621 30243
rect 11480 30212 11621 30240
rect 11480 30200 11486 30212
rect 11609 30209 11621 30212
rect 11655 30209 11667 30243
rect 11609 30203 11667 30209
rect 11698 30200 11704 30252
rect 11756 30240 11762 30252
rect 11756 30212 11801 30240
rect 11756 30200 11762 30212
rect 11882 30200 11888 30252
rect 11940 30200 11946 30252
rect 11977 30243 12035 30249
rect 11977 30209 11989 30243
rect 12023 30209 12035 30243
rect 11977 30203 12035 30209
rect 12115 30243 12173 30249
rect 12115 30209 12127 30243
rect 12161 30240 12173 30243
rect 12250 30240 12256 30252
rect 12161 30212 12256 30240
rect 12161 30209 12173 30212
rect 12115 30203 12173 30209
rect 6733 30175 6791 30181
rect 6733 30172 6745 30175
rect 4571 30144 6040 30172
rect 6564 30144 6745 30172
rect 4571 30141 4583 30144
rect 4525 30135 4583 30141
rect 6012 30104 6040 30144
rect 6733 30141 6745 30144
rect 6779 30172 6791 30175
rect 11992 30172 12020 30203
rect 12250 30200 12256 30212
rect 12308 30200 12314 30252
rect 14752 30249 14780 30280
rect 14737 30243 14795 30249
rect 14737 30209 14749 30243
rect 14783 30209 14795 30243
rect 14737 30203 14795 30209
rect 16482 30200 16488 30252
rect 16540 30240 16546 30252
rect 17681 30243 17739 30249
rect 17681 30240 17693 30243
rect 16540 30212 17693 30240
rect 16540 30200 16546 30212
rect 17681 30209 17693 30212
rect 17727 30209 17739 30243
rect 17681 30203 17739 30209
rect 18046 30200 18052 30252
rect 18104 30200 18110 30252
rect 18138 30200 18144 30252
rect 18196 30240 18202 30252
rect 18417 30243 18475 30249
rect 18417 30240 18429 30243
rect 18196 30212 18429 30240
rect 18196 30200 18202 30212
rect 18417 30209 18429 30212
rect 18463 30209 18475 30243
rect 18417 30203 18475 30209
rect 18506 30200 18512 30252
rect 18564 30200 18570 30252
rect 18598 30200 18604 30252
rect 18656 30200 18662 30252
rect 18782 30200 18788 30252
rect 18840 30200 18846 30252
rect 19076 30240 19104 30280
rect 19150 30268 19156 30320
rect 19208 30308 19214 30320
rect 19306 30308 19334 30348
rect 19208 30280 19334 30308
rect 19208 30268 19214 30280
rect 19886 30268 19892 30320
rect 19944 30268 19950 30320
rect 20070 30268 20076 30320
rect 20128 30268 20134 30320
rect 20456 30317 20484 30348
rect 23842 30336 23848 30348
rect 23900 30376 23906 30388
rect 24486 30376 24492 30388
rect 23900 30348 24492 30376
rect 23900 30336 23906 30348
rect 24486 30336 24492 30348
rect 24544 30336 24550 30388
rect 32858 30376 32864 30388
rect 25700 30348 28994 30376
rect 20441 30311 20499 30317
rect 20441 30277 20453 30311
rect 20487 30277 20499 30311
rect 20441 30271 20499 30277
rect 20622 30268 20628 30320
rect 20680 30268 20686 30320
rect 20806 30268 20812 30320
rect 20864 30308 20870 30320
rect 24210 30308 24216 30320
rect 20864 30280 24216 30308
rect 20864 30268 20870 30280
rect 24210 30268 24216 30280
rect 24268 30268 24274 30320
rect 20254 30240 20260 30252
rect 19076 30212 20260 30240
rect 20254 30200 20260 30212
rect 20312 30240 20318 30252
rect 25700 30249 25728 30348
rect 25869 30311 25927 30317
rect 25869 30277 25881 30311
rect 25915 30308 25927 30311
rect 28966 30308 28994 30348
rect 31726 30348 32864 30376
rect 30650 30308 30656 30320
rect 25915 30280 26188 30308
rect 28966 30280 30656 30308
rect 25915 30277 25927 30280
rect 25869 30271 25927 30277
rect 26160 30252 26188 30280
rect 30650 30268 30656 30280
rect 30708 30308 30714 30320
rect 31110 30308 31116 30320
rect 30708 30280 31116 30308
rect 30708 30268 30714 30280
rect 31110 30268 31116 30280
rect 31168 30268 31174 30320
rect 23385 30243 23443 30249
rect 23385 30240 23397 30243
rect 20312 30212 23397 30240
rect 20312 30200 20318 30212
rect 23385 30209 23397 30212
rect 23431 30209 23443 30243
rect 25685 30243 25743 30249
rect 25685 30240 25697 30243
rect 23385 30203 23443 30209
rect 24688 30212 25697 30240
rect 14826 30172 14832 30184
rect 6779 30144 14832 30172
rect 6779 30141 6791 30144
rect 6733 30135 6791 30141
rect 14826 30132 14832 30144
rect 14884 30172 14890 30184
rect 16666 30172 16672 30184
rect 14884 30144 16672 30172
rect 14884 30132 14890 30144
rect 16666 30132 16672 30144
rect 16724 30132 16730 30184
rect 17218 30132 17224 30184
rect 17276 30172 17282 30184
rect 17773 30175 17831 30181
rect 17773 30172 17785 30175
rect 17276 30144 17785 30172
rect 17276 30132 17282 30144
rect 17773 30141 17785 30144
rect 17819 30141 17831 30175
rect 17773 30135 17831 30141
rect 7469 30107 7527 30113
rect 7469 30104 7481 30107
rect 6012 30076 7481 30104
rect 7469 30073 7481 30076
rect 7515 30073 7527 30107
rect 9490 30104 9496 30116
rect 7469 30067 7527 30073
rect 7576 30076 9496 30104
rect 5258 29996 5264 30048
rect 5316 30036 5322 30048
rect 5718 30036 5724 30048
rect 5316 30008 5724 30036
rect 5316 29996 5322 30008
rect 5718 29996 5724 30008
rect 5776 29996 5782 30048
rect 6822 29996 6828 30048
rect 6880 30036 6886 30048
rect 7576 30036 7604 30076
rect 9490 30064 9496 30076
rect 9548 30064 9554 30116
rect 14274 30064 14280 30116
rect 14332 30104 14338 30116
rect 14734 30104 14740 30116
rect 14332 30076 14740 30104
rect 14332 30064 14338 30076
rect 14734 30064 14740 30076
rect 14792 30064 14798 30116
rect 18064 30104 18092 30200
rect 18524 30172 18552 30200
rect 18524 30144 18644 30172
rect 18616 30116 18644 30144
rect 18690 30132 18696 30184
rect 18748 30172 18754 30184
rect 24688 30172 24716 30212
rect 25685 30209 25697 30212
rect 25731 30209 25743 30243
rect 25685 30203 25743 30209
rect 25957 30243 26015 30249
rect 25957 30209 25969 30243
rect 26003 30209 26015 30243
rect 25957 30203 26015 30209
rect 26053 30243 26111 30249
rect 26053 30209 26065 30243
rect 26099 30209 26111 30243
rect 26053 30203 26111 30209
rect 18748 30144 24716 30172
rect 25133 30175 25191 30181
rect 18748 30132 18754 30144
rect 25133 30141 25145 30175
rect 25179 30172 25191 30175
rect 25590 30172 25596 30184
rect 25179 30144 25596 30172
rect 25179 30141 25191 30144
rect 25133 30135 25191 30141
rect 25590 30132 25596 30144
rect 25648 30132 25654 30184
rect 17788 30076 18092 30104
rect 6880 30008 7604 30036
rect 6880 29996 6886 30008
rect 7926 29996 7932 30048
rect 7984 30036 7990 30048
rect 8665 30039 8723 30045
rect 8665 30036 8677 30039
rect 7984 30008 8677 30036
rect 7984 29996 7990 30008
rect 8665 30005 8677 30008
rect 8711 30036 8723 30039
rect 9398 30036 9404 30048
rect 8711 30008 9404 30036
rect 8711 30005 8723 30008
rect 8665 29999 8723 30005
rect 9398 29996 9404 30008
rect 9456 29996 9462 30048
rect 12250 29996 12256 30048
rect 12308 29996 12314 30048
rect 12342 29996 12348 30048
rect 12400 30036 12406 30048
rect 13722 30036 13728 30048
rect 12400 30008 13728 30036
rect 12400 29996 12406 30008
rect 13722 29996 13728 30008
rect 13780 29996 13786 30048
rect 15010 29996 15016 30048
rect 15068 30036 15074 30048
rect 15838 30036 15844 30048
rect 15068 30008 15844 30036
rect 15068 29996 15074 30008
rect 15838 29996 15844 30008
rect 15896 29996 15902 30048
rect 16114 29996 16120 30048
rect 16172 30036 16178 30048
rect 16942 30036 16948 30048
rect 16172 30008 16948 30036
rect 16172 29996 16178 30008
rect 16942 29996 16948 30008
rect 17000 29996 17006 30048
rect 17788 30045 17816 30076
rect 18598 30064 18604 30116
rect 18656 30064 18662 30116
rect 20254 30064 20260 30116
rect 20312 30064 20318 30116
rect 20364 30076 21036 30104
rect 17773 30039 17831 30045
rect 17773 30005 17785 30039
rect 17819 30005 17831 30039
rect 17773 29999 17831 30005
rect 18046 29996 18052 30048
rect 18104 29996 18110 30048
rect 18141 30039 18199 30045
rect 18141 30005 18153 30039
rect 18187 30036 18199 30039
rect 18322 30036 18328 30048
rect 18187 30008 18328 30036
rect 18187 30005 18199 30008
rect 18141 29999 18199 30005
rect 18322 29996 18328 30008
rect 18380 29996 18386 30048
rect 19426 29996 19432 30048
rect 19484 30036 19490 30048
rect 20073 30039 20131 30045
rect 20073 30036 20085 30039
rect 19484 30008 20085 30036
rect 19484 29996 19490 30008
rect 20073 30005 20085 30008
rect 20119 30036 20131 30039
rect 20364 30036 20392 30076
rect 21008 30048 21036 30076
rect 25314 30064 25320 30116
rect 25372 30064 25378 30116
rect 25866 30064 25872 30116
rect 25924 30104 25930 30116
rect 25976 30104 26004 30203
rect 25924 30076 26004 30104
rect 25924 30064 25930 30076
rect 20119 30008 20392 30036
rect 20119 30005 20131 30008
rect 20073 29999 20131 30005
rect 20438 29996 20444 30048
rect 20496 30036 20502 30048
rect 20625 30039 20683 30045
rect 20625 30036 20637 30039
rect 20496 30008 20637 30036
rect 20496 29996 20502 30008
rect 20625 30005 20637 30008
rect 20671 30005 20683 30039
rect 20625 29999 20683 30005
rect 20806 29996 20812 30048
rect 20864 29996 20870 30048
rect 20990 29996 20996 30048
rect 21048 29996 21054 30048
rect 25332 30036 25360 30064
rect 26068 30036 26096 30203
rect 26142 30200 26148 30252
rect 26200 30200 26206 30252
rect 30377 30243 30435 30249
rect 30377 30209 30389 30243
rect 30423 30240 30435 30243
rect 31294 30240 31300 30252
rect 30423 30212 31300 30240
rect 30423 30209 30435 30212
rect 30377 30203 30435 30209
rect 31294 30200 31300 30212
rect 31352 30200 31358 30252
rect 29822 30132 29828 30184
rect 29880 30172 29886 30184
rect 30558 30172 30564 30184
rect 29880 30144 30564 30172
rect 29880 30132 29886 30144
rect 30558 30132 30564 30144
rect 30616 30132 30622 30184
rect 29089 30107 29147 30113
rect 29089 30073 29101 30107
rect 29135 30104 29147 30107
rect 30282 30104 30288 30116
rect 29135 30076 30288 30104
rect 29135 30073 29147 30076
rect 29089 30067 29147 30073
rect 30282 30064 30288 30076
rect 30340 30064 30346 30116
rect 31110 30064 31116 30116
rect 31168 30104 31174 30116
rect 31726 30104 31754 30348
rect 32858 30336 32864 30348
rect 32916 30376 32922 30388
rect 32916 30348 36032 30376
rect 32916 30336 32922 30348
rect 36004 30320 36032 30348
rect 33042 30308 33048 30320
rect 32416 30280 33048 30308
rect 32122 30200 32128 30252
rect 32180 30200 32186 30252
rect 32306 30200 32312 30252
rect 32364 30200 32370 30252
rect 32416 30249 32444 30280
rect 33042 30268 33048 30280
rect 33100 30308 33106 30320
rect 33226 30308 33232 30320
rect 33100 30280 33232 30308
rect 33100 30268 33106 30280
rect 33226 30268 33232 30280
rect 33284 30268 33290 30320
rect 35986 30268 35992 30320
rect 36044 30268 36050 30320
rect 32401 30243 32459 30249
rect 32401 30209 32413 30243
rect 32447 30209 32459 30243
rect 32401 30203 32459 30209
rect 32490 30200 32496 30252
rect 32548 30200 32554 30252
rect 31168 30076 31754 30104
rect 31168 30064 31174 30076
rect 25332 30008 26096 30036
rect 26234 29996 26240 30048
rect 26292 29996 26298 30048
rect 26602 29996 26608 30048
rect 26660 30036 26666 30048
rect 32490 30036 32496 30048
rect 26660 30008 32496 30036
rect 26660 29996 26666 30008
rect 32490 29996 32496 30008
rect 32548 29996 32554 30048
rect 32769 30039 32827 30045
rect 32769 30005 32781 30039
rect 32815 30036 32827 30039
rect 32950 30036 32956 30048
rect 32815 30008 32956 30036
rect 32815 30005 32827 30008
rect 32769 29999 32827 30005
rect 32950 29996 32956 30008
rect 33008 29996 33014 30048
rect 1104 29946 38272 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 38272 29946
rect 1104 29872 38272 29894
rect 12250 29792 12256 29844
rect 12308 29832 12314 29844
rect 15749 29835 15807 29841
rect 15749 29832 15761 29835
rect 12308 29804 12434 29832
rect 12308 29792 12314 29804
rect 8481 29767 8539 29773
rect 8481 29733 8493 29767
rect 8527 29733 8539 29767
rect 8481 29727 8539 29733
rect 6089 29699 6147 29705
rect 6089 29665 6101 29699
rect 6135 29696 6147 29699
rect 6822 29696 6828 29708
rect 6135 29668 6828 29696
rect 6135 29665 6147 29668
rect 6089 29659 6147 29665
rect 6822 29656 6828 29668
rect 6880 29656 6886 29708
rect 8496 29696 8524 29727
rect 9217 29699 9275 29705
rect 9217 29696 9229 29699
rect 8496 29668 9229 29696
rect 9217 29665 9229 29668
rect 9263 29665 9275 29699
rect 12406 29696 12434 29804
rect 14384 29804 15761 29832
rect 14384 29773 14412 29804
rect 15749 29801 15761 29804
rect 15795 29801 15807 29835
rect 15749 29795 15807 29801
rect 16574 29792 16580 29844
rect 16632 29832 16638 29844
rect 16669 29835 16727 29841
rect 16669 29832 16681 29835
rect 16632 29804 16681 29832
rect 16632 29792 16638 29804
rect 16669 29801 16681 29804
rect 16715 29801 16727 29835
rect 18690 29832 18696 29844
rect 16669 29795 16727 29801
rect 16868 29804 18696 29832
rect 13725 29767 13783 29773
rect 13725 29733 13737 29767
rect 13771 29764 13783 29767
rect 14093 29767 14151 29773
rect 14093 29764 14105 29767
rect 13771 29736 14105 29764
rect 13771 29733 13783 29736
rect 13725 29727 13783 29733
rect 14093 29733 14105 29736
rect 14139 29733 14151 29767
rect 14093 29727 14151 29733
rect 14369 29767 14427 29773
rect 14369 29733 14381 29767
rect 14415 29733 14427 29767
rect 15105 29767 15163 29773
rect 15105 29764 15117 29767
rect 14369 29727 14427 29733
rect 14476 29736 15117 29764
rect 14476 29705 14504 29736
rect 15105 29733 15117 29736
rect 15151 29733 15163 29767
rect 15105 29727 15163 29733
rect 15378 29724 15384 29776
rect 15436 29764 15442 29776
rect 15436 29736 15792 29764
rect 15436 29724 15442 29736
rect 14461 29699 14519 29705
rect 12406 29668 13492 29696
rect 9217 29659 9275 29665
rect 4157 29631 4215 29637
rect 4157 29597 4169 29631
rect 4203 29597 4215 29631
rect 4157 29591 4215 29597
rect 4172 29560 4200 29591
rect 8294 29588 8300 29640
rect 8352 29588 8358 29640
rect 8573 29631 8631 29637
rect 8573 29597 8585 29631
rect 8619 29597 8631 29631
rect 8573 29591 8631 29597
rect 8665 29631 8723 29637
rect 8665 29597 8677 29631
rect 8711 29628 8723 29631
rect 8941 29631 8999 29637
rect 8941 29628 8953 29631
rect 8711 29600 8953 29628
rect 8711 29597 8723 29600
rect 8665 29591 8723 29597
rect 8941 29597 8953 29600
rect 8987 29597 8999 29631
rect 8941 29591 8999 29597
rect 4614 29560 4620 29572
rect 4172 29532 4620 29560
rect 4614 29520 4620 29532
rect 4672 29520 4678 29572
rect 5813 29563 5871 29569
rect 5813 29529 5825 29563
rect 5859 29560 5871 29563
rect 6822 29560 6828 29572
rect 5859 29532 6828 29560
rect 5859 29529 5871 29532
rect 5813 29523 5871 29529
rect 6822 29520 6828 29532
rect 6880 29520 6886 29572
rect 4062 29452 4068 29504
rect 4120 29452 4126 29504
rect 5442 29452 5448 29504
rect 5500 29452 5506 29504
rect 5902 29452 5908 29504
rect 5960 29492 5966 29504
rect 8386 29492 8392 29504
rect 5960 29464 8392 29492
rect 5960 29452 5966 29464
rect 8386 29452 8392 29464
rect 8444 29452 8450 29504
rect 8588 29492 8616 29591
rect 10962 29588 10968 29640
rect 11020 29628 11026 29640
rect 12529 29631 12587 29637
rect 12529 29628 12541 29631
rect 11020 29600 12541 29628
rect 11020 29588 11026 29600
rect 12529 29597 12541 29600
rect 12575 29597 12587 29631
rect 12529 29591 12587 29597
rect 12710 29588 12716 29640
rect 12768 29588 12774 29640
rect 13464 29637 13492 29668
rect 14461 29665 14473 29699
rect 14507 29665 14519 29699
rect 14461 29659 14519 29665
rect 14826 29656 14832 29708
rect 14884 29696 14890 29708
rect 14884 29668 15424 29696
rect 14884 29656 14890 29668
rect 12897 29631 12955 29637
rect 12897 29597 12909 29631
rect 12943 29597 12955 29631
rect 12897 29591 12955 29597
rect 13449 29631 13507 29637
rect 13449 29597 13461 29631
rect 13495 29597 13507 29631
rect 13449 29591 13507 29597
rect 9674 29520 9680 29572
rect 9732 29520 9738 29572
rect 12912 29560 12940 29591
rect 13538 29588 13544 29640
rect 13596 29588 13602 29640
rect 13814 29588 13820 29640
rect 13872 29588 13878 29640
rect 14090 29588 14096 29640
rect 14148 29628 14154 29640
rect 14277 29631 14335 29637
rect 14277 29628 14289 29631
rect 14148 29600 14289 29628
rect 14148 29588 14154 29600
rect 14277 29597 14289 29600
rect 14323 29597 14335 29631
rect 14277 29591 14335 29597
rect 14553 29631 14611 29637
rect 14553 29597 14565 29631
rect 14599 29597 14611 29631
rect 14553 29591 14611 29597
rect 14737 29631 14795 29637
rect 14737 29597 14749 29631
rect 14783 29628 14795 29631
rect 14783 29600 14964 29628
rect 14783 29597 14795 29600
rect 14737 29591 14795 29597
rect 14568 29560 14596 29591
rect 14936 29572 14964 29600
rect 15194 29588 15200 29640
rect 15252 29628 15258 29640
rect 15396 29637 15424 29668
rect 15289 29631 15347 29637
rect 15289 29628 15301 29631
rect 15252 29600 15301 29628
rect 15252 29588 15258 29600
rect 15289 29597 15301 29600
rect 15335 29597 15347 29631
rect 15289 29591 15347 29597
rect 15381 29631 15439 29637
rect 15381 29597 15393 29631
rect 15427 29597 15439 29631
rect 15381 29591 15439 29597
rect 15473 29631 15531 29637
rect 15473 29597 15485 29631
rect 15519 29628 15531 29631
rect 15562 29628 15568 29640
rect 15519 29600 15568 29628
rect 15519 29597 15531 29600
rect 15473 29591 15531 29597
rect 15562 29588 15568 29600
rect 15620 29588 15626 29640
rect 15654 29588 15660 29640
rect 15712 29588 15718 29640
rect 14826 29560 14832 29572
rect 12912 29532 14832 29560
rect 14826 29520 14832 29532
rect 14884 29520 14890 29572
rect 14918 29520 14924 29572
rect 14976 29520 14982 29572
rect 15764 29560 15792 29736
rect 16868 29696 16896 29804
rect 18690 29792 18696 29804
rect 18748 29792 18754 29844
rect 20346 29792 20352 29844
rect 20404 29832 20410 29844
rect 20622 29832 20628 29844
rect 20404 29804 20628 29832
rect 20404 29792 20410 29804
rect 20622 29792 20628 29804
rect 20680 29792 20686 29844
rect 23106 29832 23112 29844
rect 20732 29804 23112 29832
rect 18046 29724 18052 29776
rect 18104 29764 18110 29776
rect 18104 29736 18644 29764
rect 18104 29724 18110 29736
rect 16224 29668 16896 29696
rect 15838 29588 15844 29640
rect 15896 29628 15902 29640
rect 15933 29631 15991 29637
rect 15933 29628 15945 29631
rect 15896 29600 15945 29628
rect 15896 29588 15902 29600
rect 15933 29597 15945 29600
rect 15979 29597 15991 29631
rect 15933 29591 15991 29597
rect 16022 29588 16028 29640
rect 16080 29637 16086 29640
rect 16080 29628 16091 29637
rect 16224 29628 16252 29668
rect 16080 29600 16252 29628
rect 16301 29631 16359 29637
rect 16080 29591 16091 29600
rect 16301 29597 16313 29631
rect 16347 29597 16359 29631
rect 16301 29591 16359 29597
rect 16853 29631 16911 29637
rect 16853 29597 16865 29631
rect 16899 29628 16911 29631
rect 17494 29628 17500 29640
rect 16899 29600 17500 29628
rect 16899 29597 16911 29600
rect 16853 29591 16911 29597
rect 16080 29588 16086 29591
rect 16117 29563 16175 29569
rect 16117 29560 16129 29563
rect 15764 29532 16129 29560
rect 16117 29529 16129 29532
rect 16163 29529 16175 29563
rect 16316 29560 16344 29591
rect 17494 29588 17500 29600
rect 17552 29588 17558 29640
rect 18138 29588 18144 29640
rect 18196 29628 18202 29640
rect 18233 29631 18291 29637
rect 18233 29628 18245 29631
rect 18196 29600 18245 29628
rect 18196 29588 18202 29600
rect 18233 29597 18245 29600
rect 18279 29597 18291 29631
rect 18233 29591 18291 29597
rect 18322 29588 18328 29640
rect 18380 29588 18386 29640
rect 18616 29637 18644 29736
rect 18966 29724 18972 29776
rect 19024 29764 19030 29776
rect 19978 29764 19984 29776
rect 19024 29736 19984 29764
rect 19024 29724 19030 29736
rect 19978 29724 19984 29736
rect 20036 29724 20042 29776
rect 20254 29724 20260 29776
rect 20312 29764 20318 29776
rect 20732 29764 20760 29804
rect 20312 29736 20760 29764
rect 20312 29724 20318 29736
rect 19702 29656 19708 29708
rect 19760 29696 19766 29708
rect 20272 29696 20300 29724
rect 19760 29668 20300 29696
rect 22848 29696 22876 29804
rect 23106 29792 23112 29804
rect 23164 29792 23170 29844
rect 24486 29792 24492 29844
rect 24544 29832 24550 29844
rect 24581 29835 24639 29841
rect 24581 29832 24593 29835
rect 24544 29804 24593 29832
rect 24544 29792 24550 29804
rect 24581 29801 24593 29804
rect 24627 29801 24639 29835
rect 24581 29795 24639 29801
rect 28074 29792 28080 29844
rect 28132 29832 28138 29844
rect 28132 29804 31754 29832
rect 28132 29792 28138 29804
rect 22922 29724 22928 29776
rect 22980 29764 22986 29776
rect 22980 29736 23428 29764
rect 22980 29724 22986 29736
rect 22848 29668 22922 29696
rect 19760 29656 19766 29668
rect 18601 29631 18659 29637
rect 18601 29597 18613 29631
rect 18647 29597 18659 29631
rect 18601 29591 18659 29597
rect 18690 29588 18696 29640
rect 18748 29588 18754 29640
rect 18874 29588 18880 29640
rect 18932 29588 18938 29640
rect 20625 29631 20683 29637
rect 20625 29597 20637 29631
rect 20671 29628 20683 29631
rect 20806 29628 20812 29640
rect 20671 29600 20812 29628
rect 20671 29597 20683 29600
rect 20625 29591 20683 29597
rect 20806 29588 20812 29600
rect 20864 29588 20870 29640
rect 20901 29631 20959 29637
rect 20901 29597 20913 29631
rect 20947 29628 20959 29631
rect 20990 29628 20996 29640
rect 20947 29600 20996 29628
rect 20947 29597 20959 29600
rect 20901 29591 20959 29597
rect 20990 29588 20996 29600
rect 21048 29588 21054 29640
rect 22094 29628 22100 29640
rect 21468 29600 22100 29628
rect 17221 29563 17279 29569
rect 17221 29560 17233 29563
rect 16316 29532 17233 29560
rect 16117 29523 16175 29529
rect 17221 29529 17233 29532
rect 17267 29529 17279 29563
rect 17221 29523 17279 29529
rect 9030 29492 9036 29504
rect 8588 29464 9036 29492
rect 9030 29452 9036 29464
rect 9088 29492 9094 29504
rect 9950 29492 9956 29504
rect 9088 29464 9956 29492
rect 9088 29452 9094 29464
rect 9950 29452 9956 29464
rect 10008 29452 10014 29504
rect 10686 29452 10692 29504
rect 10744 29492 10750 29504
rect 13170 29492 13176 29504
rect 10744 29464 13176 29492
rect 10744 29452 10750 29464
rect 13170 29452 13176 29464
rect 13228 29452 13234 29504
rect 13262 29452 13268 29504
rect 13320 29452 13326 29504
rect 16758 29452 16764 29504
rect 16816 29492 16822 29504
rect 16945 29495 17003 29501
rect 16945 29492 16957 29495
rect 16816 29464 16957 29492
rect 16816 29452 16822 29464
rect 16945 29461 16957 29464
rect 16991 29461 17003 29495
rect 16945 29455 17003 29461
rect 17034 29452 17040 29504
rect 17092 29452 17098 29504
rect 17236 29492 17264 29523
rect 18506 29520 18512 29572
rect 18564 29520 18570 29572
rect 18892 29560 18920 29588
rect 21468 29560 21496 29600
rect 22094 29588 22100 29600
rect 22152 29588 22158 29640
rect 22894 29637 22922 29668
rect 23216 29668 23337 29696
rect 23216 29640 23244 29668
rect 22879 29631 22937 29637
rect 22879 29597 22891 29631
rect 22925 29597 22937 29631
rect 22879 29591 22937 29597
rect 23198 29588 23204 29640
rect 23256 29588 23262 29640
rect 23309 29637 23337 29668
rect 23400 29637 23428 29736
rect 24394 29724 24400 29776
rect 24452 29764 24458 29776
rect 24762 29764 24768 29776
rect 24452 29736 24768 29764
rect 24452 29724 24458 29736
rect 24762 29724 24768 29736
rect 24820 29764 24826 29776
rect 26510 29764 26516 29776
rect 24820 29736 26516 29764
rect 24820 29724 24826 29736
rect 23474 29656 23480 29708
rect 23532 29696 23538 29708
rect 23532 29668 23796 29696
rect 23532 29656 23538 29668
rect 23768 29640 23796 29668
rect 23292 29631 23350 29637
rect 23292 29597 23304 29631
rect 23338 29597 23350 29631
rect 23292 29591 23350 29597
rect 23385 29631 23443 29637
rect 23385 29597 23397 29631
rect 23431 29597 23443 29631
rect 23385 29591 23443 29597
rect 23750 29588 23756 29640
rect 23808 29588 23814 29640
rect 24026 29588 24032 29640
rect 24084 29588 24090 29640
rect 24578 29588 24584 29640
rect 24636 29628 24642 29640
rect 24673 29631 24731 29637
rect 24673 29628 24685 29631
rect 24636 29600 24685 29628
rect 24636 29588 24642 29600
rect 24673 29597 24685 29600
rect 24719 29597 24731 29631
rect 24673 29591 24731 29597
rect 24762 29588 24768 29640
rect 24820 29588 24826 29640
rect 24854 29588 24860 29640
rect 24912 29628 24918 29640
rect 25774 29637 25780 29640
rect 25757 29631 25780 29637
rect 25757 29628 25769 29631
rect 24912 29600 25769 29628
rect 24912 29588 24918 29600
rect 25757 29597 25769 29600
rect 25757 29591 25780 29597
rect 25774 29588 25780 29591
rect 25832 29588 25838 29640
rect 25884 29637 25912 29736
rect 26510 29724 26516 29736
rect 26568 29724 26574 29776
rect 26602 29724 26608 29776
rect 26660 29764 26666 29776
rect 26660 29736 26832 29764
rect 26660 29724 26666 29736
rect 26326 29656 26332 29708
rect 26384 29696 26390 29708
rect 26384 29668 26740 29696
rect 26384 29656 26390 29668
rect 25869 29631 25927 29637
rect 25869 29597 25881 29631
rect 25915 29597 25927 29631
rect 25869 29591 25927 29597
rect 25961 29631 26019 29637
rect 25961 29597 25973 29631
rect 26007 29597 26019 29631
rect 25961 29591 26019 29597
rect 18892 29532 21496 29560
rect 21542 29520 21548 29572
rect 21600 29560 21606 29572
rect 22997 29563 23055 29569
rect 22997 29560 23009 29563
rect 21600 29532 23009 29560
rect 21600 29520 21606 29532
rect 22997 29529 23009 29532
rect 23043 29529 23055 29563
rect 22997 29523 23055 29529
rect 23106 29520 23112 29572
rect 23164 29520 23170 29572
rect 25976 29560 26004 29591
rect 26050 29588 26056 29640
rect 26108 29628 26114 29640
rect 26145 29631 26203 29637
rect 26145 29628 26157 29631
rect 26108 29600 26157 29628
rect 26108 29588 26114 29600
rect 26145 29597 26157 29600
rect 26191 29628 26203 29631
rect 26191 29600 26372 29628
rect 26191 29597 26203 29600
rect 26145 29591 26203 29597
rect 26344 29572 26372 29600
rect 26418 29588 26424 29640
rect 26476 29588 26482 29640
rect 26712 29637 26740 29668
rect 26804 29637 26832 29736
rect 26878 29724 26884 29776
rect 26936 29764 26942 29776
rect 28902 29764 28908 29776
rect 26936 29736 28908 29764
rect 26936 29724 26942 29736
rect 27448 29637 27476 29736
rect 28902 29724 28908 29736
rect 28960 29724 28966 29776
rect 29086 29724 29092 29776
rect 29144 29764 29150 29776
rect 29144 29736 30512 29764
rect 29144 29724 29150 29736
rect 27614 29656 27620 29708
rect 27672 29656 27678 29708
rect 28994 29696 29000 29708
rect 27816 29668 29000 29696
rect 27816 29637 27844 29668
rect 28994 29656 29000 29668
rect 29052 29696 29058 29708
rect 29052 29668 30420 29696
rect 29052 29656 29058 29668
rect 26513 29631 26571 29637
rect 26513 29597 26525 29631
rect 26559 29597 26571 29631
rect 26513 29591 26571 29597
rect 26697 29631 26755 29637
rect 26697 29597 26709 29631
rect 26743 29597 26755 29631
rect 26697 29591 26755 29597
rect 26789 29631 26847 29637
rect 26789 29597 26801 29631
rect 26835 29597 26847 29631
rect 26789 29591 26847 29597
rect 27433 29631 27491 29637
rect 27433 29597 27445 29631
rect 27479 29597 27491 29631
rect 27433 29591 27491 29597
rect 27801 29631 27859 29637
rect 27801 29597 27813 29631
rect 27847 29597 27859 29631
rect 28537 29631 28595 29637
rect 28537 29628 28549 29631
rect 27801 29591 27859 29597
rect 28276 29600 28549 29628
rect 26237 29563 26295 29569
rect 26237 29560 26249 29563
rect 23308 29532 25912 29560
rect 25976 29532 26249 29560
rect 18414 29492 18420 29504
rect 17236 29464 18420 29492
rect 18414 29452 18420 29464
rect 18472 29452 18478 29504
rect 18874 29452 18880 29504
rect 18932 29452 18938 29504
rect 19058 29452 19064 29504
rect 19116 29492 19122 29504
rect 20714 29492 20720 29504
rect 19116 29464 20720 29492
rect 19116 29452 19122 29464
rect 20714 29452 20720 29464
rect 20772 29492 20778 29504
rect 20809 29495 20867 29501
rect 20809 29492 20821 29495
rect 20772 29464 20821 29492
rect 20772 29452 20778 29464
rect 20809 29461 20821 29464
rect 20855 29461 20867 29495
rect 20809 29455 20867 29461
rect 20993 29495 21051 29501
rect 20993 29461 21005 29495
rect 21039 29492 21051 29495
rect 21082 29492 21088 29504
rect 21039 29464 21088 29492
rect 21039 29461 21051 29464
rect 20993 29455 21051 29461
rect 21082 29452 21088 29464
rect 21140 29452 21146 29504
rect 21174 29452 21180 29504
rect 21232 29452 21238 29504
rect 22738 29452 22744 29504
rect 22796 29452 22802 29504
rect 22830 29452 22836 29504
rect 22888 29492 22894 29504
rect 23129 29492 23157 29520
rect 23308 29504 23336 29532
rect 22888 29464 23157 29492
rect 22888 29452 22894 29464
rect 23290 29452 23296 29504
rect 23348 29452 23354 29504
rect 23566 29452 23572 29504
rect 23624 29452 23630 29504
rect 23937 29495 23995 29501
rect 23937 29461 23949 29495
rect 23983 29492 23995 29495
rect 24397 29495 24455 29501
rect 24397 29492 24409 29495
rect 23983 29464 24409 29492
rect 23983 29461 23995 29464
rect 23937 29455 23995 29461
rect 24397 29461 24409 29464
rect 24443 29461 24455 29495
rect 24397 29455 24455 29461
rect 25406 29452 25412 29504
rect 25464 29492 25470 29504
rect 25501 29495 25559 29501
rect 25501 29492 25513 29495
rect 25464 29464 25513 29492
rect 25464 29452 25470 29464
rect 25501 29461 25513 29464
rect 25547 29461 25559 29495
rect 25884 29492 25912 29532
rect 26237 29529 26249 29532
rect 26283 29529 26295 29563
rect 26237 29523 26295 29529
rect 26326 29520 26332 29572
rect 26384 29520 26390 29572
rect 26528 29560 26556 29591
rect 27816 29560 27844 29591
rect 26528 29532 27844 29560
rect 26528 29492 26556 29532
rect 25884 29464 26556 29492
rect 25501 29455 25559 29461
rect 27338 29452 27344 29504
rect 27396 29452 27402 29504
rect 27614 29452 27620 29504
rect 27672 29492 27678 29504
rect 27798 29492 27804 29504
rect 27672 29464 27804 29492
rect 27672 29452 27678 29464
rect 27798 29452 27804 29464
rect 27856 29452 27862 29504
rect 27893 29495 27951 29501
rect 27893 29461 27905 29495
rect 27939 29492 27951 29495
rect 28074 29492 28080 29504
rect 27939 29464 28080 29492
rect 27939 29461 27951 29464
rect 27893 29455 27951 29461
rect 28074 29452 28080 29464
rect 28132 29452 28138 29504
rect 28276 29501 28304 29600
rect 28537 29597 28549 29600
rect 28583 29597 28595 29631
rect 28537 29591 28595 29597
rect 28902 29588 28908 29640
rect 28960 29628 28966 29640
rect 29365 29631 29423 29637
rect 29365 29628 29377 29631
rect 28960 29600 29377 29628
rect 28960 29588 28966 29600
rect 29365 29597 29377 29600
rect 29411 29597 29423 29631
rect 29365 29591 29423 29597
rect 29822 29588 29828 29640
rect 29880 29588 29886 29640
rect 29917 29631 29975 29637
rect 29917 29597 29929 29631
rect 29963 29597 29975 29631
rect 29917 29591 29975 29597
rect 28442 29520 28448 29572
rect 28500 29560 28506 29572
rect 29840 29560 29868 29588
rect 28500 29532 29868 29560
rect 29932 29560 29960 29591
rect 30006 29588 30012 29640
rect 30064 29588 30070 29640
rect 30392 29637 30420 29668
rect 30193 29631 30251 29637
rect 30193 29597 30205 29631
rect 30239 29597 30251 29631
rect 30193 29591 30251 29597
rect 30285 29631 30343 29637
rect 30285 29597 30297 29631
rect 30331 29597 30343 29631
rect 30285 29591 30343 29597
rect 30378 29631 30436 29637
rect 30378 29597 30390 29631
rect 30424 29597 30436 29631
rect 30378 29591 30436 29597
rect 30098 29560 30104 29572
rect 29932 29532 30104 29560
rect 28500 29520 28506 29532
rect 30098 29520 30104 29532
rect 30156 29520 30162 29572
rect 28261 29495 28319 29501
rect 28261 29461 28273 29495
rect 28307 29461 28319 29495
rect 28261 29455 28319 29461
rect 28350 29452 28356 29504
rect 28408 29452 28414 29504
rect 29270 29452 29276 29504
rect 29328 29452 29334 29504
rect 29362 29452 29368 29504
rect 29420 29492 29426 29504
rect 29549 29495 29607 29501
rect 29549 29492 29561 29495
rect 29420 29464 29561 29492
rect 29420 29452 29426 29464
rect 29549 29461 29561 29464
rect 29595 29461 29607 29495
rect 30208 29492 30236 29591
rect 30300 29560 30328 29591
rect 30484 29560 30512 29736
rect 30650 29588 30656 29640
rect 30708 29588 30714 29640
rect 30834 29637 30840 29640
rect 30791 29631 30840 29637
rect 30791 29597 30803 29631
rect 30837 29597 30840 29631
rect 30791 29591 30840 29597
rect 30834 29588 30840 29591
rect 30892 29588 30898 29640
rect 31205 29631 31263 29637
rect 31205 29597 31217 29631
rect 31251 29628 31263 29631
rect 31294 29628 31300 29640
rect 31251 29600 31300 29628
rect 31251 29597 31263 29600
rect 31205 29591 31263 29597
rect 31294 29588 31300 29600
rect 31352 29588 31358 29640
rect 30300 29532 30512 29560
rect 30392 29504 30420 29532
rect 30558 29520 30564 29572
rect 30616 29520 30622 29572
rect 30282 29492 30288 29504
rect 30208 29464 30288 29492
rect 29549 29455 29607 29461
rect 30282 29452 30288 29464
rect 30340 29452 30346 29504
rect 30374 29452 30380 29504
rect 30432 29452 30438 29504
rect 30929 29495 30987 29501
rect 30929 29461 30941 29495
rect 30975 29492 30987 29495
rect 31294 29492 31300 29504
rect 30975 29464 31300 29492
rect 30975 29461 30987 29464
rect 30929 29455 30987 29461
rect 31294 29452 31300 29464
rect 31352 29452 31358 29504
rect 31726 29492 31754 29804
rect 33502 29724 33508 29776
rect 33560 29764 33566 29776
rect 34238 29764 34244 29776
rect 33560 29736 34244 29764
rect 33560 29724 33566 29736
rect 33980 29705 34008 29736
rect 34238 29724 34244 29736
rect 34296 29724 34302 29776
rect 33965 29699 34023 29705
rect 33965 29665 33977 29699
rect 34011 29665 34023 29699
rect 36817 29699 36875 29705
rect 36817 29696 36829 29699
rect 33965 29659 34023 29665
rect 34164 29668 36829 29696
rect 34164 29640 34192 29668
rect 36817 29665 36829 29668
rect 36863 29665 36875 29699
rect 36817 29659 36875 29665
rect 34146 29588 34152 29640
rect 34204 29588 34210 29640
rect 34790 29588 34796 29640
rect 34848 29588 34854 29640
rect 32953 29563 33011 29569
rect 32953 29529 32965 29563
rect 32999 29560 33011 29563
rect 34330 29560 34336 29572
rect 32999 29532 34336 29560
rect 32999 29529 33011 29532
rect 32953 29523 33011 29529
rect 34330 29520 34336 29532
rect 34388 29520 34394 29572
rect 34974 29520 34980 29572
rect 35032 29560 35038 29572
rect 35069 29563 35127 29569
rect 35069 29560 35081 29563
rect 35032 29532 35081 29560
rect 35032 29520 35038 29532
rect 35069 29529 35081 29532
rect 35115 29529 35127 29563
rect 35069 29523 35127 29529
rect 33318 29492 33324 29504
rect 31726 29464 33324 29492
rect 33318 29452 33324 29464
rect 33376 29492 33382 29504
rect 34057 29495 34115 29501
rect 34057 29492 34069 29495
rect 33376 29464 34069 29492
rect 33376 29452 33382 29464
rect 34057 29461 34069 29464
rect 34103 29461 34115 29495
rect 34057 29455 34115 29461
rect 34514 29452 34520 29504
rect 34572 29452 34578 29504
rect 35986 29452 35992 29504
rect 36044 29492 36050 29504
rect 36188 29492 36216 29614
rect 36044 29464 36216 29492
rect 36044 29452 36050 29464
rect 1104 29402 38272 29424
rect 1104 29350 4874 29402
rect 4926 29350 4938 29402
rect 4990 29350 5002 29402
rect 5054 29350 5066 29402
rect 5118 29350 5130 29402
rect 5182 29350 35594 29402
rect 35646 29350 35658 29402
rect 35710 29350 35722 29402
rect 35774 29350 35786 29402
rect 35838 29350 35850 29402
rect 35902 29350 38272 29402
rect 1104 29328 38272 29350
rect 4062 29248 4068 29300
rect 4120 29248 4126 29300
rect 5902 29248 5908 29300
rect 5960 29248 5966 29300
rect 7466 29288 7472 29300
rect 6932 29260 7472 29288
rect 4080 29220 4108 29248
rect 3896 29192 4108 29220
rect 3896 29161 3924 29192
rect 3881 29155 3939 29161
rect 3881 29121 3893 29155
rect 3927 29121 3939 29155
rect 3881 29115 3939 29121
rect 5258 29112 5264 29164
rect 5316 29152 5322 29164
rect 5920 29161 5948 29248
rect 6932 29161 6960 29260
rect 7466 29248 7472 29260
rect 7524 29248 7530 29300
rect 7558 29248 7564 29300
rect 7616 29288 7622 29300
rect 9861 29291 9919 29297
rect 9861 29288 9873 29291
rect 7616 29260 9873 29288
rect 7616 29248 7622 29260
rect 9861 29257 9873 29260
rect 9907 29257 9919 29291
rect 9861 29251 9919 29257
rect 14826 29248 14832 29300
rect 14884 29288 14890 29300
rect 14884 29260 18644 29288
rect 14884 29248 14890 29260
rect 7101 29223 7159 29229
rect 7101 29189 7113 29223
rect 7147 29220 7159 29223
rect 7926 29220 7932 29232
rect 7147 29192 7932 29220
rect 7147 29189 7159 29192
rect 7101 29183 7159 29189
rect 7926 29180 7932 29192
rect 7984 29180 7990 29232
rect 9125 29223 9183 29229
rect 9125 29189 9137 29223
rect 9171 29220 9183 29223
rect 10686 29220 10692 29232
rect 9171 29192 10692 29220
rect 9171 29189 9183 29192
rect 9125 29183 9183 29189
rect 10686 29180 10692 29192
rect 10744 29180 10750 29232
rect 11333 29223 11391 29229
rect 11333 29189 11345 29223
rect 11379 29220 11391 29223
rect 17954 29220 17960 29232
rect 11379 29192 17960 29220
rect 11379 29189 11391 29192
rect 11333 29183 11391 29189
rect 17954 29180 17960 29192
rect 18012 29180 18018 29232
rect 18616 29220 18644 29260
rect 18690 29248 18696 29300
rect 18748 29288 18754 29300
rect 18877 29291 18935 29297
rect 18877 29288 18889 29291
rect 18748 29260 18889 29288
rect 18748 29248 18754 29260
rect 18877 29257 18889 29260
rect 18923 29257 18935 29291
rect 21269 29291 21327 29297
rect 18877 29251 18935 29257
rect 19076 29260 19334 29288
rect 18966 29220 18972 29232
rect 18616 29192 18972 29220
rect 5905 29155 5963 29161
rect 5316 29124 5396 29152
rect 5316 29112 5322 29124
rect 5368 28960 5396 29124
rect 5905 29121 5917 29155
rect 5951 29121 5963 29155
rect 5905 29115 5963 29121
rect 6917 29155 6975 29161
rect 6917 29121 6929 29155
rect 6963 29121 6975 29155
rect 6917 29115 6975 29121
rect 7009 29155 7067 29161
rect 7009 29121 7021 29155
rect 7055 29121 7067 29155
rect 7009 29115 7067 29121
rect 7285 29155 7343 29161
rect 7285 29121 7297 29155
rect 7331 29152 7343 29155
rect 7653 29155 7711 29161
rect 7653 29152 7665 29155
rect 7331 29124 7665 29152
rect 7331 29121 7343 29124
rect 7285 29115 7343 29121
rect 7653 29121 7665 29124
rect 7699 29121 7711 29155
rect 7653 29115 7711 29121
rect 7760 29124 8432 29152
rect 6822 29044 6828 29096
rect 6880 29084 6886 29096
rect 7024 29084 7052 29115
rect 7760 29084 7788 29124
rect 6880 29056 7788 29084
rect 8205 29087 8263 29093
rect 6880 29044 6886 29056
rect 8205 29053 8217 29087
rect 8251 29053 8263 29087
rect 8205 29047 8263 29053
rect 4144 28951 4202 28957
rect 4144 28917 4156 28951
rect 4190 28948 4202 28951
rect 4706 28948 4712 28960
rect 4190 28920 4712 28948
rect 4190 28917 4202 28920
rect 4144 28911 4202 28917
rect 4706 28908 4712 28920
rect 4764 28908 4770 28960
rect 5350 28908 5356 28960
rect 5408 28908 5414 28960
rect 6546 28908 6552 28960
rect 6604 28948 6610 28960
rect 6733 28951 6791 28957
rect 6733 28948 6745 28951
rect 6604 28920 6745 28948
rect 6604 28908 6610 28920
rect 6733 28917 6745 28920
rect 6779 28917 6791 28951
rect 8220 28948 8248 29047
rect 8294 29044 8300 29096
rect 8352 29044 8358 29096
rect 8404 29084 8432 29124
rect 12710 29112 12716 29164
rect 12768 29152 12774 29164
rect 13081 29155 13139 29161
rect 13081 29152 13093 29155
rect 12768 29124 13093 29152
rect 12768 29112 12774 29124
rect 13081 29121 13093 29124
rect 13127 29121 13139 29155
rect 13081 29115 13139 29121
rect 13265 29155 13323 29161
rect 13265 29121 13277 29155
rect 13311 29152 13323 29155
rect 16114 29152 16120 29164
rect 13311 29124 16120 29152
rect 13311 29121 13323 29124
rect 13265 29115 13323 29121
rect 16114 29112 16120 29124
rect 16172 29112 16178 29164
rect 16850 29112 16856 29164
rect 16908 29152 16914 29164
rect 17402 29152 17408 29164
rect 16908 29124 17408 29152
rect 16908 29112 16914 29124
rect 17402 29112 17408 29124
rect 17460 29112 17466 29164
rect 18509 29155 18567 29161
rect 18509 29121 18521 29155
rect 18555 29152 18567 29155
rect 18598 29152 18604 29164
rect 18555 29124 18604 29152
rect 18555 29121 18567 29124
rect 18509 29115 18567 29121
rect 18598 29112 18604 29124
rect 18656 29112 18662 29164
rect 18708 29161 18736 29192
rect 18966 29180 18972 29192
rect 19024 29180 19030 29232
rect 18693 29155 18751 29161
rect 18693 29121 18705 29155
rect 18739 29121 18751 29155
rect 18693 29115 18751 29121
rect 9122 29084 9128 29096
rect 8404 29056 9128 29084
rect 9122 29044 9128 29056
rect 9180 29084 9186 29096
rect 9217 29087 9275 29093
rect 9217 29084 9229 29087
rect 9180 29056 9229 29084
rect 9180 29044 9186 29056
rect 9217 29053 9229 29056
rect 9263 29053 9275 29087
rect 9217 29047 9275 29053
rect 9401 29087 9459 29093
rect 9401 29053 9413 29087
rect 9447 29084 9459 29087
rect 10778 29084 10784 29096
rect 9447 29056 10784 29084
rect 9447 29053 9459 29056
rect 9401 29047 9459 29053
rect 10778 29044 10784 29056
rect 10836 29084 10842 29096
rect 10836 29056 11008 29084
rect 10836 29044 10842 29056
rect 8312 29016 8340 29044
rect 8757 29019 8815 29025
rect 8757 29016 8769 29019
rect 8312 28988 8769 29016
rect 8757 28985 8769 28988
rect 8803 28985 8815 29019
rect 8757 28979 8815 28985
rect 8294 28948 8300 28960
rect 8220 28920 8300 28948
rect 6733 28911 6791 28917
rect 8294 28908 8300 28920
rect 8352 28908 8358 28960
rect 10980 28948 11008 29056
rect 13722 29044 13728 29096
rect 13780 29084 13786 29096
rect 19076 29084 19104 29260
rect 19306 29220 19334 29260
rect 21269 29257 21281 29291
rect 21315 29288 21327 29291
rect 22462 29288 22468 29300
rect 21315 29260 22468 29288
rect 21315 29257 21327 29260
rect 21269 29251 21327 29257
rect 22462 29248 22468 29260
rect 22520 29248 22526 29300
rect 22554 29248 22560 29300
rect 22612 29248 22618 29300
rect 22738 29248 22744 29300
rect 22796 29248 22802 29300
rect 23198 29248 23204 29300
rect 23256 29288 23262 29300
rect 26418 29288 26424 29300
rect 23256 29260 25820 29288
rect 23256 29248 23262 29260
rect 21634 29220 21640 29232
rect 19306 29192 21640 29220
rect 19794 29152 19800 29164
rect 13780 29056 19104 29084
rect 19306 29124 19800 29152
rect 13780 29044 13786 29056
rect 12894 28976 12900 29028
rect 12952 28976 12958 29028
rect 13170 28976 13176 29028
rect 13228 29016 13234 29028
rect 19306 29016 19334 29124
rect 19794 29112 19800 29124
rect 19852 29152 19858 29164
rect 20717 29155 20775 29161
rect 20717 29152 20729 29155
rect 19852 29124 20729 29152
rect 19852 29112 19858 29124
rect 20717 29121 20729 29124
rect 20763 29152 20775 29155
rect 20806 29152 20812 29164
rect 20763 29124 20812 29152
rect 20763 29121 20775 29124
rect 20717 29115 20775 29121
rect 20806 29112 20812 29124
rect 20864 29112 20870 29164
rect 20898 29112 20904 29164
rect 20956 29112 20962 29164
rect 21100 29161 21128 29192
rect 21634 29180 21640 29192
rect 21692 29180 21698 29232
rect 22094 29180 22100 29232
rect 22152 29180 22158 29232
rect 20993 29155 21051 29161
rect 20993 29121 21005 29155
rect 21039 29121 21051 29155
rect 20993 29115 21051 29121
rect 21085 29155 21143 29161
rect 21085 29121 21097 29155
rect 21131 29121 21143 29155
rect 21085 29115 21143 29121
rect 21008 29084 21036 29115
rect 21174 29112 21180 29164
rect 21232 29152 21238 29164
rect 22002 29161 22008 29164
rect 21821 29155 21879 29161
rect 21821 29152 21833 29155
rect 21232 29124 21833 29152
rect 21232 29112 21238 29124
rect 21821 29121 21833 29124
rect 21867 29121 21879 29155
rect 21821 29115 21879 29121
rect 21969 29155 22008 29161
rect 21969 29121 21981 29155
rect 21969 29115 22008 29121
rect 22002 29112 22008 29115
rect 22060 29112 22066 29164
rect 22186 29112 22192 29164
rect 22244 29112 22250 29164
rect 22278 29112 22284 29164
rect 22336 29161 22342 29164
rect 22572 29161 22600 29248
rect 22336 29115 22344 29161
rect 22557 29155 22615 29161
rect 22557 29121 22569 29155
rect 22603 29121 22615 29155
rect 22756 29152 22784 29248
rect 22833 29155 22891 29161
rect 22833 29152 22845 29155
rect 22756 29124 22845 29152
rect 22557 29115 22615 29121
rect 22833 29121 22845 29124
rect 22879 29121 22891 29155
rect 22833 29115 22891 29121
rect 22336 29112 22342 29115
rect 23014 29112 23020 29164
rect 23072 29112 23078 29164
rect 23492 29161 23520 29260
rect 23658 29180 23664 29232
rect 23716 29180 23722 29232
rect 23753 29223 23811 29229
rect 23753 29189 23765 29223
rect 23799 29220 23811 29223
rect 24026 29220 24032 29232
rect 23799 29192 24032 29220
rect 23799 29189 23811 29192
rect 23753 29183 23811 29189
rect 24026 29180 24032 29192
rect 24084 29180 24090 29232
rect 23477 29155 23535 29161
rect 23477 29121 23489 29155
rect 23523 29121 23535 29155
rect 23477 29115 23535 29121
rect 23845 29155 23903 29161
rect 23845 29121 23857 29155
rect 23891 29152 23903 29155
rect 24210 29152 24216 29164
rect 23891 29124 24216 29152
rect 23891 29121 23903 29124
rect 23845 29115 23903 29121
rect 24210 29112 24216 29124
rect 24268 29112 24274 29164
rect 25501 29155 25559 29161
rect 25501 29121 25513 29155
rect 25547 29121 25559 29155
rect 25501 29115 25559 29121
rect 21542 29084 21548 29096
rect 13228 28988 19334 29016
rect 20088 29056 21548 29084
rect 13228 28976 13234 28988
rect 20088 28960 20116 29056
rect 21542 29044 21548 29056
rect 21600 29044 21606 29096
rect 22741 29087 22799 29093
rect 22741 29053 22753 29087
rect 22787 29084 22799 29087
rect 22787 29056 23428 29084
rect 22787 29053 22799 29056
rect 22741 29047 22799 29053
rect 22465 29019 22523 29025
rect 22465 28985 22477 29019
rect 22511 29016 22523 29019
rect 22925 29019 22983 29025
rect 22925 29016 22937 29019
rect 22511 28988 22937 29016
rect 22511 28985 22523 28988
rect 22465 28979 22523 28985
rect 22925 28985 22937 28988
rect 22971 28985 22983 29019
rect 22925 28979 22983 28985
rect 11514 28948 11520 28960
rect 10980 28920 11520 28948
rect 11514 28908 11520 28920
rect 11572 28908 11578 28960
rect 11606 28908 11612 28960
rect 11664 28948 11670 28960
rect 12618 28948 12624 28960
rect 11664 28920 12624 28948
rect 11664 28908 11670 28920
rect 12618 28908 12624 28920
rect 12676 28908 12682 28960
rect 14642 28908 14648 28960
rect 14700 28948 14706 28960
rect 18322 28948 18328 28960
rect 14700 28920 18328 28948
rect 14700 28908 14706 28920
rect 18322 28908 18328 28920
rect 18380 28908 18386 28960
rect 18598 28908 18604 28960
rect 18656 28948 18662 28960
rect 19150 28948 19156 28960
rect 18656 28920 19156 28948
rect 18656 28908 18662 28920
rect 19150 28908 19156 28920
rect 19208 28908 19214 28960
rect 19610 28908 19616 28960
rect 19668 28948 19674 28960
rect 19978 28948 19984 28960
rect 19668 28920 19984 28948
rect 19668 28908 19674 28920
rect 19978 28908 19984 28920
rect 20036 28908 20042 28960
rect 20070 28908 20076 28960
rect 20128 28908 20134 28960
rect 23198 28908 23204 28960
rect 23256 28908 23262 28960
rect 23400 28948 23428 29056
rect 23768 29056 24900 29084
rect 23768 29016 23796 29056
rect 24872 29028 24900 29056
rect 25038 29044 25044 29096
rect 25096 29084 25102 29096
rect 25516 29084 25544 29115
rect 25590 29112 25596 29164
rect 25648 29112 25654 29164
rect 25792 29161 25820 29260
rect 25884 29260 26424 29288
rect 25884 29161 25912 29260
rect 26418 29248 26424 29260
rect 26476 29248 26482 29300
rect 26510 29248 26516 29300
rect 26568 29248 26574 29300
rect 27338 29248 27344 29300
rect 27396 29248 27402 29300
rect 28350 29288 28356 29300
rect 27908 29260 28356 29288
rect 26053 29223 26111 29229
rect 26053 29189 26065 29223
rect 26099 29220 26111 29223
rect 26528 29220 26556 29248
rect 27356 29220 27384 29248
rect 26099 29192 26372 29220
rect 26099 29189 26111 29192
rect 26053 29183 26111 29189
rect 25777 29155 25835 29161
rect 25777 29121 25789 29155
rect 25823 29121 25835 29155
rect 25777 29115 25835 29121
rect 25869 29155 25927 29161
rect 25869 29121 25881 29155
rect 25915 29121 25927 29155
rect 25869 29115 25927 29121
rect 26145 29155 26203 29161
rect 26145 29121 26157 29155
rect 26191 29152 26203 29155
rect 26234 29152 26240 29164
rect 26191 29124 26240 29152
rect 26191 29121 26203 29124
rect 26145 29115 26203 29121
rect 25096 29056 25544 29084
rect 25792 29084 25820 29115
rect 26234 29112 26240 29124
rect 26292 29112 26298 29164
rect 26344 29161 26372 29192
rect 26436 29192 26556 29220
rect 27264 29192 27384 29220
rect 27525 29223 27583 29229
rect 26436 29161 26464 29192
rect 26329 29155 26387 29161
rect 26329 29121 26341 29155
rect 26375 29121 26387 29155
rect 26329 29115 26387 29121
rect 26421 29155 26479 29161
rect 26421 29121 26433 29155
rect 26467 29121 26479 29155
rect 26421 29115 26479 29121
rect 26510 29112 26516 29164
rect 26568 29112 26574 29164
rect 27264 29161 27292 29192
rect 27525 29189 27537 29223
rect 27571 29220 27583 29223
rect 27908 29220 27936 29260
rect 28350 29248 28356 29260
rect 28408 29248 28414 29300
rect 28994 29248 29000 29300
rect 29052 29248 29058 29300
rect 29270 29248 29276 29300
rect 29328 29248 29334 29300
rect 29822 29248 29828 29300
rect 29880 29288 29886 29300
rect 30282 29288 30288 29300
rect 29880 29260 30288 29288
rect 29880 29248 29886 29260
rect 30282 29248 30288 29260
rect 30340 29288 30346 29300
rect 30340 29260 31248 29288
rect 30340 29248 30346 29260
rect 29288 29220 29316 29248
rect 31110 29220 31116 29232
rect 27571 29192 27936 29220
rect 29196 29192 29316 29220
rect 30682 29192 31116 29220
rect 27571 29189 27583 29192
rect 27525 29183 27583 29189
rect 27249 29155 27307 29161
rect 27249 29121 27261 29155
rect 27295 29121 27307 29155
rect 27249 29115 27307 29121
rect 28626 29112 28632 29164
rect 28684 29112 28690 29164
rect 29196 29161 29224 29192
rect 31110 29180 31116 29192
rect 31168 29180 31174 29232
rect 29181 29155 29239 29161
rect 29181 29121 29193 29155
rect 29227 29121 29239 29155
rect 29181 29115 29239 29121
rect 30006 29084 30012 29096
rect 25792 29056 30012 29084
rect 25096 29044 25102 29056
rect 30006 29044 30012 29056
rect 30064 29084 30070 29096
rect 30929 29087 30987 29093
rect 30929 29084 30941 29087
rect 30064 29056 30941 29084
rect 30064 29044 30070 29056
rect 30929 29053 30941 29056
rect 30975 29053 30987 29087
rect 31220 29084 31248 29260
rect 31294 29248 31300 29300
rect 31352 29288 31358 29300
rect 31352 29260 31754 29288
rect 31352 29248 31358 29260
rect 31478 29180 31484 29232
rect 31536 29180 31542 29232
rect 31570 29180 31576 29232
rect 31628 29180 31634 29232
rect 31726 29220 31754 29260
rect 32306 29248 32312 29300
rect 32364 29248 32370 29300
rect 32490 29248 32496 29300
rect 32548 29288 32554 29300
rect 34146 29288 34152 29300
rect 32548 29260 34152 29288
rect 32548 29248 32554 29260
rect 34146 29248 34152 29260
rect 34204 29248 34210 29300
rect 34790 29248 34796 29300
rect 34848 29288 34854 29300
rect 34977 29291 35035 29297
rect 34977 29288 34989 29291
rect 34848 29260 34989 29288
rect 34848 29248 34854 29260
rect 34977 29257 34989 29260
rect 35023 29257 35035 29291
rect 34977 29251 35035 29257
rect 31726 29192 31800 29220
rect 31484 29177 31542 29180
rect 31484 29143 31496 29177
rect 31530 29143 31542 29177
rect 31772 29161 31800 29192
rect 32324 29161 32352 29248
rect 32508 29183 32536 29248
rect 32494 29177 32552 29183
rect 33226 29180 33232 29232
rect 33284 29180 33290 29232
rect 34330 29180 34336 29232
rect 34388 29220 34394 29232
rect 34388 29192 35112 29220
rect 34388 29180 34394 29192
rect 31484 29137 31542 29143
rect 31757 29155 31815 29161
rect 31757 29121 31769 29155
rect 31803 29121 31815 29155
rect 31757 29115 31815 29121
rect 31941 29155 31999 29161
rect 31941 29121 31953 29155
rect 31987 29152 31999 29155
rect 32125 29155 32183 29161
rect 32125 29152 32137 29155
rect 31987 29124 32137 29152
rect 31987 29121 31999 29124
rect 31941 29115 31999 29121
rect 32125 29121 32137 29124
rect 32171 29121 32183 29155
rect 32125 29115 32183 29121
rect 32309 29155 32367 29161
rect 32309 29121 32321 29155
rect 32355 29121 32367 29155
rect 32309 29115 32367 29121
rect 32401 29155 32459 29161
rect 32401 29121 32413 29155
rect 32447 29121 32459 29155
rect 32494 29143 32506 29177
rect 32540 29143 32552 29177
rect 32494 29137 32552 29143
rect 32401 29115 32459 29121
rect 32324 29084 32352 29115
rect 31220 29056 32352 29084
rect 32416 29084 32444 29115
rect 33042 29112 33048 29164
rect 33100 29112 33106 29164
rect 33244 29084 33272 29180
rect 34514 29112 34520 29164
rect 34572 29152 34578 29164
rect 34609 29155 34667 29161
rect 34609 29152 34621 29155
rect 34572 29124 34621 29152
rect 34572 29112 34578 29124
rect 34609 29121 34621 29124
rect 34655 29121 34667 29155
rect 34609 29115 34667 29121
rect 34974 29112 34980 29164
rect 35032 29112 35038 29164
rect 35084 29161 35112 29192
rect 35069 29155 35127 29161
rect 35069 29121 35081 29155
rect 35115 29121 35127 29155
rect 35069 29115 35127 29121
rect 36630 29112 36636 29164
rect 36688 29112 36694 29164
rect 36814 29112 36820 29164
rect 36872 29112 36878 29164
rect 32416 29056 33272 29084
rect 30929 29047 30987 29053
rect 23584 28988 23796 29016
rect 24029 29019 24087 29025
rect 23584 28948 23612 28988
rect 24029 28985 24041 29019
rect 24075 29016 24087 29019
rect 24210 29016 24216 29028
rect 24075 28988 24216 29016
rect 24075 28985 24087 28988
rect 24029 28979 24087 28985
rect 24210 28976 24216 28988
rect 24268 28976 24274 29028
rect 24854 28976 24860 29028
rect 24912 29016 24918 29028
rect 26510 29016 26516 29028
rect 24912 28988 26516 29016
rect 24912 28976 24918 28988
rect 26510 28976 26516 28988
rect 26568 28976 26574 29028
rect 26789 29019 26847 29025
rect 26789 28985 26801 29019
rect 26835 29016 26847 29019
rect 27062 29016 27068 29028
rect 26835 28988 27068 29016
rect 26835 28985 26847 28988
rect 26789 28979 26847 28985
rect 27062 28976 27068 28988
rect 27120 28976 27126 29028
rect 29086 29016 29092 29028
rect 28920 28988 29092 29016
rect 23400 28920 23612 28948
rect 23934 28908 23940 28960
rect 23992 28948 23998 28960
rect 26970 28948 26976 28960
rect 23992 28920 26976 28948
rect 23992 28908 23998 28920
rect 26970 28908 26976 28920
rect 27028 28948 27034 28960
rect 28920 28948 28948 28988
rect 29086 28976 29092 28988
rect 29144 28976 29150 29028
rect 31662 29016 31668 29028
rect 30484 28988 31668 29016
rect 27028 28920 28948 28948
rect 27028 28908 27034 28920
rect 29270 28908 29276 28960
rect 29328 28948 29334 28960
rect 29444 28951 29502 28957
rect 29444 28948 29456 28951
rect 29328 28920 29456 28948
rect 29328 28908 29334 28920
rect 29444 28917 29456 28920
rect 29490 28917 29502 28951
rect 29444 28911 29502 28917
rect 30098 28908 30104 28960
rect 30156 28948 30162 28960
rect 30484 28948 30512 28988
rect 31662 28976 31668 28988
rect 31720 29016 31726 29028
rect 32416 29016 32444 29056
rect 31720 28988 32444 29016
rect 32769 29019 32827 29025
rect 31720 28976 31726 28988
rect 32769 28985 32781 29019
rect 32815 29016 32827 29019
rect 34698 29016 34704 29028
rect 32815 28988 34704 29016
rect 32815 28985 32827 28988
rect 32769 28979 32827 28985
rect 34698 28976 34704 28988
rect 34756 28976 34762 29028
rect 34793 29019 34851 29025
rect 34793 28985 34805 29019
rect 34839 29016 34851 29019
rect 34992 29016 35020 29112
rect 34839 28988 35020 29016
rect 37001 29019 37059 29025
rect 34839 28985 34851 28988
rect 34793 28979 34851 28985
rect 37001 28985 37013 29019
rect 37047 29016 37059 29019
rect 37274 29016 37280 29028
rect 37047 28988 37280 29016
rect 37047 28985 37059 28988
rect 37001 28979 37059 28985
rect 37274 28976 37280 28988
rect 37332 28976 37338 29028
rect 30156 28920 30512 28948
rect 30156 28908 30162 28920
rect 32398 28908 32404 28960
rect 32456 28948 32462 28960
rect 32861 28951 32919 28957
rect 32861 28948 32873 28951
rect 32456 28920 32873 28948
rect 32456 28908 32462 28920
rect 32861 28917 32873 28920
rect 32907 28917 32919 28951
rect 32861 28911 32919 28917
rect 1104 28858 38272 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 38272 28858
rect 1104 28784 38272 28806
rect 4525 28747 4583 28753
rect 4525 28713 4537 28747
rect 4571 28744 4583 28747
rect 4706 28744 4712 28756
rect 4571 28716 4712 28744
rect 4571 28713 4583 28716
rect 4525 28707 4583 28713
rect 4706 28704 4712 28716
rect 4764 28704 4770 28756
rect 8018 28704 8024 28756
rect 8076 28744 8082 28756
rect 14642 28744 14648 28756
rect 8076 28716 14648 28744
rect 8076 28704 8082 28716
rect 14642 28704 14648 28716
rect 14700 28704 14706 28756
rect 20254 28744 20260 28756
rect 18156 28716 20260 28744
rect 7929 28679 7987 28685
rect 7929 28645 7941 28679
rect 7975 28676 7987 28679
rect 8294 28676 8300 28688
rect 7975 28648 8300 28676
rect 7975 28645 7987 28648
rect 7929 28639 7987 28645
rect 8294 28636 8300 28648
rect 8352 28676 8358 28688
rect 9490 28676 9496 28688
rect 8352 28648 9496 28676
rect 8352 28636 8358 28648
rect 9490 28636 9496 28648
rect 9548 28636 9554 28688
rect 11514 28636 11520 28688
rect 11572 28676 11578 28688
rect 12066 28676 12072 28688
rect 11572 28648 12072 28676
rect 11572 28636 11578 28648
rect 12066 28636 12072 28648
rect 12124 28636 12130 28688
rect 18156 28676 18184 28716
rect 20254 28704 20260 28716
rect 20312 28704 20318 28756
rect 21542 28704 21548 28756
rect 21600 28744 21606 28756
rect 23566 28744 23572 28756
rect 21600 28716 23572 28744
rect 21600 28704 21606 28716
rect 23566 28704 23572 28716
rect 23624 28704 23630 28756
rect 24302 28704 24308 28756
rect 24360 28744 24366 28756
rect 24762 28744 24768 28756
rect 24360 28716 24768 28744
rect 24360 28704 24366 28716
rect 24762 28704 24768 28716
rect 24820 28704 24826 28756
rect 25590 28704 25596 28756
rect 25648 28744 25654 28756
rect 25777 28747 25835 28753
rect 25777 28744 25789 28747
rect 25648 28716 25789 28744
rect 25648 28704 25654 28716
rect 25777 28713 25789 28716
rect 25823 28713 25835 28747
rect 29086 28744 29092 28756
rect 25777 28707 25835 28713
rect 26068 28716 29092 28744
rect 14476 28648 18184 28676
rect 5997 28611 6055 28617
rect 5997 28577 6009 28611
rect 6043 28608 6055 28611
rect 6181 28611 6239 28617
rect 6181 28608 6193 28611
rect 6043 28580 6193 28608
rect 6043 28577 6055 28580
rect 5997 28571 6055 28577
rect 6181 28577 6193 28580
rect 6227 28577 6239 28611
rect 6181 28571 6239 28577
rect 6457 28611 6515 28617
rect 6457 28577 6469 28611
rect 6503 28608 6515 28611
rect 6546 28608 6552 28620
rect 6503 28580 6552 28608
rect 6503 28577 6515 28580
rect 6457 28571 6515 28577
rect 6546 28568 6552 28580
rect 6604 28568 6610 28620
rect 14476 28608 14504 28648
rect 19334 28636 19340 28688
rect 19392 28676 19398 28688
rect 20070 28676 20076 28688
rect 19392 28648 20076 28676
rect 19392 28636 19398 28648
rect 20070 28636 20076 28648
rect 20128 28636 20134 28688
rect 22002 28636 22008 28688
rect 22060 28676 22066 28688
rect 26068 28676 26096 28716
rect 29086 28704 29092 28716
rect 29144 28704 29150 28756
rect 31404 28716 34100 28744
rect 22060 28636 22094 28676
rect 8312 28580 14504 28608
rect 16132 28580 18000 28608
rect 4341 28543 4399 28549
rect 4341 28509 4353 28543
rect 4387 28509 4399 28543
rect 4341 28503 4399 28509
rect 4709 28543 4767 28549
rect 4709 28509 4721 28543
rect 4755 28540 4767 28543
rect 5442 28540 5448 28552
rect 4755 28512 5448 28540
rect 4755 28509 4767 28512
rect 4709 28503 4767 28509
rect 4356 28472 4384 28503
rect 5442 28500 5448 28512
rect 5500 28500 5506 28552
rect 5626 28500 5632 28552
rect 5684 28500 5690 28552
rect 8312 28549 8340 28580
rect 16132 28552 16160 28580
rect 6089 28543 6147 28549
rect 6089 28509 6101 28543
rect 6135 28509 6147 28543
rect 6089 28503 6147 28509
rect 8297 28543 8355 28549
rect 8297 28509 8309 28543
rect 8343 28509 8355 28543
rect 8297 28503 8355 28509
rect 5644 28472 5672 28500
rect 4356 28444 5672 28472
rect 4246 28364 4252 28416
rect 4304 28364 4310 28416
rect 6104 28404 6132 28503
rect 7190 28432 7196 28484
rect 7248 28432 7254 28484
rect 8110 28472 8116 28484
rect 7760 28444 8116 28472
rect 7760 28404 7788 28444
rect 8110 28432 8116 28444
rect 8168 28472 8174 28484
rect 8312 28472 8340 28503
rect 9950 28500 9956 28552
rect 10008 28500 10014 28552
rect 10045 28543 10103 28549
rect 10045 28509 10057 28543
rect 10091 28540 10103 28543
rect 10229 28543 10287 28549
rect 10229 28540 10241 28543
rect 10091 28512 10241 28540
rect 10091 28509 10103 28512
rect 10045 28503 10103 28509
rect 10229 28509 10241 28512
rect 10275 28509 10287 28543
rect 10229 28503 10287 28509
rect 16114 28500 16120 28552
rect 16172 28500 16178 28552
rect 16206 28500 16212 28552
rect 16264 28540 16270 28552
rect 16301 28543 16359 28549
rect 16301 28540 16313 28543
rect 16264 28512 16313 28540
rect 16264 28500 16270 28512
rect 16301 28509 16313 28512
rect 16347 28509 16359 28543
rect 16301 28503 16359 28509
rect 16482 28500 16488 28552
rect 16540 28500 16546 28552
rect 17862 28500 17868 28552
rect 17920 28500 17926 28552
rect 17972 28540 18000 28580
rect 18322 28568 18328 28620
rect 18380 28608 18386 28620
rect 19610 28608 19616 28620
rect 18380 28580 19616 28608
rect 18380 28568 18386 28580
rect 19610 28568 19616 28580
rect 19668 28568 19674 28620
rect 19720 28580 20024 28608
rect 18046 28540 18052 28552
rect 17972 28512 18052 28540
rect 18046 28500 18052 28512
rect 18104 28500 18110 28552
rect 19720 28549 19748 28580
rect 19705 28543 19763 28549
rect 19705 28540 19717 28543
rect 19536 28512 19717 28540
rect 8168 28444 8340 28472
rect 9968 28472 9996 28500
rect 10410 28472 10416 28484
rect 9968 28444 10416 28472
rect 8168 28432 8174 28444
rect 10410 28432 10416 28444
rect 10468 28432 10474 28484
rect 10502 28432 10508 28484
rect 10560 28432 10566 28484
rect 11054 28432 11060 28484
rect 11112 28432 11118 28484
rect 16393 28475 16451 28481
rect 16393 28441 16405 28475
rect 16439 28472 16451 28475
rect 16574 28472 16580 28484
rect 16439 28444 16580 28472
rect 16439 28441 16451 28444
rect 16393 28435 16451 28441
rect 16574 28432 16580 28444
rect 16632 28432 16638 28484
rect 17880 28472 17908 28500
rect 19536 28472 19564 28512
rect 19705 28509 19717 28512
rect 19751 28509 19763 28543
rect 19705 28503 19763 28509
rect 19794 28500 19800 28552
rect 19852 28500 19858 28552
rect 17880 28444 19564 28472
rect 19610 28432 19616 28484
rect 19668 28472 19674 28484
rect 19889 28475 19947 28481
rect 19889 28472 19901 28475
rect 19668 28444 19901 28472
rect 19668 28432 19674 28444
rect 19889 28441 19901 28444
rect 19935 28441 19947 28475
rect 19996 28472 20024 28580
rect 20088 28549 20116 28636
rect 20073 28543 20131 28549
rect 20073 28509 20085 28543
rect 20119 28509 20131 28543
rect 20073 28503 20131 28509
rect 20162 28500 20168 28552
rect 20220 28540 20226 28552
rect 20809 28543 20867 28549
rect 20809 28540 20821 28543
rect 20220 28512 20821 28540
rect 20220 28500 20226 28512
rect 20809 28509 20821 28512
rect 20855 28509 20867 28543
rect 20809 28503 20867 28509
rect 20990 28500 20996 28552
rect 21048 28500 21054 28552
rect 21008 28472 21036 28500
rect 19996 28444 21036 28472
rect 22066 28472 22094 28636
rect 24688 28648 26096 28676
rect 24688 28552 24716 28648
rect 25314 28608 25320 28620
rect 24872 28580 25320 28608
rect 24872 28552 24900 28580
rect 25314 28568 25320 28580
rect 25372 28608 25378 28620
rect 25590 28608 25596 28620
rect 25372 28580 25596 28608
rect 25372 28568 25378 28580
rect 25590 28568 25596 28580
rect 25648 28608 25654 28620
rect 25648 28580 26004 28608
rect 25648 28568 25654 28580
rect 22557 28543 22615 28549
rect 22557 28509 22569 28543
rect 22603 28540 22615 28543
rect 22738 28540 22744 28552
rect 22603 28512 22744 28540
rect 22603 28509 22615 28512
rect 22557 28503 22615 28509
rect 22738 28500 22744 28512
rect 22796 28500 22802 28552
rect 24486 28500 24492 28552
rect 24544 28540 24550 28552
rect 24581 28543 24639 28549
rect 24581 28540 24593 28543
rect 24544 28512 24593 28540
rect 24544 28500 24550 28512
rect 24581 28509 24593 28512
rect 24627 28509 24639 28543
rect 24581 28503 24639 28509
rect 24670 28500 24676 28552
rect 24728 28500 24734 28552
rect 24854 28500 24860 28552
rect 24912 28500 24918 28552
rect 25976 28549 26004 28580
rect 26068 28549 26096 28648
rect 26344 28648 28994 28676
rect 26344 28549 26372 28648
rect 28966 28608 28994 28648
rect 29270 28636 29276 28688
rect 29328 28636 29334 28688
rect 29932 28648 30788 28676
rect 29932 28608 29960 28648
rect 28966 28580 29960 28608
rect 30006 28568 30012 28620
rect 30064 28568 30070 28620
rect 30193 28611 30251 28617
rect 30193 28577 30205 28611
rect 30239 28608 30251 28611
rect 30282 28608 30288 28620
rect 30239 28580 30288 28608
rect 30239 28577 30251 28580
rect 30193 28571 30251 28577
rect 30282 28568 30288 28580
rect 30340 28568 30346 28620
rect 24949 28543 25007 28549
rect 24949 28509 24961 28543
rect 24995 28540 25007 28543
rect 25961 28543 26019 28549
rect 24995 28512 25084 28540
rect 24995 28509 25007 28512
rect 24949 28503 25007 28509
rect 22066 28444 24716 28472
rect 19889 28435 19947 28441
rect 6104 28376 7788 28404
rect 8202 28364 8208 28416
rect 8260 28364 8266 28416
rect 11974 28364 11980 28416
rect 12032 28364 12038 28416
rect 16669 28407 16727 28413
rect 16669 28373 16681 28407
rect 16715 28404 16727 28407
rect 17218 28404 17224 28416
rect 16715 28376 17224 28404
rect 16715 28373 16727 28376
rect 16669 28367 16727 28373
rect 17218 28364 17224 28376
rect 17276 28364 17282 28416
rect 19426 28364 19432 28416
rect 19484 28404 19490 28416
rect 19521 28407 19579 28413
rect 19521 28404 19533 28407
rect 19484 28376 19533 28404
rect 19484 28364 19490 28376
rect 19521 28373 19533 28376
rect 19567 28373 19579 28407
rect 19521 28367 19579 28373
rect 22370 28364 22376 28416
rect 22428 28404 22434 28416
rect 23934 28404 23940 28416
rect 22428 28376 23940 28404
rect 22428 28364 22434 28376
rect 23934 28364 23940 28376
rect 23992 28364 23998 28416
rect 24394 28364 24400 28416
rect 24452 28364 24458 28416
rect 24688 28404 24716 28444
rect 24762 28432 24768 28484
rect 24820 28432 24826 28484
rect 25056 28404 25084 28512
rect 25961 28509 25973 28543
rect 26007 28509 26019 28543
rect 25961 28503 26019 28509
rect 26053 28543 26111 28549
rect 26053 28509 26065 28543
rect 26099 28509 26111 28543
rect 26053 28503 26111 28509
rect 26329 28543 26387 28549
rect 26329 28509 26341 28543
rect 26375 28509 26387 28543
rect 26329 28503 26387 28509
rect 29089 28543 29147 28549
rect 29089 28509 29101 28543
rect 29135 28540 29147 28543
rect 29135 28512 29592 28540
rect 29135 28509 29147 28512
rect 29089 28503 29147 28509
rect 26142 28432 26148 28484
rect 26200 28432 26206 28484
rect 26344 28404 26372 28503
rect 29564 28413 29592 28512
rect 30024 28472 30052 28568
rect 30760 28552 30788 28648
rect 31404 28552 31432 28716
rect 31478 28636 31484 28688
rect 31536 28636 31542 28688
rect 30374 28500 30380 28552
rect 30432 28500 30438 28552
rect 30470 28543 30528 28549
rect 30470 28509 30482 28543
rect 30516 28509 30528 28543
rect 30470 28503 30528 28509
rect 30484 28472 30512 28503
rect 30558 28500 30564 28552
rect 30616 28500 30622 28552
rect 30742 28500 30748 28552
rect 30800 28500 30806 28552
rect 30834 28500 30840 28552
rect 30892 28549 30898 28552
rect 30892 28540 30900 28549
rect 31297 28543 31355 28549
rect 31297 28540 31309 28543
rect 30892 28512 30937 28540
rect 31036 28512 31309 28540
rect 30892 28503 30900 28512
rect 30892 28500 30898 28503
rect 30024 28444 30512 28472
rect 30576 28472 30604 28500
rect 30653 28475 30711 28481
rect 30653 28472 30665 28475
rect 30576 28444 30665 28472
rect 30653 28441 30665 28444
rect 30699 28441 30711 28475
rect 30653 28435 30711 28441
rect 24688 28376 26372 28404
rect 29549 28407 29607 28413
rect 29549 28373 29561 28407
rect 29595 28373 29607 28407
rect 29549 28367 29607 28373
rect 29917 28407 29975 28413
rect 29917 28373 29929 28407
rect 29963 28404 29975 28407
rect 30190 28404 30196 28416
rect 29963 28376 30196 28404
rect 29963 28373 29975 28376
rect 29917 28367 29975 28373
rect 30190 28364 30196 28376
rect 30248 28364 30254 28416
rect 31036 28413 31064 28512
rect 31297 28509 31309 28512
rect 31343 28509 31355 28543
rect 31297 28503 31355 28509
rect 31386 28500 31392 28552
rect 31444 28500 31450 28552
rect 31496 28550 31524 28636
rect 32033 28611 32091 28617
rect 32033 28577 32045 28611
rect 32079 28608 32091 28611
rect 32398 28608 32404 28620
rect 32079 28580 32404 28608
rect 32079 28577 32091 28580
rect 32033 28571 32091 28577
rect 32398 28568 32404 28580
rect 32456 28568 32462 28620
rect 33318 28568 33324 28620
rect 33376 28608 33382 28620
rect 33873 28611 33931 28617
rect 33873 28608 33885 28611
rect 33376 28580 33885 28608
rect 33376 28568 33382 28580
rect 33873 28577 33885 28580
rect 33919 28608 33931 28611
rect 33962 28608 33968 28620
rect 33919 28580 33968 28608
rect 33919 28577 33931 28580
rect 33873 28571 33931 28577
rect 33962 28568 33968 28580
rect 34020 28568 34026 28620
rect 34072 28617 34100 28716
rect 34057 28611 34115 28617
rect 34057 28577 34069 28611
rect 34103 28608 34115 28611
rect 36449 28611 36507 28617
rect 36449 28608 36461 28611
rect 34103 28580 36461 28608
rect 34103 28577 34115 28580
rect 34057 28571 34115 28577
rect 36449 28577 36461 28580
rect 36495 28577 36507 28611
rect 36449 28571 36507 28577
rect 31557 28553 31615 28559
rect 31557 28550 31569 28553
rect 31496 28522 31569 28550
rect 31557 28519 31569 28522
rect 31603 28519 31615 28553
rect 31557 28513 31615 28519
rect 31754 28500 31760 28552
rect 31812 28500 31818 28552
rect 34698 28500 34704 28552
rect 34756 28500 34762 28552
rect 31404 28472 31432 28500
rect 31481 28475 31539 28481
rect 31481 28472 31493 28475
rect 31404 28444 31493 28472
rect 31481 28441 31493 28444
rect 31527 28441 31539 28475
rect 34054 28472 34060 28484
rect 33258 28444 34060 28472
rect 31481 28435 31539 28441
rect 34054 28432 34060 28444
rect 34112 28432 34118 28484
rect 34422 28432 34428 28484
rect 34480 28472 34486 28484
rect 34977 28475 35035 28481
rect 34977 28472 34989 28475
rect 34480 28444 34989 28472
rect 34480 28432 34486 28444
rect 34977 28441 34989 28444
rect 35023 28441 35035 28475
rect 34977 28435 35035 28441
rect 35986 28432 35992 28484
rect 36044 28432 36050 28484
rect 31021 28407 31079 28413
rect 31021 28373 31033 28407
rect 31067 28373 31079 28407
rect 31021 28367 31079 28373
rect 31110 28364 31116 28416
rect 31168 28364 31174 28416
rect 32674 28364 32680 28416
rect 32732 28404 32738 28416
rect 33505 28407 33563 28413
rect 33505 28404 33517 28407
rect 32732 28376 33517 28404
rect 32732 28364 32738 28376
rect 33505 28373 33517 28376
rect 33551 28373 33563 28407
rect 33505 28367 33563 28373
rect 34146 28364 34152 28416
rect 34204 28364 34210 28416
rect 34514 28364 34520 28416
rect 34572 28364 34578 28416
rect 1104 28314 38272 28336
rect 1104 28262 4874 28314
rect 4926 28262 4938 28314
rect 4990 28262 5002 28314
rect 5054 28262 5066 28314
rect 5118 28262 5130 28314
rect 5182 28262 35594 28314
rect 35646 28262 35658 28314
rect 35710 28262 35722 28314
rect 35774 28262 35786 28314
rect 35838 28262 35850 28314
rect 35902 28262 38272 28314
rect 1104 28240 38272 28262
rect 4246 28160 4252 28212
rect 4304 28160 4310 28212
rect 5813 28203 5871 28209
rect 5813 28169 5825 28203
rect 5859 28200 5871 28203
rect 6733 28203 6791 28209
rect 6733 28200 6745 28203
rect 5859 28172 6745 28200
rect 5859 28169 5871 28172
rect 5813 28163 5871 28169
rect 6733 28169 6745 28172
rect 6779 28200 6791 28203
rect 8018 28200 8024 28212
rect 6779 28172 8024 28200
rect 6779 28169 6791 28172
rect 6733 28163 6791 28169
rect 8018 28160 8024 28172
rect 8076 28160 8082 28212
rect 8202 28160 8208 28212
rect 8260 28160 8266 28212
rect 10502 28160 10508 28212
rect 10560 28200 10566 28212
rect 10597 28203 10655 28209
rect 10597 28200 10609 28203
rect 10560 28172 10609 28200
rect 10560 28160 10566 28172
rect 10597 28169 10609 28172
rect 10643 28169 10655 28203
rect 10597 28163 10655 28169
rect 11517 28203 11575 28209
rect 11517 28169 11529 28203
rect 11563 28169 11575 28203
rect 11517 28163 11575 28169
rect 4264 28132 4292 28160
rect 4080 28104 4292 28132
rect 4080 28073 4108 28104
rect 6822 28092 6828 28144
rect 6880 28092 6886 28144
rect 8220 28132 8248 28160
rect 7668 28104 8248 28132
rect 4065 28067 4123 28073
rect 4065 28033 4077 28067
rect 4111 28033 4123 28067
rect 4065 28027 4123 28033
rect 5442 28024 5448 28076
rect 5500 28024 5506 28076
rect 7668 28073 7696 28104
rect 9490 28092 9496 28144
rect 9548 28132 9554 28144
rect 11238 28132 11244 28144
rect 9548 28104 11244 28132
rect 9548 28092 9554 28104
rect 11238 28092 11244 28104
rect 11296 28092 11302 28144
rect 7653 28067 7711 28073
rect 7653 28033 7665 28067
rect 7699 28033 7711 28067
rect 9674 28064 9680 28076
rect 9062 28050 9680 28064
rect 7653 28027 7711 28033
rect 9048 28036 9680 28050
rect 4341 27999 4399 28005
rect 4341 27965 4353 27999
rect 4387 27996 4399 27999
rect 4706 27996 4712 28008
rect 4387 27968 4712 27996
rect 4387 27965 4399 27968
rect 4341 27959 4399 27965
rect 4706 27956 4712 27968
rect 4764 27956 4770 28008
rect 7006 27956 7012 28008
rect 7064 27956 7070 28008
rect 7929 27999 7987 28005
rect 7929 27965 7941 27999
rect 7975 27996 7987 27999
rect 8294 27996 8300 28008
rect 7975 27968 8300 27996
rect 7975 27965 7987 27968
rect 7929 27959 7987 27965
rect 8294 27956 8300 27968
rect 8352 27956 8358 28008
rect 6362 27820 6368 27872
rect 6420 27820 6426 27872
rect 7190 27820 7196 27872
rect 7248 27860 7254 27872
rect 9048 27860 9076 28036
rect 9674 28024 9680 28036
rect 9732 28024 9738 28076
rect 9766 28024 9772 28076
rect 9824 28064 9830 28076
rect 9953 28067 10011 28073
rect 9953 28064 9965 28067
rect 9824 28036 9965 28064
rect 9824 28024 9830 28036
rect 9953 28033 9965 28036
rect 9999 28033 10011 28067
rect 9953 28027 10011 28033
rect 10781 28067 10839 28073
rect 10781 28033 10793 28067
rect 10827 28064 10839 28067
rect 11532 28064 11560 28163
rect 13354 28160 13360 28212
rect 13412 28200 13418 28212
rect 13725 28203 13783 28209
rect 13725 28200 13737 28203
rect 13412 28172 13737 28200
rect 13412 28160 13418 28172
rect 13725 28169 13737 28172
rect 13771 28169 13783 28203
rect 13725 28163 13783 28169
rect 13906 28160 13912 28212
rect 13964 28200 13970 28212
rect 15746 28200 15752 28212
rect 13964 28172 15752 28200
rect 13964 28160 13970 28172
rect 15746 28160 15752 28172
rect 15804 28160 15810 28212
rect 16114 28160 16120 28212
rect 16172 28160 16178 28212
rect 17313 28203 17371 28209
rect 17313 28169 17325 28203
rect 17359 28200 17371 28203
rect 17494 28200 17500 28212
rect 17359 28172 17500 28200
rect 17359 28169 17371 28172
rect 17313 28163 17371 28169
rect 17494 28160 17500 28172
rect 17552 28160 17558 28212
rect 17586 28160 17592 28212
rect 17644 28200 17650 28212
rect 18782 28200 18788 28212
rect 17644 28172 18788 28200
rect 17644 28160 17650 28172
rect 18782 28160 18788 28172
rect 18840 28160 18846 28212
rect 22186 28200 22192 28212
rect 19076 28172 19472 28200
rect 11885 28135 11943 28141
rect 11885 28101 11897 28135
rect 11931 28132 11943 28135
rect 11974 28132 11980 28144
rect 11931 28104 11980 28132
rect 11931 28101 11943 28104
rect 11885 28095 11943 28101
rect 11974 28092 11980 28104
rect 12032 28132 12038 28144
rect 14090 28132 14096 28144
rect 12032 28104 14096 28132
rect 12032 28092 12038 28104
rect 12452 28073 12480 28104
rect 14090 28092 14096 28104
rect 14148 28092 14154 28144
rect 16132 28132 16160 28160
rect 14752 28104 16160 28132
rect 10827 28036 11560 28064
rect 12437 28067 12495 28073
rect 10827 28033 10839 28036
rect 10781 28027 10839 28033
rect 12437 28033 12449 28067
rect 12483 28033 12495 28067
rect 12437 28027 12495 28033
rect 12618 28024 12624 28076
rect 12676 28024 12682 28076
rect 12713 28067 12771 28073
rect 12713 28033 12725 28067
rect 12759 28033 12771 28067
rect 12713 28027 12771 28033
rect 12805 28067 12863 28073
rect 12805 28033 12817 28067
rect 12851 28064 12863 28067
rect 13446 28064 13452 28076
rect 12851 28036 13452 28064
rect 12851 28033 12863 28036
rect 12805 28027 12863 28033
rect 10045 27999 10103 28005
rect 10045 27965 10057 27999
rect 10091 27965 10103 27999
rect 10045 27959 10103 27965
rect 9401 27931 9459 27937
rect 9401 27897 9413 27931
rect 9447 27928 9459 27931
rect 10060 27928 10088 27959
rect 10134 27956 10140 28008
rect 10192 27956 10198 28008
rect 11974 27956 11980 28008
rect 12032 27956 12038 28008
rect 12066 27956 12072 28008
rect 12124 27956 12130 28008
rect 12728 27996 12756 28027
rect 13446 28024 13452 28036
rect 13504 28024 13510 28076
rect 13817 28067 13875 28073
rect 13817 28033 13829 28067
rect 13863 28064 13875 28067
rect 14550 28064 14556 28076
rect 13863 28036 14556 28064
rect 13863 28033 13875 28036
rect 13817 28027 13875 28033
rect 14550 28024 14556 28036
rect 14608 28024 14614 28076
rect 14642 28024 14648 28076
rect 14700 28024 14706 28076
rect 14752 28073 14780 28104
rect 16574 28092 16580 28144
rect 16632 28132 16638 28144
rect 17037 28135 17095 28141
rect 17037 28132 17049 28135
rect 16632 28104 17049 28132
rect 16632 28092 16638 28104
rect 17037 28101 17049 28104
rect 17083 28101 17095 28135
rect 17037 28095 17095 28101
rect 17402 28092 17408 28144
rect 17460 28132 17466 28144
rect 19076 28141 19104 28172
rect 19061 28135 19119 28141
rect 19061 28132 19073 28135
rect 17460 28104 19073 28132
rect 17460 28092 17466 28104
rect 19061 28101 19073 28104
rect 19107 28101 19119 28135
rect 19242 28132 19248 28144
rect 19300 28141 19306 28144
rect 19300 28135 19319 28141
rect 19061 28095 19119 28101
rect 19168 28104 19248 28132
rect 14737 28067 14795 28073
rect 14737 28033 14749 28067
rect 14783 28033 14795 28067
rect 14737 28027 14795 28033
rect 14921 28067 14979 28073
rect 14921 28033 14933 28067
rect 14967 28064 14979 28067
rect 15010 28064 15016 28076
rect 14967 28036 15016 28064
rect 14967 28033 14979 28036
rect 14921 28027 14979 28033
rect 15010 28024 15016 28036
rect 15068 28064 15074 28076
rect 16022 28064 16028 28076
rect 15068 28036 16028 28064
rect 15068 28024 15074 28036
rect 16022 28024 16028 28036
rect 16080 28024 16086 28076
rect 16666 28024 16672 28076
rect 16724 28024 16730 28076
rect 16758 28024 16764 28076
rect 16816 28064 16822 28076
rect 16945 28067 17003 28073
rect 16816 28036 16861 28064
rect 16816 28024 16822 28036
rect 16945 28033 16957 28067
rect 16991 28033 17003 28067
rect 16945 28027 17003 28033
rect 17175 28067 17233 28073
rect 17175 28033 17187 28067
rect 17221 28064 17233 28067
rect 17862 28064 17868 28076
rect 17221 28036 17868 28064
rect 17221 28033 17233 28036
rect 17175 28027 17233 28033
rect 13541 27999 13599 28005
rect 13541 27996 13553 27999
rect 12728 27968 13553 27996
rect 9447 27900 12434 27928
rect 9447 27897 9459 27900
rect 9401 27891 9459 27897
rect 7248 27832 9076 27860
rect 7248 27820 7254 27832
rect 9490 27820 9496 27872
rect 9548 27860 9554 27872
rect 9585 27863 9643 27869
rect 9585 27860 9597 27863
rect 9548 27832 9597 27860
rect 9548 27820 9554 27832
rect 9585 27829 9597 27832
rect 9631 27829 9643 27863
rect 9585 27823 9643 27829
rect 9766 27820 9772 27872
rect 9824 27860 9830 27872
rect 11974 27860 11980 27872
rect 9824 27832 11980 27860
rect 9824 27820 9830 27832
rect 11974 27820 11980 27832
rect 12032 27820 12038 27872
rect 12406 27860 12434 27900
rect 12728 27860 12756 27968
rect 13541 27965 13553 27968
rect 13587 27996 13599 27999
rect 16776 27996 16804 28024
rect 13587 27968 16804 27996
rect 16960 27996 16988 28027
rect 17862 28024 17868 28036
rect 17920 28024 17926 28076
rect 18322 28024 18328 28076
rect 18380 28064 18386 28076
rect 18874 28064 18880 28076
rect 18380 28036 18880 28064
rect 18380 28024 18386 28036
rect 18874 28024 18880 28036
rect 18932 28064 18938 28076
rect 19168 28064 19196 28104
rect 19242 28092 19248 28104
rect 19307 28101 19319 28135
rect 19444 28132 19472 28172
rect 19628 28172 22192 28200
rect 19628 28132 19656 28172
rect 19444 28104 19656 28132
rect 19719 28104 19932 28132
rect 19300 28095 19319 28101
rect 19300 28092 19306 28095
rect 19518 28064 19524 28076
rect 18932 28036 19196 28064
rect 19352 28036 19524 28064
rect 18932 28024 18938 28036
rect 19352 27996 19380 28036
rect 19518 28024 19524 28036
rect 19576 28024 19582 28076
rect 19610 28024 19616 28076
rect 19668 28024 19674 28076
rect 19719 27996 19747 28104
rect 19794 28024 19800 28076
rect 19852 28024 19858 28076
rect 19904 28073 19932 28104
rect 19978 28092 19984 28144
rect 20036 28132 20042 28144
rect 20036 28104 20945 28132
rect 20036 28092 20042 28104
rect 20548 28073 20576 28104
rect 19889 28067 19947 28073
rect 19889 28033 19901 28067
rect 19935 28033 19947 28067
rect 19889 28027 19947 28033
rect 20533 28067 20591 28073
rect 20533 28033 20545 28067
rect 20579 28033 20591 28067
rect 20533 28027 20591 28033
rect 20622 28024 20628 28076
rect 20680 28064 20686 28076
rect 20917 28073 20945 28104
rect 21082 28092 21088 28144
rect 21140 28092 21146 28144
rect 21192 28141 21220 28172
rect 22186 28160 22192 28172
rect 22244 28160 22250 28212
rect 23014 28160 23020 28212
rect 23072 28200 23078 28212
rect 23109 28203 23167 28209
rect 23109 28200 23121 28203
rect 23072 28172 23121 28200
rect 23072 28160 23078 28172
rect 23109 28169 23121 28172
rect 23155 28169 23167 28203
rect 23109 28163 23167 28169
rect 23566 28160 23572 28212
rect 23624 28200 23630 28212
rect 23845 28203 23903 28209
rect 23845 28200 23857 28203
rect 23624 28172 23857 28200
rect 23624 28160 23630 28172
rect 23845 28169 23857 28172
rect 23891 28169 23903 28203
rect 23845 28163 23903 28169
rect 24670 28160 24676 28212
rect 24728 28160 24734 28212
rect 30742 28160 30748 28212
rect 30800 28160 30806 28212
rect 31754 28160 31760 28212
rect 31812 28200 31818 28212
rect 31849 28203 31907 28209
rect 31849 28200 31861 28203
rect 31812 28172 31861 28200
rect 31812 28160 31818 28172
rect 31849 28169 31861 28172
rect 31895 28169 31907 28203
rect 31849 28163 31907 28169
rect 32585 28203 32643 28209
rect 32585 28169 32597 28203
rect 32631 28200 32643 28203
rect 32674 28200 32680 28212
rect 32631 28172 32680 28200
rect 32631 28169 32643 28172
rect 32585 28163 32643 28169
rect 21177 28135 21235 28141
rect 21177 28101 21189 28135
rect 21223 28101 21235 28135
rect 21177 28095 21235 28101
rect 21542 28092 21548 28144
rect 21600 28132 21606 28144
rect 24688 28132 24716 28160
rect 21600 28104 23520 28132
rect 21600 28092 21606 28104
rect 20809 28067 20867 28073
rect 20809 28064 20821 28067
rect 20680 28036 20821 28064
rect 20680 28024 20686 28036
rect 20809 28033 20821 28036
rect 20855 28033 20867 28067
rect 20809 28027 20867 28033
rect 20902 28067 20960 28073
rect 20902 28033 20914 28067
rect 20948 28033 20960 28067
rect 20902 28027 20960 28033
rect 21315 28067 21373 28073
rect 21315 28033 21327 28067
rect 21361 28064 21373 28067
rect 21450 28064 21456 28076
rect 21361 28036 21456 28064
rect 21361 28033 21373 28036
rect 21315 28027 21373 28033
rect 20165 27999 20223 28005
rect 20165 27996 20177 27999
rect 16960 27968 19380 27996
rect 19444 27968 19747 27996
rect 19996 27968 20177 27996
rect 13587 27965 13599 27968
rect 13541 27959 13599 27965
rect 14093 27931 14151 27937
rect 14093 27897 14105 27931
rect 14139 27928 14151 27931
rect 14553 27931 14611 27937
rect 14553 27928 14565 27931
rect 14139 27900 14565 27928
rect 14139 27897 14151 27900
rect 14093 27891 14151 27897
rect 14553 27897 14565 27900
rect 14599 27897 14611 27931
rect 14553 27891 14611 27897
rect 15562 27888 15568 27940
rect 15620 27928 15626 27940
rect 19444 27937 19472 27968
rect 19429 27931 19487 27937
rect 15620 27900 19380 27928
rect 15620 27888 15626 27900
rect 12406 27832 12756 27860
rect 12989 27863 13047 27869
rect 12989 27829 13001 27863
rect 13035 27860 13047 27863
rect 13630 27860 13636 27872
rect 13035 27832 13636 27860
rect 13035 27829 13047 27832
rect 12989 27823 13047 27829
rect 13630 27820 13636 27832
rect 13688 27820 13694 27872
rect 14182 27820 14188 27872
rect 14240 27820 14246 27872
rect 14458 27820 14464 27872
rect 14516 27860 14522 27872
rect 15470 27860 15476 27872
rect 14516 27832 15476 27860
rect 14516 27820 14522 27832
rect 15470 27820 15476 27832
rect 15528 27820 15534 27872
rect 15838 27820 15844 27872
rect 15896 27860 15902 27872
rect 19242 27860 19248 27872
rect 15896 27832 19248 27860
rect 15896 27820 15902 27832
rect 19242 27820 19248 27832
rect 19300 27820 19306 27872
rect 19352 27860 19380 27900
rect 19429 27897 19441 27931
rect 19475 27897 19487 27931
rect 19429 27891 19487 27897
rect 19705 27931 19763 27937
rect 19705 27897 19717 27931
rect 19751 27928 19763 27931
rect 19996 27928 20024 27968
rect 20165 27965 20177 27968
rect 20211 27965 20223 27999
rect 20165 27959 20223 27965
rect 20254 27956 20260 28008
rect 20312 27996 20318 28008
rect 20349 27999 20407 28005
rect 20349 27996 20361 27999
rect 20312 27968 20361 27996
rect 20312 27956 20318 27968
rect 20349 27965 20361 27968
rect 20395 27965 20407 27999
rect 20349 27959 20407 27965
rect 20438 27956 20444 28008
rect 20496 27956 20502 28008
rect 19751 27900 20024 27928
rect 20073 27931 20131 27937
rect 19751 27897 19763 27900
rect 19705 27891 19763 27897
rect 20073 27897 20085 27931
rect 20119 27928 20131 27931
rect 20119 27900 20484 27928
rect 20119 27897 20131 27900
rect 20073 27891 20131 27897
rect 20456 27872 20484 27900
rect 20346 27860 20352 27872
rect 19352 27832 20352 27860
rect 20346 27820 20352 27832
rect 20404 27820 20410 27872
rect 20438 27820 20444 27872
rect 20496 27820 20502 27872
rect 20917 27860 20945 28027
rect 21450 28024 21456 28036
rect 21508 28064 21514 28076
rect 22370 28064 22376 28076
rect 21508 28036 22376 28064
rect 21508 28024 21514 28036
rect 22370 28024 22376 28036
rect 22428 28024 22434 28076
rect 22462 28024 22468 28076
rect 22520 28024 22526 28076
rect 22833 28067 22891 28073
rect 22833 28033 22845 28067
rect 22879 28064 22891 28067
rect 23198 28064 23204 28076
rect 22879 28036 23204 28064
rect 22879 28033 22891 28036
rect 22833 28027 22891 28033
rect 23198 28024 23204 28036
rect 23256 28024 23262 28076
rect 23293 28067 23351 28073
rect 23293 28033 23305 28067
rect 23339 28033 23351 28067
rect 23293 28027 23351 28033
rect 21910 27956 21916 28008
rect 21968 27956 21974 28008
rect 22281 27999 22339 28005
rect 22281 27996 22293 27999
rect 22066 27968 22293 27996
rect 21453 27931 21511 27937
rect 21453 27897 21465 27931
rect 21499 27928 21511 27931
rect 22066 27928 22094 27968
rect 22281 27965 22293 27968
rect 22327 27965 22339 27999
rect 22281 27959 22339 27965
rect 22741 27999 22799 28005
rect 22741 27965 22753 27999
rect 22787 27965 22799 27999
rect 22741 27959 22799 27965
rect 21499 27900 22094 27928
rect 22756 27928 22784 27959
rect 22922 27956 22928 28008
rect 22980 27996 22986 28008
rect 23308 27996 23336 28027
rect 23382 28024 23388 28076
rect 23440 28024 23446 28076
rect 23492 28073 23520 28104
rect 23676 28104 24716 28132
rect 30760 28132 30788 28160
rect 32600 28132 32628 28163
rect 32674 28160 32680 28172
rect 32732 28160 32738 28212
rect 32953 28203 33011 28209
rect 32953 28169 32965 28203
rect 32999 28200 33011 28203
rect 33042 28200 33048 28212
rect 32999 28172 33048 28200
rect 32999 28169 33011 28172
rect 32953 28163 33011 28169
rect 33042 28160 33048 28172
rect 33100 28160 33106 28212
rect 34422 28160 34428 28212
rect 34480 28160 34486 28212
rect 34698 28160 34704 28212
rect 34756 28200 34762 28212
rect 34885 28203 34943 28209
rect 34885 28200 34897 28203
rect 34756 28172 34897 28200
rect 34756 28160 34762 28172
rect 34885 28169 34897 28172
rect 34931 28169 34943 28203
rect 34885 28163 34943 28169
rect 37274 28160 37280 28212
rect 37332 28160 37338 28212
rect 30760 28104 32628 28132
rect 23676 28073 23704 28104
rect 23477 28067 23535 28073
rect 23477 28033 23489 28067
rect 23523 28033 23535 28067
rect 23477 28027 23535 28033
rect 23661 28067 23719 28073
rect 23661 28033 23673 28067
rect 23707 28033 23719 28067
rect 23661 28027 23719 28033
rect 23753 28067 23811 28073
rect 23753 28033 23765 28067
rect 23799 28033 23811 28067
rect 23753 28027 23811 28033
rect 24121 28067 24179 28073
rect 24121 28033 24133 28067
rect 24167 28064 24179 28067
rect 24210 28064 24216 28076
rect 24167 28036 24216 28064
rect 24167 28033 24179 28036
rect 24121 28027 24179 28033
rect 22980 27968 23336 27996
rect 22980 27956 22986 27968
rect 23566 27956 23572 28008
rect 23624 27996 23630 28008
rect 23768 27996 23796 28027
rect 24210 28024 24216 28036
rect 24268 28024 24274 28076
rect 24394 28024 24400 28076
rect 24452 28024 24458 28076
rect 24670 28024 24676 28076
rect 24728 28064 24734 28076
rect 31846 28064 31852 28076
rect 24728 28036 31852 28064
rect 24728 28024 24734 28036
rect 31846 28024 31852 28036
rect 31904 28024 31910 28076
rect 31938 28024 31944 28076
rect 31996 28024 32002 28076
rect 32493 28067 32551 28073
rect 32493 28064 32505 28067
rect 32232 28036 32505 28064
rect 23624 27968 23796 27996
rect 23624 27956 23630 27968
rect 23750 27928 23756 27940
rect 22756 27900 23756 27928
rect 21499 27897 21511 27900
rect 21453 27891 21511 27897
rect 23750 27888 23756 27900
rect 23808 27888 23814 27940
rect 24029 27931 24087 27937
rect 24029 27897 24041 27931
rect 24075 27928 24087 27931
rect 24412 27928 24440 28024
rect 30190 27956 30196 28008
rect 30248 27996 30254 28008
rect 32232 27996 32260 28036
rect 32493 28033 32505 28036
rect 32539 28064 32551 28067
rect 34146 28064 34152 28076
rect 32539 28036 34152 28064
rect 32539 28033 32551 28036
rect 32493 28027 32551 28033
rect 34146 28024 34152 28036
rect 34204 28024 34210 28076
rect 34241 28067 34299 28073
rect 34241 28033 34253 28067
rect 34287 28064 34299 28067
rect 34514 28064 34520 28076
rect 34287 28036 34520 28064
rect 34287 28033 34299 28036
rect 34241 28027 34299 28033
rect 34514 28024 34520 28036
rect 34572 28024 34578 28076
rect 34977 28067 35035 28073
rect 34977 28033 34989 28067
rect 35023 28033 35035 28067
rect 37292 28064 37320 28160
rect 37369 28067 37427 28073
rect 37369 28064 37381 28067
rect 37292 28036 37381 28064
rect 34977 28027 35035 28033
rect 37369 28033 37381 28036
rect 37415 28033 37427 28067
rect 37369 28027 37427 28033
rect 30248 27968 32260 27996
rect 32401 27999 32459 28005
rect 30248 27956 30254 27968
rect 32401 27965 32413 27999
rect 32447 27996 32459 27999
rect 33134 27996 33140 28008
rect 32447 27968 33140 27996
rect 32447 27965 32459 27968
rect 32401 27959 32459 27965
rect 33134 27956 33140 27968
rect 33192 27996 33198 28008
rect 33870 27996 33876 28008
rect 33192 27968 33876 27996
rect 33192 27956 33198 27968
rect 33870 27956 33876 27968
rect 33928 27956 33934 28008
rect 24075 27900 24440 27928
rect 24075 27897 24087 27900
rect 24029 27891 24087 27897
rect 33686 27888 33692 27940
rect 33744 27928 33750 27940
rect 34606 27928 34612 27940
rect 33744 27900 34612 27928
rect 33744 27888 33750 27900
rect 34606 27888 34612 27900
rect 34664 27928 34670 27940
rect 34992 27928 35020 28027
rect 34664 27900 35020 27928
rect 34664 27888 34670 27900
rect 23382 27860 23388 27872
rect 20917 27832 23388 27860
rect 23382 27820 23388 27832
rect 23440 27820 23446 27872
rect 24210 27820 24216 27872
rect 24268 27820 24274 27872
rect 24486 27820 24492 27872
rect 24544 27820 24550 27872
rect 37550 27820 37556 27872
rect 37608 27820 37614 27872
rect 1104 27770 38272 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 38272 27770
rect 1104 27696 38272 27718
rect 4617 27659 4675 27665
rect 4617 27625 4629 27659
rect 4663 27656 4675 27659
rect 4706 27656 4712 27668
rect 4663 27628 4712 27656
rect 4663 27625 4675 27628
rect 4617 27619 4675 27625
rect 4706 27616 4712 27628
rect 4764 27616 4770 27668
rect 8294 27616 8300 27668
rect 8352 27616 8358 27668
rect 9490 27616 9496 27668
rect 9548 27616 9554 27668
rect 12618 27616 12624 27668
rect 12676 27656 12682 27668
rect 13170 27656 13176 27668
rect 12676 27628 13176 27656
rect 12676 27616 12682 27628
rect 13170 27616 13176 27628
rect 13228 27616 13234 27668
rect 14182 27616 14188 27668
rect 14240 27656 14246 27668
rect 14458 27656 14464 27668
rect 14240 27628 14464 27656
rect 14240 27616 14246 27628
rect 14458 27616 14464 27628
rect 14516 27616 14522 27668
rect 14642 27616 14648 27668
rect 14700 27616 14706 27668
rect 16574 27656 16580 27668
rect 14752 27628 16580 27656
rect 9508 27588 9536 27616
rect 8496 27560 9536 27588
rect 7558 27480 7564 27532
rect 7616 27480 7622 27532
rect 4801 27455 4859 27461
rect 4801 27421 4813 27455
rect 4847 27452 4859 27455
rect 6362 27452 6368 27464
rect 4847 27424 6368 27452
rect 4847 27421 4859 27424
rect 4801 27415 4859 27421
rect 6362 27412 6368 27424
rect 6420 27412 6426 27464
rect 6917 27455 6975 27461
rect 6917 27421 6929 27455
rect 6963 27452 6975 27455
rect 7576 27452 7604 27480
rect 8496 27461 8524 27560
rect 9582 27548 9588 27600
rect 9640 27548 9646 27600
rect 13906 27588 13912 27600
rect 12406 27560 13912 27588
rect 9600 27520 9628 27548
rect 9508 27492 9628 27520
rect 9508 27461 9536 27492
rect 11974 27480 11980 27532
rect 12032 27520 12038 27532
rect 12069 27523 12127 27529
rect 12069 27520 12081 27523
rect 12032 27492 12081 27520
rect 12032 27480 12038 27492
rect 12069 27489 12081 27492
rect 12115 27489 12127 27523
rect 12069 27483 12127 27489
rect 12161 27523 12219 27529
rect 12161 27489 12173 27523
rect 12207 27520 12219 27523
rect 12406 27520 12434 27560
rect 13906 27548 13912 27560
rect 13964 27548 13970 27600
rect 14090 27548 14096 27600
rect 14148 27588 14154 27600
rect 14752 27588 14780 27628
rect 16574 27616 16580 27628
rect 16632 27616 16638 27668
rect 16666 27616 16672 27668
rect 16724 27616 16730 27668
rect 21450 27656 21456 27668
rect 16776 27628 21456 27656
rect 14148 27560 14780 27588
rect 14148 27548 14154 27560
rect 15010 27548 15016 27600
rect 15068 27588 15074 27600
rect 15286 27588 15292 27600
rect 15068 27560 15292 27588
rect 15068 27548 15074 27560
rect 15286 27548 15292 27560
rect 15344 27588 15350 27600
rect 16025 27591 16083 27597
rect 15344 27560 15976 27588
rect 15344 27548 15350 27560
rect 12207 27492 12434 27520
rect 13081 27523 13139 27529
rect 12207 27489 12219 27492
rect 12161 27483 12219 27489
rect 13081 27489 13093 27523
rect 13127 27520 13139 27523
rect 13722 27520 13728 27532
rect 13127 27492 13728 27520
rect 13127 27489 13139 27492
rect 13081 27483 13139 27489
rect 6963 27424 7604 27452
rect 8481 27455 8539 27461
rect 6963 27421 6975 27424
rect 6917 27415 6975 27421
rect 8481 27421 8493 27455
rect 8527 27421 8539 27455
rect 8481 27415 8539 27421
rect 9493 27455 9551 27461
rect 9493 27421 9505 27455
rect 9539 27421 9551 27455
rect 9493 27415 9551 27421
rect 9585 27455 9643 27461
rect 9585 27421 9597 27455
rect 9631 27452 9643 27455
rect 9769 27455 9827 27461
rect 9769 27452 9781 27455
rect 9631 27424 9781 27452
rect 9631 27421 9643 27424
rect 9585 27415 9643 27421
rect 9769 27421 9781 27424
rect 9815 27421 9827 27455
rect 9769 27415 9827 27421
rect 11054 27412 11060 27464
rect 11112 27452 11118 27464
rect 12176 27452 12204 27483
rect 13722 27480 13728 27492
rect 13780 27480 13786 27532
rect 15948 27520 15976 27560
rect 16025 27557 16037 27591
rect 16071 27588 16083 27591
rect 16684 27588 16712 27616
rect 16071 27560 16712 27588
rect 16071 27557 16083 27560
rect 16025 27551 16083 27557
rect 16298 27520 16304 27532
rect 15948 27492 16304 27520
rect 16298 27480 16304 27492
rect 16356 27480 16362 27532
rect 16574 27480 16580 27532
rect 16632 27520 16638 27532
rect 16776 27520 16804 27628
rect 21450 27616 21456 27628
rect 21508 27616 21514 27668
rect 22002 27616 22008 27668
rect 22060 27656 22066 27668
rect 23566 27656 23572 27668
rect 22060 27628 23572 27656
rect 22060 27616 22066 27628
rect 23566 27616 23572 27628
rect 23624 27616 23630 27668
rect 23753 27659 23811 27665
rect 23753 27625 23765 27659
rect 23799 27656 23811 27659
rect 24210 27656 24216 27668
rect 23799 27628 24216 27656
rect 23799 27625 23811 27628
rect 23753 27619 23811 27625
rect 24210 27616 24216 27628
rect 24268 27616 24274 27668
rect 25038 27616 25044 27668
rect 25096 27656 25102 27668
rect 26602 27656 26608 27668
rect 25096 27628 26608 27656
rect 25096 27616 25102 27628
rect 26602 27616 26608 27628
rect 26660 27616 26666 27668
rect 26694 27616 26700 27668
rect 26752 27656 26758 27668
rect 27890 27656 27896 27668
rect 26752 27628 27896 27656
rect 26752 27616 26758 27628
rect 27890 27616 27896 27628
rect 27948 27616 27954 27668
rect 28442 27616 28448 27668
rect 28500 27656 28506 27668
rect 29730 27656 29736 27668
rect 28500 27628 29736 27656
rect 28500 27616 28506 27628
rect 29730 27616 29736 27628
rect 29788 27616 29794 27668
rect 18322 27588 18328 27600
rect 16632 27492 16804 27520
rect 16868 27560 18328 27588
rect 16632 27480 16638 27492
rect 11112 27424 11178 27452
rect 11440 27424 12204 27452
rect 13265 27455 13323 27461
rect 11112 27412 11118 27424
rect 10042 27344 10048 27396
rect 10100 27344 10106 27396
rect 6822 27276 6828 27328
rect 6880 27276 6886 27328
rect 9858 27276 9864 27328
rect 9916 27316 9922 27328
rect 11440 27316 11468 27424
rect 13265 27421 13277 27455
rect 13311 27452 13323 27455
rect 13446 27452 13452 27464
rect 13311 27424 13452 27452
rect 13311 27421 13323 27424
rect 13265 27415 13323 27421
rect 13446 27412 13452 27424
rect 13504 27412 13510 27464
rect 14366 27412 14372 27464
rect 14424 27452 14430 27464
rect 14461 27455 14519 27461
rect 14461 27452 14473 27455
rect 14424 27424 14473 27452
rect 14424 27412 14430 27424
rect 14461 27421 14473 27424
rect 14507 27421 14519 27455
rect 14461 27415 14519 27421
rect 14826 27412 14832 27464
rect 14884 27452 14890 27464
rect 15565 27455 15623 27461
rect 15565 27452 15577 27455
rect 14884 27424 15577 27452
rect 14884 27412 14890 27424
rect 15565 27421 15577 27424
rect 15611 27421 15623 27455
rect 15565 27415 15623 27421
rect 15657 27455 15715 27461
rect 15657 27421 15669 27455
rect 15703 27421 15715 27455
rect 15657 27415 15715 27421
rect 11977 27387 12035 27393
rect 11977 27384 11989 27387
rect 11532 27356 11989 27384
rect 11532 27325 11560 27356
rect 11977 27353 11989 27356
rect 12023 27384 12035 27387
rect 12342 27384 12348 27396
rect 12023 27356 12348 27384
rect 12023 27353 12035 27356
rect 11977 27347 12035 27353
rect 12342 27344 12348 27356
rect 12400 27384 12406 27396
rect 14844 27384 14872 27412
rect 12400 27356 14872 27384
rect 15672 27384 15700 27415
rect 15838 27412 15844 27464
rect 15896 27452 15902 27464
rect 16206 27452 16212 27464
rect 15896 27424 16212 27452
rect 15896 27412 15902 27424
rect 16206 27412 16212 27424
rect 16264 27412 16270 27464
rect 16666 27412 16672 27464
rect 16724 27412 16730 27464
rect 16758 27412 16764 27464
rect 16816 27412 16822 27464
rect 16868 27384 16896 27560
rect 18322 27548 18328 27560
rect 18380 27548 18386 27600
rect 18506 27548 18512 27600
rect 18564 27588 18570 27600
rect 23658 27588 23664 27600
rect 18564 27560 23664 27588
rect 18564 27548 18570 27560
rect 23658 27548 23664 27560
rect 23716 27548 23722 27600
rect 25498 27548 25504 27600
rect 25556 27548 25562 27600
rect 28994 27548 29000 27600
rect 29052 27548 29058 27600
rect 31846 27588 31852 27600
rect 31726 27560 31852 27588
rect 18690 27520 18696 27532
rect 16960 27492 17264 27520
rect 16960 27461 16988 27492
rect 16945 27455 17003 27461
rect 16945 27421 16957 27455
rect 16991 27421 17003 27455
rect 16945 27415 17003 27421
rect 17126 27412 17132 27464
rect 17184 27461 17190 27464
rect 17184 27415 17192 27461
rect 17236 27452 17264 27492
rect 17696 27492 18696 27520
rect 17310 27452 17316 27464
rect 17236 27424 17316 27452
rect 17184 27412 17190 27415
rect 17310 27412 17316 27424
rect 17368 27412 17374 27464
rect 17402 27412 17408 27464
rect 17460 27412 17466 27464
rect 17494 27412 17500 27464
rect 17552 27452 17558 27464
rect 17696 27461 17724 27492
rect 18690 27480 18696 27492
rect 18748 27480 18754 27532
rect 20346 27480 20352 27532
rect 20404 27520 20410 27532
rect 21542 27520 21548 27532
rect 20404 27492 21548 27520
rect 20404 27480 20410 27492
rect 21542 27480 21548 27492
rect 21600 27480 21606 27532
rect 23382 27520 23388 27532
rect 22940 27492 23388 27520
rect 17589 27455 17647 27461
rect 17589 27452 17601 27455
rect 17552 27424 17601 27452
rect 17552 27412 17558 27424
rect 17589 27421 17601 27424
rect 17635 27421 17647 27455
rect 17589 27415 17647 27421
rect 17681 27455 17739 27461
rect 17681 27421 17693 27455
rect 17727 27421 17739 27455
rect 17681 27415 17739 27421
rect 17773 27455 17831 27461
rect 17773 27421 17785 27455
rect 17819 27421 17831 27455
rect 18138 27452 18144 27464
rect 17773 27415 17831 27421
rect 17972 27424 18144 27452
rect 15672 27356 16896 27384
rect 17037 27387 17095 27393
rect 12400 27344 12406 27356
rect 17037 27353 17049 27387
rect 17083 27384 17095 27387
rect 17788 27384 17816 27415
rect 17972 27396 18000 27424
rect 18138 27412 18144 27424
rect 18196 27412 18202 27464
rect 18325 27455 18383 27461
rect 18325 27421 18337 27455
rect 18371 27421 18383 27455
rect 18325 27415 18383 27421
rect 18417 27455 18475 27461
rect 18417 27421 18429 27455
rect 18463 27421 18475 27455
rect 18417 27415 18475 27421
rect 18601 27455 18659 27461
rect 18601 27421 18613 27455
rect 18647 27452 18659 27455
rect 18966 27452 18972 27464
rect 18647 27424 18972 27452
rect 18647 27421 18659 27424
rect 18601 27415 18659 27421
rect 17083 27356 17816 27384
rect 17083 27353 17095 27356
rect 17037 27347 17095 27353
rect 9916 27288 11468 27316
rect 11517 27319 11575 27325
rect 9916 27276 9922 27288
rect 11517 27285 11529 27319
rect 11563 27285 11575 27319
rect 11517 27279 11575 27285
rect 11606 27276 11612 27328
rect 11664 27276 11670 27328
rect 13354 27276 13360 27328
rect 13412 27316 13418 27328
rect 14090 27316 14096 27328
rect 13412 27288 14096 27316
rect 13412 27276 13418 27288
rect 14090 27276 14096 27288
rect 14148 27316 14154 27328
rect 14277 27319 14335 27325
rect 14277 27316 14289 27319
rect 14148 27288 14289 27316
rect 14148 27276 14154 27288
rect 14277 27285 14289 27288
rect 14323 27285 14335 27319
rect 14277 27279 14335 27285
rect 14369 27319 14427 27325
rect 14369 27285 14381 27319
rect 14415 27316 14427 27319
rect 14550 27316 14556 27328
rect 14415 27288 14556 27316
rect 14415 27285 14427 27288
rect 14369 27279 14427 27285
rect 14550 27276 14556 27288
rect 14608 27276 14614 27328
rect 15378 27276 15384 27328
rect 15436 27316 15442 27328
rect 17052 27316 17080 27347
rect 17954 27344 17960 27396
rect 18012 27344 18018 27396
rect 18049 27387 18107 27393
rect 18049 27353 18061 27387
rect 18095 27384 18107 27387
rect 18340 27384 18368 27415
rect 18095 27356 18368 27384
rect 18095 27353 18107 27356
rect 18049 27347 18107 27353
rect 15436 27288 17080 27316
rect 15436 27276 15442 27288
rect 17310 27276 17316 27328
rect 17368 27276 17374 27328
rect 17770 27276 17776 27328
rect 17828 27316 17834 27328
rect 18432 27316 18460 27415
rect 18966 27412 18972 27424
rect 19024 27412 19030 27464
rect 21266 27412 21272 27464
rect 21324 27452 21330 27464
rect 22940 27461 22968 27492
rect 23382 27480 23388 27492
rect 23440 27480 23446 27532
rect 23492 27492 25084 27520
rect 22925 27455 22983 27461
rect 21324 27424 22876 27452
rect 21324 27412 21330 27424
rect 18506 27344 18512 27396
rect 18564 27344 18570 27396
rect 20622 27384 20628 27396
rect 18616 27356 20628 27384
rect 18616 27316 18644 27356
rect 20622 27344 20628 27356
rect 20680 27384 20686 27396
rect 21818 27384 21824 27396
rect 20680 27356 21824 27384
rect 20680 27344 20686 27356
rect 21818 27344 21824 27356
rect 21876 27344 21882 27396
rect 22741 27387 22799 27393
rect 22741 27384 22753 27387
rect 22066 27356 22753 27384
rect 17828 27288 18644 27316
rect 17828 27276 17834 27288
rect 18782 27276 18788 27328
rect 18840 27276 18846 27328
rect 20162 27276 20168 27328
rect 20220 27316 20226 27328
rect 22066 27316 22094 27356
rect 22741 27353 22753 27356
rect 22787 27353 22799 27387
rect 22848 27384 22876 27424
rect 22925 27421 22937 27455
rect 22971 27421 22983 27455
rect 23201 27455 23259 27461
rect 23201 27452 23213 27455
rect 22925 27415 22983 27421
rect 23032 27424 23213 27452
rect 23032 27384 23060 27424
rect 23201 27421 23213 27424
rect 23247 27452 23259 27455
rect 23492 27452 23520 27492
rect 25056 27464 25084 27492
rect 23247 27424 23520 27452
rect 23247 27421 23259 27424
rect 23201 27415 23259 27421
rect 23566 27412 23572 27464
rect 23624 27452 23630 27464
rect 24118 27452 24124 27464
rect 23624 27424 24124 27452
rect 23624 27412 23630 27424
rect 24118 27412 24124 27424
rect 24176 27412 24182 27464
rect 25038 27412 25044 27464
rect 25096 27412 25102 27464
rect 25516 27461 25544 27548
rect 26418 27480 26424 27532
rect 26476 27520 26482 27532
rect 27525 27523 27583 27529
rect 27525 27520 27537 27523
rect 26476 27492 27537 27520
rect 26476 27480 26482 27492
rect 27525 27489 27537 27492
rect 27571 27489 27583 27523
rect 29012 27520 29040 27548
rect 31726 27520 31754 27560
rect 31846 27548 31852 27560
rect 31904 27548 31910 27600
rect 33778 27548 33784 27600
rect 33836 27548 33842 27600
rect 34330 27548 34336 27600
rect 34388 27548 34394 27600
rect 27525 27483 27583 27489
rect 27908 27492 29592 27520
rect 27908 27461 27936 27492
rect 25501 27455 25559 27461
rect 25501 27421 25513 27455
rect 25547 27421 25559 27455
rect 25501 27415 25559 27421
rect 25593 27455 25651 27461
rect 25593 27421 25605 27455
rect 25639 27452 25651 27455
rect 25777 27455 25835 27461
rect 25777 27452 25789 27455
rect 25639 27424 25789 27452
rect 25639 27421 25651 27424
rect 25593 27415 25651 27421
rect 25777 27421 25789 27424
rect 25823 27421 25835 27455
rect 25777 27415 25835 27421
rect 27893 27455 27951 27461
rect 27893 27421 27905 27455
rect 27939 27421 27951 27455
rect 27893 27415 27951 27421
rect 28166 27412 28172 27464
rect 28224 27412 28230 27464
rect 29564 27461 29592 27492
rect 29656 27492 31754 27520
rect 29549 27455 29607 27461
rect 29549 27421 29561 27455
rect 29595 27421 29607 27455
rect 29549 27415 29607 27421
rect 22848 27356 23060 27384
rect 23109 27387 23167 27393
rect 22741 27347 22799 27353
rect 23109 27353 23121 27387
rect 23155 27384 23167 27387
rect 23385 27387 23443 27393
rect 23385 27384 23397 27387
rect 23155 27356 23397 27384
rect 23155 27353 23167 27356
rect 23109 27347 23167 27353
rect 23385 27353 23397 27356
rect 23431 27353 23443 27387
rect 23385 27347 23443 27353
rect 23477 27387 23535 27393
rect 23477 27353 23489 27387
rect 23523 27353 23535 27387
rect 23477 27347 23535 27353
rect 20220 27288 22094 27316
rect 20220 27276 20226 27288
rect 22186 27276 22192 27328
rect 22244 27316 22250 27328
rect 23492 27316 23520 27347
rect 25682 27344 25688 27396
rect 25740 27344 25746 27396
rect 26053 27387 26111 27393
rect 26053 27353 26065 27387
rect 26099 27384 26111 27387
rect 26326 27384 26332 27396
rect 26099 27356 26332 27384
rect 26099 27353 26111 27356
rect 26053 27347 26111 27353
rect 26326 27344 26332 27356
rect 26384 27344 26390 27396
rect 26786 27344 26792 27396
rect 26844 27344 26850 27396
rect 29656 27384 29684 27492
rect 30006 27412 30012 27464
rect 30064 27412 30070 27464
rect 30374 27412 30380 27464
rect 30432 27412 30438 27464
rect 30470 27455 30528 27461
rect 30470 27421 30482 27455
rect 30516 27421 30528 27455
rect 30470 27415 30528 27421
rect 30484 27384 30512 27415
rect 30558 27412 30564 27464
rect 30616 27452 30622 27464
rect 30653 27455 30711 27461
rect 30653 27452 30665 27455
rect 30616 27424 30665 27452
rect 30616 27412 30622 27424
rect 30653 27421 30665 27424
rect 30699 27421 30711 27455
rect 30653 27415 30711 27421
rect 30745 27455 30803 27461
rect 30745 27421 30757 27455
rect 30791 27421 30803 27455
rect 30745 27415 30803 27421
rect 27356 27356 29684 27384
rect 30116 27356 30512 27384
rect 22244 27288 23520 27316
rect 25700 27316 25728 27344
rect 27356 27316 27384 27356
rect 30116 27328 30144 27356
rect 30760 27328 30788 27415
rect 30834 27412 30840 27464
rect 30892 27461 30898 27464
rect 30892 27455 30941 27461
rect 30892 27421 30895 27455
rect 30929 27452 30941 27455
rect 31018 27452 31024 27464
rect 30929 27424 31024 27452
rect 30929 27421 30941 27424
rect 30892 27415 30941 27421
rect 30892 27412 30898 27415
rect 31018 27412 31024 27424
rect 31076 27412 31082 27464
rect 31938 27412 31944 27464
rect 31996 27452 32002 27464
rect 33686 27452 33692 27464
rect 31996 27424 33692 27452
rect 31996 27412 32002 27424
rect 33686 27412 33692 27424
rect 33744 27412 33750 27464
rect 33965 27455 34023 27461
rect 33965 27421 33977 27455
rect 34011 27452 34023 27455
rect 34348 27452 34376 27548
rect 34011 27424 34376 27452
rect 34011 27421 34023 27424
rect 33965 27415 34023 27421
rect 25700 27288 27384 27316
rect 22244 27276 22250 27288
rect 27798 27276 27804 27328
rect 27856 27276 27862 27328
rect 27890 27276 27896 27328
rect 27948 27316 27954 27328
rect 27985 27319 28043 27325
rect 27985 27316 27997 27319
rect 27948 27288 27997 27316
rect 27948 27276 27954 27288
rect 27985 27285 27997 27288
rect 28031 27285 28043 27319
rect 27985 27279 28043 27285
rect 29638 27276 29644 27328
rect 29696 27276 29702 27328
rect 29822 27276 29828 27328
rect 29880 27276 29886 27328
rect 30098 27276 30104 27328
rect 30156 27276 30162 27328
rect 30742 27276 30748 27328
rect 30800 27276 30806 27328
rect 31021 27319 31079 27325
rect 31021 27285 31033 27319
rect 31067 27316 31079 27319
rect 31754 27316 31760 27328
rect 31067 27288 31760 27316
rect 31067 27285 31079 27288
rect 31021 27279 31079 27285
rect 31754 27276 31760 27288
rect 31812 27276 31818 27328
rect 33594 27276 33600 27328
rect 33652 27276 33658 27328
rect 1104 27226 38272 27248
rect 1104 27174 4874 27226
rect 4926 27174 4938 27226
rect 4990 27174 5002 27226
rect 5054 27174 5066 27226
rect 5118 27174 5130 27226
rect 5182 27174 35594 27226
rect 35646 27174 35658 27226
rect 35710 27174 35722 27226
rect 35774 27174 35786 27226
rect 35838 27174 35850 27226
rect 35902 27174 38272 27226
rect 1104 27152 38272 27174
rect 6822 27072 6828 27124
rect 6880 27072 6886 27124
rect 7006 27072 7012 27124
rect 7064 27112 7070 27124
rect 9858 27112 9864 27124
rect 7064 27084 9864 27112
rect 7064 27072 7070 27084
rect 9858 27072 9864 27084
rect 9916 27072 9922 27124
rect 10042 27072 10048 27124
rect 10100 27112 10106 27124
rect 10229 27115 10287 27121
rect 10229 27112 10241 27115
rect 10100 27084 10241 27112
rect 10100 27072 10106 27084
rect 10229 27081 10241 27084
rect 10275 27081 10287 27115
rect 10229 27075 10287 27081
rect 11606 27072 11612 27124
rect 11664 27072 11670 27124
rect 12250 27072 12256 27124
rect 12308 27112 12314 27124
rect 16574 27112 16580 27124
rect 12308 27084 12802 27112
rect 12308 27072 12314 27084
rect 6840 27044 6868 27072
rect 6656 27016 6868 27044
rect 6656 26985 6684 27016
rect 7190 27004 7196 27056
rect 7248 27044 7254 27056
rect 7248 27016 7406 27044
rect 7248 27004 7254 27016
rect 6641 26979 6699 26985
rect 6641 26945 6653 26979
rect 6687 26945 6699 26979
rect 6641 26939 6699 26945
rect 10413 26979 10471 26985
rect 10413 26945 10425 26979
rect 10459 26976 10471 26979
rect 11624 26976 11652 27072
rect 12242 26979 12300 26985
rect 12242 26976 12254 26979
rect 10459 26948 11652 26976
rect 12176 26948 12254 26976
rect 10459 26945 10471 26948
rect 10413 26939 10471 26945
rect 6914 26868 6920 26920
rect 6972 26868 6978 26920
rect 11422 26868 11428 26920
rect 11480 26908 11486 26920
rect 11974 26908 11980 26920
rect 11480 26880 11980 26908
rect 11480 26868 11486 26880
rect 11974 26868 11980 26880
rect 12032 26908 12038 26920
rect 12176 26908 12204 26948
rect 12242 26945 12254 26948
rect 12288 26945 12300 26979
rect 12242 26939 12300 26945
rect 12342 26936 12348 26988
rect 12400 26976 12406 26988
rect 12774 26985 12802 27084
rect 14384 27084 16580 27112
rect 12529 26979 12587 26985
rect 12400 26948 12445 26976
rect 12400 26936 12406 26948
rect 12529 26945 12541 26979
rect 12575 26945 12587 26979
rect 12529 26939 12587 26945
rect 12621 26979 12679 26985
rect 12621 26945 12633 26979
rect 12667 26945 12679 26979
rect 12621 26939 12679 26945
rect 12759 26979 12817 26985
rect 12759 26945 12771 26979
rect 12805 26976 12817 26979
rect 14384 26976 14412 27084
rect 16574 27072 16580 27084
rect 16632 27072 16638 27124
rect 16666 27072 16672 27124
rect 16724 27072 16730 27124
rect 16942 27072 16948 27124
rect 17000 27072 17006 27124
rect 17218 27072 17224 27124
rect 17276 27072 17282 27124
rect 17310 27072 17316 27124
rect 17368 27072 17374 27124
rect 18049 27115 18107 27121
rect 18049 27081 18061 27115
rect 18095 27112 18107 27115
rect 18506 27112 18512 27124
rect 18095 27084 18512 27112
rect 18095 27081 18107 27084
rect 18049 27075 18107 27081
rect 18506 27072 18512 27084
rect 18564 27072 18570 27124
rect 18690 27072 18696 27124
rect 18748 27072 18754 27124
rect 18785 27115 18843 27121
rect 18785 27081 18797 27115
rect 18831 27112 18843 27115
rect 18966 27112 18972 27124
rect 18831 27084 18972 27112
rect 18831 27081 18843 27084
rect 18785 27075 18843 27081
rect 18966 27072 18972 27084
rect 19024 27072 19030 27124
rect 22480 27084 26288 27112
rect 12805 26948 14412 26976
rect 14449 27001 14507 27007
rect 15470 27004 15476 27056
rect 15528 27004 15534 27056
rect 14449 26967 14461 27001
rect 14495 26988 14507 27001
rect 14449 26961 14464 26967
rect 12805 26945 12817 26948
rect 12759 26939 12817 26945
rect 12032 26880 12204 26908
rect 12032 26868 12038 26880
rect 8570 26840 8576 26852
rect 7944 26812 8576 26840
rect 7650 26732 7656 26784
rect 7708 26772 7714 26784
rect 7944 26772 7972 26812
rect 8570 26800 8576 26812
rect 8628 26800 8634 26852
rect 11882 26800 11888 26852
rect 11940 26840 11946 26852
rect 12342 26840 12348 26852
rect 11940 26812 12348 26840
rect 11940 26800 11946 26812
rect 12342 26800 12348 26812
rect 12400 26840 12406 26852
rect 12544 26840 12572 26939
rect 12400 26812 12572 26840
rect 12636 26908 12664 26939
rect 14458 26936 14464 26961
rect 14516 26936 14522 26988
rect 14918 26936 14924 26988
rect 14976 26936 14982 26988
rect 15654 26936 15660 26988
rect 15712 26936 15718 26988
rect 16853 26979 16911 26985
rect 16853 26945 16865 26979
rect 16899 26945 16911 26979
rect 16853 26939 16911 26945
rect 12636 26880 14412 26908
rect 12400 26800 12406 26812
rect 7708 26744 7972 26772
rect 7708 26732 7714 26744
rect 8386 26732 8392 26784
rect 8444 26772 8450 26784
rect 12636 26772 12664 26880
rect 8444 26744 12664 26772
rect 8444 26732 8450 26744
rect 12894 26732 12900 26784
rect 12952 26732 12958 26784
rect 14274 26732 14280 26784
rect 14332 26732 14338 26784
rect 14384 26772 14412 26880
rect 14642 26868 14648 26920
rect 14700 26868 14706 26920
rect 14734 26868 14740 26920
rect 14792 26868 14798 26920
rect 14553 26843 14611 26849
rect 14553 26809 14565 26843
rect 14599 26840 14611 26843
rect 15102 26840 15108 26852
rect 14599 26812 15108 26840
rect 14599 26809 14611 26812
rect 14553 26803 14611 26809
rect 15102 26800 15108 26812
rect 15160 26800 15166 26852
rect 15378 26800 15384 26852
rect 15436 26800 15442 26852
rect 16868 26840 16896 26939
rect 17034 26936 17040 26988
rect 17092 26936 17098 26988
rect 17236 26976 17264 27072
rect 17328 27044 17356 27072
rect 17328 27016 17816 27044
rect 17788 26985 17816 27016
rect 17681 26979 17739 26985
rect 17681 26976 17693 26979
rect 17236 26948 17693 26976
rect 17681 26945 17693 26948
rect 17727 26945 17739 26979
rect 17681 26939 17739 26945
rect 17773 26979 17831 26985
rect 17773 26945 17785 26979
rect 17819 26945 17831 26979
rect 18708 26976 18736 27072
rect 22480 27053 22508 27084
rect 22465 27047 22523 27053
rect 22465 27044 22477 27047
rect 21744 27016 22477 27044
rect 21744 26988 21772 27016
rect 22465 27013 22477 27016
rect 22511 27013 22523 27047
rect 23474 27044 23480 27056
rect 22465 27007 22523 27013
rect 22664 27016 23480 27044
rect 19153 26979 19211 26985
rect 19153 26976 19165 26979
rect 18708 26948 19165 26976
rect 17773 26939 17831 26945
rect 19153 26945 19165 26948
rect 19199 26945 19211 26979
rect 19153 26939 19211 26945
rect 21726 26936 21732 26988
rect 21784 26936 21790 26988
rect 22370 26936 22376 26988
rect 22428 26936 22434 26988
rect 22557 26979 22615 26985
rect 22557 26945 22569 26979
rect 22603 26976 22615 26979
rect 22664 26976 22692 27016
rect 23474 27004 23480 27016
rect 23532 27004 23538 27056
rect 26260 27044 26288 27084
rect 26326 27072 26332 27124
rect 26384 27112 26390 27124
rect 26973 27115 27031 27121
rect 26973 27112 26985 27115
rect 26384 27084 26985 27112
rect 26384 27072 26390 27084
rect 26973 27081 26985 27084
rect 27019 27081 27031 27115
rect 26973 27075 27031 27081
rect 27798 27072 27804 27124
rect 27856 27072 27862 27124
rect 28626 27072 28632 27124
rect 28684 27112 28690 27124
rect 28684 27084 28948 27112
rect 28684 27072 28690 27084
rect 26418 27044 26424 27056
rect 26260 27016 26424 27044
rect 26418 27004 26424 27016
rect 26476 27004 26482 27056
rect 27816 27044 27844 27072
rect 27540 27016 27844 27044
rect 22603 26948 22692 26976
rect 22741 26979 22799 26985
rect 22603 26945 22615 26948
rect 22557 26939 22615 26945
rect 22741 26945 22753 26979
rect 22787 26976 22799 26979
rect 24946 26976 24952 26988
rect 22787 26948 24952 26976
rect 22787 26945 22799 26948
rect 22741 26939 22799 26945
rect 16942 26868 16948 26920
rect 17000 26908 17006 26920
rect 18506 26908 18512 26920
rect 17000 26880 18512 26908
rect 17000 26868 17006 26880
rect 18506 26868 18512 26880
rect 18564 26868 18570 26920
rect 18966 26868 18972 26920
rect 19024 26908 19030 26920
rect 19061 26911 19119 26917
rect 19061 26908 19073 26911
rect 19024 26880 19073 26908
rect 19024 26868 19030 26880
rect 19061 26877 19073 26880
rect 19107 26877 19119 26911
rect 19061 26871 19119 26877
rect 20070 26868 20076 26920
rect 20128 26908 20134 26920
rect 22756 26908 22784 26939
rect 24946 26936 24952 26948
rect 25004 26936 25010 26988
rect 26694 26976 26700 26988
rect 26160 26948 26700 26976
rect 20128 26880 22784 26908
rect 20128 26868 20134 26880
rect 24854 26868 24860 26920
rect 24912 26908 24918 26920
rect 26160 26917 26188 26948
rect 26694 26936 26700 26948
rect 26752 26936 26758 26988
rect 27540 26985 27568 27016
rect 27157 26979 27215 26985
rect 27157 26976 27169 26979
rect 26804 26948 27169 26976
rect 26145 26911 26203 26917
rect 26145 26908 26157 26911
rect 24912 26880 26157 26908
rect 24912 26868 24918 26880
rect 26145 26877 26157 26880
rect 26191 26877 26203 26911
rect 26145 26871 26203 26877
rect 26329 26911 26387 26917
rect 26329 26877 26341 26911
rect 26375 26877 26387 26911
rect 26329 26871 26387 26877
rect 17126 26840 17132 26852
rect 16868 26812 17132 26840
rect 17126 26800 17132 26812
rect 17184 26800 17190 26852
rect 17218 26800 17224 26852
rect 17276 26840 17282 26852
rect 21910 26840 21916 26852
rect 17276 26812 21916 26840
rect 17276 26800 17282 26812
rect 21910 26800 21916 26812
rect 21968 26800 21974 26852
rect 15396 26772 15424 26800
rect 14384 26744 15424 26772
rect 17678 26732 17684 26784
rect 17736 26732 17742 26784
rect 18138 26732 18144 26784
rect 18196 26772 18202 26784
rect 18598 26772 18604 26784
rect 18196 26744 18604 26772
rect 18196 26732 18202 26744
rect 18598 26732 18604 26744
rect 18656 26772 18662 26784
rect 18969 26775 19027 26781
rect 18969 26772 18981 26775
rect 18656 26744 18981 26772
rect 18656 26732 18662 26744
rect 18969 26741 18981 26744
rect 19015 26741 19027 26775
rect 18969 26735 19027 26741
rect 19610 26732 19616 26784
rect 19668 26772 19674 26784
rect 20714 26772 20720 26784
rect 19668 26744 20720 26772
rect 19668 26732 19674 26744
rect 20714 26732 20720 26744
rect 20772 26732 20778 26784
rect 22186 26732 22192 26784
rect 22244 26732 22250 26784
rect 26344 26772 26372 26871
rect 26804 26849 26832 26948
rect 27157 26945 27169 26948
rect 27203 26945 27215 26979
rect 27157 26939 27215 26945
rect 27525 26979 27583 26985
rect 27525 26945 27537 26979
rect 27571 26945 27583 26979
rect 27525 26939 27583 26945
rect 27801 26911 27859 26917
rect 27801 26877 27813 26911
rect 27847 26908 27859 26911
rect 27890 26908 27896 26920
rect 27847 26880 27896 26908
rect 27847 26877 27859 26880
rect 27801 26871 27859 26877
rect 27890 26868 27896 26880
rect 27948 26868 27954 26920
rect 28920 26908 28948 27084
rect 29638 27072 29644 27124
rect 29696 27072 29702 27124
rect 29822 27112 29828 27124
rect 29748 27084 29828 27112
rect 29656 27044 29684 27072
rect 29748 27053 29776 27084
rect 29822 27072 29828 27084
rect 29880 27072 29886 27124
rect 31570 27112 31576 27124
rect 30852 27084 31576 27112
rect 29472 27016 29684 27044
rect 29733 27047 29791 27053
rect 29472 26985 29500 27016
rect 29733 27013 29745 27047
rect 29779 27013 29791 27047
rect 29733 27007 29791 27013
rect 29457 26979 29515 26985
rect 29457 26945 29469 26979
rect 29503 26945 29515 26979
rect 29457 26939 29515 26945
rect 30852 26908 30880 27084
rect 31570 27072 31576 27084
rect 31628 27112 31634 27124
rect 34054 27112 34060 27124
rect 31628 27084 34060 27112
rect 31628 27072 31634 27084
rect 34054 27072 34060 27084
rect 34112 27112 34118 27124
rect 34112 27084 34836 27112
rect 34112 27072 34118 27084
rect 33594 27044 33600 27056
rect 33428 27016 33600 27044
rect 31665 26979 31723 26985
rect 31665 26945 31677 26979
rect 31711 26976 31723 26979
rect 32122 26976 32128 26988
rect 31711 26948 32128 26976
rect 31711 26945 31723 26948
rect 31665 26939 31723 26945
rect 32122 26936 32128 26948
rect 32180 26936 32186 26988
rect 33134 26936 33140 26988
rect 33192 26936 33198 26988
rect 33428 26985 33456 27016
rect 33594 27004 33600 27016
rect 33652 27004 33658 27056
rect 33413 26979 33471 26985
rect 33413 26945 33425 26979
rect 33459 26945 33471 26979
rect 34808 26976 34836 27084
rect 35986 26976 35992 26988
rect 34808 26962 35992 26976
rect 34822 26948 35992 26962
rect 33413 26939 33471 26945
rect 35986 26936 35992 26948
rect 36044 26936 36050 26988
rect 33689 26911 33747 26917
rect 33689 26908 33701 26911
rect 28920 26880 30880 26908
rect 33336 26880 33701 26908
rect 29472 26852 29500 26880
rect 26789 26843 26847 26849
rect 26789 26809 26801 26843
rect 26835 26809 26847 26843
rect 26789 26803 26847 26809
rect 29454 26800 29460 26852
rect 29512 26800 29518 26852
rect 33336 26849 33364 26880
rect 33689 26877 33701 26880
rect 33735 26877 33747 26911
rect 33689 26871 33747 26877
rect 35434 26868 35440 26920
rect 35492 26868 35498 26920
rect 33321 26843 33379 26849
rect 33321 26809 33333 26843
rect 33367 26809 33379 26843
rect 33321 26803 33379 26809
rect 27338 26772 27344 26784
rect 26344 26744 27344 26772
rect 27338 26732 27344 26744
rect 27396 26732 27402 26784
rect 28258 26732 28264 26784
rect 28316 26772 28322 26784
rect 29273 26775 29331 26781
rect 29273 26772 29285 26775
rect 28316 26744 29285 26772
rect 28316 26732 28322 26744
rect 29273 26741 29285 26744
rect 29319 26741 29331 26775
rect 29273 26735 29331 26741
rect 30098 26732 30104 26784
rect 30156 26772 30162 26784
rect 31205 26775 31263 26781
rect 31205 26772 31217 26775
rect 30156 26744 31217 26772
rect 30156 26732 30162 26744
rect 31205 26741 31217 26744
rect 31251 26741 31263 26775
rect 31205 26735 31263 26741
rect 31386 26732 31392 26784
rect 31444 26772 31450 26784
rect 31481 26775 31539 26781
rect 31481 26772 31493 26775
rect 31444 26744 31493 26772
rect 31444 26732 31450 26744
rect 31481 26741 31493 26744
rect 31527 26741 31539 26775
rect 31481 26735 31539 26741
rect 1104 26682 38272 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 38272 26682
rect 1104 26608 38272 26630
rect 6914 26528 6920 26580
rect 6972 26568 6978 26580
rect 7745 26571 7803 26577
rect 7745 26568 7757 26571
rect 6972 26540 7757 26568
rect 6972 26528 6978 26540
rect 7745 26537 7757 26540
rect 7791 26537 7803 26571
rect 11146 26568 11152 26580
rect 7745 26531 7803 26537
rect 7852 26540 11152 26568
rect 7650 26460 7656 26512
rect 7708 26460 7714 26512
rect 7561 26435 7619 26441
rect 7561 26401 7573 26435
rect 7607 26432 7619 26435
rect 7668 26432 7696 26460
rect 7607 26404 7696 26432
rect 7607 26401 7619 26404
rect 7561 26395 7619 26401
rect 4522 26324 4528 26376
rect 4580 26324 4586 26376
rect 4617 26367 4675 26373
rect 4617 26333 4629 26367
rect 4663 26364 4675 26367
rect 4801 26367 4859 26373
rect 4801 26364 4813 26367
rect 4663 26336 4813 26364
rect 4663 26333 4675 26336
rect 4617 26327 4675 26333
rect 4801 26333 4813 26336
rect 4847 26333 4859 26367
rect 4801 26327 4859 26333
rect 6825 26367 6883 26373
rect 6825 26333 6837 26367
rect 6871 26364 6883 26367
rect 7285 26367 7343 26373
rect 7285 26364 7297 26367
rect 6871 26336 7297 26364
rect 6871 26333 6883 26336
rect 6825 26327 6883 26333
rect 7285 26333 7297 26336
rect 7331 26364 7343 26367
rect 7852 26364 7880 26540
rect 11146 26528 11152 26540
rect 11204 26528 11210 26580
rect 12894 26528 12900 26580
rect 12952 26528 12958 26580
rect 13817 26571 13875 26577
rect 13817 26537 13829 26571
rect 13863 26568 13875 26571
rect 14274 26568 14280 26580
rect 13863 26540 14280 26568
rect 13863 26537 13875 26540
rect 13817 26531 13875 26537
rect 14274 26528 14280 26540
rect 14332 26528 14338 26580
rect 14461 26571 14519 26577
rect 14461 26537 14473 26571
rect 14507 26568 14519 26571
rect 14642 26568 14648 26580
rect 14507 26540 14648 26568
rect 14507 26537 14519 26540
rect 14461 26531 14519 26537
rect 14642 26528 14648 26540
rect 14700 26528 14706 26580
rect 15102 26528 15108 26580
rect 15160 26528 15166 26580
rect 15286 26528 15292 26580
rect 15344 26568 15350 26580
rect 17405 26571 17463 26577
rect 15344 26540 17356 26568
rect 15344 26528 15350 26540
rect 8021 26503 8079 26509
rect 8021 26469 8033 26503
rect 8067 26469 8079 26503
rect 8021 26463 8079 26469
rect 7331 26336 7880 26364
rect 7929 26367 7987 26373
rect 7331 26333 7343 26336
rect 7285 26327 7343 26333
rect 7929 26333 7941 26367
rect 7975 26364 7987 26367
rect 8036 26364 8064 26463
rect 8386 26460 8392 26512
rect 8444 26460 8450 26512
rect 9582 26460 9588 26512
rect 9640 26460 9646 26512
rect 8404 26373 8432 26460
rect 8570 26392 8576 26444
rect 8628 26392 8634 26444
rect 7975 26336 8064 26364
rect 8389 26367 8447 26373
rect 7975 26333 7987 26336
rect 7929 26327 7987 26333
rect 8389 26333 8401 26367
rect 8435 26333 8447 26367
rect 8389 26327 8447 26333
rect 9125 26367 9183 26373
rect 9125 26333 9137 26367
rect 9171 26364 9183 26367
rect 9600 26364 9628 26460
rect 9171 26336 9628 26364
rect 9171 26333 9183 26336
rect 9125 26327 9183 26333
rect 12342 26324 12348 26376
rect 12400 26364 12406 26376
rect 12618 26364 12624 26376
rect 12400 26336 12624 26364
rect 12400 26324 12406 26336
rect 12618 26324 12624 26336
rect 12676 26324 12682 26376
rect 12912 26364 12940 26528
rect 17218 26500 17224 26512
rect 15028 26472 17224 26500
rect 14274 26392 14280 26444
rect 14332 26432 14338 26444
rect 14332 26404 14688 26432
rect 14332 26392 14338 26404
rect 13541 26367 13599 26373
rect 13541 26364 13553 26367
rect 12912 26336 13553 26364
rect 13541 26333 13553 26336
rect 13587 26333 13599 26367
rect 13541 26327 13599 26333
rect 13630 26324 13636 26376
rect 13688 26324 13694 26376
rect 13814 26324 13820 26376
rect 13872 26364 13878 26376
rect 14660 26373 14688 26404
rect 14826 26392 14832 26444
rect 14884 26392 14890 26444
rect 13909 26367 13967 26373
rect 13909 26364 13921 26367
rect 13872 26336 13921 26364
rect 13872 26324 13878 26336
rect 13909 26333 13921 26336
rect 13955 26364 13967 26367
rect 14645 26367 14703 26373
rect 13955 26336 14596 26364
rect 13955 26333 13967 26336
rect 13909 26327 13967 26333
rect 5077 26299 5135 26305
rect 5077 26265 5089 26299
rect 5123 26296 5135 26299
rect 5350 26296 5356 26308
rect 5123 26268 5356 26296
rect 5123 26265 5135 26268
rect 5077 26259 5135 26265
rect 5350 26256 5356 26268
rect 5408 26256 5414 26308
rect 5534 26296 5540 26308
rect 5460 26268 5540 26296
rect 3878 26188 3884 26240
rect 3936 26228 3942 26240
rect 5460 26228 5488 26268
rect 5534 26256 5540 26268
rect 5592 26256 5598 26308
rect 7190 26296 7196 26308
rect 6840 26268 7196 26296
rect 5994 26228 6000 26240
rect 3936 26200 6000 26228
rect 3936 26188 3942 26200
rect 5994 26188 6000 26200
rect 6052 26228 6058 26240
rect 6840 26228 6868 26268
rect 7190 26256 7196 26268
rect 7248 26256 7254 26308
rect 7377 26299 7435 26305
rect 7377 26265 7389 26299
rect 7423 26296 7435 26299
rect 7423 26268 8432 26296
rect 7423 26265 7435 26268
rect 7377 26259 7435 26265
rect 6052 26200 6868 26228
rect 6052 26188 6058 26200
rect 6914 26188 6920 26240
rect 6972 26188 6978 26240
rect 8404 26228 8432 26268
rect 8478 26256 8484 26308
rect 8536 26256 8542 26308
rect 11146 26296 11152 26308
rect 8588 26268 11152 26296
rect 8588 26228 8616 26268
rect 11146 26256 11152 26268
rect 11204 26256 11210 26308
rect 13357 26299 13415 26305
rect 13357 26265 13369 26299
rect 13403 26296 13415 26299
rect 14458 26296 14464 26308
rect 13403 26268 14464 26296
rect 13403 26265 13415 26268
rect 13357 26259 13415 26265
rect 14458 26256 14464 26268
rect 14516 26256 14522 26308
rect 14568 26296 14596 26336
rect 14645 26333 14657 26367
rect 14691 26333 14703 26367
rect 14645 26327 14703 26333
rect 14737 26367 14795 26373
rect 14737 26333 14749 26367
rect 14783 26364 14795 26367
rect 14844 26364 14872 26392
rect 15028 26373 15056 26472
rect 17218 26460 17224 26472
rect 17276 26460 17282 26512
rect 17328 26500 17356 26540
rect 17405 26537 17417 26571
rect 17451 26568 17463 26571
rect 17678 26568 17684 26580
rect 17451 26540 17684 26568
rect 17451 26537 17463 26540
rect 17405 26531 17463 26537
rect 17678 26528 17684 26540
rect 17736 26528 17742 26580
rect 18046 26528 18052 26580
rect 18104 26568 18110 26580
rect 27801 26571 27859 26577
rect 18104 26540 27752 26568
rect 18104 26528 18110 26540
rect 17586 26500 17592 26512
rect 17328 26472 17592 26500
rect 17586 26460 17592 26472
rect 17644 26460 17650 26512
rect 18322 26460 18328 26512
rect 18380 26500 18386 26512
rect 19334 26500 19340 26512
rect 18380 26472 19340 26500
rect 18380 26460 18386 26472
rect 19334 26460 19340 26472
rect 19392 26460 19398 26512
rect 20898 26460 20904 26512
rect 20956 26460 20962 26512
rect 21361 26503 21419 26509
rect 21361 26469 21373 26503
rect 21407 26500 21419 26503
rect 22646 26500 22652 26512
rect 21407 26472 22652 26500
rect 21407 26469 21419 26472
rect 21361 26463 21419 26469
rect 22646 26460 22652 26472
rect 22704 26460 22710 26512
rect 15102 26392 15108 26444
rect 15160 26432 15166 26444
rect 15160 26404 15332 26432
rect 15160 26392 15166 26404
rect 15304 26373 15332 26404
rect 15378 26392 15384 26444
rect 15436 26392 15442 26444
rect 20346 26432 20352 26444
rect 15672 26404 20352 26432
rect 15013 26367 15071 26373
rect 14783 26336 14964 26364
rect 14783 26333 14795 26336
rect 14737 26327 14795 26333
rect 14829 26299 14887 26305
rect 14568 26268 14688 26296
rect 14660 26240 14688 26268
rect 14829 26265 14841 26299
rect 14875 26265 14887 26299
rect 14936 26296 14964 26336
rect 15013 26333 15025 26367
rect 15059 26333 15071 26367
rect 15013 26327 15071 26333
rect 15289 26367 15347 26373
rect 15289 26333 15301 26367
rect 15335 26333 15347 26367
rect 15289 26327 15347 26333
rect 15396 26305 15424 26392
rect 15473 26367 15531 26373
rect 15473 26333 15485 26367
rect 15519 26364 15531 26367
rect 15562 26364 15568 26376
rect 15519 26336 15568 26364
rect 15519 26333 15531 26336
rect 15473 26327 15531 26333
rect 15562 26324 15568 26336
rect 15620 26324 15626 26376
rect 15672 26373 15700 26404
rect 15657 26367 15715 26373
rect 15657 26333 15669 26367
rect 15703 26333 15715 26367
rect 16209 26367 16267 26373
rect 16209 26364 16221 26367
rect 15657 26327 15715 26333
rect 15764 26336 16221 26364
rect 15381 26299 15439 26305
rect 14936 26268 15240 26296
rect 14829 26259 14887 26265
rect 8404 26200 8616 26228
rect 8662 26188 8668 26240
rect 8720 26228 8726 26240
rect 9033 26231 9091 26237
rect 9033 26228 9045 26231
rect 8720 26200 9045 26228
rect 8720 26188 8726 26200
rect 9033 26197 9045 26200
rect 9079 26197 9091 26231
rect 9033 26191 9091 26197
rect 14642 26188 14648 26240
rect 14700 26188 14706 26240
rect 14844 26228 14872 26259
rect 15102 26228 15108 26240
rect 14844 26200 15108 26228
rect 15102 26188 15108 26200
rect 15160 26188 15166 26240
rect 15212 26228 15240 26268
rect 15381 26265 15393 26299
rect 15427 26265 15439 26299
rect 15381 26259 15439 26265
rect 15764 26228 15792 26336
rect 16209 26333 16221 26336
rect 16255 26333 16267 26367
rect 16209 26327 16267 26333
rect 16850 26324 16856 26376
rect 16908 26324 16914 26376
rect 17144 26373 17172 26404
rect 20346 26392 20352 26404
rect 20404 26392 20410 26444
rect 20916 26432 20944 26460
rect 21266 26432 21272 26444
rect 20548 26404 20944 26432
rect 21105 26404 21272 26432
rect 17129 26367 17187 26373
rect 17129 26333 17141 26367
rect 17175 26333 17187 26367
rect 17129 26327 17187 26333
rect 17218 26324 17224 26376
rect 17276 26324 17282 26376
rect 18690 26324 18696 26376
rect 18748 26364 18754 26376
rect 18966 26364 18972 26376
rect 18748 26336 18972 26364
rect 18748 26324 18754 26336
rect 18966 26324 18972 26336
rect 19024 26364 19030 26376
rect 19242 26364 19248 26376
rect 19024 26336 19248 26364
rect 19024 26324 19030 26336
rect 19242 26324 19248 26336
rect 19300 26324 19306 26376
rect 19334 26324 19340 26376
rect 19392 26364 19398 26376
rect 19702 26364 19708 26376
rect 19392 26336 19708 26364
rect 19392 26324 19398 26336
rect 19702 26324 19708 26336
rect 19760 26324 19766 26376
rect 16025 26299 16083 26305
rect 16025 26265 16037 26299
rect 16071 26265 16083 26299
rect 16025 26259 16083 26265
rect 16393 26299 16451 26305
rect 16393 26265 16405 26299
rect 16439 26296 16451 26299
rect 17037 26299 17095 26305
rect 17037 26296 17049 26299
rect 16439 26268 17049 26296
rect 16439 26265 16451 26268
rect 16393 26259 16451 26265
rect 17037 26265 17049 26268
rect 17083 26265 17095 26299
rect 20162 26296 20168 26308
rect 17037 26259 17095 26265
rect 17236 26268 20168 26296
rect 15212 26200 15792 26228
rect 16040 26228 16068 26259
rect 16482 26228 16488 26240
rect 16040 26200 16488 26228
rect 16482 26188 16488 26200
rect 16540 26228 16546 26240
rect 16758 26228 16764 26240
rect 16540 26200 16764 26228
rect 16540 26188 16546 26200
rect 16758 26188 16764 26200
rect 16816 26228 16822 26240
rect 17236 26228 17264 26268
rect 20162 26256 20168 26268
rect 20220 26296 20226 26308
rect 20257 26299 20315 26305
rect 20257 26296 20269 26299
rect 20220 26268 20269 26296
rect 20220 26256 20226 26268
rect 20257 26265 20269 26268
rect 20303 26265 20315 26299
rect 20257 26259 20315 26265
rect 20346 26256 20352 26308
rect 20404 26296 20410 26308
rect 20441 26299 20499 26305
rect 20441 26296 20453 26299
rect 20404 26268 20453 26296
rect 20404 26256 20410 26268
rect 20441 26265 20453 26268
rect 20487 26265 20499 26299
rect 20441 26259 20499 26265
rect 16816 26200 17264 26228
rect 16816 26188 16822 26200
rect 18966 26188 18972 26240
rect 19024 26228 19030 26240
rect 20548 26228 20576 26404
rect 20809 26367 20867 26373
rect 20809 26333 20821 26367
rect 20855 26364 20867 26367
rect 21105 26364 21133 26404
rect 21266 26392 21272 26404
rect 21324 26392 21330 26444
rect 20855 26336 21133 26364
rect 21177 26367 21235 26373
rect 20855 26333 20867 26336
rect 20809 26327 20867 26333
rect 21177 26333 21189 26367
rect 21223 26364 21235 26367
rect 22002 26364 22008 26376
rect 21223 26336 22008 26364
rect 21223 26333 21235 26336
rect 21177 26327 21235 26333
rect 22002 26324 22008 26336
rect 22060 26324 22066 26376
rect 22370 26324 22376 26376
rect 22428 26364 22434 26376
rect 23569 26367 23627 26373
rect 23569 26364 23581 26367
rect 22428 26336 23581 26364
rect 22428 26324 22434 26336
rect 23569 26333 23581 26336
rect 23615 26364 23627 26367
rect 23750 26364 23756 26376
rect 23615 26336 23756 26364
rect 23615 26333 23627 26336
rect 23569 26327 23627 26333
rect 23750 26324 23756 26336
rect 23808 26324 23814 26376
rect 23845 26367 23903 26373
rect 23845 26333 23857 26367
rect 23891 26364 23903 26367
rect 24486 26364 24492 26376
rect 23891 26336 24492 26364
rect 23891 26333 23903 26336
rect 23845 26327 23903 26333
rect 24486 26324 24492 26336
rect 24544 26324 24550 26376
rect 24578 26324 24584 26376
rect 24636 26364 24642 26376
rect 25332 26364 25360 26540
rect 25961 26503 26019 26509
rect 25961 26469 25973 26503
rect 26007 26469 26019 26503
rect 25961 26463 26019 26469
rect 25498 26392 25504 26444
rect 25556 26432 25562 26444
rect 25976 26432 26004 26463
rect 26786 26460 26792 26512
rect 26844 26500 26850 26512
rect 27522 26500 27528 26512
rect 26844 26472 27528 26500
rect 26844 26460 26850 26472
rect 27522 26460 27528 26472
rect 27580 26460 27586 26512
rect 27724 26500 27752 26540
rect 27801 26537 27813 26571
rect 27847 26568 27859 26571
rect 28166 26568 28172 26580
rect 27847 26540 28172 26568
rect 27847 26537 27859 26540
rect 27801 26531 27859 26537
rect 28166 26528 28172 26540
rect 28224 26528 28230 26580
rect 30006 26528 30012 26580
rect 30064 26568 30070 26580
rect 30285 26571 30343 26577
rect 30285 26568 30297 26571
rect 30064 26540 30297 26568
rect 30064 26528 30070 26540
rect 30285 26537 30297 26540
rect 30331 26537 30343 26571
rect 30285 26531 30343 26537
rect 31128 26540 33088 26568
rect 30742 26500 30748 26512
rect 27724 26472 30748 26500
rect 30742 26460 30748 26472
rect 30800 26500 30806 26512
rect 31128 26500 31156 26540
rect 30800 26472 31156 26500
rect 33060 26500 33088 26540
rect 33134 26528 33140 26580
rect 33192 26568 33198 26580
rect 33229 26571 33287 26577
rect 33229 26568 33241 26571
rect 33192 26540 33241 26568
rect 33192 26528 33198 26540
rect 33229 26537 33241 26540
rect 33275 26537 33287 26571
rect 35434 26568 35440 26580
rect 33229 26531 33287 26537
rect 33704 26540 35440 26568
rect 33704 26500 33732 26540
rect 35434 26528 35440 26540
rect 35492 26528 35498 26580
rect 33060 26472 33732 26500
rect 30800 26460 30806 26472
rect 25556 26404 25820 26432
rect 25976 26404 26556 26432
rect 25556 26392 25562 26404
rect 25409 26367 25467 26373
rect 25409 26364 25421 26367
rect 24636 26336 24992 26364
rect 25332 26336 25421 26364
rect 24636 26324 24642 26336
rect 20625 26299 20683 26305
rect 20625 26265 20637 26299
rect 20671 26296 20683 26299
rect 20993 26299 21051 26305
rect 20993 26296 21005 26299
rect 20671 26268 21005 26296
rect 20671 26265 20683 26268
rect 20625 26259 20683 26265
rect 20993 26265 21005 26268
rect 21039 26265 21051 26299
rect 20993 26259 21051 26265
rect 21085 26299 21143 26305
rect 21085 26265 21097 26299
rect 21131 26265 21143 26299
rect 21085 26259 21143 26265
rect 19024 26200 20576 26228
rect 19024 26188 19030 26200
rect 20806 26188 20812 26240
rect 20864 26228 20870 26240
rect 21100 26228 21128 26259
rect 23014 26256 23020 26308
rect 23072 26296 23078 26308
rect 23385 26299 23443 26305
rect 23385 26296 23397 26299
rect 23072 26268 23397 26296
rect 23072 26256 23078 26268
rect 23385 26265 23397 26268
rect 23431 26265 23443 26299
rect 23385 26259 23443 26265
rect 24854 26256 24860 26308
rect 24912 26256 24918 26308
rect 24964 26296 24992 26336
rect 25409 26333 25421 26336
rect 25455 26333 25467 26367
rect 25682 26364 25688 26376
rect 25409 26327 25467 26333
rect 25516 26336 25688 26364
rect 25516 26296 25544 26336
rect 25682 26324 25688 26336
rect 25740 26324 25746 26376
rect 25792 26373 25820 26404
rect 25777 26367 25835 26373
rect 25777 26333 25789 26367
rect 25823 26333 25835 26367
rect 25777 26327 25835 26333
rect 26240 26345 26298 26351
rect 26240 26311 26252 26345
rect 26286 26311 26298 26345
rect 26326 26324 26332 26376
rect 26384 26324 26390 26376
rect 26528 26373 26556 26404
rect 27614 26392 27620 26444
rect 27672 26432 27678 26444
rect 27982 26432 27988 26444
rect 27672 26404 27988 26432
rect 27672 26392 27678 26404
rect 27982 26392 27988 26404
rect 28040 26432 28046 26444
rect 28353 26435 28411 26441
rect 28353 26432 28365 26435
rect 28040 26404 28365 26432
rect 28040 26392 28046 26404
rect 28353 26401 28365 26404
rect 28399 26432 28411 26435
rect 29641 26435 29699 26441
rect 29641 26432 29653 26435
rect 28399 26404 29653 26432
rect 28399 26401 28411 26404
rect 28353 26395 28411 26401
rect 29641 26401 29653 26404
rect 29687 26432 29699 26435
rect 30282 26432 30288 26444
rect 29687 26404 30288 26432
rect 29687 26401 29699 26404
rect 29641 26395 29699 26401
rect 30282 26392 30288 26404
rect 30340 26392 30346 26444
rect 30466 26392 30472 26444
rect 30524 26392 30530 26444
rect 31297 26435 31355 26441
rect 31297 26401 31309 26435
rect 31343 26432 31355 26435
rect 31386 26432 31392 26444
rect 31343 26404 31392 26432
rect 31343 26401 31355 26404
rect 31297 26395 31355 26401
rect 31386 26392 31392 26404
rect 31444 26392 31450 26444
rect 31846 26392 31852 26444
rect 31904 26432 31910 26444
rect 33045 26435 33103 26441
rect 33045 26432 33057 26435
rect 31904 26404 33057 26432
rect 31904 26392 31910 26404
rect 33045 26401 33057 26404
rect 33091 26401 33103 26435
rect 33045 26395 33103 26401
rect 26513 26367 26571 26373
rect 26513 26333 26525 26367
rect 26559 26333 26571 26367
rect 26513 26327 26571 26333
rect 26602 26324 26608 26376
rect 26660 26324 26666 26376
rect 29825 26367 29883 26373
rect 29825 26364 29837 26367
rect 26712 26336 29837 26364
rect 26240 26308 26298 26311
rect 24964 26268 25544 26296
rect 25593 26299 25651 26305
rect 25593 26265 25605 26299
rect 25639 26296 25651 26299
rect 26142 26296 26148 26308
rect 25639 26268 26148 26296
rect 25639 26265 25651 26268
rect 25593 26259 25651 26265
rect 21542 26228 21548 26240
rect 20864 26200 21548 26228
rect 20864 26188 20870 26200
rect 21542 26188 21548 26200
rect 21600 26188 21606 26240
rect 23750 26188 23756 26240
rect 23808 26188 23814 26240
rect 24872 26228 24900 26256
rect 25608 26228 25636 26259
rect 26142 26256 26148 26268
rect 26200 26256 26206 26308
rect 26234 26256 26240 26308
rect 26292 26256 26298 26308
rect 26344 26296 26372 26324
rect 26712 26296 26740 26336
rect 29825 26333 29837 26336
rect 29871 26364 29883 26367
rect 30098 26364 30104 26376
rect 29871 26336 30104 26364
rect 29871 26333 29883 26336
rect 29825 26327 29883 26333
rect 30098 26324 30104 26336
rect 30156 26324 30162 26376
rect 30484 26364 30512 26392
rect 30745 26367 30803 26373
rect 30745 26364 30757 26367
rect 30484 26336 30757 26364
rect 30745 26333 30757 26336
rect 30791 26333 30803 26367
rect 30745 26327 30803 26333
rect 30837 26367 30895 26373
rect 30837 26333 30849 26367
rect 30883 26364 30895 26367
rect 31021 26367 31079 26373
rect 31021 26364 31033 26367
rect 30883 26336 31033 26364
rect 30883 26333 30895 26336
rect 30837 26327 30895 26333
rect 31021 26333 31033 26336
rect 31067 26333 31079 26367
rect 31021 26327 31079 26333
rect 33597 26367 33655 26373
rect 33597 26333 33609 26367
rect 33643 26364 33655 26367
rect 33704 26364 33732 26472
rect 34885 26503 34943 26509
rect 34885 26469 34897 26503
rect 34931 26469 34943 26503
rect 34885 26463 34943 26469
rect 33870 26392 33876 26444
rect 33928 26392 33934 26444
rect 34900 26432 34928 26463
rect 35253 26435 35311 26441
rect 35253 26432 35265 26435
rect 34900 26404 35265 26432
rect 35253 26401 35265 26404
rect 35299 26401 35311 26435
rect 35253 26395 35311 26401
rect 33643 26336 33732 26364
rect 33643 26333 33655 26336
rect 33597 26327 33655 26333
rect 34698 26324 34704 26376
rect 34756 26324 34762 26376
rect 34974 26324 34980 26376
rect 35032 26324 35038 26376
rect 26344 26268 26740 26296
rect 28258 26256 28264 26308
rect 28316 26256 28322 26308
rect 29917 26299 29975 26305
rect 29917 26265 29929 26299
rect 29963 26265 29975 26299
rect 29917 26259 29975 26265
rect 25682 26228 25688 26240
rect 24872 26200 25688 26228
rect 25682 26188 25688 26200
rect 25740 26188 25746 26240
rect 26050 26188 26056 26240
rect 26108 26188 26114 26240
rect 27338 26188 27344 26240
rect 27396 26228 27402 26240
rect 28166 26228 28172 26240
rect 27396 26200 28172 26228
rect 27396 26188 27402 26200
rect 28166 26188 28172 26200
rect 28224 26188 28230 26240
rect 29086 26188 29092 26240
rect 29144 26228 29150 26240
rect 29932 26228 29960 26259
rect 31570 26256 31576 26308
rect 31628 26296 31634 26308
rect 31628 26268 31786 26296
rect 31628 26256 31634 26268
rect 35986 26256 35992 26308
rect 36044 26256 36050 26308
rect 36630 26256 36636 26308
rect 36688 26296 36694 26308
rect 37001 26299 37059 26305
rect 37001 26296 37013 26299
rect 36688 26268 37013 26296
rect 36688 26256 36694 26268
rect 37001 26265 37013 26268
rect 37047 26265 37059 26299
rect 37001 26259 37059 26265
rect 30006 26228 30012 26240
rect 29144 26200 30012 26228
rect 29144 26188 29150 26200
rect 30006 26188 30012 26200
rect 30064 26188 30070 26240
rect 30282 26188 30288 26240
rect 30340 26228 30346 26240
rect 31662 26228 31668 26240
rect 30340 26200 31668 26228
rect 30340 26188 30346 26200
rect 31662 26188 31668 26200
rect 31720 26228 31726 26240
rect 33226 26228 33232 26240
rect 31720 26200 33232 26228
rect 31720 26188 31726 26200
rect 33226 26188 33232 26200
rect 33284 26188 33290 26240
rect 33686 26188 33692 26240
rect 33744 26188 33750 26240
rect 1104 26138 38272 26160
rect 1104 26086 4874 26138
rect 4926 26086 4938 26138
rect 4990 26086 5002 26138
rect 5054 26086 5066 26138
rect 5118 26086 5130 26138
rect 5182 26086 35594 26138
rect 35646 26086 35658 26138
rect 35710 26086 35722 26138
rect 35774 26086 35786 26138
rect 35838 26086 35850 26138
rect 35902 26086 38272 26138
rect 1104 26064 38272 26086
rect 5350 25984 5356 26036
rect 5408 26024 5414 26036
rect 5445 26027 5503 26033
rect 5445 26024 5457 26027
rect 5408 25996 5457 26024
rect 5408 25984 5414 25996
rect 5445 25993 5457 25996
rect 5491 25993 5503 26027
rect 5445 25987 5503 25993
rect 6914 25984 6920 26036
rect 6972 25984 6978 26036
rect 14734 25984 14740 26036
rect 14792 25984 14798 26036
rect 15562 25984 15568 26036
rect 15620 26024 15626 26036
rect 15930 26024 15936 26036
rect 15620 25996 15936 26024
rect 15620 25984 15626 25996
rect 15930 25984 15936 25996
rect 15988 25984 15994 26036
rect 16393 26027 16451 26033
rect 16393 25993 16405 26027
rect 16439 26024 16451 26027
rect 17126 26024 17132 26036
rect 16439 25996 17132 26024
rect 16439 25993 16451 25996
rect 16393 25987 16451 25993
rect 17126 25984 17132 25996
rect 17184 25984 17190 26036
rect 19061 26027 19119 26033
rect 19061 25993 19073 26027
rect 19107 26024 19119 26027
rect 19426 26024 19432 26036
rect 19107 25996 19432 26024
rect 19107 25993 19119 25996
rect 19061 25987 19119 25993
rect 19426 25984 19432 25996
rect 19484 25984 19490 26036
rect 20070 26024 20076 26036
rect 19637 25996 20076 26024
rect 3878 25956 3884 25968
rect 3252 25928 3884 25956
rect 3252 25900 3280 25928
rect 3878 25916 3884 25928
rect 3936 25956 3942 25968
rect 3936 25928 4094 25956
rect 3936 25916 3942 25928
rect 1762 25848 1768 25900
rect 1820 25848 1826 25900
rect 3050 25848 3056 25900
rect 3108 25848 3114 25900
rect 3234 25848 3240 25900
rect 3292 25848 3298 25900
rect 5629 25891 5687 25897
rect 5629 25857 5641 25891
rect 5675 25888 5687 25891
rect 6932 25888 6960 25984
rect 14752 25956 14780 25984
rect 18322 25956 18328 25968
rect 14752 25928 18328 25956
rect 18322 25916 18328 25928
rect 18380 25956 18386 25968
rect 18785 25959 18843 25965
rect 18785 25956 18797 25959
rect 18380 25928 18797 25956
rect 18380 25916 18386 25928
rect 18785 25925 18797 25928
rect 18831 25925 18843 25959
rect 18785 25919 18843 25925
rect 18877 25959 18935 25965
rect 18877 25925 18889 25959
rect 18923 25956 18935 25959
rect 18966 25956 18972 25968
rect 18923 25928 18972 25956
rect 18923 25925 18935 25928
rect 18877 25919 18935 25925
rect 18966 25916 18972 25928
rect 19024 25916 19030 25968
rect 19150 25916 19156 25968
rect 19208 25916 19214 25968
rect 19521 25959 19579 25965
rect 19521 25925 19533 25959
rect 19567 25925 19579 25959
rect 19521 25919 19579 25925
rect 5675 25860 6960 25888
rect 5675 25857 5687 25860
rect 5629 25851 5687 25857
rect 10042 25848 10048 25900
rect 10100 25848 10106 25900
rect 13814 25848 13820 25900
rect 13872 25888 13878 25900
rect 16209 25891 16267 25897
rect 16209 25888 16221 25891
rect 13872 25860 16221 25888
rect 13872 25848 13878 25860
rect 16209 25857 16221 25860
rect 16255 25857 16267 25891
rect 16209 25851 16267 25857
rect 17126 25848 17132 25900
rect 17184 25888 17190 25900
rect 17862 25888 17868 25900
rect 17184 25860 17868 25888
rect 17184 25848 17190 25860
rect 17862 25848 17868 25860
rect 17920 25848 17926 25900
rect 18046 25848 18052 25900
rect 18104 25888 18110 25900
rect 18690 25888 18696 25900
rect 18104 25860 18696 25888
rect 18104 25848 18110 25860
rect 18690 25848 18696 25860
rect 18748 25848 18754 25900
rect 1854 25780 1860 25832
rect 1912 25820 1918 25832
rect 3329 25823 3387 25829
rect 3329 25820 3341 25823
rect 1912 25792 3341 25820
rect 1912 25780 1918 25792
rect 3329 25789 3341 25792
rect 3375 25789 3387 25823
rect 3329 25783 3387 25789
rect 3602 25780 3608 25832
rect 3660 25780 3666 25832
rect 8662 25780 8668 25832
rect 8720 25780 8726 25832
rect 8938 25780 8944 25832
rect 8996 25780 9002 25832
rect 11974 25780 11980 25832
rect 12032 25820 12038 25832
rect 13538 25820 13544 25832
rect 12032 25792 13544 25820
rect 12032 25780 12038 25792
rect 13538 25780 13544 25792
rect 13596 25780 13602 25832
rect 14642 25780 14648 25832
rect 14700 25820 14706 25832
rect 17402 25820 17408 25832
rect 14700 25792 17408 25820
rect 14700 25780 14706 25792
rect 17402 25780 17408 25792
rect 17460 25780 17466 25832
rect 18984 25820 19012 25916
rect 18616 25792 19012 25820
rect 19168 25820 19196 25916
rect 19334 25897 19340 25900
rect 19291 25891 19340 25897
rect 19291 25857 19303 25891
rect 19337 25857 19340 25891
rect 19291 25851 19340 25857
rect 19334 25848 19340 25851
rect 19392 25848 19398 25900
rect 19426 25848 19432 25900
rect 19484 25848 19490 25900
rect 19525 25820 19553 25919
rect 19637 25897 19665 25996
rect 20070 25984 20076 25996
rect 20128 25984 20134 26036
rect 20806 26024 20812 26036
rect 20180 25996 20812 26024
rect 20180 25968 20208 25996
rect 20806 25984 20812 25996
rect 20864 25984 20870 26036
rect 23106 25984 23112 26036
rect 23164 25984 23170 26036
rect 23750 25984 23756 26036
rect 23808 26024 23814 26036
rect 23937 26027 23995 26033
rect 23937 26024 23949 26027
rect 23808 25996 23949 26024
rect 23808 25984 23814 25996
rect 23937 25993 23949 25996
rect 23983 25993 23995 26027
rect 23937 25987 23995 25993
rect 25225 26027 25283 26033
rect 25225 25993 25237 26027
rect 25271 26024 25283 26027
rect 25314 26024 25320 26036
rect 25271 25996 25320 26024
rect 25271 25993 25283 25996
rect 25225 25987 25283 25993
rect 25314 25984 25320 25996
rect 25372 25984 25378 26036
rect 25866 25984 25872 26036
rect 25924 25984 25930 26036
rect 26142 25984 26148 26036
rect 26200 25984 26206 26036
rect 32030 26024 32036 26036
rect 26528 25996 32036 26024
rect 20162 25916 20168 25968
rect 20220 25916 20226 25968
rect 20622 25916 20628 25968
rect 20680 25916 20686 25968
rect 20898 25916 20904 25968
rect 20956 25956 20962 25968
rect 23124 25956 23152 25984
rect 25884 25956 25912 25984
rect 26160 25956 26188 25984
rect 20956 25928 23060 25956
rect 23124 25928 23428 25956
rect 20956 25916 20962 25928
rect 19637 25891 19707 25897
rect 19637 25860 19661 25891
rect 19649 25857 19661 25860
rect 19695 25857 19707 25891
rect 19649 25851 19707 25857
rect 19794 25848 19800 25900
rect 19852 25848 19858 25900
rect 19886 25848 19892 25900
rect 19944 25888 19950 25900
rect 20346 25888 20352 25900
rect 19944 25860 20352 25888
rect 19944 25848 19950 25860
rect 20346 25848 20352 25860
rect 20404 25888 20410 25900
rect 20441 25891 20499 25897
rect 20441 25888 20453 25891
rect 20404 25860 20453 25888
rect 20404 25848 20410 25860
rect 20441 25857 20453 25860
rect 20487 25857 20499 25891
rect 20441 25851 20499 25857
rect 20717 25891 20775 25897
rect 20717 25857 20729 25891
rect 20763 25857 20775 25891
rect 20717 25851 20775 25857
rect 20809 25891 20867 25897
rect 20809 25857 20821 25891
rect 20855 25888 20867 25891
rect 20990 25888 20996 25900
rect 20855 25860 20996 25888
rect 20855 25857 20867 25860
rect 20809 25851 20867 25857
rect 19168 25792 19553 25820
rect 18616 25764 18644 25792
rect 20070 25780 20076 25832
rect 20128 25820 20134 25832
rect 20732 25820 20760 25851
rect 20990 25848 20996 25860
rect 21048 25848 21054 25900
rect 22186 25848 22192 25900
rect 22244 25888 22250 25900
rect 22465 25891 22523 25897
rect 22465 25888 22477 25891
rect 22244 25860 22477 25888
rect 22244 25848 22250 25860
rect 22465 25857 22477 25860
rect 22511 25857 22523 25891
rect 22465 25851 22523 25857
rect 22646 25848 22652 25900
rect 22704 25848 22710 25900
rect 22741 25891 22799 25897
rect 22741 25857 22753 25891
rect 22787 25857 22799 25891
rect 22741 25851 22799 25857
rect 20128 25792 20760 25820
rect 21008 25820 21036 25848
rect 21008 25792 22692 25820
rect 20128 25780 20134 25792
rect 14826 25712 14832 25764
rect 14884 25752 14890 25764
rect 18230 25752 18236 25764
rect 14884 25724 18236 25752
rect 14884 25712 14890 25724
rect 18230 25712 18236 25724
rect 18288 25712 18294 25764
rect 18509 25755 18567 25761
rect 18509 25721 18521 25755
rect 18555 25721 18567 25755
rect 18509 25715 18567 25721
rect 934 25644 940 25696
rect 992 25684 998 25696
rect 1489 25687 1547 25693
rect 1489 25684 1501 25687
rect 992 25656 1501 25684
rect 992 25644 998 25656
rect 1489 25653 1501 25656
rect 1535 25653 1547 25687
rect 1489 25647 1547 25653
rect 2866 25644 2872 25696
rect 2924 25644 2930 25696
rect 4706 25644 4712 25696
rect 4764 25684 4770 25696
rect 5077 25687 5135 25693
rect 5077 25684 5089 25687
rect 4764 25656 5089 25684
rect 4764 25644 4770 25656
rect 5077 25653 5089 25656
rect 5123 25653 5135 25687
rect 5077 25647 5135 25653
rect 9674 25644 9680 25696
rect 9732 25684 9738 25696
rect 10413 25687 10471 25693
rect 10413 25684 10425 25687
rect 9732 25656 10425 25684
rect 9732 25644 9738 25656
rect 10413 25653 10425 25656
rect 10459 25684 10471 25687
rect 12986 25684 12992 25696
rect 10459 25656 12992 25684
rect 10459 25653 10471 25656
rect 10413 25647 10471 25653
rect 12986 25644 12992 25656
rect 13044 25644 13050 25696
rect 15010 25644 15016 25696
rect 15068 25684 15074 25696
rect 18524 25684 18552 25715
rect 18598 25712 18604 25764
rect 18656 25712 18662 25764
rect 19334 25752 19340 25764
rect 18708 25724 19340 25752
rect 18708 25684 18736 25724
rect 19334 25712 19340 25724
rect 19392 25712 19398 25764
rect 20732 25752 20760 25792
rect 22664 25764 22692 25792
rect 21174 25752 21180 25764
rect 20732 25724 21180 25752
rect 21174 25712 21180 25724
rect 21232 25712 21238 25764
rect 22554 25712 22560 25764
rect 22612 25712 22618 25764
rect 22646 25712 22652 25764
rect 22704 25712 22710 25764
rect 22756 25752 22784 25851
rect 23032 25820 23060 25928
rect 23400 25900 23428 25928
rect 24596 25928 26004 25956
rect 26160 25928 26280 25956
rect 23106 25848 23112 25900
rect 23164 25848 23170 25900
rect 23382 25848 23388 25900
rect 23440 25848 23446 25900
rect 23845 25891 23903 25897
rect 23845 25857 23857 25891
rect 23891 25888 23903 25891
rect 24302 25888 24308 25900
rect 23891 25860 24308 25888
rect 23891 25857 23903 25860
rect 23845 25851 23903 25857
rect 24302 25848 24308 25860
rect 24360 25848 24366 25900
rect 24596 25897 24624 25928
rect 24581 25891 24639 25897
rect 24581 25857 24593 25891
rect 24627 25888 24639 25891
rect 24670 25888 24676 25900
rect 24627 25860 24676 25888
rect 24627 25857 24639 25860
rect 24581 25851 24639 25857
rect 24670 25848 24676 25860
rect 24728 25848 24734 25900
rect 24762 25848 24768 25900
rect 24820 25848 24826 25900
rect 24857 25891 24915 25897
rect 24857 25857 24869 25891
rect 24903 25857 24915 25891
rect 24857 25851 24915 25857
rect 24949 25891 25007 25897
rect 24949 25857 24961 25891
rect 24995 25857 25007 25891
rect 24949 25851 25007 25857
rect 23753 25823 23811 25829
rect 23753 25820 23765 25823
rect 23032 25792 23765 25820
rect 23753 25789 23765 25792
rect 23799 25789 23811 25823
rect 23753 25783 23811 25789
rect 23477 25755 23535 25761
rect 23477 25752 23489 25755
rect 22756 25724 23489 25752
rect 23477 25721 23489 25724
rect 23523 25721 23535 25755
rect 23768 25752 23796 25783
rect 24026 25780 24032 25832
rect 24084 25820 24090 25832
rect 24213 25823 24271 25829
rect 24213 25820 24225 25823
rect 24084 25792 24225 25820
rect 24084 25780 24090 25792
rect 24213 25789 24225 25792
rect 24259 25789 24271 25823
rect 24320 25820 24348 25848
rect 24872 25820 24900 25851
rect 24320 25792 24900 25820
rect 24213 25783 24271 25789
rect 24486 25752 24492 25764
rect 23768 25724 24492 25752
rect 23477 25715 23535 25721
rect 24486 25712 24492 25724
rect 24544 25752 24550 25764
rect 24964 25752 24992 25851
rect 25314 25848 25320 25900
rect 25372 25888 25378 25900
rect 25498 25888 25504 25900
rect 25372 25860 25504 25888
rect 25372 25848 25378 25860
rect 25498 25848 25504 25860
rect 25556 25848 25562 25900
rect 25593 25891 25651 25897
rect 25593 25857 25605 25891
rect 25639 25857 25651 25891
rect 25593 25851 25651 25857
rect 25608 25820 25636 25851
rect 25682 25848 25688 25900
rect 25740 25848 25746 25900
rect 25976 25897 26004 25928
rect 25869 25891 25927 25897
rect 25869 25857 25881 25891
rect 25915 25857 25927 25891
rect 25869 25851 25927 25857
rect 25961 25891 26019 25897
rect 25961 25857 25973 25891
rect 26007 25857 26019 25891
rect 25961 25851 26019 25857
rect 24544 25724 24992 25752
rect 25240 25792 25636 25820
rect 25884 25820 25912 25851
rect 26050 25848 26056 25900
rect 26108 25888 26114 25900
rect 26252 25897 26280 25928
rect 26528 25900 26556 25996
rect 32030 25984 32036 25996
rect 32088 25984 32094 26036
rect 32122 25984 32128 26036
rect 32180 25984 32186 26036
rect 32674 25984 32680 26036
rect 32732 26024 32738 26036
rect 33318 26024 33324 26036
rect 32732 25996 33324 26024
rect 32732 25984 32738 25996
rect 33318 25984 33324 25996
rect 33376 25984 33382 26036
rect 34330 25984 34336 26036
rect 34388 25984 34394 26036
rect 34698 25984 34704 26036
rect 34756 26024 34762 26036
rect 34793 26027 34851 26033
rect 34793 26024 34805 26027
rect 34756 25996 34805 26024
rect 34756 25984 34762 25996
rect 34793 25993 34805 25996
rect 34839 25993 34851 26027
rect 34793 25987 34851 25993
rect 34974 25984 34980 26036
rect 35032 26024 35038 26036
rect 35253 26027 35311 26033
rect 35253 26024 35265 26027
rect 35032 25996 35265 26024
rect 35032 25984 35038 25996
rect 35253 25993 35265 25996
rect 35299 25993 35311 26027
rect 35253 25987 35311 25993
rect 30006 25916 30012 25968
rect 30064 25956 30070 25968
rect 31941 25959 31999 25965
rect 30064 25928 31892 25956
rect 30064 25916 30070 25928
rect 26145 25891 26203 25897
rect 26145 25888 26157 25891
rect 26108 25860 26157 25888
rect 26108 25848 26114 25860
rect 26145 25857 26157 25860
rect 26191 25857 26203 25891
rect 26145 25851 26203 25857
rect 26237 25891 26295 25897
rect 26237 25857 26249 25891
rect 26283 25857 26295 25891
rect 26237 25851 26295 25857
rect 26329 25891 26387 25897
rect 26329 25857 26341 25891
rect 26375 25888 26387 25891
rect 26510 25888 26516 25900
rect 26375 25860 26516 25888
rect 26375 25857 26387 25860
rect 26329 25851 26387 25857
rect 26510 25848 26516 25860
rect 26568 25848 26574 25900
rect 27890 25848 27896 25900
rect 27948 25888 27954 25900
rect 31481 25891 31539 25897
rect 31481 25888 31493 25891
rect 27948 25860 31493 25888
rect 27948 25848 27954 25860
rect 31481 25857 31493 25860
rect 31527 25857 31539 25891
rect 31481 25851 31539 25857
rect 31573 25891 31631 25897
rect 31573 25857 31585 25891
rect 31619 25857 31631 25891
rect 31573 25851 31631 25857
rect 26418 25820 26424 25832
rect 25884 25792 26424 25820
rect 24544 25712 24550 25724
rect 15068 25656 18736 25684
rect 15068 25644 15074 25656
rect 19150 25644 19156 25696
rect 19208 25644 19214 25696
rect 19426 25644 19432 25696
rect 19484 25684 19490 25696
rect 20162 25684 20168 25696
rect 19484 25656 20168 25684
rect 19484 25644 19490 25656
rect 20162 25644 20168 25656
rect 20220 25644 20226 25696
rect 20990 25644 20996 25696
rect 21048 25644 21054 25696
rect 21082 25644 21088 25696
rect 21140 25684 21146 25696
rect 21634 25684 21640 25696
rect 21140 25656 21640 25684
rect 21140 25644 21146 25656
rect 21634 25644 21640 25656
rect 21692 25644 21698 25696
rect 22278 25644 22284 25696
rect 22336 25644 22342 25696
rect 23842 25644 23848 25696
rect 23900 25684 23906 25696
rect 24121 25687 24179 25693
rect 24121 25684 24133 25687
rect 23900 25656 24133 25684
rect 23900 25644 23906 25656
rect 24121 25653 24133 25656
rect 24167 25653 24179 25687
rect 24121 25647 24179 25653
rect 24302 25644 24308 25696
rect 24360 25684 24366 25696
rect 25240 25684 25268 25792
rect 25608 25752 25636 25792
rect 26418 25780 26424 25792
rect 26476 25780 26482 25832
rect 31588 25820 31616 25851
rect 31754 25848 31760 25900
rect 31812 25848 31818 25900
rect 31864 25888 31892 25928
rect 31941 25925 31953 25959
rect 31987 25956 31999 25959
rect 33686 25956 33692 25968
rect 31987 25928 32996 25956
rect 31987 25925 31999 25928
rect 31941 25919 31999 25925
rect 32968 25897 32996 25928
rect 33060 25928 33692 25956
rect 32493 25891 32551 25897
rect 32493 25888 32505 25891
rect 31864 25860 32505 25888
rect 32493 25857 32505 25860
rect 32539 25888 32551 25891
rect 32953 25891 33011 25897
rect 32539 25860 32904 25888
rect 32539 25857 32551 25860
rect 32493 25851 32551 25857
rect 31846 25820 31852 25832
rect 31588 25792 31852 25820
rect 31846 25780 31852 25792
rect 31904 25820 31910 25832
rect 32585 25823 32643 25829
rect 32585 25820 32597 25823
rect 31904 25792 32597 25820
rect 31904 25780 31910 25792
rect 32585 25789 32597 25792
rect 32631 25789 32643 25823
rect 32585 25783 32643 25789
rect 32674 25780 32680 25832
rect 32732 25780 32738 25832
rect 32876 25820 32904 25860
rect 32953 25857 32965 25891
rect 32999 25857 33011 25891
rect 32953 25851 33011 25857
rect 33060 25820 33088 25928
rect 33686 25916 33692 25928
rect 33744 25916 33750 25968
rect 34348 25956 34376 25984
rect 34348 25928 35112 25956
rect 33137 25891 33195 25897
rect 33137 25857 33149 25891
rect 33183 25857 33195 25891
rect 33137 25851 33195 25857
rect 32876 25792 33088 25820
rect 26326 25752 26332 25764
rect 25608 25724 26332 25752
rect 26326 25712 26332 25724
rect 26384 25712 26390 25764
rect 29086 25752 29092 25764
rect 26528 25724 29092 25752
rect 24360 25656 25268 25684
rect 24360 25644 24366 25656
rect 25314 25644 25320 25696
rect 25372 25644 25378 25696
rect 25498 25644 25504 25696
rect 25556 25684 25562 25696
rect 26528 25684 26556 25724
rect 29086 25712 29092 25724
rect 29144 25712 29150 25764
rect 33152 25752 33180 25851
rect 33226 25848 33232 25900
rect 33284 25848 33290 25900
rect 33321 25891 33379 25897
rect 33321 25857 33333 25891
rect 33367 25888 33379 25891
rect 33704 25888 33732 25916
rect 35084 25897 35112 25928
rect 34333 25891 34391 25897
rect 34333 25888 34345 25891
rect 33367 25860 33640 25888
rect 33704 25860 34345 25888
rect 33367 25857 33379 25860
rect 33321 25851 33379 25857
rect 33612 25752 33640 25860
rect 34333 25857 34345 25860
rect 34379 25857 34391 25891
rect 34333 25851 34391 25857
rect 34425 25891 34483 25897
rect 34425 25857 34437 25891
rect 34471 25857 34483 25891
rect 34425 25851 34483 25857
rect 35069 25891 35127 25897
rect 35069 25857 35081 25891
rect 35115 25888 35127 25891
rect 35161 25891 35219 25897
rect 35161 25888 35173 25891
rect 35115 25860 35173 25888
rect 35115 25857 35127 25860
rect 35069 25851 35127 25857
rect 35161 25857 35173 25860
rect 35207 25857 35219 25891
rect 35161 25851 35219 25857
rect 34146 25780 34152 25832
rect 34204 25780 34210 25832
rect 34440 25820 34468 25851
rect 36630 25848 36636 25900
rect 36688 25848 36694 25900
rect 36648 25820 36676 25848
rect 34440 25792 36676 25820
rect 34440 25752 34468 25792
rect 31312 25724 33180 25752
rect 33244 25724 34468 25752
rect 31312 25696 31340 25724
rect 25556 25656 26556 25684
rect 25556 25644 25562 25656
rect 26602 25644 26608 25696
rect 26660 25644 26666 25696
rect 27798 25644 27804 25696
rect 27856 25684 27862 25696
rect 28718 25684 28724 25696
rect 27856 25656 28724 25684
rect 27856 25644 27862 25656
rect 28718 25644 28724 25656
rect 28776 25644 28782 25696
rect 31294 25644 31300 25696
rect 31352 25644 31358 25696
rect 32030 25644 32036 25696
rect 32088 25684 32094 25696
rect 33244 25684 33272 25724
rect 34698 25712 34704 25764
rect 34756 25752 34762 25764
rect 34977 25755 35035 25761
rect 34977 25752 34989 25755
rect 34756 25724 34989 25752
rect 34756 25712 34762 25724
rect 34977 25721 34989 25724
rect 35023 25721 35035 25755
rect 34977 25715 35035 25721
rect 32088 25656 33272 25684
rect 33597 25687 33655 25693
rect 32088 25644 32094 25656
rect 33597 25653 33609 25687
rect 33643 25684 33655 25687
rect 34790 25684 34796 25696
rect 33643 25656 34796 25684
rect 33643 25653 33655 25656
rect 33597 25647 33655 25653
rect 34790 25644 34796 25656
rect 34848 25644 34854 25696
rect 1104 25594 38272 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 38272 25594
rect 1104 25520 38272 25542
rect 3602 25440 3608 25492
rect 3660 25480 3666 25492
rect 3881 25483 3939 25489
rect 3881 25480 3893 25483
rect 3660 25452 3893 25480
rect 3660 25440 3666 25452
rect 3881 25449 3893 25452
rect 3927 25449 3939 25483
rect 3881 25443 3939 25449
rect 8938 25440 8944 25492
rect 8996 25480 9002 25492
rect 9033 25483 9091 25489
rect 9033 25480 9045 25483
rect 8996 25452 9045 25480
rect 8996 25440 9002 25452
rect 9033 25449 9045 25452
rect 9079 25449 9091 25483
rect 9033 25443 9091 25449
rect 9674 25440 9680 25492
rect 9732 25440 9738 25492
rect 12986 25440 12992 25492
rect 13044 25440 13050 25492
rect 17218 25440 17224 25492
rect 17276 25480 17282 25492
rect 18785 25483 18843 25489
rect 18785 25480 18797 25483
rect 17276 25452 18797 25480
rect 17276 25440 17282 25452
rect 18785 25449 18797 25452
rect 18831 25480 18843 25483
rect 18831 25452 22508 25480
rect 18831 25449 18843 25452
rect 18785 25443 18843 25449
rect 2133 25347 2191 25353
rect 2133 25313 2145 25347
rect 2179 25344 2191 25347
rect 2866 25344 2872 25356
rect 2179 25316 2872 25344
rect 2179 25313 2191 25316
rect 2133 25307 2191 25313
rect 2866 25304 2872 25316
rect 2924 25304 2930 25356
rect 1394 25236 1400 25288
rect 1452 25276 1458 25288
rect 1854 25276 1860 25288
rect 1452 25248 1860 25276
rect 1452 25236 1458 25248
rect 1854 25236 1860 25248
rect 1912 25236 1918 25288
rect 3234 25236 3240 25288
rect 3292 25236 3298 25288
rect 4065 25279 4123 25285
rect 4065 25245 4077 25279
rect 4111 25276 4123 25279
rect 4338 25276 4344 25288
rect 4111 25248 4344 25276
rect 4111 25245 4123 25248
rect 4065 25239 4123 25245
rect 4338 25236 4344 25248
rect 4396 25236 4402 25288
rect 7558 25236 7564 25288
rect 7616 25276 7622 25288
rect 8662 25276 8668 25288
rect 7616 25248 8668 25276
rect 7616 25236 7622 25248
rect 8662 25236 8668 25248
rect 8720 25236 8726 25288
rect 9692 25285 9720 25440
rect 12066 25372 12072 25424
rect 12124 25412 12130 25424
rect 12342 25412 12348 25424
rect 12124 25384 12348 25412
rect 12124 25372 12130 25384
rect 12342 25372 12348 25384
rect 12400 25412 12406 25424
rect 13004 25412 13032 25440
rect 18966 25412 18972 25424
rect 12400 25372 12434 25412
rect 9858 25304 9864 25356
rect 9916 25304 9922 25356
rect 11885 25347 11943 25353
rect 11885 25313 11897 25347
rect 11931 25313 11943 25347
rect 12406 25344 12434 25372
rect 13004 25384 18972 25412
rect 12529 25347 12587 25353
rect 12529 25344 12541 25347
rect 12406 25316 12541 25344
rect 11885 25307 11943 25313
rect 12529 25313 12541 25316
rect 12575 25313 12587 25347
rect 13004 25344 13032 25384
rect 18966 25372 18972 25384
rect 19024 25412 19030 25424
rect 19886 25412 19892 25424
rect 19024 25384 19892 25412
rect 19024 25372 19030 25384
rect 19886 25372 19892 25384
rect 19944 25372 19950 25424
rect 20901 25415 20959 25421
rect 20901 25381 20913 25415
rect 20947 25412 20959 25415
rect 21085 25415 21143 25421
rect 21085 25412 21097 25415
rect 20947 25384 21097 25412
rect 20947 25381 20959 25384
rect 20901 25375 20959 25381
rect 21085 25381 21097 25384
rect 21131 25381 21143 25415
rect 21085 25375 21143 25381
rect 13722 25344 13728 25356
rect 13004 25316 13124 25344
rect 12529 25307 12587 25313
rect 9217 25279 9275 25285
rect 9217 25245 9229 25279
rect 9263 25276 9275 25279
rect 9677 25279 9735 25285
rect 9263 25248 9352 25276
rect 9263 25245 9275 25248
rect 9217 25239 9275 25245
rect 2958 25100 2964 25152
rect 3016 25140 3022 25152
rect 3252 25140 3280 25236
rect 3016 25112 3280 25140
rect 3605 25143 3663 25149
rect 3016 25100 3022 25112
rect 3605 25109 3617 25143
rect 3651 25140 3663 25143
rect 4614 25140 4620 25152
rect 3651 25112 4620 25140
rect 3651 25109 3663 25112
rect 3605 25103 3663 25109
rect 4614 25100 4620 25112
rect 4672 25100 4678 25152
rect 7282 25100 7288 25152
rect 7340 25140 7346 25152
rect 9324 25149 9352 25248
rect 9677 25245 9689 25279
rect 9723 25245 9735 25279
rect 9677 25239 9735 25245
rect 10134 25236 10140 25288
rect 10192 25236 10198 25288
rect 11900 25276 11928 25307
rect 12345 25279 12403 25285
rect 12345 25276 12357 25279
rect 11900 25248 12357 25276
rect 12345 25245 12357 25248
rect 12391 25276 12403 25279
rect 12391 25248 12572 25276
rect 12391 25245 12403 25248
rect 12345 25239 12403 25245
rect 10413 25211 10471 25217
rect 10413 25177 10425 25211
rect 10459 25208 10471 25211
rect 10502 25208 10508 25220
rect 10459 25180 10508 25208
rect 10459 25177 10471 25180
rect 10413 25171 10471 25177
rect 10502 25168 10508 25180
rect 10560 25168 10566 25220
rect 11054 25168 11060 25220
rect 11112 25168 11118 25220
rect 11790 25168 11796 25220
rect 11848 25208 11854 25220
rect 12437 25211 12495 25217
rect 12437 25208 12449 25211
rect 11848 25180 12449 25208
rect 11848 25168 11854 25180
rect 12437 25177 12449 25180
rect 12483 25177 12495 25211
rect 12544 25208 12572 25248
rect 12618 25236 12624 25288
rect 12676 25276 12682 25288
rect 13096 25285 13124 25316
rect 13188 25316 13728 25344
rect 13188 25288 13216 25316
rect 13722 25304 13728 25316
rect 13780 25344 13786 25356
rect 13780 25316 14596 25344
rect 13780 25304 13786 25316
rect 12943 25279 13001 25285
rect 12943 25276 12955 25279
rect 12676 25248 12955 25276
rect 12676 25236 12682 25248
rect 12943 25245 12955 25248
rect 12989 25245 13001 25279
rect 12943 25239 13001 25245
rect 13081 25279 13139 25285
rect 13081 25245 13093 25279
rect 13127 25245 13139 25279
rect 13081 25239 13139 25245
rect 13170 25236 13176 25288
rect 13228 25236 13234 25288
rect 13356 25279 13414 25285
rect 13356 25276 13368 25279
rect 13335 25248 13368 25276
rect 13356 25245 13368 25248
rect 13402 25245 13414 25279
rect 13356 25239 13414 25245
rect 13449 25279 13507 25285
rect 13449 25245 13461 25279
rect 13495 25276 13507 25279
rect 13538 25276 13544 25288
rect 13495 25248 13544 25276
rect 13495 25245 13507 25248
rect 13449 25239 13507 25245
rect 13372 25208 13400 25239
rect 13538 25236 13544 25248
rect 13596 25236 13602 25288
rect 14568 25285 14596 25316
rect 14826 25304 14832 25356
rect 14884 25304 14890 25356
rect 15654 25304 15660 25356
rect 15712 25344 15718 25356
rect 17405 25347 17463 25353
rect 15712 25316 17264 25344
rect 15712 25304 15718 25316
rect 14553 25279 14611 25285
rect 14553 25245 14565 25279
rect 14599 25245 14611 25279
rect 14553 25239 14611 25245
rect 15010 25236 15016 25288
rect 15068 25236 15074 25288
rect 15930 25236 15936 25288
rect 15988 25236 15994 25288
rect 16022 25236 16028 25288
rect 16080 25236 16086 25288
rect 17236 25285 17264 25316
rect 17405 25313 17417 25347
rect 17451 25344 17463 25347
rect 19058 25344 19064 25356
rect 17451 25316 19064 25344
rect 17451 25313 17463 25316
rect 17405 25307 17463 25313
rect 19058 25304 19064 25316
rect 19116 25304 19122 25356
rect 20990 25304 20996 25356
rect 21048 25304 21054 25356
rect 21105 25316 22416 25344
rect 16761 25279 16819 25285
rect 16668 25257 16726 25263
rect 15028 25208 15056 25236
rect 12544 25180 15056 25208
rect 16040 25208 16068 25236
rect 16668 25223 16680 25257
rect 16714 25223 16726 25257
rect 16761 25245 16773 25279
rect 16807 25245 16819 25279
rect 16761 25239 16819 25245
rect 16853 25279 16911 25285
rect 16853 25245 16865 25279
rect 16899 25276 16911 25279
rect 17037 25279 17095 25285
rect 16899 25248 16988 25276
rect 16899 25245 16911 25248
rect 16853 25239 16911 25245
rect 16668 25217 16726 25223
rect 16393 25211 16451 25217
rect 16393 25208 16405 25211
rect 16040 25180 16405 25208
rect 12437 25171 12495 25177
rect 16393 25177 16405 25180
rect 16439 25177 16451 25211
rect 16393 25171 16451 25177
rect 7469 25143 7527 25149
rect 7469 25140 7481 25143
rect 7340 25112 7481 25140
rect 7340 25100 7346 25112
rect 7469 25109 7481 25112
rect 7515 25109 7527 25143
rect 7469 25103 7527 25109
rect 9309 25143 9367 25149
rect 9309 25109 9321 25143
rect 9355 25109 9367 25143
rect 9309 25103 9367 25109
rect 9582 25100 9588 25152
rect 9640 25140 9646 25152
rect 9769 25143 9827 25149
rect 9769 25140 9781 25143
rect 9640 25112 9781 25140
rect 9640 25100 9646 25112
rect 9769 25109 9781 25112
rect 9815 25140 9827 25143
rect 11808 25140 11836 25168
rect 16683 25152 16711 25217
rect 16776 25208 16804 25239
rect 16776 25180 16896 25208
rect 16868 25152 16896 25180
rect 9815 25112 11836 25140
rect 9815 25109 9827 25112
rect 9769 25103 9827 25109
rect 11974 25100 11980 25152
rect 12032 25100 12038 25152
rect 12802 25100 12808 25152
rect 12860 25100 12866 25152
rect 16117 25143 16175 25149
rect 16117 25109 16129 25143
rect 16163 25140 16175 25143
rect 16666 25140 16672 25152
rect 16163 25112 16672 25140
rect 16163 25109 16175 25112
rect 16117 25103 16175 25109
rect 16666 25100 16672 25112
rect 16724 25100 16730 25152
rect 16850 25100 16856 25152
rect 16908 25100 16914 25152
rect 16960 25140 16988 25248
rect 17037 25245 17049 25279
rect 17083 25245 17095 25279
rect 17037 25239 17095 25245
rect 17221 25279 17279 25285
rect 17221 25245 17233 25279
rect 17267 25245 17279 25279
rect 17221 25239 17279 25245
rect 17052 25208 17080 25239
rect 17310 25236 17316 25288
rect 17368 25276 17374 25288
rect 17368 25248 18000 25276
rect 17368 25236 17374 25248
rect 17972 25208 18000 25248
rect 18414 25236 18420 25288
rect 18472 25236 18478 25288
rect 18506 25236 18512 25288
rect 18564 25236 18570 25288
rect 18601 25279 18659 25285
rect 18601 25245 18613 25279
rect 18647 25276 18659 25279
rect 19334 25276 19340 25288
rect 18647 25248 19340 25276
rect 18647 25245 18659 25248
rect 18601 25239 18659 25245
rect 18616 25208 18644 25239
rect 19334 25236 19340 25248
rect 19392 25276 19398 25288
rect 20254 25276 20260 25288
rect 19392 25248 20260 25276
rect 19392 25236 19398 25248
rect 20254 25236 20260 25248
rect 20312 25236 20318 25288
rect 20714 25236 20720 25288
rect 20772 25236 20778 25288
rect 21105 25276 21133 25316
rect 21266 25285 21272 25288
rect 21264 25276 21272 25285
rect 20916 25248 21133 25276
rect 21227 25248 21272 25276
rect 20916 25220 20944 25248
rect 21264 25239 21272 25248
rect 21266 25236 21272 25239
rect 21324 25236 21330 25288
rect 21450 25236 21456 25288
rect 21508 25236 21514 25288
rect 21542 25236 21548 25288
rect 21600 25285 21606 25288
rect 21600 25279 21639 25285
rect 21627 25245 21639 25279
rect 21600 25239 21639 25245
rect 21729 25279 21787 25285
rect 21729 25245 21741 25279
rect 21775 25276 21787 25279
rect 21818 25276 21824 25288
rect 21775 25248 21824 25276
rect 21775 25245 21787 25248
rect 21729 25239 21787 25245
rect 21600 25236 21606 25239
rect 21818 25236 21824 25248
rect 21876 25236 21882 25288
rect 22002 25236 22008 25288
rect 22060 25236 22066 25288
rect 22186 25236 22192 25288
rect 22244 25236 22250 25288
rect 22282 25279 22340 25285
rect 22282 25245 22294 25279
rect 22328 25245 22340 25279
rect 22282 25239 22340 25245
rect 17052 25180 17724 25208
rect 17972 25180 18644 25208
rect 17696 25152 17724 25180
rect 19518 25168 19524 25220
rect 19576 25208 19582 25220
rect 19576 25180 20852 25208
rect 19576 25168 19582 25180
rect 17494 25140 17500 25152
rect 16960 25112 17500 25140
rect 17494 25100 17500 25112
rect 17552 25100 17558 25152
rect 17678 25100 17684 25152
rect 17736 25100 17742 25152
rect 17954 25100 17960 25152
rect 18012 25140 18018 25152
rect 19426 25140 19432 25152
rect 18012 25112 19432 25140
rect 18012 25100 18018 25112
rect 19426 25100 19432 25112
rect 19484 25100 19490 25152
rect 20533 25143 20591 25149
rect 20533 25109 20545 25143
rect 20579 25140 20591 25143
rect 20622 25140 20628 25152
rect 20579 25112 20628 25140
rect 20579 25109 20591 25112
rect 20533 25103 20591 25109
rect 20622 25100 20628 25112
rect 20680 25100 20686 25152
rect 20824 25140 20852 25180
rect 20898 25168 20904 25220
rect 20956 25168 20962 25220
rect 21361 25211 21419 25217
rect 21361 25177 21373 25211
rect 21407 25208 21419 25211
rect 22020 25208 22048 25236
rect 22296 25208 22324 25239
rect 21407 25180 22324 25208
rect 22388 25208 22416 25316
rect 22480 25276 22508 25452
rect 22554 25440 22560 25492
rect 22612 25480 22618 25492
rect 22833 25483 22891 25489
rect 22833 25480 22845 25483
rect 22612 25452 22845 25480
rect 22612 25440 22618 25452
rect 22833 25449 22845 25452
rect 22879 25449 22891 25483
rect 22833 25443 22891 25449
rect 24946 25440 24952 25492
rect 25004 25440 25010 25492
rect 25130 25440 25136 25492
rect 25188 25440 25194 25492
rect 25314 25440 25320 25492
rect 25372 25480 25378 25492
rect 31018 25480 31024 25492
rect 25372 25452 25544 25480
rect 25372 25440 25378 25452
rect 22646 25372 22652 25424
rect 22704 25412 22710 25424
rect 22704 25384 24900 25412
rect 22704 25372 22710 25384
rect 22922 25304 22928 25356
rect 22980 25344 22986 25356
rect 22980 25316 23060 25344
rect 22980 25304 22986 25316
rect 23032 25285 23060 25316
rect 23658 25304 23664 25356
rect 23716 25304 23722 25356
rect 22654 25279 22712 25285
rect 22654 25276 22666 25279
rect 22480 25248 22666 25276
rect 22654 25245 22666 25248
rect 22700 25276 22712 25279
rect 23017 25279 23075 25285
rect 22700 25248 22968 25276
rect 22700 25245 22712 25248
rect 22654 25239 22712 25245
rect 22465 25211 22523 25217
rect 22465 25208 22477 25211
rect 22388 25180 22477 25208
rect 21407 25177 21419 25180
rect 21361 25171 21419 25177
rect 22465 25177 22477 25180
rect 22511 25177 22523 25211
rect 22465 25171 22523 25177
rect 21726 25140 21732 25152
rect 20824 25112 21732 25140
rect 21726 25100 21732 25112
rect 21784 25100 21790 25152
rect 22480 25140 22508 25171
rect 22554 25168 22560 25220
rect 22612 25168 22618 25220
rect 22940 25208 22968 25248
rect 23017 25245 23029 25279
rect 23063 25245 23075 25279
rect 24394 25276 24400 25288
rect 23017 25239 23075 25245
rect 23493 25248 24400 25276
rect 23493 25208 23521 25248
rect 24394 25236 24400 25248
rect 24452 25236 24458 25288
rect 24762 25236 24768 25288
rect 24820 25236 24826 25288
rect 24872 25276 24900 25384
rect 24964 25344 24992 25440
rect 25148 25412 25176 25440
rect 25148 25384 25452 25412
rect 24964 25316 25084 25344
rect 24946 25276 24952 25288
rect 24872 25248 24952 25276
rect 24946 25236 24952 25248
rect 25004 25236 25010 25288
rect 25056 25285 25084 25316
rect 25041 25279 25099 25285
rect 25041 25245 25053 25279
rect 25087 25245 25099 25279
rect 25041 25239 25099 25245
rect 25225 25279 25283 25285
rect 25225 25245 25237 25279
rect 25271 25245 25283 25279
rect 25225 25239 25283 25245
rect 25317 25279 25375 25285
rect 25317 25245 25329 25279
rect 25363 25276 25375 25279
rect 25424 25276 25452 25384
rect 25363 25248 25452 25276
rect 25363 25245 25375 25248
rect 25317 25239 25375 25245
rect 22940 25180 23521 25208
rect 23934 25168 23940 25220
rect 23992 25168 23998 25220
rect 25240 25208 25268 25239
rect 25516 25208 25544 25452
rect 27448 25452 31024 25480
rect 26418 25236 26424 25288
rect 26476 25236 26482 25288
rect 26970 25236 26976 25288
rect 27028 25276 27034 25288
rect 27448 25285 27476 25452
rect 31018 25440 31024 25452
rect 31076 25440 31082 25492
rect 27798 25372 27804 25424
rect 27856 25372 27862 25424
rect 30558 25412 30564 25424
rect 28736 25384 30564 25412
rect 28736 25344 28764 25384
rect 30558 25372 30564 25384
rect 30616 25372 30622 25424
rect 34698 25372 34704 25424
rect 34756 25372 34762 25424
rect 28368 25316 28764 25344
rect 28905 25347 28963 25353
rect 27157 25279 27215 25285
rect 27157 25276 27169 25279
rect 27028 25248 27169 25276
rect 27028 25236 27034 25248
rect 27157 25245 27169 25248
rect 27203 25245 27215 25279
rect 27157 25239 27215 25245
rect 27250 25279 27308 25285
rect 27250 25245 27262 25279
rect 27296 25245 27308 25279
rect 27250 25239 27308 25245
rect 27433 25279 27491 25285
rect 27433 25245 27445 25279
rect 27479 25245 27491 25279
rect 27433 25239 27491 25245
rect 27622 25279 27680 25285
rect 27622 25245 27634 25279
rect 27668 25276 27680 25279
rect 27890 25276 27896 25288
rect 27668 25248 27896 25276
rect 27668 25245 27680 25248
rect 27622 25239 27680 25245
rect 25240 25180 25544 25208
rect 26436 25208 26464 25236
rect 27265 25208 27293 25239
rect 26436 25180 27293 25208
rect 27338 25168 27344 25220
rect 27396 25208 27402 25220
rect 27525 25211 27583 25217
rect 27525 25208 27537 25211
rect 27396 25180 27537 25208
rect 27396 25168 27402 25180
rect 27525 25177 27537 25180
rect 27571 25177 27583 25211
rect 27525 25171 27583 25177
rect 23566 25140 23572 25152
rect 22480 25112 23572 25140
rect 23566 25100 23572 25112
rect 23624 25100 23630 25152
rect 23952 25140 23980 25168
rect 27632 25140 27660 25239
rect 27890 25236 27896 25248
rect 27948 25236 27954 25288
rect 28368 25276 28396 25316
rect 28905 25313 28917 25347
rect 28951 25344 28963 25347
rect 28951 25316 30052 25344
rect 28951 25313 28963 25316
rect 28905 25307 28963 25313
rect 28445 25279 28503 25285
rect 28445 25276 28457 25279
rect 28368 25248 28457 25276
rect 28445 25245 28457 25248
rect 28491 25245 28503 25279
rect 28445 25239 28503 25245
rect 28718 25236 28724 25288
rect 28776 25236 28782 25288
rect 28994 25236 29000 25288
rect 29052 25276 29058 25288
rect 29181 25279 29239 25285
rect 29181 25276 29193 25279
rect 29052 25248 29193 25276
rect 29052 25236 29058 25248
rect 29181 25245 29193 25248
rect 29227 25245 29239 25279
rect 29181 25239 29239 25245
rect 29730 25236 29736 25288
rect 29788 25236 29794 25288
rect 30024 25285 30052 25316
rect 30009 25279 30067 25285
rect 30009 25245 30021 25279
rect 30055 25245 30067 25279
rect 30009 25239 30067 25245
rect 30193 25279 30251 25285
rect 30193 25245 30205 25279
rect 30239 25245 30251 25279
rect 30193 25239 30251 25245
rect 27798 25168 27804 25220
rect 27856 25208 27862 25220
rect 29748 25208 29776 25236
rect 30208 25208 30236 25239
rect 30282 25236 30288 25288
rect 30340 25236 30346 25288
rect 30374 25236 30380 25288
rect 30432 25236 30438 25288
rect 34330 25236 34336 25288
rect 34388 25236 34394 25288
rect 34716 25285 34744 25372
rect 34701 25279 34759 25285
rect 34701 25245 34713 25279
rect 34747 25245 34759 25279
rect 34701 25239 34759 25245
rect 34977 25211 35035 25217
rect 34977 25208 34989 25211
rect 27856 25180 29224 25208
rect 29748 25180 30236 25208
rect 30300 25180 31432 25208
rect 27856 25168 27862 25180
rect 23952 25112 27660 25140
rect 28258 25100 28264 25152
rect 28316 25140 28322 25152
rect 28537 25143 28595 25149
rect 28537 25140 28549 25143
rect 28316 25112 28549 25140
rect 28316 25100 28322 25112
rect 28537 25109 28549 25112
rect 28583 25109 28595 25143
rect 28537 25103 28595 25109
rect 29086 25100 29092 25152
rect 29144 25100 29150 25152
rect 29196 25140 29224 25180
rect 30300 25140 30328 25180
rect 31404 25152 31432 25180
rect 34532 25180 34989 25208
rect 29196 25112 30328 25140
rect 30650 25100 30656 25152
rect 30708 25100 30714 25152
rect 31386 25100 31392 25152
rect 31444 25100 31450 25152
rect 34532 25149 34560 25180
rect 34977 25177 34989 25180
rect 35023 25177 35035 25211
rect 34977 25171 35035 25177
rect 35986 25168 35992 25220
rect 36044 25168 36050 25220
rect 36722 25168 36728 25220
rect 36780 25168 36786 25220
rect 34517 25143 34575 25149
rect 34517 25109 34529 25143
rect 34563 25109 34575 25143
rect 34517 25103 34575 25109
rect 1104 25050 38272 25072
rect 1104 24998 4874 25050
rect 4926 24998 4938 25050
rect 4990 24998 5002 25050
rect 5054 24998 5066 25050
rect 5118 24998 5130 25050
rect 5182 24998 35594 25050
rect 35646 24998 35658 25050
rect 35710 24998 35722 25050
rect 35774 24998 35786 25050
rect 35838 24998 35850 25050
rect 35902 24998 38272 25050
rect 1104 24976 38272 24998
rect 4338 24896 4344 24948
rect 4396 24896 4402 24948
rect 4706 24896 4712 24948
rect 4764 24936 4770 24948
rect 5810 24936 5816 24948
rect 4764 24908 5816 24936
rect 4764 24896 4770 24908
rect 5810 24896 5816 24908
rect 5868 24896 5874 24948
rect 9582 24896 9588 24948
rect 9640 24896 9646 24948
rect 10134 24896 10140 24948
rect 10192 24936 10198 24948
rect 10321 24939 10379 24945
rect 10321 24936 10333 24939
rect 10192 24908 10333 24936
rect 10192 24896 10198 24908
rect 10321 24905 10333 24908
rect 10367 24905 10379 24939
rect 10321 24899 10379 24905
rect 10502 24896 10508 24948
rect 10560 24936 10566 24948
rect 10597 24939 10655 24945
rect 10597 24936 10609 24939
rect 10560 24908 10609 24936
rect 10560 24896 10566 24908
rect 10597 24905 10609 24908
rect 10643 24905 10655 24939
rect 10597 24899 10655 24905
rect 11974 24896 11980 24948
rect 12032 24896 12038 24948
rect 12434 24936 12440 24948
rect 12176 24908 12440 24936
rect 9674 24828 9680 24880
rect 9732 24868 9738 24880
rect 10042 24868 10048 24880
rect 9732 24840 10048 24868
rect 9732 24828 9738 24840
rect 10042 24828 10048 24840
rect 10100 24828 10106 24880
rect 2958 24800 2964 24812
rect 2806 24772 2964 24800
rect 2958 24760 2964 24772
rect 3016 24760 3022 24812
rect 5902 24760 5908 24812
rect 5960 24760 5966 24812
rect 9692 24800 9720 24828
rect 8588 24772 9720 24800
rect 1394 24692 1400 24744
rect 1452 24692 1458 24744
rect 1670 24692 1676 24744
rect 1728 24692 1734 24744
rect 4798 24692 4804 24744
rect 4856 24692 4862 24744
rect 4985 24735 5043 24741
rect 4985 24701 4997 24735
rect 5031 24701 5043 24735
rect 4985 24695 5043 24701
rect 2682 24556 2688 24608
rect 2740 24596 2746 24608
rect 3145 24599 3203 24605
rect 3145 24596 3157 24599
rect 2740 24568 3157 24596
rect 2740 24556 2746 24568
rect 3145 24565 3157 24568
rect 3191 24565 3203 24599
rect 3145 24559 3203 24565
rect 3970 24556 3976 24608
rect 4028 24596 4034 24608
rect 5000 24596 5028 24695
rect 7282 24692 7288 24744
rect 7340 24692 7346 24744
rect 7561 24735 7619 24741
rect 7561 24701 7573 24735
rect 7607 24732 7619 24735
rect 7926 24732 7932 24744
rect 7607 24704 7932 24732
rect 7607 24701 7619 24704
rect 7561 24695 7619 24701
rect 7926 24692 7932 24704
rect 7984 24692 7990 24744
rect 4028 24568 5028 24596
rect 4028 24556 4034 24568
rect 5626 24556 5632 24608
rect 5684 24596 5690 24608
rect 5721 24599 5779 24605
rect 5721 24596 5733 24599
rect 5684 24568 5733 24596
rect 5684 24556 5690 24568
rect 5721 24565 5733 24568
rect 5767 24565 5779 24599
rect 5721 24559 5779 24565
rect 7282 24556 7288 24608
rect 7340 24596 7346 24608
rect 8588 24596 8616 24772
rect 10410 24760 10416 24812
rect 10468 24760 10474 24812
rect 10781 24803 10839 24809
rect 10781 24769 10793 24803
rect 10827 24800 10839 24803
rect 11992 24800 12020 24896
rect 12176 24809 12204 24908
rect 12434 24896 12440 24908
rect 12492 24896 12498 24948
rect 12802 24896 12808 24948
rect 12860 24936 12866 24948
rect 12860 24908 13032 24936
rect 12860 24896 12866 24908
rect 12250 24828 12256 24880
rect 12308 24868 12314 24880
rect 13004 24877 13032 24908
rect 13722 24896 13728 24948
rect 13780 24936 13786 24948
rect 14277 24939 14335 24945
rect 14277 24936 14289 24939
rect 13780 24908 14289 24936
rect 13780 24896 13786 24908
rect 14277 24905 14289 24908
rect 14323 24905 14335 24939
rect 15010 24936 15016 24948
rect 14277 24899 14335 24905
rect 14384 24908 15016 24936
rect 12345 24871 12403 24877
rect 12345 24868 12357 24871
rect 12308 24840 12357 24868
rect 12308 24828 12314 24840
rect 12345 24837 12357 24840
rect 12391 24837 12403 24871
rect 12989 24871 13047 24877
rect 12345 24831 12403 24837
rect 12544 24840 12940 24868
rect 12544 24809 12572 24840
rect 10827 24772 12020 24800
rect 12161 24803 12219 24809
rect 10827 24769 10839 24772
rect 10781 24763 10839 24769
rect 12161 24769 12173 24803
rect 12207 24769 12219 24803
rect 12161 24763 12219 24769
rect 12437 24803 12495 24809
rect 12437 24769 12449 24803
rect 12483 24769 12495 24803
rect 12437 24763 12495 24769
rect 12529 24803 12587 24809
rect 12529 24769 12541 24803
rect 12575 24769 12587 24803
rect 12805 24803 12863 24809
rect 12805 24800 12817 24803
rect 12529 24763 12587 24769
rect 12728 24772 12817 24800
rect 9033 24735 9091 24741
rect 9033 24701 9045 24735
rect 9079 24732 9091 24735
rect 9677 24735 9735 24741
rect 9677 24732 9689 24735
rect 9079 24704 9689 24732
rect 9079 24701 9091 24704
rect 9033 24695 9091 24701
rect 9677 24701 9689 24704
rect 9723 24701 9735 24735
rect 9677 24695 9735 24701
rect 7340 24568 8616 24596
rect 7340 24556 7346 24568
rect 9214 24556 9220 24608
rect 9272 24556 9278 24608
rect 9692 24596 9720 24695
rect 9858 24692 9864 24744
rect 9916 24692 9922 24744
rect 12452 24732 12480 24763
rect 12406 24704 12480 24732
rect 12406 24596 12434 24704
rect 12728 24673 12756 24772
rect 12805 24769 12817 24772
rect 12851 24769 12863 24803
rect 12912 24800 12940 24840
rect 12989 24837 13001 24871
rect 13035 24837 13047 24871
rect 12989 24831 13047 24837
rect 13446 24800 13452 24812
rect 12912 24772 13452 24800
rect 12805 24763 12863 24769
rect 13446 24760 13452 24772
rect 13504 24800 13510 24812
rect 14182 24800 14188 24812
rect 13504 24772 14188 24800
rect 13504 24760 13510 24772
rect 14182 24760 14188 24772
rect 14240 24760 14246 24812
rect 14277 24803 14335 24809
rect 14277 24769 14289 24803
rect 14323 24800 14335 24803
rect 14384 24800 14412 24908
rect 15010 24896 15016 24908
rect 15068 24936 15074 24948
rect 15838 24936 15844 24948
rect 15068 24908 15844 24936
rect 15068 24896 15074 24908
rect 15838 24896 15844 24908
rect 15896 24936 15902 24948
rect 17678 24936 17684 24948
rect 15896 24908 17684 24936
rect 15896 24896 15902 24908
rect 17678 24896 17684 24908
rect 17736 24896 17742 24948
rect 18138 24896 18144 24948
rect 18196 24936 18202 24948
rect 18196 24908 21036 24936
rect 18196 24896 18202 24908
rect 17310 24868 17316 24880
rect 16132 24840 17316 24868
rect 16132 24812 16160 24840
rect 14323 24772 14412 24800
rect 14323 24769 14335 24772
rect 14277 24763 14335 24769
rect 14918 24760 14924 24812
rect 14976 24760 14982 24812
rect 15378 24760 15384 24812
rect 15436 24760 15442 24812
rect 16114 24760 16120 24812
rect 16172 24760 16178 24812
rect 16209 24803 16267 24809
rect 16209 24769 16221 24803
rect 16255 24800 16267 24803
rect 16574 24800 16580 24812
rect 16255 24772 16580 24800
rect 16255 24769 16267 24772
rect 16209 24763 16267 24769
rect 16574 24760 16580 24772
rect 16632 24760 16638 24812
rect 16850 24760 16856 24812
rect 16908 24760 16914 24812
rect 17236 24809 17264 24840
rect 17310 24828 17316 24840
rect 17368 24868 17374 24880
rect 18046 24868 18052 24880
rect 17368 24840 18052 24868
rect 17368 24828 17374 24840
rect 18046 24828 18052 24840
rect 18104 24828 18110 24880
rect 18506 24828 18512 24880
rect 18564 24828 18570 24880
rect 20898 24868 20904 24880
rect 19076 24840 20904 24868
rect 17221 24803 17279 24809
rect 17221 24769 17233 24803
rect 17267 24769 17279 24803
rect 17221 24763 17279 24769
rect 17586 24760 17592 24812
rect 17644 24800 17650 24812
rect 17865 24803 17923 24809
rect 17865 24800 17877 24803
rect 17644 24772 17877 24800
rect 17644 24760 17650 24772
rect 17865 24769 17877 24772
rect 17911 24769 17923 24803
rect 17865 24763 17923 24769
rect 18601 24803 18659 24809
rect 18601 24769 18613 24803
rect 18647 24800 18659 24803
rect 18782 24800 18788 24812
rect 18647 24772 18788 24800
rect 18647 24769 18659 24772
rect 18601 24763 18659 24769
rect 18782 24760 18788 24772
rect 18840 24760 18846 24812
rect 19076 24809 19104 24840
rect 20898 24828 20904 24840
rect 20956 24828 20962 24880
rect 19061 24803 19119 24809
rect 19061 24769 19073 24803
rect 19107 24769 19119 24803
rect 19061 24763 19119 24769
rect 19242 24760 19248 24812
rect 19300 24800 19306 24812
rect 20070 24800 20076 24812
rect 19300 24772 20076 24800
rect 19300 24760 19306 24772
rect 20070 24760 20076 24772
rect 20128 24760 20134 24812
rect 14366 24692 14372 24744
rect 14424 24732 14430 24744
rect 15013 24735 15071 24741
rect 15013 24732 15025 24735
rect 14424 24704 15025 24732
rect 14424 24692 14430 24704
rect 15013 24701 15025 24704
rect 15059 24701 15071 24735
rect 15013 24695 15071 24701
rect 16666 24692 16672 24744
rect 16724 24692 16730 24744
rect 16868 24732 16896 24760
rect 17313 24735 17371 24741
rect 16868 24704 17264 24732
rect 17236 24676 17264 24704
rect 17313 24701 17325 24735
rect 17359 24732 17371 24735
rect 17494 24732 17500 24744
rect 17359 24704 17500 24732
rect 17359 24701 17371 24704
rect 17313 24695 17371 24701
rect 17494 24692 17500 24704
rect 17552 24692 17558 24744
rect 21008 24732 21036 24908
rect 21450 24896 21456 24948
rect 21508 24896 21514 24948
rect 21818 24896 21824 24948
rect 21876 24936 21882 24948
rect 22922 24936 22928 24948
rect 21876 24908 22928 24936
rect 21876 24896 21882 24908
rect 22922 24896 22928 24908
rect 22980 24896 22986 24948
rect 23382 24896 23388 24948
rect 23440 24896 23446 24948
rect 26973 24939 27031 24945
rect 26973 24905 26985 24939
rect 27019 24905 27031 24939
rect 26973 24899 27031 24905
rect 21085 24871 21143 24877
rect 21085 24837 21097 24871
rect 21131 24868 21143 24871
rect 21174 24868 21180 24880
rect 21131 24840 21180 24868
rect 21131 24837 21143 24840
rect 21085 24831 21143 24837
rect 21174 24828 21180 24840
rect 21232 24828 21238 24880
rect 21361 24871 21419 24877
rect 21361 24837 21373 24871
rect 21407 24837 21419 24871
rect 21634 24868 21640 24880
rect 21361 24831 21419 24837
rect 21560 24840 21640 24868
rect 21269 24803 21327 24809
rect 21269 24769 21281 24803
rect 21315 24769 21327 24803
rect 21376 24800 21404 24831
rect 21560 24800 21588 24840
rect 21634 24828 21640 24840
rect 21692 24828 21698 24880
rect 22554 24828 22560 24880
rect 22612 24868 22618 24880
rect 24302 24868 24308 24880
rect 22612 24840 24308 24868
rect 22612 24828 22618 24840
rect 24302 24828 24308 24840
rect 24360 24828 24366 24880
rect 24486 24828 24492 24880
rect 24544 24868 24550 24880
rect 26878 24868 26884 24880
rect 24544 24840 26884 24868
rect 24544 24828 24550 24840
rect 26878 24828 26884 24840
rect 26936 24828 26942 24880
rect 21376 24772 21588 24800
rect 21269 24763 21327 24769
rect 21284 24732 21312 24763
rect 23474 24760 23480 24812
rect 23532 24760 23538 24812
rect 23658 24760 23664 24812
rect 23716 24760 23722 24812
rect 23842 24760 23848 24812
rect 23900 24760 23906 24812
rect 25869 24803 25927 24809
rect 25869 24769 25881 24803
rect 25915 24769 25927 24803
rect 25869 24763 25927 24769
rect 26145 24803 26203 24809
rect 26145 24769 26157 24803
rect 26191 24800 26203 24803
rect 26988 24800 27016 24899
rect 29086 24896 29092 24948
rect 29144 24896 29150 24948
rect 29822 24896 29828 24948
rect 29880 24936 29886 24948
rect 31294 24936 31300 24948
rect 29880 24908 31300 24936
rect 29880 24896 29886 24908
rect 31294 24896 31300 24908
rect 31352 24896 31358 24948
rect 31386 24896 31392 24948
rect 31444 24936 31450 24948
rect 34241 24939 34299 24945
rect 31444 24908 31984 24936
rect 31444 24896 31450 24908
rect 27341 24871 27399 24877
rect 27341 24837 27353 24871
rect 27387 24837 27399 24871
rect 29104 24868 29132 24896
rect 27341 24831 27399 24837
rect 28920 24840 29132 24868
rect 26191 24772 27016 24800
rect 26191 24769 26203 24772
rect 26145 24763 26203 24769
rect 17604 24704 20945 24732
rect 21008 24704 21312 24732
rect 23676 24732 23704 24760
rect 24118 24732 24124 24744
rect 23676 24704 24124 24732
rect 12713 24667 12771 24673
rect 12713 24633 12725 24667
rect 12759 24633 12771 24667
rect 17126 24664 17132 24676
rect 12713 24627 12771 24633
rect 13096 24636 17132 24664
rect 13096 24596 13124 24636
rect 17126 24624 17132 24636
rect 17184 24624 17190 24676
rect 17218 24624 17224 24676
rect 17276 24624 17282 24676
rect 9692 24568 13124 24596
rect 13170 24556 13176 24608
rect 13228 24556 13234 24608
rect 14182 24556 14188 24608
rect 14240 24596 14246 24608
rect 15194 24596 15200 24608
rect 14240 24568 15200 24596
rect 14240 24556 14246 24568
rect 15194 24556 15200 24568
rect 15252 24596 15258 24608
rect 17604 24596 17632 24704
rect 17678 24624 17684 24676
rect 17736 24664 17742 24676
rect 19886 24664 19892 24676
rect 17736 24636 19892 24664
rect 17736 24624 17742 24636
rect 19886 24624 19892 24636
rect 19944 24624 19950 24676
rect 20917 24664 20945 24704
rect 24118 24692 24124 24704
rect 24176 24692 24182 24744
rect 25884 24732 25912 24763
rect 27154 24760 27160 24812
rect 27212 24800 27218 24812
rect 27356 24800 27384 24831
rect 28166 24800 28172 24812
rect 27212 24772 28172 24800
rect 27212 24760 27218 24772
rect 28166 24760 28172 24772
rect 28224 24760 28230 24812
rect 28626 24760 28632 24812
rect 28684 24760 28690 24812
rect 28920 24809 28948 24840
rect 29454 24828 29460 24880
rect 29512 24868 29518 24880
rect 29512 24840 29670 24868
rect 29512 24828 29518 24840
rect 30466 24828 30472 24880
rect 30524 24868 30530 24880
rect 30929 24871 30987 24877
rect 30929 24868 30941 24871
rect 30524 24840 30941 24868
rect 30524 24828 30530 24840
rect 30929 24837 30941 24840
rect 30975 24837 30987 24871
rect 30929 24831 30987 24837
rect 28905 24803 28963 24809
rect 28905 24769 28917 24803
rect 28951 24769 28963 24803
rect 28905 24763 28963 24769
rect 31110 24760 31116 24812
rect 31168 24760 31174 24812
rect 31312 24809 31340 24896
rect 31956 24868 31984 24908
rect 34241 24905 34253 24939
rect 34287 24936 34299 24939
rect 34330 24936 34336 24948
rect 34287 24908 34336 24936
rect 34287 24905 34299 24908
rect 34241 24899 34299 24905
rect 34330 24896 34336 24908
rect 34388 24896 34394 24948
rect 34609 24939 34667 24945
rect 34609 24905 34621 24939
rect 34655 24936 34667 24939
rect 36722 24936 36728 24948
rect 34655 24908 36728 24936
rect 34655 24905 34667 24908
rect 34609 24899 34667 24905
rect 34624 24868 34652 24899
rect 36722 24896 36728 24908
rect 36780 24896 36786 24948
rect 31956 24840 34652 24868
rect 31297 24803 31355 24809
rect 31297 24769 31309 24803
rect 31343 24769 31355 24803
rect 31297 24763 31355 24769
rect 31570 24760 31576 24812
rect 31628 24760 31634 24812
rect 31956 24809 31984 24840
rect 31941 24803 31999 24809
rect 31941 24769 31953 24803
rect 31987 24769 31999 24803
rect 31941 24763 31999 24769
rect 33042 24760 33048 24812
rect 33100 24760 33106 24812
rect 33134 24760 33140 24812
rect 33192 24800 33198 24812
rect 33229 24803 33287 24809
rect 33229 24800 33241 24803
rect 33192 24772 33241 24800
rect 33192 24760 33198 24772
rect 33229 24769 33241 24772
rect 33275 24800 33287 24803
rect 33505 24803 33563 24809
rect 33505 24800 33517 24803
rect 33275 24772 33517 24800
rect 33275 24769 33287 24772
rect 33229 24763 33287 24769
rect 33505 24769 33517 24772
rect 33551 24800 33563 24803
rect 33778 24800 33784 24812
rect 33551 24772 33784 24800
rect 33551 24769 33563 24772
rect 33505 24763 33563 24769
rect 33778 24760 33784 24772
rect 33836 24760 33842 24812
rect 26694 24732 26700 24744
rect 25884 24704 26700 24732
rect 26694 24692 26700 24704
rect 26752 24692 26758 24744
rect 27338 24692 27344 24744
rect 27396 24732 27402 24744
rect 27433 24735 27491 24741
rect 27433 24732 27445 24735
rect 27396 24704 27445 24732
rect 27396 24692 27402 24704
rect 27433 24701 27445 24704
rect 27479 24701 27491 24735
rect 27433 24695 27491 24701
rect 27525 24735 27583 24741
rect 27525 24701 27537 24735
rect 27571 24701 27583 24735
rect 29181 24735 29239 24741
rect 29181 24732 29193 24735
rect 27525 24695 27583 24701
rect 28828 24704 29193 24732
rect 23934 24664 23940 24676
rect 20917 24636 23940 24664
rect 23934 24624 23940 24636
rect 23992 24624 23998 24676
rect 27540 24664 27568 24695
rect 28828 24673 28856 24704
rect 29181 24701 29193 24704
rect 29227 24701 29239 24735
rect 29181 24695 29239 24701
rect 29270 24692 29276 24744
rect 29328 24732 29334 24744
rect 30190 24732 30196 24744
rect 29328 24704 30196 24732
rect 29328 24692 29334 24704
rect 30190 24692 30196 24704
rect 30248 24732 30254 24744
rect 34701 24735 34759 24741
rect 34701 24732 34713 24735
rect 30248 24704 30880 24732
rect 30248 24692 30254 24704
rect 24044 24636 26924 24664
rect 24044 24608 24072 24636
rect 15252 24568 17632 24596
rect 18325 24599 18383 24605
rect 15252 24556 15258 24568
rect 18325 24565 18337 24599
rect 18371 24596 18383 24599
rect 18414 24596 18420 24608
rect 18371 24568 18420 24596
rect 18371 24565 18383 24568
rect 18325 24559 18383 24565
rect 18414 24556 18420 24568
rect 18472 24556 18478 24608
rect 18874 24556 18880 24608
rect 18932 24596 18938 24608
rect 20806 24596 20812 24608
rect 18932 24568 20812 24596
rect 18932 24556 18938 24568
rect 20806 24556 20812 24568
rect 20864 24556 20870 24608
rect 21637 24599 21695 24605
rect 21637 24565 21649 24599
rect 21683 24596 21695 24599
rect 22186 24596 22192 24608
rect 21683 24568 22192 24596
rect 21683 24565 21695 24568
rect 21637 24559 21695 24565
rect 22186 24556 22192 24568
rect 22244 24556 22250 24608
rect 24026 24556 24032 24608
rect 24084 24556 24090 24608
rect 25682 24556 25688 24608
rect 25740 24596 25746 24608
rect 25777 24599 25835 24605
rect 25777 24596 25789 24599
rect 25740 24568 25789 24596
rect 25740 24556 25746 24568
rect 25777 24565 25789 24568
rect 25823 24565 25835 24599
rect 25777 24559 25835 24565
rect 25958 24556 25964 24608
rect 26016 24556 26022 24608
rect 26896 24596 26924 24636
rect 27448 24636 27568 24664
rect 28813 24667 28871 24673
rect 27448 24596 27476 24636
rect 28813 24633 28825 24667
rect 28859 24633 28871 24667
rect 30852 24664 30880 24704
rect 31036 24704 34713 24732
rect 31036 24664 31064 24704
rect 34701 24701 34713 24704
rect 34747 24701 34759 24735
rect 34701 24695 34759 24701
rect 34793 24735 34851 24741
rect 34793 24701 34805 24735
rect 34839 24701 34851 24735
rect 34793 24695 34851 24701
rect 30852 24636 31064 24664
rect 31128 24636 31754 24664
rect 28813 24627 28871 24633
rect 31128 24596 31156 24636
rect 26896 24568 31156 24596
rect 31202 24556 31208 24608
rect 31260 24556 31266 24608
rect 31726 24596 31754 24636
rect 33226 24624 33232 24676
rect 33284 24664 33290 24676
rect 33413 24667 33471 24673
rect 33413 24664 33425 24667
rect 33284 24636 33425 24664
rect 33284 24624 33290 24636
rect 33413 24633 33425 24636
rect 33459 24633 33471 24667
rect 33413 24627 33471 24633
rect 33594 24624 33600 24676
rect 33652 24664 33658 24676
rect 34146 24664 34152 24676
rect 33652 24636 34152 24664
rect 33652 24624 33658 24636
rect 34146 24624 34152 24636
rect 34204 24664 34210 24676
rect 34808 24664 34836 24695
rect 34204 24636 34836 24664
rect 34204 24624 34210 24636
rect 32674 24596 32680 24608
rect 31726 24568 32680 24596
rect 32674 24556 32680 24568
rect 32732 24556 32738 24608
rect 33137 24599 33195 24605
rect 33137 24565 33149 24599
rect 33183 24596 33195 24599
rect 33318 24596 33324 24608
rect 33183 24568 33324 24596
rect 33183 24565 33195 24568
rect 33137 24559 33195 24565
rect 33318 24556 33324 24568
rect 33376 24556 33382 24608
rect 1104 24506 38272 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 38272 24506
rect 1104 24432 38272 24454
rect 1670 24352 1676 24404
rect 1728 24392 1734 24404
rect 1765 24395 1823 24401
rect 1765 24392 1777 24395
rect 1728 24364 1777 24392
rect 1728 24352 1734 24364
rect 1765 24361 1777 24364
rect 1811 24361 1823 24395
rect 1765 24355 1823 24361
rect 3050 24352 3056 24404
rect 3108 24392 3114 24404
rect 3789 24395 3847 24401
rect 3789 24392 3801 24395
rect 3108 24364 3801 24392
rect 3108 24352 3114 24364
rect 3789 24361 3801 24364
rect 3835 24361 3847 24395
rect 3789 24355 3847 24361
rect 4062 24352 4068 24404
rect 4120 24392 4126 24404
rect 7834 24392 7840 24404
rect 4120 24364 7840 24392
rect 4120 24352 4126 24364
rect 7834 24352 7840 24364
rect 7892 24352 7898 24404
rect 7926 24352 7932 24404
rect 7984 24352 7990 24404
rect 9214 24352 9220 24404
rect 9272 24352 9278 24404
rect 13725 24395 13783 24401
rect 13725 24361 13737 24395
rect 13771 24361 13783 24395
rect 13725 24355 13783 24361
rect 13909 24395 13967 24401
rect 13909 24361 13921 24395
rect 13955 24392 13967 24395
rect 15378 24392 15384 24404
rect 13955 24364 15384 24392
rect 13955 24361 13967 24364
rect 13909 24355 13967 24361
rect 1394 24284 1400 24336
rect 1452 24324 1458 24336
rect 1452 24296 5304 24324
rect 1452 24284 1458 24296
rect 2961 24259 3019 24265
rect 2961 24225 2973 24259
rect 3007 24256 3019 24259
rect 4062 24256 4068 24268
rect 3007 24228 4068 24256
rect 3007 24225 3019 24228
rect 2961 24219 3019 24225
rect 4062 24216 4068 24228
rect 4120 24256 4126 24268
rect 5276 24265 5304 24296
rect 6638 24284 6644 24336
rect 6696 24324 6702 24336
rect 7009 24327 7067 24333
rect 7009 24324 7021 24327
rect 6696 24296 7021 24324
rect 6696 24284 6702 24296
rect 7009 24293 7021 24296
rect 7055 24293 7067 24327
rect 9232 24324 9260 24352
rect 7009 24287 7067 24293
rect 8128 24296 9260 24324
rect 13740 24324 13768 24355
rect 15378 24352 15384 24364
rect 15436 24352 15442 24404
rect 15746 24352 15752 24404
rect 15804 24392 15810 24404
rect 15804 24364 17356 24392
rect 15804 24352 15810 24364
rect 14918 24324 14924 24336
rect 13740 24296 14924 24324
rect 4341 24259 4399 24265
rect 4341 24256 4353 24259
rect 4120 24228 4353 24256
rect 4120 24216 4126 24228
rect 4341 24225 4353 24228
rect 4387 24225 4399 24259
rect 4341 24219 4399 24225
rect 5261 24259 5319 24265
rect 5261 24225 5273 24259
rect 5307 24225 5319 24259
rect 5261 24219 5319 24225
rect 5537 24259 5595 24265
rect 5537 24225 5549 24259
rect 5583 24256 5595 24259
rect 5626 24256 5632 24268
rect 5583 24228 5632 24256
rect 5583 24225 5595 24228
rect 5537 24219 5595 24225
rect 5626 24216 5632 24228
rect 5684 24216 5690 24268
rect 1949 24191 2007 24197
rect 1949 24157 1961 24191
rect 1995 24188 2007 24191
rect 4157 24191 4215 24197
rect 1995 24160 2360 24188
rect 1995 24157 2007 24160
rect 1949 24151 2007 24157
rect 2332 24061 2360 24160
rect 4157 24157 4169 24191
rect 4203 24188 4215 24191
rect 4614 24188 4620 24200
rect 4203 24160 4620 24188
rect 4203 24157 4215 24160
rect 4157 24151 4215 24157
rect 4614 24148 4620 24160
rect 4672 24148 4678 24200
rect 8128 24197 8156 24296
rect 14918 24284 14924 24296
rect 14976 24284 14982 24336
rect 15194 24284 15200 24336
rect 15252 24284 15258 24336
rect 8662 24216 8668 24268
rect 8720 24256 8726 24268
rect 8720 24228 9168 24256
rect 8720 24216 8726 24228
rect 9140 24200 9168 24228
rect 12710 24216 12716 24268
rect 12768 24256 12774 24268
rect 12768 24228 12848 24256
rect 12768 24216 12774 24228
rect 8113 24191 8171 24197
rect 8113 24157 8125 24191
rect 8159 24157 8171 24191
rect 8113 24151 8171 24157
rect 9122 24148 9128 24200
rect 9180 24148 9186 24200
rect 12820 24197 12848 24228
rect 12986 24216 12992 24268
rect 13044 24216 13050 24268
rect 14090 24216 14096 24268
rect 14148 24256 14154 24268
rect 14550 24256 14556 24268
rect 14148 24228 14556 24256
rect 14148 24216 14154 24228
rect 14550 24216 14556 24228
rect 14608 24256 14614 24268
rect 14608 24228 15148 24256
rect 14608 24216 14614 24228
rect 12805 24191 12863 24197
rect 12805 24157 12817 24191
rect 12851 24157 12863 24191
rect 14366 24188 14372 24200
rect 13772 24163 14372 24188
rect 12805 24151 12863 24157
rect 13771 24160 14372 24163
rect 13771 24157 13829 24160
rect 5994 24080 6000 24132
rect 6052 24080 6058 24132
rect 13541 24123 13599 24129
rect 13541 24089 13553 24123
rect 13587 24089 13599 24123
rect 13771 24123 13783 24157
rect 13817 24123 13829 24157
rect 14366 24148 14372 24160
rect 14424 24148 14430 24200
rect 14737 24191 14795 24197
rect 14737 24157 14749 24191
rect 14783 24188 14795 24191
rect 14918 24188 14924 24200
rect 14783 24160 14924 24188
rect 14783 24157 14795 24160
rect 14737 24151 14795 24157
rect 14918 24148 14924 24160
rect 14976 24148 14982 24200
rect 15120 24197 15148 24228
rect 15470 24216 15476 24268
rect 15528 24216 15534 24268
rect 15764 24256 15792 24352
rect 16390 24284 16396 24336
rect 16448 24284 16454 24336
rect 17218 24324 17224 24336
rect 16500 24296 17224 24324
rect 16500 24256 16528 24296
rect 17218 24284 17224 24296
rect 17276 24284 17282 24336
rect 15764 24228 15976 24256
rect 15105 24191 15163 24197
rect 15105 24157 15117 24191
rect 15151 24188 15163 24191
rect 15378 24188 15384 24200
rect 15151 24160 15384 24188
rect 15151 24157 15163 24160
rect 15105 24151 15163 24157
rect 15378 24148 15384 24160
rect 15436 24148 15442 24200
rect 13771 24117 13829 24123
rect 13541 24083 13599 24089
rect 2317 24055 2375 24061
rect 2317 24021 2329 24055
rect 2363 24021 2375 24055
rect 2317 24015 2375 24021
rect 2498 24012 2504 24064
rect 2556 24052 2562 24064
rect 2682 24052 2688 24064
rect 2556 24024 2688 24052
rect 2556 24012 2562 24024
rect 2682 24012 2688 24024
rect 2740 24012 2746 24064
rect 2774 24012 2780 24064
rect 2832 24012 2838 24064
rect 4249 24055 4307 24061
rect 4249 24021 4261 24055
rect 4295 24052 4307 24055
rect 4614 24052 4620 24064
rect 4295 24024 4620 24052
rect 4295 24021 4307 24024
rect 4249 24015 4307 24021
rect 4614 24012 4620 24024
rect 4672 24012 4678 24064
rect 9030 24012 9036 24064
rect 9088 24012 9094 24064
rect 12618 24012 12624 24064
rect 12676 24012 12682 24064
rect 13556 24052 13584 24083
rect 15010 24080 15016 24132
rect 15068 24080 15074 24132
rect 15488 24120 15516 24216
rect 15749 24191 15807 24197
rect 15749 24157 15761 24191
rect 15795 24188 15807 24191
rect 15838 24188 15844 24200
rect 15795 24160 15844 24188
rect 15795 24157 15807 24160
rect 15749 24151 15807 24157
rect 15838 24148 15844 24160
rect 15896 24148 15902 24200
rect 15948 24197 15976 24228
rect 16040 24228 16528 24256
rect 16040 24197 16068 24228
rect 15933 24191 15991 24197
rect 15933 24157 15945 24191
rect 15979 24157 15991 24191
rect 15933 24151 15991 24157
rect 16025 24191 16083 24197
rect 16025 24157 16037 24191
rect 16071 24157 16083 24191
rect 16025 24151 16083 24157
rect 16151 24191 16209 24197
rect 16151 24157 16163 24191
rect 16197 24188 16209 24191
rect 16666 24188 16672 24200
rect 16197 24160 16672 24188
rect 16197 24157 16209 24160
rect 16151 24151 16209 24157
rect 16666 24148 16672 24160
rect 16724 24188 16730 24200
rect 17095 24191 17153 24197
rect 17095 24188 17107 24191
rect 16724 24160 17107 24188
rect 16724 24148 16730 24160
rect 17095 24157 17107 24160
rect 17141 24157 17153 24191
rect 17095 24151 17153 24157
rect 17218 24148 17224 24200
rect 17276 24148 17282 24200
rect 17328 24197 17356 24364
rect 17402 24352 17408 24404
rect 17460 24392 17466 24404
rect 18601 24395 18659 24401
rect 18601 24392 18613 24395
rect 17460 24364 18613 24392
rect 17460 24352 17466 24364
rect 18601 24361 18613 24364
rect 18647 24361 18659 24395
rect 18601 24355 18659 24361
rect 18785 24395 18843 24401
rect 18785 24361 18797 24395
rect 18831 24392 18843 24395
rect 19150 24392 19156 24404
rect 18831 24364 19156 24392
rect 18831 24361 18843 24364
rect 18785 24355 18843 24361
rect 19150 24352 19156 24364
rect 19208 24352 19214 24404
rect 19889 24395 19947 24401
rect 19889 24361 19901 24395
rect 19935 24392 19947 24395
rect 19935 24364 20392 24392
rect 19935 24361 19947 24364
rect 19889 24355 19947 24361
rect 20364 24336 20392 24364
rect 20530 24352 20536 24404
rect 20588 24392 20594 24404
rect 21450 24392 21456 24404
rect 20588 24364 21456 24392
rect 20588 24352 20594 24364
rect 21450 24352 21456 24364
rect 21508 24352 21514 24404
rect 22097 24395 22155 24401
rect 22097 24361 22109 24395
rect 22143 24392 22155 24395
rect 22186 24392 22192 24404
rect 22143 24364 22192 24392
rect 22143 24361 22155 24364
rect 22097 24355 22155 24361
rect 22186 24352 22192 24364
rect 22244 24352 22250 24404
rect 23658 24392 23664 24404
rect 23400 24364 23664 24392
rect 17862 24284 17868 24336
rect 17920 24324 17926 24336
rect 20254 24324 20260 24336
rect 17920 24296 20260 24324
rect 17920 24284 17926 24296
rect 17402 24216 17408 24268
rect 17460 24216 17466 24268
rect 17678 24216 17684 24268
rect 17736 24256 17742 24268
rect 19996 24265 20024 24296
rect 20254 24284 20260 24296
rect 20312 24284 20318 24336
rect 20346 24284 20352 24336
rect 20404 24324 20410 24336
rect 20717 24327 20775 24333
rect 20717 24324 20729 24327
rect 20404 24296 20729 24324
rect 20404 24284 20410 24296
rect 20717 24293 20729 24296
rect 20763 24293 20775 24327
rect 20717 24287 20775 24293
rect 21082 24284 21088 24336
rect 21140 24324 21146 24336
rect 21358 24324 21364 24336
rect 21140 24296 21364 24324
rect 21140 24284 21146 24296
rect 21358 24284 21364 24296
rect 21416 24324 21422 24336
rect 21416 24296 22692 24324
rect 21416 24284 21422 24296
rect 19981 24259 20039 24265
rect 17736 24228 19748 24256
rect 17736 24216 17742 24228
rect 17313 24191 17371 24197
rect 17313 24157 17325 24191
rect 17359 24157 17371 24191
rect 17420 24188 17448 24216
rect 17497 24191 17555 24197
rect 17497 24188 17509 24191
rect 17420 24160 17509 24188
rect 17313 24151 17371 24157
rect 17497 24157 17509 24160
rect 17543 24157 17555 24191
rect 17497 24151 17555 24157
rect 16853 24123 16911 24129
rect 16853 24120 16865 24123
rect 15488 24092 16865 24120
rect 16853 24089 16865 24092
rect 16899 24089 16911 24123
rect 17328 24120 17356 24151
rect 17586 24148 17592 24200
rect 17644 24188 17650 24200
rect 17865 24191 17923 24197
rect 17865 24188 17877 24191
rect 17644 24160 17877 24188
rect 17644 24148 17650 24160
rect 17865 24157 17877 24160
rect 17911 24157 17923 24191
rect 17865 24151 17923 24157
rect 18141 24191 18199 24197
rect 18141 24157 18153 24191
rect 18187 24188 18199 24191
rect 18414 24188 18420 24200
rect 18187 24160 18420 24188
rect 18187 24157 18199 24160
rect 18141 24151 18199 24157
rect 18414 24148 18420 24160
rect 18472 24148 18478 24200
rect 18690 24148 18696 24200
rect 18748 24148 18754 24200
rect 18874 24148 18880 24200
rect 18932 24148 18938 24200
rect 19058 24148 19064 24200
rect 19116 24148 19122 24200
rect 19518 24148 19524 24200
rect 19576 24148 19582 24200
rect 19720 24197 19748 24228
rect 19981 24225 19993 24259
rect 20027 24225 20039 24259
rect 19981 24219 20039 24225
rect 20070 24216 20076 24268
rect 20128 24216 20134 24268
rect 22554 24256 22560 24268
rect 20456 24228 22560 24256
rect 19705 24191 19763 24197
rect 19705 24157 19717 24191
rect 19751 24157 19763 24191
rect 20088 24188 20116 24216
rect 20349 24191 20407 24197
rect 20088 24160 20208 24188
rect 19705 24151 19763 24157
rect 17954 24120 17960 24132
rect 17328 24092 17960 24120
rect 16853 24083 16911 24089
rect 17954 24080 17960 24092
rect 18012 24080 18018 24132
rect 18892 24120 18920 24148
rect 18064 24092 18920 24120
rect 15028 24052 15056 24080
rect 13556 24024 15056 24052
rect 15562 24012 15568 24064
rect 15620 24052 15626 24064
rect 18064 24052 18092 24092
rect 19150 24080 19156 24132
rect 19208 24120 19214 24132
rect 20073 24123 20131 24129
rect 20073 24120 20085 24123
rect 19208 24092 20085 24120
rect 19208 24080 19214 24092
rect 20073 24089 20085 24092
rect 20119 24089 20131 24123
rect 20180 24120 20208 24160
rect 20349 24157 20361 24191
rect 20395 24188 20407 24191
rect 20456 24188 20484 24228
rect 22554 24216 22560 24228
rect 22612 24216 22618 24268
rect 20395 24160 20484 24188
rect 20395 24157 20407 24160
rect 20349 24151 20407 24157
rect 20714 24148 20720 24200
rect 20772 24188 20778 24200
rect 20809 24191 20867 24197
rect 20809 24188 20821 24191
rect 20772 24160 20821 24188
rect 20772 24148 20778 24160
rect 20809 24157 20821 24160
rect 20855 24157 20867 24191
rect 20809 24151 20867 24157
rect 22097 24191 22155 24197
rect 22097 24157 22109 24191
rect 22143 24188 22155 24191
rect 22143 24160 22232 24188
rect 22143 24157 22155 24160
rect 22097 24151 22155 24157
rect 20441 24123 20499 24129
rect 20441 24120 20453 24123
rect 20180 24092 20453 24120
rect 20073 24083 20131 24089
rect 20441 24089 20453 24092
rect 20487 24089 20499 24123
rect 20441 24083 20499 24089
rect 22204 24064 22232 24160
rect 15620 24024 18092 24052
rect 15620 24012 15626 24024
rect 18138 24012 18144 24064
rect 18196 24012 18202 24064
rect 18325 24055 18383 24061
rect 18325 24021 18337 24055
rect 18371 24052 18383 24055
rect 19058 24052 19064 24064
rect 18371 24024 19064 24052
rect 18371 24021 18383 24024
rect 18325 24015 18383 24021
rect 19058 24012 19064 24024
rect 19116 24012 19122 24064
rect 19242 24012 19248 24064
rect 19300 24012 19306 24064
rect 19613 24055 19671 24061
rect 19613 24021 19625 24055
rect 19659 24052 19671 24055
rect 19886 24052 19892 24064
rect 19659 24024 19892 24052
rect 19659 24021 19671 24024
rect 19613 24015 19671 24021
rect 19886 24012 19892 24024
rect 19944 24012 19950 24064
rect 19978 24012 19984 24064
rect 20036 24052 20042 24064
rect 20533 24055 20591 24061
rect 20533 24052 20545 24055
rect 20036 24024 20545 24052
rect 20036 24012 20042 24024
rect 20533 24021 20545 24024
rect 20579 24021 20591 24055
rect 20533 24015 20591 24021
rect 22186 24012 22192 24064
rect 22244 24012 22250 24064
rect 22664 24052 22692 24296
rect 23106 24216 23112 24268
rect 23164 24256 23170 24268
rect 23293 24259 23351 24265
rect 23293 24256 23305 24259
rect 23164 24228 23305 24256
rect 23164 24216 23170 24228
rect 23293 24225 23305 24228
rect 23339 24256 23351 24259
rect 23400 24256 23428 24364
rect 23658 24352 23664 24364
rect 23716 24392 23722 24404
rect 23716 24364 24716 24392
rect 23716 24352 23722 24364
rect 24688 24336 24716 24364
rect 25682 24352 25688 24404
rect 25740 24352 25746 24404
rect 26326 24352 26332 24404
rect 26384 24392 26390 24404
rect 27338 24392 27344 24404
rect 26384 24364 27344 24392
rect 26384 24352 26390 24364
rect 27338 24352 27344 24364
rect 27396 24352 27402 24404
rect 31202 24352 31208 24404
rect 31260 24392 31266 24404
rect 31757 24395 31815 24401
rect 31260 24364 31708 24392
rect 31260 24352 31266 24364
rect 24026 24284 24032 24336
rect 24084 24284 24090 24336
rect 24670 24284 24676 24336
rect 24728 24284 24734 24336
rect 23339 24228 23428 24256
rect 23492 24228 24808 24256
rect 23339 24225 23351 24228
rect 23293 24219 23351 24225
rect 23492 24200 23520 24228
rect 22925 24191 22983 24197
rect 22925 24157 22937 24191
rect 22971 24157 22983 24191
rect 22925 24151 22983 24157
rect 22940 24120 22968 24151
rect 23474 24148 23480 24200
rect 23532 24148 23538 24200
rect 23661 24191 23719 24197
rect 23661 24157 23673 24191
rect 23707 24188 23719 24191
rect 23750 24188 23756 24200
rect 23707 24160 23756 24188
rect 23707 24157 23719 24160
rect 23661 24151 23719 24157
rect 23750 24148 23756 24160
rect 23808 24148 23814 24200
rect 23934 24148 23940 24200
rect 23992 24148 23998 24200
rect 24780 24197 24808 24228
rect 24854 24216 24860 24268
rect 24912 24216 24918 24268
rect 25593 24259 25651 24265
rect 25593 24225 25605 24259
rect 25639 24256 25651 24259
rect 25700 24256 25728 24352
rect 26878 24284 26884 24336
rect 26936 24324 26942 24336
rect 28718 24324 28724 24336
rect 26936 24296 28724 24324
rect 26936 24284 26942 24296
rect 28718 24284 28724 24296
rect 28776 24324 28782 24336
rect 30374 24324 30380 24336
rect 28776 24296 30380 24324
rect 28776 24284 28782 24296
rect 30374 24284 30380 24296
rect 30432 24284 30438 24336
rect 31570 24324 31576 24336
rect 31312 24296 31576 24324
rect 25639 24228 25728 24256
rect 25869 24259 25927 24265
rect 25639 24225 25651 24228
rect 25593 24219 25651 24225
rect 25869 24225 25881 24259
rect 25915 24256 25927 24259
rect 25958 24256 25964 24268
rect 25915 24228 25964 24256
rect 25915 24225 25927 24228
rect 25869 24219 25927 24225
rect 25958 24216 25964 24228
rect 26016 24216 26022 24268
rect 26418 24216 26424 24268
rect 26476 24256 26482 24268
rect 27154 24256 27160 24268
rect 26476 24228 27160 24256
rect 26476 24216 26482 24228
rect 27154 24216 27160 24228
rect 27212 24216 27218 24268
rect 28261 24259 28319 24265
rect 28261 24225 28273 24259
rect 28307 24256 28319 24259
rect 30282 24256 30288 24268
rect 28307 24228 29684 24256
rect 28307 24225 28319 24228
rect 28261 24219 28319 24225
rect 24765 24191 24823 24197
rect 24765 24157 24777 24191
rect 24811 24157 24823 24191
rect 24765 24151 24823 24157
rect 25314 24148 25320 24200
rect 25372 24148 25378 24200
rect 27890 24148 27896 24200
rect 27948 24188 27954 24200
rect 28169 24191 28227 24197
rect 28169 24188 28181 24191
rect 27948 24160 28181 24188
rect 27948 24148 27954 24160
rect 28169 24157 28181 24160
rect 28215 24157 28227 24191
rect 28169 24151 28227 24157
rect 28350 24148 28356 24200
rect 28408 24188 28414 24200
rect 28445 24191 28503 24197
rect 28445 24188 28457 24191
rect 28408 24160 28457 24188
rect 28408 24148 28414 24160
rect 28445 24157 28457 24160
rect 28491 24157 28503 24191
rect 28445 24151 28503 24157
rect 29546 24148 29552 24200
rect 29604 24148 29610 24200
rect 29656 24188 29684 24228
rect 29840 24228 30288 24256
rect 29840 24200 29868 24228
rect 30282 24216 30288 24228
rect 30340 24256 30346 24268
rect 31312 24256 31340 24296
rect 31570 24284 31576 24296
rect 31628 24284 31634 24336
rect 31680 24324 31708 24364
rect 31757 24361 31769 24395
rect 31803 24361 31815 24395
rect 32950 24392 32956 24404
rect 31757 24355 31815 24361
rect 32784 24364 32956 24392
rect 31772 24324 31800 24355
rect 31680 24296 31800 24324
rect 31680 24256 31708 24296
rect 30340 24228 31340 24256
rect 31404 24228 32444 24256
rect 30340 24216 30346 24228
rect 29730 24197 29736 24200
rect 29728 24188 29736 24197
rect 29656 24160 29736 24188
rect 29728 24151 29736 24160
rect 29730 24148 29736 24151
rect 29788 24148 29794 24200
rect 29822 24148 29828 24200
rect 29880 24148 29886 24200
rect 29914 24148 29920 24200
rect 29972 24148 29978 24200
rect 31404 24197 31432 24228
rect 32416 24197 32444 24228
rect 32784 24197 32812 24364
rect 32950 24352 32956 24364
rect 33008 24392 33014 24404
rect 33008 24364 34468 24392
rect 33008 24352 33014 24364
rect 33042 24284 33048 24336
rect 33100 24324 33106 24336
rect 33100 24296 33456 24324
rect 33100 24284 33106 24296
rect 33428 24256 33456 24296
rect 33502 24284 33508 24336
rect 33560 24284 33566 24336
rect 34440 24333 34468 24364
rect 33689 24327 33747 24333
rect 33689 24293 33701 24327
rect 33735 24324 33747 24327
rect 34425 24327 34483 24333
rect 33735 24296 34192 24324
rect 33735 24293 33747 24296
rect 33689 24287 33747 24293
rect 33428 24228 34100 24256
rect 31389 24191 31447 24197
rect 31389 24157 31401 24191
rect 31435 24157 31447 24191
rect 31389 24151 31447 24157
rect 31573 24191 31631 24197
rect 31573 24157 31585 24191
rect 31619 24188 31631 24191
rect 31665 24191 31723 24197
rect 31665 24188 31677 24191
rect 31619 24160 31677 24188
rect 31619 24157 31631 24160
rect 31573 24151 31631 24157
rect 31665 24157 31677 24160
rect 31711 24188 31723 24191
rect 32217 24191 32275 24197
rect 32217 24188 32229 24191
rect 31711 24160 32229 24188
rect 31711 24157 31723 24160
rect 31665 24151 31723 24157
rect 32217 24157 32229 24160
rect 32263 24157 32275 24191
rect 32217 24151 32275 24157
rect 32401 24191 32459 24197
rect 32401 24157 32413 24191
rect 32447 24157 32459 24191
rect 32401 24151 32459 24157
rect 32769 24191 32827 24197
rect 32769 24157 32781 24191
rect 32815 24157 32827 24191
rect 32769 24151 32827 24157
rect 23952 24120 23980 24148
rect 22940 24092 23980 24120
rect 26878 24080 26884 24132
rect 26936 24080 26942 24132
rect 27614 24080 27620 24132
rect 27672 24120 27678 24132
rect 31680 24120 31708 24151
rect 32858 24148 32864 24200
rect 32916 24148 32922 24200
rect 33134 24148 33140 24200
rect 33192 24148 33198 24200
rect 33229 24191 33287 24197
rect 33229 24157 33241 24191
rect 33275 24157 33287 24191
rect 33229 24151 33287 24157
rect 33244 24120 33272 24151
rect 33318 24148 33324 24200
rect 33376 24188 33382 24200
rect 33597 24191 33655 24197
rect 33428 24188 33548 24190
rect 33597 24188 33609 24191
rect 33376 24162 33609 24188
rect 33376 24160 33456 24162
rect 33520 24160 33609 24162
rect 33376 24148 33382 24160
rect 33597 24157 33609 24160
rect 33643 24157 33655 24191
rect 33597 24151 33655 24157
rect 33778 24148 33784 24200
rect 33836 24188 33842 24200
rect 34072 24197 34100 24228
rect 34164 24197 34192 24296
rect 34425 24293 34437 24327
rect 34471 24293 34483 24327
rect 34425 24287 34483 24293
rect 33873 24191 33931 24197
rect 33873 24188 33885 24191
rect 33836 24160 33885 24188
rect 33836 24148 33842 24160
rect 33873 24157 33885 24160
rect 33919 24157 33931 24191
rect 33873 24151 33931 24157
rect 34057 24191 34115 24197
rect 34057 24157 34069 24191
rect 34103 24157 34115 24191
rect 34057 24151 34115 24157
rect 34149 24191 34207 24197
rect 34149 24157 34161 24191
rect 34195 24157 34207 24191
rect 34149 24151 34207 24157
rect 34333 24191 34391 24197
rect 34333 24157 34345 24191
rect 34379 24157 34391 24191
rect 34333 24151 34391 24157
rect 27672 24092 31708 24120
rect 32140 24092 33272 24120
rect 33505 24123 33563 24129
rect 27672 24080 27678 24092
rect 29822 24052 29828 24064
rect 22664 24024 29828 24052
rect 29822 24012 29828 24024
rect 29880 24012 29886 24064
rect 30190 24012 30196 24064
rect 30248 24012 30254 24064
rect 31478 24012 31484 24064
rect 31536 24012 31542 24064
rect 32140 24061 32168 24092
rect 33152 24064 33180 24092
rect 33505 24089 33517 24123
rect 33551 24120 33563 24123
rect 33965 24123 34023 24129
rect 33965 24120 33977 24123
rect 33551 24092 33977 24120
rect 33551 24089 33563 24092
rect 33505 24083 33563 24089
rect 33965 24089 33977 24092
rect 34011 24120 34023 24123
rect 34348 24120 34376 24151
rect 34011 24092 34376 24120
rect 34011 24089 34023 24092
rect 33965 24083 34023 24089
rect 32125 24055 32183 24061
rect 32125 24021 32137 24055
rect 32171 24021 32183 24055
rect 32125 24015 32183 24021
rect 32398 24012 32404 24064
rect 32456 24012 32462 24064
rect 32582 24012 32588 24064
rect 32640 24012 32646 24064
rect 33134 24012 33140 24064
rect 33192 24012 33198 24064
rect 1104 23962 38272 23984
rect 1104 23910 4874 23962
rect 4926 23910 4938 23962
rect 4990 23910 5002 23962
rect 5054 23910 5066 23962
rect 5118 23910 5130 23962
rect 5182 23910 35594 23962
rect 35646 23910 35658 23962
rect 35710 23910 35722 23962
rect 35774 23910 35786 23962
rect 35838 23910 35850 23962
rect 35902 23910 38272 23962
rect 1104 23888 38272 23910
rect 1946 23808 1952 23860
rect 2004 23808 2010 23860
rect 5902 23808 5908 23860
rect 5960 23848 5966 23860
rect 6365 23851 6423 23857
rect 6365 23848 6377 23851
rect 5960 23820 6377 23848
rect 5960 23808 5966 23820
rect 6365 23817 6377 23820
rect 6411 23817 6423 23851
rect 12713 23851 12771 23857
rect 12713 23848 12725 23851
rect 6365 23811 6423 23817
rect 7576 23820 12725 23848
rect 1964 23780 1992 23808
rect 7576 23780 7604 23820
rect 12713 23817 12725 23820
rect 12759 23817 12771 23851
rect 12713 23811 12771 23817
rect 12894 23808 12900 23860
rect 12952 23808 12958 23860
rect 14660 23820 15240 23848
rect 9030 23780 9036 23792
rect 1964 23752 7604 23780
rect 8680 23752 9036 23780
rect 5626 23672 5632 23724
rect 5684 23672 5690 23724
rect 6638 23672 6644 23724
rect 6696 23712 6702 23724
rect 6733 23715 6791 23721
rect 6733 23712 6745 23715
rect 6696 23684 6745 23712
rect 6696 23672 6702 23684
rect 6733 23681 6745 23684
rect 6779 23681 6791 23715
rect 6733 23675 6791 23681
rect 6825 23715 6883 23721
rect 6825 23681 6837 23715
rect 6871 23712 6883 23715
rect 7006 23712 7012 23724
rect 6871 23684 7012 23712
rect 6871 23681 6883 23684
rect 6825 23675 6883 23681
rect 7006 23672 7012 23684
rect 7064 23672 7070 23724
rect 8680 23721 8708 23752
rect 9030 23740 9036 23752
rect 9088 23740 9094 23792
rect 9674 23740 9680 23792
rect 9732 23740 9738 23792
rect 12912 23780 12940 23808
rect 12406 23752 12940 23780
rect 13449 23783 13507 23789
rect 8665 23715 8723 23721
rect 8665 23681 8677 23715
rect 8711 23681 8723 23715
rect 8665 23675 8723 23681
rect 11241 23715 11299 23721
rect 11241 23681 11253 23715
rect 11287 23712 11299 23715
rect 12406 23712 12434 23752
rect 13449 23749 13461 23783
rect 13495 23780 13507 23783
rect 13538 23780 13544 23792
rect 13495 23752 13544 23780
rect 13495 23749 13507 23752
rect 13449 23743 13507 23749
rect 13538 23740 13544 23752
rect 13596 23740 13602 23792
rect 14274 23740 14280 23792
rect 14332 23740 14338 23792
rect 14458 23740 14464 23792
rect 14516 23780 14522 23792
rect 14660 23789 14688 23820
rect 14645 23783 14703 23789
rect 14645 23780 14657 23783
rect 14516 23752 14657 23780
rect 14516 23740 14522 23752
rect 14645 23749 14657 23752
rect 14691 23749 14703 23783
rect 14645 23743 14703 23749
rect 15010 23740 15016 23792
rect 15068 23740 15074 23792
rect 11287 23684 12434 23712
rect 11287 23681 11299 23684
rect 11241 23675 11299 23681
rect 4062 23604 4068 23656
rect 4120 23644 4126 23656
rect 6917 23647 6975 23653
rect 6917 23644 6929 23647
rect 4120 23616 6929 23644
rect 4120 23604 4126 23616
rect 6917 23613 6929 23616
rect 6963 23613 6975 23647
rect 6917 23607 6975 23613
rect 8941 23647 8999 23653
rect 8941 23613 8953 23647
rect 8987 23644 8999 23647
rect 9306 23644 9312 23656
rect 8987 23616 9312 23644
rect 8987 23613 8999 23616
rect 8941 23607 8999 23613
rect 9306 23604 9312 23616
rect 9364 23604 9370 23656
rect 10413 23647 10471 23653
rect 10413 23613 10425 23647
rect 10459 23644 10471 23647
rect 11256 23644 11284 23675
rect 12710 23672 12716 23724
rect 12768 23712 12774 23724
rect 12894 23712 12900 23724
rect 12768 23684 12900 23712
rect 12768 23672 12774 23684
rect 12894 23672 12900 23684
rect 12952 23672 12958 23724
rect 13078 23672 13084 23724
rect 13136 23672 13142 23724
rect 14182 23672 14188 23724
rect 14240 23672 14246 23724
rect 14366 23672 14372 23724
rect 14424 23712 14430 23724
rect 14737 23715 14795 23721
rect 14737 23712 14749 23715
rect 14424 23684 14749 23712
rect 14424 23672 14430 23684
rect 14737 23681 14749 23684
rect 14783 23681 14795 23715
rect 14737 23675 14795 23681
rect 14829 23715 14887 23721
rect 14829 23681 14841 23715
rect 14875 23712 14887 23715
rect 14918 23712 14924 23724
rect 14875 23684 14924 23712
rect 14875 23681 14887 23684
rect 14829 23675 14887 23681
rect 14918 23672 14924 23684
rect 14976 23672 14982 23724
rect 10459 23616 11284 23644
rect 15212 23644 15240 23820
rect 15654 23808 15660 23860
rect 15712 23848 15718 23860
rect 15749 23851 15807 23857
rect 15749 23848 15761 23851
rect 15712 23820 15761 23848
rect 15712 23808 15718 23820
rect 15749 23817 15761 23820
rect 15795 23817 15807 23851
rect 18598 23848 18604 23860
rect 15749 23811 15807 23817
rect 16500 23820 18604 23848
rect 16022 23780 16028 23792
rect 15304 23752 16028 23780
rect 15304 23721 15332 23752
rect 16022 23740 16028 23752
rect 16080 23740 16086 23792
rect 15289 23715 15347 23721
rect 15289 23681 15301 23715
rect 15335 23681 15347 23715
rect 15289 23675 15347 23681
rect 15473 23715 15531 23721
rect 15473 23681 15485 23715
rect 15519 23712 15531 23715
rect 15562 23712 15568 23724
rect 15519 23684 15568 23712
rect 15519 23681 15531 23684
rect 15473 23675 15531 23681
rect 15562 23672 15568 23684
rect 15620 23672 15626 23724
rect 15657 23715 15715 23721
rect 15657 23681 15669 23715
rect 15703 23712 15715 23715
rect 16500 23712 16528 23820
rect 17862 23780 17868 23792
rect 17328 23752 17868 23780
rect 17328 23721 17356 23752
rect 17862 23740 17868 23752
rect 17920 23740 17926 23792
rect 18524 23789 18552 23820
rect 18598 23808 18604 23820
rect 18656 23808 18662 23860
rect 18690 23808 18696 23860
rect 18748 23808 18754 23860
rect 18966 23808 18972 23860
rect 19024 23808 19030 23860
rect 19242 23808 19248 23860
rect 19300 23808 19306 23860
rect 19886 23808 19892 23860
rect 19944 23808 19950 23860
rect 20162 23808 20168 23860
rect 20220 23848 20226 23860
rect 20220 23820 28028 23848
rect 20220 23808 20226 23820
rect 18509 23783 18567 23789
rect 18509 23749 18521 23783
rect 18555 23749 18567 23783
rect 18509 23743 18567 23749
rect 17313 23715 17371 23721
rect 17313 23712 17325 23715
rect 15703 23684 16528 23712
rect 16684 23684 17325 23712
rect 15703 23681 15715 23684
rect 15657 23675 15715 23681
rect 15672 23644 15700 23675
rect 16684 23656 16712 23684
rect 17313 23681 17325 23684
rect 17359 23681 17371 23715
rect 17313 23675 17371 23681
rect 17405 23715 17463 23721
rect 17405 23681 17417 23715
rect 17451 23712 17463 23715
rect 17957 23715 18015 23721
rect 17957 23712 17969 23715
rect 17451 23684 17969 23712
rect 17451 23681 17463 23684
rect 17405 23675 17463 23681
rect 17696 23656 17724 23684
rect 17957 23681 17969 23684
rect 18003 23681 18015 23715
rect 17957 23675 18015 23681
rect 18049 23715 18107 23721
rect 18049 23681 18061 23715
rect 18095 23681 18107 23715
rect 18049 23675 18107 23681
rect 16025 23647 16083 23653
rect 16025 23644 16037 23647
rect 15212 23616 15700 23644
rect 15764 23616 16037 23644
rect 10459 23613 10471 23616
rect 10413 23607 10471 23613
rect 5994 23536 6000 23588
rect 6052 23576 6058 23588
rect 7282 23576 7288 23588
rect 6052 23548 7288 23576
rect 6052 23536 6058 23548
rect 7282 23536 7288 23548
rect 7340 23536 7346 23588
rect 9968 23548 12434 23576
rect 5258 23468 5264 23520
rect 5316 23508 5322 23520
rect 5537 23511 5595 23517
rect 5537 23508 5549 23511
rect 5316 23480 5549 23508
rect 5316 23468 5322 23480
rect 5537 23477 5549 23480
rect 5583 23477 5595 23511
rect 5537 23471 5595 23477
rect 7466 23468 7472 23520
rect 7524 23508 7530 23520
rect 9968 23508 9996 23548
rect 7524 23480 9996 23508
rect 7524 23468 7530 23480
rect 10042 23468 10048 23520
rect 10100 23508 10106 23520
rect 10597 23511 10655 23517
rect 10597 23508 10609 23511
rect 10100 23480 10609 23508
rect 10100 23468 10106 23480
rect 10597 23477 10609 23480
rect 10643 23477 10655 23511
rect 12406 23508 12434 23548
rect 15378 23536 15384 23588
rect 15436 23576 15442 23588
rect 15764 23576 15792 23616
rect 16025 23613 16037 23616
rect 16071 23644 16083 23647
rect 16114 23644 16120 23656
rect 16071 23616 16120 23644
rect 16071 23613 16083 23616
rect 16025 23607 16083 23613
rect 16114 23604 16120 23616
rect 16172 23604 16178 23656
rect 16666 23604 16672 23656
rect 16724 23604 16730 23656
rect 17218 23604 17224 23656
rect 17276 23604 17282 23656
rect 17497 23647 17555 23653
rect 17497 23644 17509 23647
rect 17328 23616 17509 23644
rect 15436 23548 15792 23576
rect 15841 23579 15899 23585
rect 15436 23536 15442 23548
rect 15841 23545 15853 23579
rect 15887 23576 15899 23579
rect 17236 23576 17264 23604
rect 15887 23548 17264 23576
rect 17328 23576 17356 23616
rect 17497 23613 17509 23616
rect 17543 23613 17555 23647
rect 17497 23607 17555 23613
rect 17678 23604 17684 23656
rect 17736 23604 17742 23656
rect 18064 23644 18092 23675
rect 17972 23616 18092 23644
rect 18984 23644 19012 23808
rect 19260 23780 19288 23808
rect 19803 23783 19861 23789
rect 19803 23780 19815 23783
rect 19076 23752 19288 23780
rect 19628 23752 19815 23780
rect 19076 23721 19104 23752
rect 19061 23715 19119 23721
rect 19061 23681 19073 23715
rect 19107 23681 19119 23715
rect 19061 23675 19119 23681
rect 19150 23672 19156 23724
rect 19208 23672 19214 23724
rect 19245 23715 19303 23721
rect 19245 23681 19257 23715
rect 19291 23681 19303 23715
rect 19245 23675 19303 23681
rect 19260 23644 19288 23675
rect 19426 23672 19432 23724
rect 19484 23672 19490 23724
rect 18984 23616 19288 23644
rect 17972 23576 18000 23616
rect 17328 23548 18000 23576
rect 18969 23579 19027 23585
rect 15887 23545 15899 23548
rect 15841 23539 15899 23545
rect 17328 23520 17356 23548
rect 18969 23545 18981 23579
rect 19015 23576 19027 23579
rect 19521 23579 19579 23585
rect 19521 23576 19533 23579
rect 19015 23548 19533 23576
rect 19015 23545 19027 23548
rect 18969 23539 19027 23545
rect 19521 23545 19533 23548
rect 19567 23545 19579 23579
rect 19521 23539 19579 23545
rect 12802 23508 12808 23520
rect 12406 23480 12808 23508
rect 10597 23471 10655 23477
rect 12802 23468 12808 23480
rect 12860 23508 12866 23520
rect 13722 23508 13728 23520
rect 12860 23480 13728 23508
rect 12860 23468 12866 23480
rect 13722 23468 13728 23480
rect 13780 23468 13786 23520
rect 15102 23468 15108 23520
rect 15160 23468 15166 23520
rect 15930 23468 15936 23520
rect 15988 23508 15994 23520
rect 16206 23508 16212 23520
rect 15988 23480 16212 23508
rect 15988 23468 15994 23480
rect 16206 23468 16212 23480
rect 16264 23468 16270 23520
rect 17310 23468 17316 23520
rect 17368 23468 17374 23520
rect 17494 23468 17500 23520
rect 17552 23508 17558 23520
rect 17681 23511 17739 23517
rect 17681 23508 17693 23511
rect 17552 23480 17693 23508
rect 17552 23468 17558 23480
rect 17681 23477 17693 23480
rect 17727 23477 17739 23511
rect 17681 23471 17739 23477
rect 17773 23511 17831 23517
rect 17773 23477 17785 23511
rect 17819 23508 17831 23511
rect 17862 23508 17868 23520
rect 17819 23480 17868 23508
rect 17819 23477 17831 23480
rect 17773 23471 17831 23477
rect 17862 23468 17868 23480
rect 17920 23468 17926 23520
rect 18046 23468 18052 23520
rect 18104 23508 18110 23520
rect 19628 23508 19656 23752
rect 19803 23749 19815 23752
rect 19849 23780 19861 23783
rect 19849 23752 21042 23780
rect 19849 23749 19861 23752
rect 19803 23743 19861 23749
rect 19978 23672 19984 23724
rect 20036 23672 20042 23724
rect 20254 23672 20260 23724
rect 20312 23712 20318 23724
rect 20714 23712 20720 23724
rect 20312 23684 20720 23712
rect 20312 23672 20318 23684
rect 20714 23672 20720 23684
rect 20772 23672 20778 23724
rect 20806 23672 20812 23724
rect 20864 23672 20870 23724
rect 21014 23712 21042 23752
rect 21082 23740 21088 23792
rect 21140 23740 21146 23792
rect 23106 23780 23112 23792
rect 22388 23752 23112 23780
rect 22002 23712 22008 23724
rect 21014 23684 22008 23712
rect 22002 23672 22008 23684
rect 22060 23672 22066 23724
rect 22388 23721 22416 23752
rect 23106 23740 23112 23752
rect 23164 23740 23170 23792
rect 24486 23780 24492 23792
rect 24136 23752 24492 23780
rect 24136 23724 24164 23752
rect 24486 23740 24492 23752
rect 24544 23740 24550 23792
rect 25314 23780 25320 23792
rect 24688 23752 25320 23780
rect 22373 23715 22431 23721
rect 22373 23681 22385 23715
rect 22419 23681 22431 23715
rect 22373 23675 22431 23681
rect 22557 23715 22615 23721
rect 22557 23681 22569 23715
rect 22603 23712 22615 23715
rect 22922 23712 22928 23724
rect 22603 23684 22928 23712
rect 22603 23681 22615 23684
rect 22557 23675 22615 23681
rect 22922 23672 22928 23684
rect 22980 23672 22986 23724
rect 23293 23715 23351 23721
rect 23293 23681 23305 23715
rect 23339 23712 23351 23715
rect 23382 23712 23388 23724
rect 23339 23684 23388 23712
rect 23339 23681 23351 23684
rect 23293 23675 23351 23681
rect 23382 23672 23388 23684
rect 23440 23672 23446 23724
rect 23661 23715 23719 23721
rect 23661 23681 23673 23715
rect 23707 23712 23719 23715
rect 23750 23712 23756 23724
rect 23707 23684 23756 23712
rect 23707 23681 23719 23684
rect 23661 23675 23719 23681
rect 23750 23672 23756 23684
rect 23808 23672 23814 23724
rect 23845 23715 23903 23721
rect 23845 23681 23857 23715
rect 23891 23712 23903 23715
rect 24118 23712 24124 23724
rect 23891 23684 24124 23712
rect 23891 23681 23903 23684
rect 23845 23675 23903 23681
rect 21450 23604 21456 23656
rect 21508 23644 21514 23656
rect 22649 23647 22707 23653
rect 22649 23644 22661 23647
rect 21508 23616 22661 23644
rect 21508 23604 21514 23616
rect 22649 23613 22661 23616
rect 22695 23613 22707 23647
rect 22649 23607 22707 23613
rect 23201 23647 23259 23653
rect 23201 23613 23213 23647
rect 23247 23613 23259 23647
rect 23201 23607 23259 23613
rect 20165 23579 20223 23585
rect 20165 23545 20177 23579
rect 20211 23576 20223 23579
rect 20346 23576 20352 23588
rect 20211 23548 20352 23576
rect 20211 23545 20223 23548
rect 20165 23539 20223 23545
rect 20346 23536 20352 23548
rect 20404 23536 20410 23588
rect 22186 23536 22192 23588
rect 22244 23576 22250 23588
rect 23216 23576 23244 23607
rect 23566 23604 23572 23656
rect 23624 23644 23630 23656
rect 23860 23644 23888 23675
rect 24118 23672 24124 23684
rect 24176 23672 24182 23724
rect 24688 23721 24716 23752
rect 25314 23740 25320 23752
rect 25372 23780 25378 23792
rect 25869 23783 25927 23789
rect 25869 23780 25881 23783
rect 25372 23752 25881 23780
rect 25372 23740 25378 23752
rect 25869 23749 25881 23752
rect 25915 23749 25927 23783
rect 25869 23743 25927 23749
rect 26970 23740 26976 23792
rect 27028 23780 27034 23792
rect 28000 23789 28028 23820
rect 28166 23808 28172 23860
rect 28224 23808 28230 23860
rect 28626 23808 28632 23860
rect 28684 23848 28690 23860
rect 29089 23851 29147 23857
rect 29089 23848 29101 23851
rect 28684 23820 29101 23848
rect 28684 23808 28690 23820
rect 29089 23817 29101 23820
rect 29135 23817 29147 23851
rect 29089 23811 29147 23817
rect 31478 23808 31484 23860
rect 31536 23848 31542 23860
rect 32217 23851 32275 23857
rect 31536 23820 31754 23848
rect 31536 23808 31542 23820
rect 27249 23783 27307 23789
rect 27249 23780 27261 23783
rect 27028 23752 27261 23780
rect 27028 23740 27034 23752
rect 27249 23749 27261 23752
rect 27295 23780 27307 23783
rect 27893 23783 27951 23789
rect 27893 23780 27905 23783
rect 27295 23752 27905 23780
rect 27295 23749 27307 23752
rect 27249 23743 27307 23749
rect 27893 23749 27905 23752
rect 27939 23749 27951 23783
rect 27893 23743 27951 23749
rect 27985 23783 28043 23789
rect 27985 23749 27997 23783
rect 28031 23749 28043 23783
rect 27985 23743 28043 23749
rect 24673 23715 24731 23721
rect 24673 23681 24685 23715
rect 24719 23681 24731 23715
rect 24673 23675 24731 23681
rect 24762 23672 24768 23724
rect 24820 23712 24826 23724
rect 25041 23715 25099 23721
rect 25041 23712 25053 23715
rect 24820 23684 25053 23712
rect 24820 23672 24826 23684
rect 25041 23681 25053 23684
rect 25087 23681 25099 23715
rect 25041 23675 25099 23681
rect 25130 23672 25136 23724
rect 25188 23672 25194 23724
rect 26050 23672 26056 23724
rect 26108 23672 26114 23724
rect 27062 23672 27068 23724
rect 27120 23672 27126 23724
rect 27341 23715 27399 23721
rect 27341 23681 27353 23715
rect 27387 23681 27399 23715
rect 27341 23675 27399 23681
rect 23624 23616 23888 23644
rect 24400 23656 24452 23662
rect 23624 23604 23630 23616
rect 26237 23647 26295 23653
rect 26237 23613 26249 23647
rect 26283 23613 26295 23647
rect 26237 23607 26295 23613
rect 24400 23598 24452 23604
rect 22244 23548 23244 23576
rect 22244 23536 22250 23548
rect 24302 23536 24308 23588
rect 24360 23536 24366 23588
rect 24486 23536 24492 23588
rect 24544 23576 24550 23588
rect 26252 23576 26280 23607
rect 26694 23576 26700 23588
rect 24544 23548 26700 23576
rect 24544 23536 24550 23548
rect 26694 23536 26700 23548
rect 26752 23536 26758 23588
rect 18104 23480 19656 23508
rect 18104 23468 18110 23480
rect 19702 23468 19708 23520
rect 19760 23508 19766 23520
rect 27356 23508 27384 23675
rect 27430 23672 27436 23724
rect 27488 23672 27494 23724
rect 27706 23672 27712 23724
rect 27764 23672 27770 23724
rect 28077 23715 28135 23721
rect 28077 23681 28089 23715
rect 28123 23681 28135 23715
rect 28184 23712 28212 23808
rect 28718 23740 28724 23792
rect 28776 23740 28782 23792
rect 28629 23715 28687 23721
rect 28629 23712 28641 23715
rect 28184 23684 28641 23712
rect 28077 23675 28135 23681
rect 28629 23681 28641 23684
rect 28675 23681 28687 23715
rect 31726 23712 31754 23820
rect 32217 23817 32229 23851
rect 32263 23848 32275 23851
rect 32858 23848 32864 23860
rect 32263 23820 32864 23848
rect 32263 23817 32275 23820
rect 32217 23811 32275 23817
rect 32858 23808 32864 23820
rect 32916 23808 32922 23860
rect 33134 23808 33140 23860
rect 33192 23808 33198 23860
rect 34606 23808 34612 23860
rect 34664 23848 34670 23860
rect 34664 23820 35572 23848
rect 34664 23808 34670 23820
rect 33152 23721 33180 23808
rect 35544 23724 35572 23820
rect 32125 23715 32183 23721
rect 32125 23712 32137 23715
rect 31726 23684 32137 23712
rect 28629 23675 28687 23681
rect 32125 23681 32137 23684
rect 32171 23681 32183 23715
rect 32125 23675 32183 23681
rect 33137 23715 33195 23721
rect 33137 23681 33149 23715
rect 33183 23681 33195 23715
rect 33137 23675 33195 23681
rect 27448 23644 27476 23672
rect 27890 23644 27896 23656
rect 27448 23616 27896 23644
rect 27890 23604 27896 23616
rect 27948 23644 27954 23656
rect 28092 23644 28120 23675
rect 35526 23672 35532 23724
rect 35584 23672 35590 23724
rect 28445 23647 28503 23653
rect 28445 23644 28457 23647
rect 27948 23616 28120 23644
rect 28184 23616 28457 23644
rect 27948 23604 27954 23616
rect 27522 23536 27528 23588
rect 27580 23536 27586 23588
rect 27614 23536 27620 23588
rect 27672 23536 27678 23588
rect 19760 23480 27384 23508
rect 27540 23508 27568 23536
rect 28184 23508 28212 23616
rect 28445 23613 28457 23616
rect 28491 23644 28503 23647
rect 33594 23644 33600 23656
rect 28491 23616 33600 23644
rect 28491 23613 28503 23616
rect 28445 23607 28503 23613
rect 33594 23604 33600 23616
rect 33652 23604 33658 23656
rect 34698 23604 34704 23656
rect 34756 23644 34762 23656
rect 34885 23647 34943 23653
rect 34885 23644 34897 23647
rect 34756 23616 34897 23644
rect 34756 23604 34762 23616
rect 34885 23613 34897 23616
rect 34931 23613 34943 23647
rect 34885 23607 34943 23613
rect 35621 23647 35679 23653
rect 35621 23613 35633 23647
rect 35667 23613 35679 23647
rect 35621 23607 35679 23613
rect 28261 23579 28319 23585
rect 28261 23545 28273 23579
rect 28307 23576 28319 23579
rect 33042 23576 33048 23588
rect 28307 23548 33048 23576
rect 28307 23545 28319 23548
rect 28261 23539 28319 23545
rect 33042 23536 33048 23548
rect 33100 23536 33106 23588
rect 35434 23536 35440 23588
rect 35492 23576 35498 23588
rect 35636 23576 35664 23607
rect 35492 23548 35664 23576
rect 35492 23536 35498 23548
rect 27540 23480 28212 23508
rect 19760 23468 19766 23480
rect 33226 23468 33232 23520
rect 33284 23468 33290 23520
rect 1104 23418 38272 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 38272 23418
rect 1104 23344 38272 23366
rect 1762 23264 1768 23316
rect 1820 23304 1826 23316
rect 2225 23307 2283 23313
rect 2225 23304 2237 23307
rect 1820 23276 2237 23304
rect 1820 23264 1826 23276
rect 2225 23273 2237 23276
rect 2271 23273 2283 23307
rect 2225 23267 2283 23273
rect 2774 23264 2780 23316
rect 2832 23304 2838 23316
rect 2961 23307 3019 23313
rect 2961 23304 2973 23307
rect 2832 23276 2973 23304
rect 2832 23264 2838 23276
rect 2961 23273 2973 23276
rect 3007 23273 3019 23307
rect 2961 23267 3019 23273
rect 4249 23307 4307 23313
rect 4249 23273 4261 23307
rect 4295 23304 4307 23307
rect 4614 23304 4620 23316
rect 4295 23276 4620 23304
rect 4295 23273 4307 23276
rect 4249 23267 4307 23273
rect 4614 23264 4620 23276
rect 4672 23264 4678 23316
rect 4798 23264 4804 23316
rect 4856 23304 4862 23316
rect 4985 23307 5043 23313
rect 4985 23304 4997 23307
rect 4856 23276 4997 23304
rect 4856 23264 4862 23276
rect 4985 23273 4997 23276
rect 5031 23273 5043 23307
rect 4985 23267 5043 23273
rect 5626 23264 5632 23316
rect 5684 23304 5690 23316
rect 6273 23307 6331 23313
rect 6273 23304 6285 23307
rect 5684 23276 6285 23304
rect 5684 23264 5690 23276
rect 6273 23273 6285 23276
rect 6319 23273 6331 23307
rect 6454 23304 6460 23316
rect 6512 23313 6518 23316
rect 6273 23267 6331 23273
rect 6380 23276 6460 23304
rect 5810 23196 5816 23248
rect 5868 23236 5874 23248
rect 6380 23236 6408 23276
rect 6454 23264 6460 23276
rect 6512 23267 6524 23313
rect 6512 23264 6518 23267
rect 7006 23264 7012 23316
rect 7064 23264 7070 23316
rect 7650 23264 7656 23316
rect 7708 23304 7714 23316
rect 7708 23276 8156 23304
rect 7708 23264 7714 23276
rect 8018 23236 8024 23248
rect 5868 23208 6408 23236
rect 6932 23208 8024 23236
rect 5868 23196 5874 23208
rect 5721 23171 5779 23177
rect 5721 23168 5733 23171
rect 5276 23140 5733 23168
rect 5186 23113 5244 23119
rect 1946 23060 1952 23112
rect 2004 23060 2010 23112
rect 2498 23060 2504 23112
rect 2556 23060 2562 23112
rect 2593 23103 2651 23109
rect 2593 23069 2605 23103
rect 2639 23069 2651 23103
rect 2593 23063 2651 23069
rect 1765 22967 1823 22973
rect 1765 22933 1777 22967
rect 1811 22964 1823 22967
rect 1854 22964 1860 22976
rect 1811 22936 1860 22964
rect 1811 22933 1823 22936
rect 1765 22927 1823 22933
rect 1854 22924 1860 22936
rect 1912 22924 1918 22976
rect 2608 22964 2636 23063
rect 2682 23060 2688 23112
rect 2740 23060 2746 23112
rect 2869 23103 2927 23109
rect 2869 23069 2881 23103
rect 2915 23100 2927 23103
rect 3050 23100 3056 23112
rect 2915 23072 3056 23100
rect 2915 23069 2927 23072
rect 2869 23063 2927 23069
rect 3050 23060 3056 23072
rect 3108 23060 3114 23112
rect 3142 23060 3148 23112
rect 3200 23060 3206 23112
rect 3602 23060 3608 23112
rect 3660 23060 3666 23112
rect 4430 23060 4436 23112
rect 4488 23060 4494 23112
rect 4890 23060 4896 23112
rect 4948 23060 4954 23112
rect 5186 23079 5198 23113
rect 5232 23110 5244 23113
rect 5276 23110 5304 23140
rect 5721 23137 5733 23140
rect 5767 23137 5779 23171
rect 5828 23168 5856 23196
rect 6638 23168 6644 23180
rect 5828 23140 5948 23168
rect 5721 23131 5779 23137
rect 5232 23082 5304 23110
rect 5232 23079 5244 23082
rect 5186 23073 5244 23079
rect 5350 23060 5356 23112
rect 5408 23060 5414 23112
rect 5629 23103 5687 23109
rect 5629 23069 5641 23103
rect 5675 23100 5687 23103
rect 5810 23100 5816 23112
rect 5675 23072 5816 23100
rect 5675 23069 5687 23072
rect 5629 23063 5687 23069
rect 5810 23060 5816 23072
rect 5868 23060 5874 23112
rect 5920 23109 5948 23140
rect 6104 23140 6644 23168
rect 6104 23109 6132 23140
rect 6630 23128 6644 23140
rect 6696 23168 6702 23180
rect 6932 23168 6960 23208
rect 8018 23196 8024 23208
rect 8076 23196 8082 23248
rect 8128 23236 8156 23276
rect 9306 23264 9312 23316
rect 9364 23264 9370 23316
rect 14093 23307 14151 23313
rect 9646 23276 12204 23304
rect 9646 23236 9674 23276
rect 8128 23208 9674 23236
rect 12176 23236 12204 23276
rect 14093 23273 14105 23307
rect 14139 23304 14151 23307
rect 14182 23304 14188 23316
rect 14139 23276 14188 23304
rect 14139 23273 14151 23276
rect 14093 23267 14151 23273
rect 14182 23264 14188 23276
rect 14240 23264 14246 23316
rect 20162 23304 20168 23316
rect 14384 23276 20168 23304
rect 14384 23236 14412 23276
rect 20162 23264 20168 23276
rect 20220 23264 20226 23316
rect 20625 23307 20683 23313
rect 20625 23273 20637 23307
rect 20671 23304 20683 23307
rect 20714 23304 20720 23316
rect 20671 23276 20720 23304
rect 20671 23273 20683 23276
rect 20625 23267 20683 23273
rect 20714 23264 20720 23276
rect 20772 23264 20778 23316
rect 20806 23264 20812 23316
rect 20864 23264 20870 23316
rect 23290 23264 23296 23316
rect 23348 23304 23354 23316
rect 23845 23307 23903 23313
rect 23845 23304 23857 23307
rect 23348 23276 23857 23304
rect 23348 23264 23354 23276
rect 23845 23273 23857 23276
rect 23891 23304 23903 23307
rect 26050 23304 26056 23316
rect 23891 23276 26056 23304
rect 23891 23273 23903 23276
rect 23845 23267 23903 23273
rect 26050 23264 26056 23276
rect 26108 23264 26114 23316
rect 26326 23264 26332 23316
rect 26384 23304 26390 23316
rect 29178 23304 29184 23316
rect 26384 23276 29184 23304
rect 26384 23264 26390 23276
rect 29178 23264 29184 23276
rect 29236 23264 29242 23316
rect 30466 23264 30472 23316
rect 30524 23304 30530 23316
rect 35434 23304 35440 23316
rect 30524 23276 35440 23304
rect 30524 23264 30530 23276
rect 35434 23264 35440 23276
rect 35492 23304 35498 23316
rect 35713 23307 35771 23313
rect 35713 23304 35725 23307
rect 35492 23276 35725 23304
rect 35492 23264 35498 23276
rect 35713 23273 35725 23276
rect 35759 23273 35771 23307
rect 35713 23267 35771 23273
rect 19702 23236 19708 23248
rect 12176 23208 14412 23236
rect 14568 23208 19708 23236
rect 8113 23171 8171 23177
rect 8113 23168 8125 23171
rect 6696 23140 6960 23168
rect 6696 23128 6702 23140
rect 5905 23103 5963 23109
rect 5905 23069 5917 23103
rect 5951 23069 5963 23103
rect 5905 23063 5963 23069
rect 6089 23103 6147 23109
rect 6089 23069 6101 23103
rect 6135 23069 6147 23103
rect 6089 23063 6147 23069
rect 6181 23103 6239 23109
rect 6181 23069 6193 23103
rect 6227 23069 6239 23103
rect 6181 23063 6239 23069
rect 3237 23035 3295 23041
rect 3237 23001 3249 23035
rect 3283 23001 3295 23035
rect 3237 22995 3295 23001
rect 2866 22964 2872 22976
rect 2608 22936 2872 22964
rect 2866 22924 2872 22936
rect 2924 22924 2930 22976
rect 3252 22964 3280 22995
rect 3326 22992 3332 23044
rect 3384 22992 3390 23044
rect 3467 23035 3525 23041
rect 3467 23001 3479 23035
rect 3513 23032 3525 23035
rect 4338 23032 4344 23044
rect 3513 23004 4344 23032
rect 3513 23001 3525 23004
rect 3467 22995 3525 23001
rect 4338 22992 4344 23004
rect 4396 22992 4402 23044
rect 4522 22992 4528 23044
rect 4580 22992 4586 23044
rect 4614 22992 4620 23044
rect 4672 22992 4678 23044
rect 4735 23035 4793 23041
rect 4735 23032 4747 23035
rect 4724 23001 4747 23032
rect 4781 23001 4793 23035
rect 4724 22995 4793 23001
rect 3970 22964 3976 22976
rect 3252 22936 3976 22964
rect 3970 22924 3976 22936
rect 4028 22924 4034 22976
rect 4356 22964 4384 22992
rect 4724 22964 4752 22995
rect 5258 22992 5264 23044
rect 5316 22992 5322 23044
rect 5471 23035 5529 23041
rect 5471 23001 5483 23035
rect 5517 23001 5529 23035
rect 6196 23032 6224 23063
rect 6630 23041 6658 23128
rect 6932 23109 6960 23140
rect 7208 23140 8125 23168
rect 7208 23109 7236 23140
rect 8113 23137 8125 23140
rect 8159 23137 8171 23171
rect 8113 23131 8171 23137
rect 9122 23128 9128 23180
rect 9180 23168 9186 23180
rect 9180 23140 10548 23168
rect 9180 23128 9186 23140
rect 6733 23103 6791 23109
rect 6733 23069 6745 23103
rect 6779 23069 6791 23103
rect 6733 23063 6791 23069
rect 6917 23103 6975 23109
rect 6917 23069 6929 23103
rect 6963 23069 6975 23103
rect 6917 23063 6975 23069
rect 7193 23103 7251 23109
rect 7193 23069 7205 23103
rect 7239 23069 7251 23103
rect 7193 23063 7251 23069
rect 7653 23103 7711 23109
rect 7653 23069 7665 23103
rect 7699 23100 7711 23103
rect 7699 23072 8984 23100
rect 7699 23069 7711 23072
rect 7653 23063 7711 23069
rect 6425 23035 6483 23041
rect 6425 23032 6437 23035
rect 5471 22995 5529 23001
rect 5736 23004 6437 23032
rect 5486 22964 5514 22995
rect 5736 22976 5764 23004
rect 6425 23001 6437 23004
rect 6471 23001 6483 23035
rect 6630 23035 6699 23041
rect 6630 23004 6653 23035
rect 6425 22995 6483 23001
rect 6641 23001 6653 23004
rect 6687 23001 6699 23035
rect 6641 22995 6699 23001
rect 4356 22936 5514 22964
rect 5718 22924 5724 22976
rect 5776 22924 5782 22976
rect 6440 22964 6468 22995
rect 6748 22964 6776 23063
rect 6825 23035 6883 23041
rect 6825 23001 6837 23035
rect 6871 23032 6883 23035
rect 7285 23035 7343 23041
rect 7285 23032 7297 23035
rect 6871 23004 7297 23032
rect 6871 23001 6883 23004
rect 6825 22995 6883 23001
rect 7285 23001 7297 23004
rect 7331 23001 7343 23035
rect 7285 22995 7343 23001
rect 7374 22992 7380 23044
rect 7432 22992 7438 23044
rect 7466 22992 7472 23044
rect 7524 23041 7530 23044
rect 7524 23035 7553 23041
rect 7541 23001 7553 23035
rect 7524 22995 7553 23001
rect 7745 23035 7803 23041
rect 7745 23001 7757 23035
rect 7791 23001 7803 23035
rect 7745 22995 7803 23001
rect 7929 23035 7987 23041
rect 7929 23001 7941 23035
rect 7975 23032 7987 23035
rect 8018 23032 8024 23044
rect 7975 23004 8024 23032
rect 7975 23001 7987 23004
rect 7929 22995 7987 23001
rect 7524 22992 7530 22995
rect 7760 22964 7788 22995
rect 8018 22992 8024 23004
rect 8076 22992 8082 23044
rect 8956 22976 8984 23072
rect 9398 23060 9404 23112
rect 9456 23100 9462 23112
rect 9493 23103 9551 23109
rect 9493 23100 9505 23103
rect 9456 23072 9505 23100
rect 9456 23060 9462 23072
rect 9493 23069 9505 23072
rect 9539 23069 9551 23103
rect 9493 23063 9551 23069
rect 9585 23103 9643 23109
rect 9585 23069 9597 23103
rect 9631 23100 9643 23103
rect 9631 23072 9812 23100
rect 9631 23069 9643 23072
rect 9585 23063 9643 23069
rect 9674 22992 9680 23044
rect 9732 22992 9738 23044
rect 9784 23032 9812 23072
rect 9858 23060 9864 23112
rect 9916 23060 9922 23112
rect 10042 23060 10048 23112
rect 10100 23060 10106 23112
rect 10520 23109 10548 23140
rect 12434 23128 12440 23180
rect 12492 23168 12498 23180
rect 12805 23171 12863 23177
rect 12805 23168 12817 23171
rect 12492 23140 12817 23168
rect 12492 23128 12498 23140
rect 12805 23137 12817 23140
rect 12851 23168 12863 23171
rect 13906 23168 13912 23180
rect 12851 23140 13912 23168
rect 12851 23137 12863 23140
rect 12805 23131 12863 23137
rect 13906 23128 13912 23140
rect 13964 23128 13970 23180
rect 10505 23103 10563 23109
rect 10505 23069 10517 23103
rect 10551 23069 10563 23103
rect 10505 23063 10563 23069
rect 10597 23103 10655 23109
rect 10597 23069 10609 23103
rect 10643 23100 10655 23103
rect 10781 23103 10839 23109
rect 10781 23100 10793 23103
rect 10643 23072 10793 23100
rect 10643 23069 10655 23072
rect 10597 23063 10655 23069
rect 10781 23069 10793 23072
rect 10827 23069 10839 23103
rect 10781 23063 10839 23069
rect 10060 23032 10088 23060
rect 9784 23004 10088 23032
rect 11054 22992 11060 23044
rect 11112 22992 11118 23044
rect 11146 22992 11152 23044
rect 11204 23032 11210 23044
rect 11514 23032 11520 23044
rect 11204 23004 11520 23032
rect 11204 22992 11210 23004
rect 11514 22992 11520 23004
rect 11572 22992 11578 23044
rect 14274 22992 14280 23044
rect 14332 22992 14338 23044
rect 14458 22992 14464 23044
rect 14516 22992 14522 23044
rect 6440 22936 7788 22964
rect 8938 22924 8944 22976
rect 8996 22964 9002 22976
rect 14568 22964 14596 23208
rect 19702 23196 19708 23208
rect 19760 23196 19766 23248
rect 20070 23196 20076 23248
rect 20128 23236 20134 23248
rect 20128 23208 20576 23236
rect 20128 23196 20134 23208
rect 14734 23128 14740 23180
rect 14792 23128 14798 23180
rect 15473 23171 15531 23177
rect 15473 23137 15485 23171
rect 15519 23168 15531 23171
rect 16209 23171 16267 23177
rect 15519 23140 15976 23168
rect 15519 23137 15531 23140
rect 15473 23131 15531 23137
rect 15948 23112 15976 23140
rect 16209 23137 16221 23171
rect 16255 23168 16267 23171
rect 16298 23168 16304 23180
rect 16255 23140 16304 23168
rect 16255 23137 16267 23140
rect 16209 23131 16267 23137
rect 16298 23128 16304 23140
rect 16356 23128 16362 23180
rect 16684 23140 17632 23168
rect 15378 23060 15384 23112
rect 15436 23060 15442 23112
rect 15749 23103 15807 23109
rect 15749 23069 15761 23103
rect 15795 23069 15807 23103
rect 15749 23063 15807 23069
rect 15286 22992 15292 23044
rect 15344 23032 15350 23044
rect 15764 23032 15792 23063
rect 15838 23060 15844 23112
rect 15896 23060 15902 23112
rect 15930 23060 15936 23112
rect 15988 23060 15994 23112
rect 16684 23109 16712 23140
rect 17604 23112 17632 23140
rect 17954 23128 17960 23180
rect 18012 23168 18018 23180
rect 18693 23171 18751 23177
rect 18693 23168 18705 23171
rect 18012 23140 18705 23168
rect 18012 23128 18018 23140
rect 18693 23137 18705 23140
rect 18739 23168 18751 23171
rect 19978 23168 19984 23180
rect 18739 23140 19984 23168
rect 18739 23137 18751 23140
rect 18693 23131 18751 23137
rect 19978 23128 19984 23140
rect 20036 23128 20042 23180
rect 20548 23177 20576 23208
rect 23474 23196 23480 23248
rect 23532 23196 23538 23248
rect 27522 23196 27528 23248
rect 27580 23236 27586 23248
rect 34793 23239 34851 23245
rect 27580 23208 34752 23236
rect 27580 23196 27586 23208
rect 20533 23171 20591 23177
rect 20533 23137 20545 23171
rect 20579 23137 20591 23171
rect 20533 23131 20591 23137
rect 22005 23171 22063 23177
rect 22005 23137 22017 23171
rect 22051 23168 22063 23171
rect 22370 23168 22376 23180
rect 22051 23140 22376 23168
rect 22051 23137 22063 23140
rect 22005 23131 22063 23137
rect 22370 23128 22376 23140
rect 22428 23128 22434 23180
rect 22462 23128 22468 23180
rect 22520 23168 22526 23180
rect 22520 23140 23796 23168
rect 22520 23128 22526 23140
rect 16669 23103 16727 23109
rect 16669 23069 16681 23103
rect 16715 23069 16727 23103
rect 17037 23103 17095 23109
rect 17037 23100 17049 23103
rect 16669 23063 16727 23069
rect 16960 23072 17049 23100
rect 16960 23044 16988 23072
rect 17037 23069 17049 23072
rect 17083 23069 17095 23103
rect 17037 23063 17095 23069
rect 17126 23060 17132 23112
rect 17184 23060 17190 23112
rect 17310 23060 17316 23112
rect 17368 23060 17374 23112
rect 17586 23060 17592 23112
rect 17644 23060 17650 23112
rect 17678 23060 17684 23112
rect 17736 23060 17742 23112
rect 17862 23060 17868 23112
rect 17920 23100 17926 23112
rect 18049 23103 18107 23109
rect 18049 23100 18061 23103
rect 17920 23072 18061 23100
rect 17920 23060 17926 23072
rect 18049 23069 18061 23072
rect 18095 23069 18107 23103
rect 18049 23063 18107 23069
rect 18601 23103 18659 23109
rect 18601 23069 18613 23103
rect 18647 23100 18659 23103
rect 20346 23100 20352 23112
rect 18647 23072 20352 23100
rect 18647 23069 18659 23072
rect 18601 23063 18659 23069
rect 15344 23004 16160 23032
rect 15344 22992 15350 23004
rect 16132 22976 16160 23004
rect 16942 22992 16948 23044
rect 17000 22992 17006 23044
rect 17218 22992 17224 23044
rect 17276 23032 17282 23044
rect 18616 23032 18644 23063
rect 20346 23060 20352 23072
rect 20404 23100 20410 23112
rect 20441 23103 20499 23109
rect 20441 23100 20453 23103
rect 20404 23072 20453 23100
rect 20404 23060 20410 23072
rect 20441 23069 20453 23072
rect 20487 23069 20499 23103
rect 20441 23063 20499 23069
rect 20622 23060 20628 23112
rect 20680 23100 20686 23112
rect 21177 23103 21235 23109
rect 21177 23100 21189 23103
rect 20680 23072 21189 23100
rect 20680 23060 20686 23072
rect 21177 23069 21189 23072
rect 21223 23069 21235 23103
rect 21177 23063 21235 23069
rect 21729 23103 21787 23109
rect 21729 23069 21741 23103
rect 21775 23100 21787 23103
rect 22278 23100 22284 23112
rect 21775 23072 22284 23100
rect 21775 23069 21787 23072
rect 21729 23063 21787 23069
rect 22278 23060 22284 23072
rect 22336 23060 22342 23112
rect 22741 23103 22799 23109
rect 22741 23069 22753 23103
rect 22787 23069 22799 23103
rect 22741 23063 22799 23069
rect 17276 23004 18644 23032
rect 17276 22992 17282 23004
rect 19886 22992 19892 23044
rect 19944 23032 19950 23044
rect 20993 23035 21051 23041
rect 20993 23032 21005 23035
rect 19944 23004 21005 23032
rect 19944 22992 19950 23004
rect 20993 23001 21005 23004
rect 21039 23001 21051 23035
rect 20993 22995 21051 23001
rect 22646 22992 22652 23044
rect 22704 23032 22710 23044
rect 22756 23032 22784 23063
rect 22922 23060 22928 23112
rect 22980 23060 22986 23112
rect 23106 23060 23112 23112
rect 23164 23100 23170 23112
rect 23382 23100 23388 23112
rect 23164 23072 23388 23100
rect 23164 23060 23170 23072
rect 23382 23060 23388 23072
rect 23440 23060 23446 23112
rect 23566 23060 23572 23112
rect 23624 23060 23630 23112
rect 23768 23109 23796 23140
rect 23842 23128 23848 23180
rect 23900 23168 23906 23180
rect 25130 23168 25136 23180
rect 23900 23140 25136 23168
rect 23900 23128 23906 23140
rect 25130 23128 25136 23140
rect 25188 23168 25194 23180
rect 27614 23168 27620 23180
rect 25188 23140 25268 23168
rect 25188 23128 25194 23140
rect 23753 23103 23811 23109
rect 23753 23069 23765 23103
rect 23799 23069 23811 23103
rect 23753 23063 23811 23069
rect 23584 23032 23612 23060
rect 22704 23004 23612 23032
rect 22704 22992 22710 23004
rect 8996 22936 14596 22964
rect 8996 22924 9002 22936
rect 16114 22924 16120 22976
rect 16172 22924 16178 22976
rect 22002 22924 22008 22976
rect 22060 22964 22066 22976
rect 22278 22964 22284 22976
rect 22060 22936 22284 22964
rect 22060 22924 22066 22936
rect 22278 22924 22284 22936
rect 22336 22924 22342 22976
rect 22830 22924 22836 22976
rect 22888 22964 22894 22976
rect 23860 22964 23888 23128
rect 23937 23103 23995 23109
rect 23937 23069 23949 23103
rect 23983 23069 23995 23103
rect 23937 23063 23995 23069
rect 23952 23032 23980 23063
rect 24026 23060 24032 23112
rect 24084 23100 24090 23112
rect 24394 23100 24400 23112
rect 24084 23072 24400 23100
rect 24084 23060 24090 23072
rect 24394 23060 24400 23072
rect 24452 23100 24458 23112
rect 25240 23109 25268 23140
rect 25608 23140 27620 23168
rect 24949 23103 25007 23109
rect 24949 23100 24961 23103
rect 24452 23072 24961 23100
rect 24452 23060 24458 23072
rect 24949 23069 24961 23072
rect 24995 23069 25007 23103
rect 24949 23063 25007 23069
rect 25225 23103 25283 23109
rect 25225 23069 25237 23103
rect 25271 23069 25283 23103
rect 25225 23063 25283 23069
rect 23952 23004 24164 23032
rect 24136 22976 24164 23004
rect 22888 22936 23888 22964
rect 22888 22924 22894 22936
rect 24118 22924 24124 22976
rect 24176 22924 24182 22976
rect 25409 22967 25467 22973
rect 25409 22933 25421 22967
rect 25455 22964 25467 22967
rect 25608 22964 25636 23140
rect 27614 23128 27620 23140
rect 27672 23128 27678 23180
rect 34724 23168 34752 23208
rect 34793 23205 34805 23239
rect 34839 23236 34851 23239
rect 35158 23236 35164 23248
rect 34839 23208 35164 23236
rect 34839 23205 34851 23208
rect 34793 23199 34851 23205
rect 35158 23196 35164 23208
rect 35216 23196 35222 23248
rect 32416 23140 32904 23168
rect 34724 23140 35020 23168
rect 32416 23112 32444 23140
rect 25682 23060 25688 23112
rect 25740 23060 25746 23112
rect 26053 23103 26111 23109
rect 26053 23069 26065 23103
rect 26099 23100 26111 23103
rect 26142 23100 26148 23112
rect 26099 23072 26148 23100
rect 26099 23069 26111 23072
rect 26053 23063 26111 23069
rect 26142 23060 26148 23072
rect 26200 23060 26206 23112
rect 26970 23060 26976 23112
rect 27028 23060 27034 23112
rect 29730 23060 29736 23112
rect 29788 23060 29794 23112
rect 29914 23060 29920 23112
rect 29972 23060 29978 23112
rect 32306 23060 32312 23112
rect 32364 23060 32370 23112
rect 32398 23060 32404 23112
rect 32456 23060 32462 23112
rect 32490 23060 32496 23112
rect 32548 23060 32554 23112
rect 32766 23060 32772 23112
rect 32824 23060 32830 23112
rect 32876 23109 32904 23140
rect 34992 23112 35020 23140
rect 32861 23103 32919 23109
rect 32861 23069 32873 23103
rect 32907 23069 32919 23103
rect 32861 23063 32919 23069
rect 33045 23103 33103 23109
rect 33045 23069 33057 23103
rect 33091 23069 33103 23103
rect 33045 23063 33103 23069
rect 25869 23035 25927 23041
rect 25869 23001 25881 23035
rect 25915 23001 25927 23035
rect 25869 22995 25927 23001
rect 25455 22936 25636 22964
rect 25884 22964 25912 22995
rect 25958 22992 25964 23044
rect 26016 22992 26022 23044
rect 26988 23032 27016 23060
rect 27154 23032 27160 23044
rect 26068 23004 27160 23032
rect 26068 22976 26096 23004
rect 27154 22992 27160 23004
rect 27212 22992 27218 23044
rect 30006 22992 30012 23044
rect 30064 22992 30070 23044
rect 32324 23032 32352 23060
rect 32784 23032 32812 23060
rect 33060 23032 33088 23063
rect 34606 23060 34612 23112
rect 34664 23102 34670 23112
rect 34701 23103 34759 23109
rect 34701 23102 34713 23103
rect 34664 23074 34713 23102
rect 34664 23060 34670 23074
rect 34701 23069 34713 23074
rect 34747 23069 34759 23103
rect 34701 23063 34759 23069
rect 34974 23060 34980 23112
rect 35032 23060 35038 23112
rect 35345 23103 35403 23109
rect 35345 23069 35357 23103
rect 35391 23102 35403 23103
rect 35452 23102 35480 23264
rect 35529 23239 35587 23245
rect 35529 23205 35541 23239
rect 35575 23236 35587 23239
rect 35575 23208 35940 23236
rect 35575 23205 35587 23208
rect 35529 23199 35587 23205
rect 35621 23171 35679 23177
rect 35621 23168 35633 23171
rect 35544 23140 35633 23168
rect 35544 23112 35572 23140
rect 35621 23137 35633 23140
rect 35667 23137 35679 23171
rect 35621 23131 35679 23137
rect 35391 23074 35480 23102
rect 35391 23069 35403 23074
rect 35345 23063 35403 23069
rect 32324 23004 32720 23032
rect 32784 23004 33088 23032
rect 33229 23035 33287 23041
rect 26050 22964 26056 22976
rect 25884 22936 26056 22964
rect 25455 22933 25467 22936
rect 25409 22927 25467 22933
rect 26050 22924 26056 22936
rect 26108 22924 26114 22976
rect 26234 22924 26240 22976
rect 26292 22924 26298 22976
rect 31846 22924 31852 22976
rect 31904 22964 31910 22976
rect 32692 22973 32720 23004
rect 33229 23001 33241 23035
rect 33275 23032 33287 23035
rect 33318 23032 33324 23044
rect 33275 23004 33324 23032
rect 33275 23001 33287 23004
rect 33229 22995 33287 23001
rect 33318 22992 33324 23004
rect 33376 22992 33382 23044
rect 35161 23035 35219 23041
rect 35161 23001 35173 23035
rect 35207 23001 35219 23035
rect 35161 22995 35219 23001
rect 32309 22967 32367 22973
rect 32309 22964 32321 22967
rect 31904 22936 32321 22964
rect 31904 22924 31910 22936
rect 32309 22933 32321 22936
rect 32355 22933 32367 22967
rect 32309 22927 32367 22933
rect 32677 22967 32735 22973
rect 32677 22933 32689 22967
rect 32723 22964 32735 22967
rect 34790 22964 34796 22976
rect 32723 22936 34796 22964
rect 32723 22933 32735 22936
rect 32677 22927 32735 22933
rect 34790 22924 34796 22936
rect 34848 22924 34854 22976
rect 34882 22924 34888 22976
rect 34940 22964 34946 22976
rect 35176 22964 35204 22995
rect 35250 22992 35256 23044
rect 35308 22992 35314 23044
rect 35452 23032 35480 23074
rect 35526 23060 35532 23112
rect 35584 23060 35590 23112
rect 35912 23109 35940 23208
rect 36078 23196 36084 23248
rect 36136 23236 36142 23248
rect 36136 23208 36400 23236
rect 36136 23196 36142 23208
rect 35986 23128 35992 23180
rect 36044 23168 36050 23180
rect 36265 23171 36323 23177
rect 36265 23168 36277 23171
rect 36044 23140 36277 23168
rect 36044 23128 36050 23140
rect 36265 23137 36277 23140
rect 36311 23137 36323 23171
rect 36265 23131 36323 23137
rect 36372 23109 36400 23208
rect 35897 23103 35955 23109
rect 35897 23069 35909 23103
rect 35943 23069 35955 23103
rect 35897 23063 35955 23069
rect 36173 23103 36231 23109
rect 36173 23069 36185 23103
rect 36219 23069 36231 23103
rect 36173 23063 36231 23069
rect 36357 23103 36415 23109
rect 36357 23069 36369 23103
rect 36403 23069 36415 23103
rect 36357 23063 36415 23069
rect 36188 23032 36216 23063
rect 35452 23004 36216 23032
rect 35434 22964 35440 22976
rect 34940 22936 35440 22964
rect 34940 22924 34946 22936
rect 35434 22924 35440 22936
rect 35492 22924 35498 22976
rect 36078 22924 36084 22976
rect 36136 22924 36142 22976
rect 1104 22874 38272 22896
rect 1104 22822 4874 22874
rect 4926 22822 4938 22874
rect 4990 22822 5002 22874
rect 5054 22822 5066 22874
rect 5118 22822 5130 22874
rect 5182 22822 35594 22874
rect 35646 22822 35658 22874
rect 35710 22822 35722 22874
rect 35774 22822 35786 22874
rect 35838 22822 35850 22874
rect 35902 22822 38272 22874
rect 1104 22800 38272 22822
rect 2682 22720 2688 22772
rect 2740 22760 2746 22772
rect 2869 22763 2927 22769
rect 2869 22760 2881 22763
rect 2740 22732 2881 22760
rect 2740 22720 2746 22732
rect 2869 22729 2881 22732
rect 2915 22729 2927 22763
rect 2869 22723 2927 22729
rect 3142 22720 3148 22772
rect 3200 22760 3206 22772
rect 3421 22763 3479 22769
rect 3421 22760 3433 22763
rect 3200 22732 3433 22760
rect 3200 22720 3206 22732
rect 3421 22729 3433 22732
rect 3467 22729 3479 22763
rect 3421 22723 3479 22729
rect 3970 22720 3976 22772
rect 4028 22720 4034 22772
rect 4430 22720 4436 22772
rect 4488 22760 4494 22772
rect 5077 22763 5135 22769
rect 5077 22760 5089 22763
rect 4488 22732 5089 22760
rect 4488 22720 4494 22732
rect 5077 22729 5089 22732
rect 5123 22729 5135 22763
rect 5537 22763 5595 22769
rect 5537 22760 5549 22763
rect 5077 22723 5135 22729
rect 5184 22732 5549 22760
rect 2498 22652 2504 22704
rect 2556 22692 2562 22704
rect 2556 22664 3648 22692
rect 2556 22652 2562 22664
rect 2777 22627 2835 22633
rect 2777 22593 2789 22627
rect 2823 22593 2835 22627
rect 2777 22587 2835 22593
rect 2792 22556 2820 22587
rect 2958 22584 2964 22636
rect 3016 22584 3022 22636
rect 3620 22633 3648 22664
rect 4522 22652 4528 22704
rect 4580 22692 4586 22704
rect 4798 22692 4804 22704
rect 4580 22664 4804 22692
rect 4580 22652 4586 22664
rect 4798 22652 4804 22664
rect 4856 22692 4862 22704
rect 5184 22692 5212 22732
rect 5537 22729 5549 22732
rect 5583 22729 5595 22763
rect 5537 22723 5595 22729
rect 5626 22720 5632 22772
rect 5684 22720 5690 22772
rect 9493 22763 9551 22769
rect 9493 22729 9505 22763
rect 9539 22760 9551 22763
rect 9858 22760 9864 22772
rect 9539 22732 9864 22760
rect 9539 22729 9551 22732
rect 9493 22723 9551 22729
rect 9858 22720 9864 22732
rect 9916 22720 9922 22772
rect 11054 22720 11060 22772
rect 11112 22720 11118 22772
rect 11885 22763 11943 22769
rect 11885 22729 11897 22763
rect 11931 22760 11943 22763
rect 12434 22760 12440 22772
rect 11931 22732 12440 22760
rect 11931 22729 11943 22732
rect 11885 22723 11943 22729
rect 12434 22720 12440 22732
rect 12492 22720 12498 22772
rect 12526 22720 12532 22772
rect 12584 22760 12590 22772
rect 12989 22763 13047 22769
rect 12989 22760 13001 22763
rect 12584 22732 13001 22760
rect 12584 22720 12590 22732
rect 12989 22729 13001 22732
rect 13035 22729 13047 22763
rect 15286 22760 15292 22772
rect 12989 22723 13047 22729
rect 13372 22732 15292 22760
rect 4856 22664 5212 22692
rect 5445 22695 5503 22701
rect 4856 22652 4862 22664
rect 5445 22661 5457 22695
rect 5491 22692 5503 22695
rect 5644 22692 5672 22720
rect 5491 22664 5672 22692
rect 5491 22661 5503 22664
rect 5445 22655 5503 22661
rect 3605 22627 3663 22633
rect 3605 22593 3617 22627
rect 3651 22624 3663 22627
rect 3789 22627 3847 22633
rect 3651 22596 3740 22624
rect 3651 22593 3663 22596
rect 3605 22587 3663 22593
rect 3712 22568 3740 22596
rect 3789 22593 3801 22627
rect 3835 22624 3847 22627
rect 3878 22624 3884 22636
rect 3835 22596 3884 22624
rect 3835 22593 3847 22596
rect 3789 22587 3847 22593
rect 3878 22584 3884 22596
rect 3936 22584 3942 22636
rect 4065 22627 4123 22633
rect 4065 22593 4077 22627
rect 4111 22593 4123 22627
rect 4065 22587 4123 22593
rect 2866 22556 2872 22568
rect 2792 22528 2872 22556
rect 2866 22516 2872 22528
rect 2924 22516 2930 22568
rect 3694 22516 3700 22568
rect 3752 22556 3758 22568
rect 4080 22556 4108 22587
rect 4706 22584 4712 22636
rect 4764 22624 4770 22636
rect 5258 22624 5264 22636
rect 4764 22596 5264 22624
rect 4764 22584 4770 22596
rect 5258 22584 5264 22596
rect 5316 22624 5322 22636
rect 5537 22627 5595 22633
rect 5537 22624 5549 22627
rect 5316 22596 5549 22624
rect 5316 22584 5322 22596
rect 5537 22593 5549 22596
rect 5583 22593 5595 22627
rect 5644 22624 5672 22664
rect 6365 22695 6423 22701
rect 6365 22661 6377 22695
rect 6411 22692 6423 22695
rect 7742 22692 7748 22704
rect 6411 22664 7748 22692
rect 6411 22661 6423 22664
rect 6365 22655 6423 22661
rect 7742 22652 7748 22664
rect 7800 22692 7806 22704
rect 7837 22695 7895 22701
rect 7837 22692 7849 22695
rect 7800 22664 7849 22692
rect 7800 22652 7806 22664
rect 7837 22661 7849 22664
rect 7883 22661 7895 22695
rect 7837 22655 7895 22661
rect 7944 22664 12572 22692
rect 5721 22627 5779 22633
rect 5721 22624 5733 22627
rect 5644 22596 5733 22624
rect 5537 22587 5595 22593
rect 5721 22593 5733 22596
rect 5767 22593 5779 22627
rect 5721 22587 5779 22593
rect 6454 22584 6460 22636
rect 6512 22624 6518 22636
rect 6549 22627 6607 22633
rect 6549 22624 6561 22627
rect 6512 22596 6561 22624
rect 6512 22584 6518 22596
rect 6549 22593 6561 22596
rect 6595 22593 6607 22627
rect 6549 22587 6607 22593
rect 6733 22627 6791 22633
rect 6733 22593 6745 22627
rect 6779 22624 6791 22627
rect 7944 22624 7972 22664
rect 6779 22596 7972 22624
rect 6779 22593 6791 22596
rect 6733 22587 6791 22593
rect 8018 22584 8024 22636
rect 8076 22584 8082 22636
rect 8570 22584 8576 22636
rect 8628 22624 8634 22636
rect 9677 22627 9735 22633
rect 9677 22624 9689 22627
rect 8628 22596 9689 22624
rect 8628 22584 8634 22596
rect 9677 22593 9689 22596
rect 9723 22624 9735 22627
rect 11241 22627 11299 22633
rect 9723 22596 10088 22624
rect 9723 22593 9735 22596
rect 9677 22587 9735 22593
rect 3752 22528 4108 22556
rect 3752 22516 3758 22528
rect 5350 22516 5356 22568
rect 5408 22556 5414 22568
rect 7374 22556 7380 22568
rect 5408 22528 7380 22556
rect 5408 22516 5414 22528
rect 7374 22516 7380 22528
rect 7432 22516 7438 22568
rect 9953 22559 10011 22565
rect 9953 22525 9965 22559
rect 9999 22525 10011 22559
rect 10060 22556 10088 22596
rect 11241 22593 11253 22627
rect 11287 22624 11299 22627
rect 11422 22624 11428 22636
rect 11287 22596 11428 22624
rect 11287 22593 11299 22596
rect 11241 22587 11299 22593
rect 11422 22584 11428 22596
rect 11480 22584 11486 22636
rect 12544 22633 12572 22664
rect 12345 22627 12403 22633
rect 11900 22596 12112 22624
rect 11900 22556 11928 22596
rect 12084 22568 12112 22596
rect 12345 22593 12357 22627
rect 12391 22593 12403 22627
rect 12345 22587 12403 22593
rect 12529 22627 12587 22633
rect 12529 22593 12541 22627
rect 12575 22593 12587 22627
rect 12529 22587 12587 22593
rect 10060 22528 11928 22556
rect 9953 22519 10011 22525
rect 3326 22448 3332 22500
rect 3384 22488 3390 22500
rect 4614 22488 4620 22500
rect 3384 22460 4620 22488
rect 3384 22448 3390 22460
rect 4614 22448 4620 22460
rect 4672 22448 4678 22500
rect 8202 22448 8208 22500
rect 8260 22448 8266 22500
rect 9968 22488 9996 22519
rect 11974 22516 11980 22568
rect 12032 22516 12038 22568
rect 12066 22516 12072 22568
rect 12124 22516 12130 22568
rect 10042 22488 10048 22500
rect 9968 22460 10048 22488
rect 10042 22448 10048 22460
rect 10100 22448 10106 22500
rect 11422 22448 11428 22500
rect 11480 22488 11486 22500
rect 11517 22491 11575 22497
rect 11517 22488 11529 22491
rect 11480 22460 11529 22488
rect 11480 22448 11486 22460
rect 11517 22457 11529 22460
rect 11563 22457 11575 22491
rect 11517 22451 11575 22457
rect 11606 22448 11612 22500
rect 11664 22488 11670 22500
rect 12360 22488 12388 22587
rect 12618 22584 12624 22636
rect 12676 22584 12682 22636
rect 13372 22633 13400 22732
rect 15286 22720 15292 22732
rect 15344 22720 15350 22772
rect 15473 22763 15531 22769
rect 15473 22729 15485 22763
rect 15519 22760 15531 22763
rect 15746 22760 15752 22772
rect 15519 22732 15752 22760
rect 15519 22729 15531 22732
rect 15473 22723 15531 22729
rect 15746 22720 15752 22732
rect 15804 22720 15810 22772
rect 17957 22763 18015 22769
rect 17957 22729 17969 22763
rect 18003 22760 18015 22763
rect 18506 22760 18512 22772
rect 18003 22732 18512 22760
rect 18003 22729 18015 22732
rect 17957 22723 18015 22729
rect 18506 22720 18512 22732
rect 18564 22720 18570 22772
rect 22097 22763 22155 22769
rect 22097 22729 22109 22763
rect 22143 22760 22155 22763
rect 22922 22760 22928 22772
rect 22143 22732 22928 22760
rect 22143 22729 22155 22732
rect 22097 22723 22155 22729
rect 22922 22720 22928 22732
rect 22980 22720 22986 22772
rect 23750 22720 23756 22772
rect 23808 22760 23814 22772
rect 24397 22763 24455 22769
rect 24397 22760 24409 22763
rect 23808 22732 24409 22760
rect 23808 22720 23814 22732
rect 24397 22729 24409 22732
rect 24443 22729 24455 22763
rect 24397 22723 24455 22729
rect 25866 22720 25872 22772
rect 25924 22720 25930 22772
rect 26234 22720 26240 22772
rect 26292 22720 26298 22772
rect 27522 22720 27528 22772
rect 27580 22720 27586 22772
rect 27982 22720 27988 22772
rect 28040 22720 28046 22772
rect 29914 22720 29920 22772
rect 29972 22760 29978 22772
rect 30285 22763 30343 22769
rect 30285 22760 30297 22763
rect 29972 22732 30297 22760
rect 29972 22720 29978 22732
rect 30285 22729 30297 22732
rect 30331 22729 30343 22763
rect 30285 22723 30343 22729
rect 32217 22763 32275 22769
rect 32217 22729 32229 22763
rect 32263 22760 32275 22763
rect 32490 22760 32496 22772
rect 32263 22732 32496 22760
rect 32263 22729 32275 22732
rect 32217 22723 32275 22729
rect 32490 22720 32496 22732
rect 32548 22720 32554 22772
rect 34698 22720 34704 22772
rect 34756 22760 34762 22772
rect 35342 22760 35348 22772
rect 34756 22732 35348 22760
rect 34756 22720 34762 22732
rect 35342 22720 35348 22732
rect 35400 22720 35406 22772
rect 35434 22720 35440 22772
rect 35492 22760 35498 22772
rect 37369 22763 37427 22769
rect 37369 22760 37381 22763
rect 35492 22732 36216 22760
rect 35492 22720 35498 22732
rect 13633 22695 13691 22701
rect 13633 22661 13645 22695
rect 13679 22692 13691 22695
rect 14274 22692 14280 22704
rect 13679 22664 14280 22692
rect 13679 22661 13691 22664
rect 13633 22655 13691 22661
rect 12713 22627 12771 22633
rect 12713 22593 12725 22627
rect 12759 22593 12771 22627
rect 12713 22587 12771 22593
rect 13357 22627 13415 22633
rect 13357 22593 13369 22627
rect 13403 22593 13415 22627
rect 13357 22587 13415 22593
rect 12728 22556 12756 22587
rect 13538 22584 13544 22636
rect 13596 22584 13602 22636
rect 14200 22633 14228 22664
rect 14274 22652 14280 22664
rect 14332 22652 14338 22704
rect 14384 22664 17448 22692
rect 14185 22627 14243 22633
rect 14185 22593 14197 22627
rect 14231 22593 14243 22627
rect 14185 22587 14243 22593
rect 14384 22556 14412 22664
rect 14458 22584 14464 22636
rect 14516 22624 14522 22636
rect 14553 22627 14611 22633
rect 14553 22624 14565 22627
rect 14516 22596 14565 22624
rect 14516 22584 14522 22596
rect 14553 22593 14565 22596
rect 14599 22593 14611 22627
rect 14553 22587 14611 22593
rect 12728 22528 14412 22556
rect 11664 22460 12388 22488
rect 11664 22448 11670 22460
rect 14090 22448 14096 22500
rect 14148 22488 14154 22500
rect 14568 22488 14596 22587
rect 15194 22584 15200 22636
rect 15252 22624 15258 22636
rect 15411 22627 15469 22633
rect 15411 22624 15423 22627
rect 15252 22596 15423 22624
rect 15252 22584 15258 22596
rect 15411 22593 15423 22596
rect 15457 22593 15469 22627
rect 15411 22587 15469 22593
rect 16114 22584 16120 22636
rect 16172 22584 16178 22636
rect 16301 22627 16359 22633
rect 16301 22593 16313 22627
rect 16347 22624 16359 22627
rect 16666 22624 16672 22636
rect 16347 22596 16672 22624
rect 16347 22593 16359 22596
rect 16301 22587 16359 22593
rect 16666 22584 16672 22596
rect 16724 22584 16730 22636
rect 16850 22584 16856 22636
rect 16908 22624 16914 22636
rect 17126 22624 17132 22636
rect 16908 22596 17132 22624
rect 16908 22584 16914 22596
rect 17126 22584 17132 22596
rect 17184 22584 17190 22636
rect 17313 22627 17371 22633
rect 17313 22593 17325 22627
rect 17359 22593 17371 22627
rect 17313 22587 17371 22593
rect 14642 22516 14648 22568
rect 14700 22516 14706 22568
rect 15930 22516 15936 22568
rect 15988 22556 15994 22568
rect 16390 22556 16396 22568
rect 15988 22528 16396 22556
rect 15988 22516 15994 22528
rect 16390 22516 16396 22528
rect 16448 22516 16454 22568
rect 16485 22559 16543 22565
rect 16485 22525 16497 22559
rect 16531 22556 16543 22559
rect 16942 22556 16948 22568
rect 16531 22528 16948 22556
rect 16531 22525 16543 22528
rect 16485 22519 16543 22525
rect 16942 22516 16948 22528
rect 17000 22556 17006 22568
rect 17328 22556 17356 22587
rect 17000 22528 17356 22556
rect 17420 22556 17448 22664
rect 20346 22652 20352 22704
rect 20404 22652 20410 22704
rect 22020 22664 22600 22692
rect 17586 22584 17592 22636
rect 17644 22624 17650 22636
rect 17865 22627 17923 22633
rect 17865 22624 17877 22627
rect 17644 22596 17877 22624
rect 17644 22584 17650 22596
rect 17865 22593 17877 22596
rect 17911 22593 17923 22627
rect 17865 22587 17923 22593
rect 20714 22584 20720 22636
rect 20772 22584 20778 22636
rect 21910 22584 21916 22636
rect 21968 22624 21974 22636
rect 22020 22633 22048 22664
rect 22005 22627 22063 22633
rect 22005 22624 22017 22627
rect 21968 22596 22017 22624
rect 21968 22584 21974 22596
rect 22005 22593 22017 22596
rect 22051 22593 22063 22627
rect 22005 22587 22063 22593
rect 22186 22584 22192 22636
rect 22244 22624 22250 22636
rect 22462 22624 22468 22636
rect 22244 22596 22468 22624
rect 22244 22584 22250 22596
rect 22462 22584 22468 22596
rect 22520 22584 22526 22636
rect 22572 22633 22600 22664
rect 22940 22664 24532 22692
rect 22940 22636 22968 22664
rect 22557 22627 22615 22633
rect 22557 22593 22569 22627
rect 22603 22593 22615 22627
rect 22557 22587 22615 22593
rect 22649 22627 22707 22633
rect 22649 22593 22661 22627
rect 22695 22624 22707 22627
rect 22830 22624 22836 22636
rect 22695 22596 22836 22624
rect 22695 22593 22707 22596
rect 22649 22587 22707 22593
rect 22572 22556 22600 22587
rect 22830 22584 22836 22596
rect 22888 22584 22894 22636
rect 22922 22584 22928 22636
rect 22980 22584 22986 22636
rect 23290 22584 23296 22636
rect 23348 22584 23354 22636
rect 23658 22584 23664 22636
rect 23716 22584 23722 22636
rect 24026 22584 24032 22636
rect 24084 22584 24090 22636
rect 24504 22633 24532 22664
rect 24305 22627 24363 22633
rect 24305 22593 24317 22627
rect 24351 22593 24363 22627
rect 24305 22587 24363 22593
rect 24489 22627 24547 22633
rect 24489 22593 24501 22627
rect 24535 22593 24547 22627
rect 24489 22587 24547 22593
rect 24118 22556 24124 22568
rect 17420 22528 19334 22556
rect 22572 22528 24124 22556
rect 17000 22516 17006 22528
rect 15841 22491 15899 22497
rect 15841 22488 15853 22491
rect 14148 22460 14596 22488
rect 14844 22460 15853 22488
rect 14148 22448 14154 22460
rect 14844 22432 14872 22460
rect 15841 22457 15853 22460
rect 15887 22488 15899 22491
rect 18138 22488 18144 22500
rect 15887 22460 18144 22488
rect 15887 22457 15899 22460
rect 15841 22451 15899 22457
rect 18138 22448 18144 22460
rect 18196 22448 18202 22500
rect 4338 22380 4344 22432
rect 4396 22420 4402 22432
rect 4706 22420 4712 22432
rect 4396 22392 4712 22420
rect 4396 22380 4402 22392
rect 4706 22380 4712 22392
rect 4764 22380 4770 22432
rect 5810 22380 5816 22432
rect 5868 22420 5874 22432
rect 7650 22420 7656 22432
rect 5868 22392 7656 22420
rect 5868 22380 5874 22392
rect 7650 22380 7656 22392
rect 7708 22380 7714 22432
rect 9861 22423 9919 22429
rect 9861 22389 9873 22423
rect 9907 22420 9919 22423
rect 10134 22420 10140 22432
rect 9907 22392 10140 22420
rect 9907 22389 9919 22392
rect 9861 22383 9919 22389
rect 10134 22380 10140 22392
rect 10192 22380 10198 22432
rect 14826 22380 14832 22432
rect 14884 22380 14890 22432
rect 15010 22380 15016 22432
rect 15068 22420 15074 22432
rect 15289 22423 15347 22429
rect 15289 22420 15301 22423
rect 15068 22392 15301 22420
rect 15068 22380 15074 22392
rect 15289 22389 15301 22392
rect 15335 22389 15347 22423
rect 19306 22420 19334 22528
rect 24118 22516 24124 22528
rect 24176 22556 24182 22568
rect 24320 22556 24348 22587
rect 25406 22584 25412 22636
rect 25464 22584 25470 22636
rect 25593 22627 25651 22633
rect 25593 22593 25605 22627
rect 25639 22624 25651 22627
rect 25884 22624 25912 22720
rect 26252 22692 26280 22720
rect 26252 22664 30696 22692
rect 26510 22624 26516 22636
rect 25639 22596 26516 22624
rect 25639 22593 25651 22596
rect 25593 22587 25651 22593
rect 26510 22584 26516 22596
rect 26568 22584 26574 22636
rect 26602 22584 26608 22636
rect 26660 22624 26666 22636
rect 26973 22627 27031 22633
rect 26973 22624 26985 22627
rect 26660 22596 26985 22624
rect 26660 22584 26666 22596
rect 26973 22593 26985 22596
rect 27019 22593 27031 22627
rect 26973 22587 27031 22593
rect 27154 22584 27160 22636
rect 27212 22584 27218 22636
rect 27249 22627 27307 22633
rect 27249 22593 27261 22627
rect 27295 22593 27307 22627
rect 27249 22587 27307 22593
rect 24176 22528 24348 22556
rect 25424 22556 25452 22584
rect 25774 22556 25780 22568
rect 25424 22528 25780 22556
rect 24176 22516 24182 22528
rect 25774 22516 25780 22528
rect 25832 22516 25838 22568
rect 26142 22516 26148 22568
rect 26200 22516 26206 22568
rect 26234 22516 26240 22568
rect 26292 22556 26298 22568
rect 27264 22556 27292 22587
rect 27338 22584 27344 22636
rect 27396 22584 27402 22636
rect 27430 22584 27436 22636
rect 27488 22624 27494 22636
rect 29656 22633 29684 22664
rect 27709 22627 27767 22633
rect 27709 22624 27721 22627
rect 27488 22596 27721 22624
rect 27488 22584 27494 22596
rect 27709 22593 27721 22596
rect 27755 22593 27767 22627
rect 27709 22587 27767 22593
rect 29641 22627 29699 22633
rect 29641 22593 29653 22627
rect 29687 22593 29699 22627
rect 29641 22587 29699 22593
rect 29825 22627 29883 22633
rect 29825 22593 29837 22627
rect 29871 22624 29883 22627
rect 29917 22627 29975 22633
rect 29917 22624 29929 22627
rect 29871 22596 29929 22624
rect 29871 22593 29883 22596
rect 29825 22587 29883 22593
rect 29917 22593 29929 22596
rect 29963 22624 29975 22627
rect 30190 22624 30196 22636
rect 29963 22596 30196 22624
rect 29963 22593 29975 22596
rect 29917 22587 29975 22593
rect 30190 22584 30196 22596
rect 30248 22584 30254 22636
rect 30392 22633 30420 22664
rect 30668 22633 30696 22664
rect 32398 22652 32404 22704
rect 32456 22652 32462 22704
rect 33689 22695 33747 22701
rect 33689 22692 33701 22695
rect 32784 22664 33701 22692
rect 30377 22627 30435 22633
rect 30377 22593 30389 22627
rect 30423 22593 30435 22627
rect 30377 22587 30435 22593
rect 30469 22627 30527 22633
rect 30469 22593 30481 22627
rect 30515 22593 30527 22627
rect 30469 22587 30527 22593
rect 30653 22627 30711 22633
rect 30653 22593 30665 22627
rect 30699 22593 30711 22627
rect 30653 22587 30711 22593
rect 26292 22528 27292 22556
rect 26292 22516 26298 22528
rect 23934 22448 23940 22500
rect 23992 22448 23998 22500
rect 26160 22488 26188 22516
rect 27356 22488 27384 22584
rect 30009 22559 30067 22565
rect 30009 22525 30021 22559
rect 30055 22556 30067 22559
rect 30484 22556 30512 22587
rect 31938 22584 31944 22636
rect 31996 22624 32002 22636
rect 32125 22627 32183 22633
rect 32125 22624 32137 22627
rect 31996 22596 32137 22624
rect 31996 22584 32002 22596
rect 32125 22593 32137 22596
rect 32171 22593 32183 22627
rect 32125 22587 32183 22593
rect 32309 22627 32367 22633
rect 32309 22593 32321 22627
rect 32355 22624 32367 22627
rect 32416 22624 32444 22652
rect 32355 22596 32444 22624
rect 32355 22593 32367 22596
rect 32309 22587 32367 22593
rect 32490 22584 32496 22636
rect 32548 22624 32554 22636
rect 32784 22633 32812 22664
rect 33689 22661 33701 22664
rect 33735 22661 33747 22695
rect 33689 22655 33747 22661
rect 35161 22695 35219 22701
rect 35161 22661 35173 22695
rect 35207 22692 35219 22695
rect 35986 22692 35992 22704
rect 35207 22664 35992 22692
rect 35207 22661 35219 22664
rect 35161 22655 35219 22661
rect 35986 22652 35992 22664
rect 36044 22652 36050 22704
rect 32769 22627 32827 22633
rect 32769 22624 32781 22627
rect 32548 22596 32781 22624
rect 32548 22584 32554 22596
rect 32769 22593 32781 22596
rect 32815 22593 32827 22627
rect 32769 22587 32827 22593
rect 32858 22584 32864 22636
rect 32916 22584 32922 22636
rect 33137 22627 33195 22633
rect 33137 22593 33149 22627
rect 33183 22593 33195 22627
rect 33137 22587 33195 22593
rect 30055 22528 30512 22556
rect 30055 22525 30067 22528
rect 30009 22519 30067 22525
rect 31846 22516 31852 22568
rect 31904 22556 31910 22568
rect 32677 22559 32735 22565
rect 32677 22556 32689 22559
rect 31904 22528 32689 22556
rect 31904 22516 31910 22528
rect 32677 22525 32689 22528
rect 32723 22525 32735 22559
rect 32677 22519 32735 22525
rect 32950 22516 32956 22568
rect 33008 22516 33014 22568
rect 24964 22460 26096 22488
rect 26160 22460 27384 22488
rect 24964 22432 24992 22460
rect 24946 22420 24952 22432
rect 19306 22392 24952 22420
rect 15289 22383 15347 22389
rect 24946 22380 24952 22392
rect 25004 22380 25010 22432
rect 25406 22380 25412 22432
rect 25464 22380 25470 22432
rect 26068 22420 26096 22460
rect 31938 22448 31944 22500
rect 31996 22488 32002 22500
rect 33152 22488 33180 22587
rect 33226 22584 33232 22636
rect 33284 22584 33290 22636
rect 33318 22584 33324 22636
rect 33376 22624 33382 22636
rect 33413 22627 33471 22633
rect 33413 22624 33425 22627
rect 33376 22596 33425 22624
rect 33376 22584 33382 22596
rect 33413 22593 33425 22596
rect 33459 22593 33471 22627
rect 33413 22587 33471 22593
rect 33505 22627 33563 22633
rect 33505 22593 33517 22627
rect 33551 22624 33563 22627
rect 34422 22624 34428 22636
rect 33551 22596 34428 22624
rect 33551 22593 33563 22596
rect 33505 22587 33563 22593
rect 34422 22584 34428 22596
rect 34480 22584 34486 22636
rect 34974 22584 34980 22636
rect 35032 22584 35038 22636
rect 35434 22584 35440 22636
rect 35492 22584 35498 22636
rect 36081 22627 36139 22633
rect 36081 22593 36093 22627
rect 36127 22593 36139 22627
rect 36081 22587 36139 22593
rect 34992 22556 35020 22584
rect 36096 22556 36124 22587
rect 34992 22528 36124 22556
rect 36188 22556 36216 22732
rect 36280 22732 37381 22760
rect 36280 22633 36308 22732
rect 37369 22729 37381 22732
rect 37415 22729 37427 22763
rect 37369 22723 37427 22729
rect 36817 22695 36875 22701
rect 36817 22692 36829 22695
rect 36464 22664 36829 22692
rect 36265 22627 36323 22633
rect 36265 22593 36277 22627
rect 36311 22593 36323 22627
rect 36265 22587 36323 22593
rect 36357 22627 36415 22633
rect 36357 22593 36369 22627
rect 36403 22624 36415 22627
rect 36464 22624 36492 22664
rect 36817 22661 36829 22664
rect 36863 22692 36875 22695
rect 36863 22664 37320 22692
rect 36863 22661 36875 22664
rect 36817 22655 36875 22661
rect 37292 22633 37320 22664
rect 36403 22596 36492 22624
rect 36541 22627 36599 22633
rect 36403 22593 36415 22596
rect 36357 22587 36415 22593
rect 36541 22593 36553 22627
rect 36587 22624 36599 22627
rect 36633 22627 36691 22633
rect 36633 22624 36645 22627
rect 36587 22596 36645 22624
rect 36587 22593 36599 22596
rect 36541 22587 36599 22593
rect 36633 22593 36645 22596
rect 36679 22593 36691 22627
rect 36633 22587 36691 22593
rect 37277 22627 37335 22633
rect 37277 22593 37289 22627
rect 37323 22593 37335 22627
rect 37277 22587 37335 22593
rect 36372 22556 36400 22587
rect 36188 22528 36400 22556
rect 31996 22460 33180 22488
rect 36096 22488 36124 22528
rect 36556 22488 36584 22587
rect 37550 22584 37556 22636
rect 37608 22624 37614 22636
rect 37645 22627 37703 22633
rect 37645 22624 37657 22627
rect 37608 22596 37657 22624
rect 37608 22584 37614 22596
rect 37645 22593 37657 22596
rect 37691 22593 37703 22627
rect 37645 22587 37703 22593
rect 36096 22460 36584 22488
rect 31996 22448 32002 22460
rect 37826 22448 37832 22500
rect 37884 22448 37890 22500
rect 28166 22420 28172 22432
rect 26068 22392 28172 22420
rect 28166 22380 28172 22392
rect 28224 22380 28230 22432
rect 29457 22423 29515 22429
rect 29457 22389 29469 22423
rect 29503 22420 29515 22423
rect 29730 22420 29736 22432
rect 29503 22392 29736 22420
rect 29503 22389 29515 22392
rect 29457 22383 29515 22389
rect 29730 22380 29736 22392
rect 29788 22380 29794 22432
rect 30650 22380 30656 22432
rect 30708 22380 30714 22432
rect 32030 22380 32036 22432
rect 32088 22420 32094 22432
rect 32398 22420 32404 22432
rect 32088 22392 32404 22420
rect 32088 22380 32094 22392
rect 32398 22380 32404 22392
rect 32456 22380 32462 22432
rect 32490 22380 32496 22432
rect 32548 22380 32554 22432
rect 34790 22380 34796 22432
rect 34848 22420 34854 22432
rect 35161 22423 35219 22429
rect 35161 22420 35173 22423
rect 34848 22392 35173 22420
rect 34848 22380 34854 22392
rect 35161 22389 35173 22392
rect 35207 22389 35219 22423
rect 35161 22383 35219 22389
rect 36078 22380 36084 22432
rect 36136 22380 36142 22432
rect 36446 22380 36452 22432
rect 36504 22380 36510 22432
rect 36998 22380 37004 22432
rect 37056 22380 37062 22432
rect 1104 22330 38272 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 38272 22330
rect 1104 22256 38272 22278
rect 3602 22176 3608 22228
rect 3660 22216 3666 22228
rect 3973 22219 4031 22225
rect 3973 22216 3985 22219
rect 3660 22188 3985 22216
rect 3660 22176 3666 22188
rect 3973 22185 3985 22188
rect 4019 22185 4031 22219
rect 3973 22179 4031 22185
rect 9674 22176 9680 22228
rect 9732 22216 9738 22228
rect 10321 22219 10379 22225
rect 10321 22216 10333 22219
rect 9732 22188 10333 22216
rect 9732 22176 9738 22188
rect 10321 22185 10333 22188
rect 10367 22185 10379 22219
rect 10321 22179 10379 22185
rect 11974 22176 11980 22228
rect 12032 22216 12038 22228
rect 12161 22219 12219 22225
rect 12161 22216 12173 22219
rect 12032 22188 12173 22216
rect 12032 22176 12038 22188
rect 12161 22185 12173 22188
rect 12207 22185 12219 22219
rect 26234 22216 26240 22228
rect 12161 22179 12219 22185
rect 12406 22188 26240 22216
rect 3050 22108 3056 22160
rect 3108 22148 3114 22160
rect 3418 22148 3424 22160
rect 3108 22120 3424 22148
rect 3108 22108 3114 22120
rect 3418 22108 3424 22120
rect 3476 22148 3482 22160
rect 6178 22148 6184 22160
rect 3476 22120 6184 22148
rect 3476 22108 3482 22120
rect 6178 22108 6184 22120
rect 6236 22108 6242 22160
rect 12406 22148 12434 22188
rect 26234 22176 26240 22188
rect 26292 22176 26298 22228
rect 27154 22176 27160 22228
rect 27212 22216 27218 22228
rect 27706 22216 27712 22228
rect 27212 22188 27712 22216
rect 27212 22176 27218 22188
rect 27706 22176 27712 22188
rect 27764 22176 27770 22228
rect 29181 22219 29239 22225
rect 29181 22185 29193 22219
rect 29227 22216 29239 22219
rect 29270 22216 29276 22228
rect 29227 22188 29276 22216
rect 29227 22185 29239 22188
rect 29181 22179 29239 22185
rect 29270 22176 29276 22188
rect 29328 22176 29334 22228
rect 32858 22176 32864 22228
rect 32916 22176 32922 22228
rect 36262 22216 36268 22228
rect 35728 22188 36268 22216
rect 9646 22120 12434 22148
rect 3786 22040 3792 22092
rect 3844 22080 3850 22092
rect 6270 22080 6276 22092
rect 3844 22052 6276 22080
rect 3844 22040 3850 22052
rect 6270 22040 6276 22052
rect 6328 22080 6334 22092
rect 9646 22080 9674 22120
rect 14550 22108 14556 22160
rect 14608 22108 14614 22160
rect 14642 22108 14648 22160
rect 14700 22148 14706 22160
rect 16022 22148 16028 22160
rect 14700 22120 16028 22148
rect 14700 22108 14706 22120
rect 16022 22108 16028 22120
rect 16080 22108 16086 22160
rect 16298 22108 16304 22160
rect 16356 22148 16362 22160
rect 16356 22120 16528 22148
rect 16356 22108 16362 22120
rect 6328 22052 9674 22080
rect 6328 22040 6334 22052
rect 10042 22040 10048 22092
rect 10100 22080 10106 22092
rect 11609 22083 11667 22089
rect 11609 22080 11621 22083
rect 10100 22052 11621 22080
rect 10100 22040 10106 22052
rect 1946 21972 1952 22024
rect 2004 21972 2010 22024
rect 4249 22015 4307 22021
rect 4249 22012 4261 22015
rect 4172 21984 4261 22012
rect 3786 21904 3792 21956
rect 3844 21904 3850 21956
rect 1762 21836 1768 21888
rect 1820 21836 1826 21888
rect 3878 21836 3884 21888
rect 3936 21876 3942 21888
rect 4172 21885 4200 21984
rect 4249 21981 4261 21984
rect 4295 22012 4307 22015
rect 5718 22012 5724 22024
rect 4295 21984 5724 22012
rect 4295 21981 4307 21984
rect 4249 21975 4307 21981
rect 5718 21972 5724 21984
rect 5776 21972 5782 22024
rect 5810 21972 5816 22024
rect 5868 22012 5874 22024
rect 10244 22021 10272 22052
rect 11609 22049 11621 22052
rect 11655 22049 11667 22083
rect 11609 22043 11667 22049
rect 7745 22015 7803 22021
rect 7745 22012 7757 22015
rect 5868 21984 7757 22012
rect 5868 21972 5874 21984
rect 7745 21981 7757 21984
rect 7791 21981 7803 22015
rect 7745 21975 7803 21981
rect 10229 22015 10287 22021
rect 10229 21981 10241 22015
rect 10275 21981 10287 22015
rect 10229 21975 10287 21981
rect 10410 21972 10416 22024
rect 10468 21972 10474 22024
rect 6178 21904 6184 21956
rect 6236 21944 6242 21956
rect 11624 21944 11652 22043
rect 12066 22040 12072 22092
rect 12124 22080 12130 22092
rect 12253 22083 12311 22089
rect 12253 22080 12265 22083
rect 12124 22052 12265 22080
rect 12124 22040 12130 22052
rect 12253 22049 12265 22052
rect 12299 22049 12311 22083
rect 12253 22043 12311 22049
rect 15470 22040 15476 22092
rect 15528 22080 15534 22092
rect 16500 22080 16528 22120
rect 16758 22108 16764 22160
rect 16816 22148 16822 22160
rect 17037 22151 17095 22157
rect 17037 22148 17049 22151
rect 16816 22120 17049 22148
rect 16816 22108 16822 22120
rect 17037 22117 17049 22120
rect 17083 22117 17095 22151
rect 17037 22111 17095 22117
rect 19334 22108 19340 22160
rect 19392 22108 19398 22160
rect 22370 22148 22376 22160
rect 22020 22120 22376 22148
rect 15528 22052 16436 22080
rect 16500 22052 17540 22080
rect 15528 22040 15534 22052
rect 16408 22024 16436 22052
rect 12802 21972 12808 22024
rect 12860 21972 12866 22024
rect 13538 21972 13544 22024
rect 13596 22012 13602 22024
rect 14550 22012 14556 22024
rect 13596 21984 14556 22012
rect 13596 21972 13602 21984
rect 14550 21972 14556 21984
rect 14608 22012 14614 22024
rect 14826 22012 14832 22024
rect 14608 21984 14832 22012
rect 14608 21972 14614 21984
rect 14826 21972 14832 21984
rect 14884 21972 14890 22024
rect 15013 22015 15071 22021
rect 15013 21981 15025 22015
rect 15059 21981 15071 22015
rect 15013 21975 15071 21981
rect 6236 21916 10180 21944
rect 11624 21916 12204 21944
rect 6236 21904 6242 21916
rect 3989 21879 4047 21885
rect 3989 21876 4001 21879
rect 3936 21848 4001 21876
rect 3936 21836 3942 21848
rect 3989 21845 4001 21848
rect 4035 21845 4047 21879
rect 3989 21839 4047 21845
rect 4157 21879 4215 21885
rect 4157 21845 4169 21879
rect 4203 21845 4215 21879
rect 4157 21839 4215 21845
rect 4338 21836 4344 21888
rect 4396 21836 4402 21888
rect 7742 21836 7748 21888
rect 7800 21876 7806 21888
rect 8202 21876 8208 21888
rect 7800 21848 8208 21876
rect 7800 21836 7806 21848
rect 8202 21836 8208 21848
rect 8260 21836 8266 21888
rect 8478 21836 8484 21888
rect 8536 21876 8542 21888
rect 9401 21879 9459 21885
rect 9401 21876 9413 21879
rect 8536 21848 9413 21876
rect 8536 21836 8542 21848
rect 9401 21845 9413 21848
rect 9447 21845 9459 21879
rect 9401 21839 9459 21845
rect 9766 21836 9772 21888
rect 9824 21836 9830 21888
rect 9858 21836 9864 21888
rect 9916 21836 9922 21888
rect 10152 21876 10180 21916
rect 12176 21888 12204 21916
rect 12434 21904 12440 21956
rect 12492 21904 12498 21956
rect 15028 21944 15056 21975
rect 15194 21972 15200 22024
rect 15252 22012 15258 22024
rect 15565 22015 15623 22021
rect 15565 22012 15577 22015
rect 15252 21984 15577 22012
rect 15252 21972 15258 21984
rect 15565 21981 15577 21984
rect 15611 21981 15623 22015
rect 15565 21975 15623 21981
rect 15746 21972 15752 22024
rect 15804 21972 15810 22024
rect 15838 21972 15844 22024
rect 15896 21972 15902 22024
rect 16025 22015 16083 22021
rect 16025 21981 16037 22015
rect 16071 21981 16083 22015
rect 16025 21975 16083 21981
rect 15028 21916 15516 21944
rect 15488 21888 15516 21916
rect 16040 21888 16068 21975
rect 16390 21972 16396 22024
rect 16448 21972 16454 22024
rect 16482 21972 16488 22024
rect 16540 22012 16546 22024
rect 16577 22015 16635 22021
rect 16577 22012 16589 22015
rect 16540 21984 16589 22012
rect 16540 21972 16546 21984
rect 16577 21981 16589 21984
rect 16623 21981 16635 22015
rect 16577 21975 16635 21981
rect 16758 21972 16764 22024
rect 16816 21972 16822 22024
rect 16853 22015 16911 22021
rect 16853 21981 16865 22015
rect 16899 22012 16911 22015
rect 16942 22012 16948 22024
rect 16899 21984 16948 22012
rect 16899 21981 16911 21984
rect 16853 21975 16911 21981
rect 16942 21972 16948 21984
rect 17000 21972 17006 22024
rect 17034 21972 17040 22024
rect 17092 21972 17098 22024
rect 17512 22021 17540 22052
rect 17862 22040 17868 22092
rect 17920 22080 17926 22092
rect 22020 22080 22048 22120
rect 22370 22108 22376 22120
rect 22428 22108 22434 22160
rect 22649 22151 22707 22157
rect 22649 22117 22661 22151
rect 22695 22148 22707 22151
rect 23106 22148 23112 22160
rect 22695 22120 23112 22148
rect 22695 22117 22707 22120
rect 22649 22111 22707 22117
rect 23106 22108 23112 22120
rect 23164 22108 23170 22160
rect 25700 22120 26556 22148
rect 17920 22052 22048 22080
rect 23661 22083 23719 22089
rect 17920 22040 17926 22052
rect 23661 22049 23673 22083
rect 23707 22080 23719 22083
rect 24026 22080 24032 22092
rect 23707 22052 24032 22080
rect 23707 22049 23719 22052
rect 23661 22043 23719 22049
rect 24026 22040 24032 22052
rect 24084 22040 24090 22092
rect 25314 22040 25320 22092
rect 25372 22040 25378 22092
rect 17497 22015 17555 22021
rect 17497 21981 17509 22015
rect 17543 21981 17555 22015
rect 17497 21975 17555 21981
rect 18046 21972 18052 22024
rect 18104 22012 18110 22024
rect 19242 22012 19248 22024
rect 18104 21984 19248 22012
rect 18104 21972 18110 21984
rect 19242 21972 19248 21984
rect 19300 22012 19306 22024
rect 19429 22015 19487 22021
rect 19429 22012 19441 22015
rect 19300 21984 19441 22012
rect 19300 21972 19306 21984
rect 19429 21981 19441 21984
rect 19475 21981 19487 22015
rect 19429 21975 19487 21981
rect 19702 21972 19708 22024
rect 19760 21972 19766 22024
rect 19794 21972 19800 22024
rect 19852 22012 19858 22024
rect 19981 22015 20039 22021
rect 19981 22012 19993 22015
rect 19852 21984 19993 22012
rect 19852 21972 19858 21984
rect 19981 21981 19993 21984
rect 20027 21981 20039 22015
rect 19981 21975 20039 21981
rect 20070 21972 20076 22024
rect 20128 21972 20134 22024
rect 22002 21972 22008 22024
rect 22060 22012 22066 22024
rect 22189 22015 22247 22021
rect 22189 22012 22201 22015
rect 22060 21984 22201 22012
rect 22060 21972 22066 21984
rect 22189 21981 22201 21984
rect 22235 21981 22247 22015
rect 22189 21975 22247 21981
rect 22373 22015 22431 22021
rect 22373 21981 22385 22015
rect 22419 22012 22431 22015
rect 22646 22012 22652 22024
rect 22419 21984 22652 22012
rect 22419 21981 22431 21984
rect 22373 21975 22431 21981
rect 16206 21904 16212 21956
rect 16264 21944 16270 21956
rect 16669 21947 16727 21953
rect 16669 21944 16681 21947
rect 16264 21916 16681 21944
rect 16264 21904 16270 21916
rect 16669 21913 16681 21916
rect 16715 21913 16727 21947
rect 16776 21944 16804 21972
rect 22204 21944 22232 21975
rect 22646 21972 22652 21984
rect 22704 21972 22710 22024
rect 22738 21972 22744 22024
rect 22796 22012 22802 22024
rect 22925 22015 22983 22021
rect 22925 22012 22937 22015
rect 22796 21984 22937 22012
rect 22796 21972 22802 21984
rect 22925 21981 22937 21984
rect 22971 21981 22983 22015
rect 23569 22015 23627 22021
rect 23569 22012 23581 22015
rect 22925 21975 22983 21981
rect 23124 21984 23581 22012
rect 23124 21956 23152 21984
rect 23569 21981 23581 21984
rect 23615 21981 23627 22015
rect 23569 21975 23627 21981
rect 23750 21972 23756 22024
rect 23808 22012 23814 22024
rect 23845 22015 23903 22021
rect 23845 22012 23857 22015
rect 23808 21984 23857 22012
rect 23808 21972 23814 21984
rect 23845 21981 23857 21984
rect 23891 21981 23903 22015
rect 23845 21975 23903 21981
rect 24578 21972 24584 22024
rect 24636 22012 24642 22024
rect 24673 22015 24731 22021
rect 24673 22012 24685 22015
rect 24636 21984 24685 22012
rect 24636 21972 24642 21984
rect 24673 21981 24685 21984
rect 24719 21981 24731 22015
rect 24673 21975 24731 21981
rect 24762 21972 24768 22024
rect 24820 22012 24826 22024
rect 24857 22015 24915 22021
rect 24857 22012 24869 22015
rect 24820 21984 24869 22012
rect 24820 21972 24826 21984
rect 24857 21981 24869 21984
rect 24903 21981 24915 22015
rect 24857 21975 24915 21981
rect 24949 22015 25007 22021
rect 24949 21981 24961 22015
rect 24995 21981 25007 22015
rect 24949 21975 25007 21981
rect 25041 22015 25099 22021
rect 25041 21981 25053 22015
rect 25087 22012 25099 22015
rect 25700 22012 25728 22120
rect 25087 21984 25728 22012
rect 25087 21981 25099 21984
rect 25041 21975 25099 21981
rect 23106 21944 23112 21956
rect 16776 21916 16896 21944
rect 22204 21916 23112 21944
rect 16669 21907 16727 21913
rect 11606 21876 11612 21888
rect 10152 21848 11612 21876
rect 11606 21836 11612 21848
rect 11664 21836 11670 21888
rect 11698 21836 11704 21888
rect 11756 21836 11762 21888
rect 11790 21836 11796 21888
rect 11848 21836 11854 21888
rect 12158 21836 12164 21888
rect 12216 21876 12222 21888
rect 12529 21879 12587 21885
rect 12529 21876 12541 21879
rect 12216 21848 12541 21876
rect 12216 21836 12222 21848
rect 12529 21845 12541 21848
rect 12575 21845 12587 21879
rect 12529 21839 12587 21845
rect 12618 21836 12624 21888
rect 12676 21836 12682 21888
rect 15470 21836 15476 21888
rect 15528 21836 15534 21888
rect 16022 21836 16028 21888
rect 16080 21836 16086 21888
rect 16868 21876 16896 21916
rect 23106 21904 23112 21916
rect 23164 21904 23170 21956
rect 23290 21904 23296 21956
rect 23348 21944 23354 21956
rect 24964 21944 24992 21975
rect 23348 21916 24992 21944
rect 23348 21904 23354 21916
rect 22370 21876 22376 21888
rect 16868 21848 22376 21876
rect 22370 21836 22376 21848
rect 22428 21836 22434 21888
rect 24670 21836 24676 21888
rect 24728 21876 24734 21888
rect 25056 21876 25084 21975
rect 25774 21974 25780 22026
rect 25832 21974 25838 22026
rect 26234 22021 26240 22024
rect 26053 22015 26111 22021
rect 26053 22012 26065 22015
rect 25881 21984 26065 22012
rect 25130 21904 25136 21956
rect 25188 21944 25194 21956
rect 25881 21944 25909 21984
rect 26053 21981 26065 21984
rect 26099 21981 26111 22015
rect 26053 21975 26111 21981
rect 26197 22015 26240 22021
rect 26197 21981 26209 22015
rect 26197 21975 26240 21981
rect 26234 21972 26240 21975
rect 26292 21972 26298 22024
rect 26528 22012 26556 22120
rect 28258 22108 28264 22160
rect 28316 22148 28322 22160
rect 30745 22151 30803 22157
rect 30745 22148 30757 22151
rect 28316 22120 28948 22148
rect 28316 22108 28322 22120
rect 26602 22040 26608 22092
rect 26660 22080 26666 22092
rect 27249 22083 27307 22089
rect 27249 22080 27261 22083
rect 26660 22052 27261 22080
rect 26660 22040 26666 22052
rect 27249 22049 27261 22052
rect 27295 22049 27307 22083
rect 27249 22043 27307 22049
rect 27356 22052 28856 22080
rect 27356 22012 27384 22052
rect 28828 22024 28856 22052
rect 26528 21984 27384 22012
rect 27433 22015 27491 22021
rect 27433 21981 27445 22015
rect 27479 21981 27491 22015
rect 27433 21975 27491 21981
rect 25188 21916 25909 21944
rect 25961 21947 26019 21953
rect 25188 21904 25194 21916
rect 25961 21913 25973 21947
rect 26007 21944 26019 21947
rect 26007 21916 26096 21944
rect 26007 21913 26019 21916
rect 25961 21907 26019 21913
rect 26068 21888 26096 21916
rect 26510 21904 26516 21956
rect 26568 21944 26574 21956
rect 27448 21944 27476 21975
rect 27706 21972 27712 22024
rect 27764 21972 27770 22024
rect 27985 22015 28043 22021
rect 27985 21981 27997 22015
rect 28031 21981 28043 22015
rect 27985 21975 28043 21981
rect 27801 21947 27859 21953
rect 27801 21944 27813 21947
rect 26568 21916 27813 21944
rect 26568 21904 26574 21916
rect 27801 21913 27813 21916
rect 27847 21913 27859 21947
rect 27801 21907 27859 21913
rect 24728 21848 25084 21876
rect 24728 21836 24734 21848
rect 26050 21836 26056 21888
rect 26108 21836 26114 21888
rect 26346 21879 26404 21885
rect 26346 21845 26358 21879
rect 26392 21876 26404 21879
rect 27522 21876 27528 21888
rect 26392 21848 27528 21876
rect 26392 21845 26404 21848
rect 26346 21839 26404 21845
rect 27522 21836 27528 21848
rect 27580 21836 27586 21888
rect 27614 21836 27620 21888
rect 27672 21836 27678 21888
rect 27890 21836 27896 21888
rect 27948 21876 27954 21888
rect 28000 21876 28028 21975
rect 28350 21972 28356 22024
rect 28408 21972 28414 22024
rect 28629 22015 28687 22021
rect 28629 21981 28641 22015
rect 28675 21981 28687 22015
rect 28629 21975 28687 21981
rect 28166 21904 28172 21956
rect 28224 21904 28230 21956
rect 28258 21904 28264 21956
rect 28316 21904 28322 21956
rect 28644 21944 28672 21975
rect 28810 21972 28816 22024
rect 28868 21972 28874 22024
rect 28920 22021 28948 22120
rect 30484 22120 30757 22148
rect 29012 22052 29868 22080
rect 29012 22021 29040 22052
rect 29840 22024 29868 22052
rect 30006 22040 30012 22092
rect 30064 22080 30070 22092
rect 30377 22083 30435 22089
rect 30377 22080 30389 22083
rect 30064 22052 30389 22080
rect 30064 22040 30070 22052
rect 30377 22049 30389 22052
rect 30423 22049 30435 22083
rect 30377 22043 30435 22049
rect 28905 22015 28963 22021
rect 28905 21981 28917 22015
rect 28951 21981 28963 22015
rect 28905 21975 28963 21981
rect 28997 22015 29055 22021
rect 28997 21981 29009 22015
rect 29043 21981 29055 22015
rect 28997 21975 29055 21981
rect 29822 21972 29828 22024
rect 29880 21972 29886 22024
rect 30484 21998 30512 22120
rect 30745 22117 30757 22120
rect 30791 22117 30803 22151
rect 32217 22151 32275 22157
rect 32217 22148 32229 22151
rect 30745 22111 30803 22117
rect 31588 22120 32229 22148
rect 30558 22040 30564 22092
rect 30616 22080 30622 22092
rect 31202 22080 31208 22092
rect 30616 22052 31208 22080
rect 30616 22040 30622 22052
rect 31202 22040 31208 22052
rect 31260 22040 31266 22092
rect 31389 22083 31447 22089
rect 31389 22049 31401 22083
rect 31435 22080 31447 22083
rect 31478 22080 31484 22092
rect 31435 22052 31484 22080
rect 31435 22049 31447 22052
rect 31389 22043 31447 22049
rect 31478 22040 31484 22052
rect 31536 22040 31542 22092
rect 31110 21972 31116 22024
rect 31168 22012 31174 22024
rect 31588 22012 31616 22120
rect 32217 22117 32229 22120
rect 32263 22117 32275 22151
rect 32217 22111 32275 22117
rect 32398 22108 32404 22160
rect 32456 22108 32462 22160
rect 32493 22151 32551 22157
rect 32493 22117 32505 22151
rect 32539 22117 32551 22151
rect 32876 22148 32904 22176
rect 32493 22111 32551 22117
rect 32784 22120 33272 22148
rect 31168 21984 31616 22012
rect 31168 21972 31174 21984
rect 31846 21972 31852 22024
rect 31904 21972 31910 22024
rect 31941 22015 31999 22021
rect 31941 21981 31953 22015
rect 31987 22006 31999 22015
rect 32030 22006 32036 22024
rect 31987 21981 32036 22006
rect 31941 21978 32036 21981
rect 31941 21975 31999 21978
rect 32030 21972 32036 21978
rect 32088 21972 32094 22024
rect 32416 22021 32444 22108
rect 32508 22080 32536 22111
rect 32784 22080 32812 22120
rect 32508 22052 32812 22080
rect 32401 22015 32459 22021
rect 32125 21981 32183 21987
rect 28368 21916 28672 21944
rect 29549 21947 29607 21953
rect 28368 21876 28396 21916
rect 29549 21913 29561 21947
rect 29595 21913 29607 21947
rect 32125 21947 32137 21981
rect 32171 21978 32183 21981
rect 32401 21981 32413 22015
rect 32447 21981 32459 22015
rect 32171 21950 32260 21978
rect 32401 21975 32459 21981
rect 32171 21947 32183 21950
rect 32125 21941 32183 21947
rect 32232 21944 32260 21950
rect 32508 21944 32536 22052
rect 32858 22040 32864 22092
rect 32916 22040 32922 22092
rect 33045 22083 33103 22089
rect 33045 22049 33057 22083
rect 33091 22049 33103 22083
rect 33045 22043 33103 22049
rect 32585 22015 32643 22021
rect 32585 21981 32597 22015
rect 32631 21981 32643 22015
rect 32585 21975 32643 21981
rect 32232 21916 32536 21944
rect 29549 21907 29607 21913
rect 27948 21848 28396 21876
rect 27948 21836 27954 21848
rect 28534 21836 28540 21888
rect 28592 21836 28598 21888
rect 29564 21876 29592 21907
rect 29822 21876 29828 21888
rect 29564 21848 29828 21876
rect 29822 21836 29828 21848
rect 29880 21836 29886 21888
rect 32026 21879 32084 21885
rect 32026 21845 32038 21879
rect 32072 21876 32084 21879
rect 32214 21876 32220 21888
rect 32072 21848 32220 21876
rect 32072 21845 32084 21848
rect 32026 21839 32084 21845
rect 32214 21836 32220 21848
rect 32272 21836 32278 21888
rect 32600 21876 32628 21975
rect 32674 21972 32680 22024
rect 32732 21972 32738 22024
rect 33060 21944 33088 22043
rect 33134 22040 33140 22092
rect 33192 22040 33198 22092
rect 33244 22089 33272 22120
rect 33229 22083 33287 22089
rect 33229 22049 33241 22083
rect 33275 22049 33287 22083
rect 33229 22043 33287 22049
rect 35158 22040 35164 22092
rect 35216 22040 35222 22092
rect 35250 22040 35256 22092
rect 35308 22040 35314 22092
rect 35728 22089 35756 22188
rect 36262 22176 36268 22188
rect 36320 22176 36326 22228
rect 35820 22120 36400 22148
rect 35820 22089 35848 22120
rect 35713 22083 35771 22089
rect 35713 22049 35725 22083
rect 35759 22049 35771 22083
rect 35713 22043 35771 22049
rect 35805 22083 35863 22089
rect 35805 22049 35817 22083
rect 35851 22049 35863 22083
rect 35805 22043 35863 22049
rect 35989 22083 36047 22089
rect 35989 22049 36001 22083
rect 36035 22080 36047 22083
rect 36078 22080 36084 22092
rect 36035 22052 36084 22080
rect 36035 22049 36047 22052
rect 35989 22043 36047 22049
rect 36078 22040 36084 22052
rect 36136 22040 36142 22092
rect 33321 22015 33379 22021
rect 33321 21981 33333 22015
rect 33367 22012 33379 22015
rect 33502 22012 33508 22024
rect 33367 21984 33508 22012
rect 33367 21981 33379 21984
rect 33321 21975 33379 21981
rect 33502 21972 33508 21984
rect 33560 21972 33566 22024
rect 34790 21972 34796 22024
rect 34848 22012 34854 22024
rect 35069 22015 35127 22021
rect 35069 22012 35081 22015
rect 34848 21984 35081 22012
rect 34848 21972 34854 21984
rect 35069 21981 35081 21984
rect 35115 21981 35127 22015
rect 35176 22012 35204 22040
rect 35897 22015 35955 22021
rect 35897 22012 35909 22015
rect 35176 21984 35909 22012
rect 35069 21975 35127 21981
rect 35897 21981 35909 21984
rect 35943 21981 35955 22015
rect 35897 21975 35955 21981
rect 34422 21944 34428 21956
rect 33060 21916 34428 21944
rect 34422 21904 34428 21916
rect 34480 21944 34486 21956
rect 35161 21947 35219 21953
rect 35161 21944 35173 21947
rect 34480 21916 35173 21944
rect 34480 21904 34486 21916
rect 35161 21913 35173 21916
rect 35207 21913 35219 21947
rect 35161 21907 35219 21913
rect 33318 21876 33324 21888
rect 32600 21848 33324 21876
rect 33318 21836 33324 21848
rect 33376 21836 33382 21888
rect 34698 21836 34704 21888
rect 34756 21836 34762 21888
rect 35176 21876 35204 21907
rect 36372 21888 36400 22120
rect 36446 22040 36452 22092
rect 36504 22080 36510 22092
rect 37001 22083 37059 22089
rect 37001 22080 37013 22083
rect 36504 22052 37013 22080
rect 36504 22040 36510 22052
rect 37001 22049 37013 22052
rect 37047 22049 37059 22083
rect 37001 22043 37059 22049
rect 36817 22015 36875 22021
rect 36817 21981 36829 22015
rect 36863 22012 36875 22015
rect 36906 22012 36912 22024
rect 36863 21984 36912 22012
rect 36863 21981 36875 21984
rect 36817 21975 36875 21981
rect 36906 21972 36912 21984
rect 36964 21972 36970 22024
rect 35529 21879 35587 21885
rect 35529 21876 35541 21879
rect 35176 21848 35541 21876
rect 35529 21845 35541 21848
rect 35575 21845 35587 21879
rect 35529 21839 35587 21845
rect 36354 21836 36360 21888
rect 36412 21876 36418 21888
rect 36633 21879 36691 21885
rect 36633 21876 36645 21879
rect 36412 21848 36645 21876
rect 36412 21836 36418 21848
rect 36633 21845 36645 21848
rect 36679 21845 36691 21879
rect 36633 21839 36691 21845
rect 1104 21786 38272 21808
rect 1104 21734 4874 21786
rect 4926 21734 4938 21786
rect 4990 21734 5002 21786
rect 5054 21734 5066 21786
rect 5118 21734 5130 21786
rect 5182 21734 35594 21786
rect 35646 21734 35658 21786
rect 35710 21734 35722 21786
rect 35774 21734 35786 21786
rect 35838 21734 35850 21786
rect 35902 21734 38272 21786
rect 1104 21712 38272 21734
rect 1762 21672 1768 21684
rect 1688 21644 1768 21672
rect 1688 21613 1716 21644
rect 1762 21632 1768 21644
rect 1820 21632 1826 21684
rect 1946 21632 1952 21684
rect 2004 21672 2010 21684
rect 3237 21675 3295 21681
rect 3237 21672 3249 21675
rect 2004 21644 3249 21672
rect 2004 21632 2010 21644
rect 3237 21641 3249 21644
rect 3283 21641 3295 21675
rect 3237 21635 3295 21641
rect 4338 21632 4344 21684
rect 4396 21632 4402 21684
rect 4706 21632 4712 21684
rect 4764 21632 4770 21684
rect 8846 21632 8852 21684
rect 8904 21672 8910 21684
rect 9125 21675 9183 21681
rect 9125 21672 9137 21675
rect 8904 21644 9137 21672
rect 8904 21632 8910 21644
rect 9125 21641 9137 21644
rect 9171 21641 9183 21675
rect 9125 21635 9183 21641
rect 9582 21632 9588 21684
rect 9640 21672 9646 21684
rect 9769 21675 9827 21681
rect 9769 21672 9781 21675
rect 9640 21644 9781 21672
rect 9640 21632 9646 21644
rect 9769 21641 9781 21644
rect 9815 21641 9827 21675
rect 9769 21635 9827 21641
rect 11146 21632 11152 21684
rect 11204 21672 11210 21684
rect 11517 21675 11575 21681
rect 11517 21672 11529 21675
rect 11204 21644 11529 21672
rect 11204 21632 11210 21644
rect 11517 21641 11529 21644
rect 11563 21641 11575 21675
rect 11517 21635 11575 21641
rect 14918 21632 14924 21684
rect 14976 21632 14982 21684
rect 15102 21632 15108 21684
rect 15160 21672 15166 21684
rect 16298 21672 16304 21684
rect 15160 21644 16304 21672
rect 15160 21632 15166 21644
rect 16298 21632 16304 21644
rect 16356 21632 16362 21684
rect 17310 21632 17316 21684
rect 17368 21632 17374 21684
rect 17862 21632 17868 21684
rect 17920 21632 17926 21684
rect 17972 21644 20392 21672
rect 1673 21607 1731 21613
rect 1673 21573 1685 21607
rect 1719 21573 1731 21607
rect 1673 21567 1731 21573
rect 2774 21496 2780 21548
rect 2832 21496 2838 21548
rect 3602 21536 3608 21548
rect 3160 21508 3608 21536
rect 1394 21428 1400 21480
rect 1452 21428 1458 21480
rect 3160 21477 3188 21508
rect 3602 21496 3608 21508
rect 3660 21496 3666 21548
rect 4356 21545 4384 21632
rect 4571 21607 4629 21613
rect 4571 21573 4583 21607
rect 4617 21604 4629 21607
rect 4724 21604 4752 21632
rect 4617 21576 4752 21604
rect 4617 21573 4629 21576
rect 4571 21567 4629 21573
rect 5166 21564 5172 21616
rect 5224 21564 5230 21616
rect 7282 21564 7288 21616
rect 7340 21564 7346 21616
rect 17880 21604 17908 21632
rect 8404 21576 17908 21604
rect 3697 21539 3755 21545
rect 3697 21505 3709 21539
rect 3743 21536 3755 21539
rect 4065 21539 4123 21545
rect 4065 21536 4077 21539
rect 3743 21508 4077 21536
rect 3743 21505 3755 21508
rect 3697 21499 3755 21505
rect 4065 21505 4077 21508
rect 4111 21505 4123 21539
rect 4065 21499 4123 21505
rect 4249 21539 4307 21545
rect 4249 21505 4261 21539
rect 4295 21505 4307 21539
rect 4249 21499 4307 21505
rect 4341 21539 4399 21545
rect 4341 21505 4353 21539
rect 4387 21505 4399 21539
rect 4341 21499 4399 21505
rect 4433 21539 4491 21545
rect 4433 21505 4445 21539
rect 4479 21505 4491 21539
rect 4433 21499 4491 21505
rect 4709 21539 4767 21545
rect 4709 21505 4721 21539
rect 4755 21536 4767 21539
rect 4890 21536 4896 21548
rect 4755 21508 4896 21536
rect 4755 21505 4767 21508
rect 4709 21499 4767 21505
rect 3145 21471 3203 21477
rect 3145 21437 3157 21471
rect 3191 21437 3203 21471
rect 3145 21431 3203 21437
rect 3881 21471 3939 21477
rect 3881 21437 3893 21471
rect 3927 21468 3939 21471
rect 3970 21468 3976 21480
rect 3927 21440 3976 21468
rect 3927 21437 3939 21440
rect 3881 21431 3939 21437
rect 3050 21292 3056 21344
rect 3108 21332 3114 21344
rect 3896 21332 3924 21431
rect 3970 21428 3976 21440
rect 4028 21428 4034 21480
rect 4264 21400 4292 21499
rect 4448 21468 4476 21499
rect 4890 21496 4896 21508
rect 4948 21496 4954 21548
rect 4985 21539 5043 21545
rect 4985 21505 4997 21539
rect 5031 21505 5043 21539
rect 4985 21499 5043 21505
rect 4522 21468 4528 21480
rect 4448 21440 4528 21468
rect 4522 21428 4528 21440
rect 4580 21468 4586 21480
rect 5000 21468 5028 21499
rect 5718 21496 5724 21548
rect 5776 21496 5782 21548
rect 5810 21496 5816 21548
rect 5868 21496 5874 21548
rect 5905 21539 5963 21545
rect 5905 21505 5917 21539
rect 5951 21505 5963 21539
rect 5905 21499 5963 21505
rect 6089 21539 6147 21545
rect 6089 21505 6101 21539
rect 6135 21536 6147 21539
rect 6178 21536 6184 21548
rect 6135 21508 6184 21536
rect 6135 21505 6147 21508
rect 6089 21499 6147 21505
rect 5258 21468 5264 21480
rect 4580 21440 4752 21468
rect 5000 21440 5264 21468
rect 4580 21428 4586 21440
rect 4614 21400 4620 21412
rect 4264 21372 4620 21400
rect 4614 21360 4620 21372
rect 4672 21360 4678 21412
rect 4724 21400 4752 21440
rect 5258 21428 5264 21440
rect 5316 21428 5322 21480
rect 5353 21471 5411 21477
rect 5353 21437 5365 21471
rect 5399 21468 5411 21471
rect 5920 21468 5948 21499
rect 6178 21496 6184 21508
rect 6236 21496 6242 21548
rect 8404 21536 8432 21576
rect 8312 21508 8432 21536
rect 9309 21539 9367 21545
rect 5399 21440 5948 21468
rect 6549 21471 6607 21477
rect 5399 21437 5411 21440
rect 5353 21431 5411 21437
rect 6549 21437 6561 21471
rect 6595 21468 6607 21471
rect 6595 21440 6684 21468
rect 6595 21437 6607 21440
rect 6549 21431 6607 21437
rect 4724 21372 5396 21400
rect 5368 21344 5396 21372
rect 6656 21344 6684 21440
rect 6822 21428 6828 21480
rect 6880 21428 6886 21480
rect 8312 21409 8340 21508
rect 9309 21505 9321 21539
rect 9355 21505 9367 21539
rect 9309 21499 9367 21505
rect 9324 21468 9352 21499
rect 9398 21496 9404 21548
rect 9456 21496 9462 21548
rect 9493 21539 9551 21545
rect 9493 21505 9505 21539
rect 9539 21536 9551 21539
rect 9582 21536 9588 21548
rect 9539 21508 9588 21536
rect 9539 21505 9551 21508
rect 9493 21499 9551 21505
rect 9582 21496 9588 21508
rect 9640 21496 9646 21548
rect 9674 21496 9680 21548
rect 9732 21496 9738 21548
rect 9953 21539 10011 21545
rect 9953 21505 9965 21539
rect 9999 21505 10011 21539
rect 9953 21499 10011 21505
rect 9968 21468 9996 21499
rect 10042 21496 10048 21548
rect 10100 21496 10106 21548
rect 10137 21539 10195 21545
rect 10137 21505 10149 21539
rect 10183 21536 10195 21539
rect 10226 21536 10232 21548
rect 10183 21508 10232 21536
rect 10183 21505 10195 21508
rect 10137 21499 10195 21505
rect 10226 21496 10232 21508
rect 10284 21496 10290 21548
rect 10318 21496 10324 21548
rect 10376 21496 10382 21548
rect 11882 21496 11888 21548
rect 11940 21496 11946 21548
rect 13357 21539 13415 21545
rect 13357 21505 13369 21539
rect 13403 21505 13415 21539
rect 13357 21499 13415 21505
rect 15100 21539 15158 21545
rect 15100 21505 15112 21539
rect 15146 21505 15158 21539
rect 15100 21499 15158 21505
rect 15197 21539 15255 21545
rect 15197 21505 15209 21539
rect 15243 21505 15255 21539
rect 15197 21499 15255 21505
rect 9324 21440 9996 21468
rect 9968 21412 9996 21440
rect 11974 21428 11980 21480
rect 12032 21428 12038 21480
rect 12158 21428 12164 21480
rect 12216 21428 12222 21480
rect 12802 21428 12808 21480
rect 12860 21468 12866 21480
rect 13081 21471 13139 21477
rect 13081 21468 13093 21471
rect 12860 21440 13093 21468
rect 12860 21428 12866 21440
rect 13081 21437 13093 21440
rect 13127 21437 13139 21471
rect 13081 21431 13139 21437
rect 13372 21468 13400 21499
rect 13998 21468 14004 21480
rect 13372 21440 14004 21468
rect 8297 21403 8355 21409
rect 8297 21400 8309 21403
rect 7944 21372 8309 21400
rect 7944 21344 7972 21372
rect 8297 21369 8309 21372
rect 8343 21369 8355 21403
rect 8297 21363 8355 21369
rect 9950 21360 9956 21412
rect 10008 21400 10014 21412
rect 13372 21400 13400 21440
rect 13998 21428 14004 21440
rect 14056 21428 14062 21480
rect 14277 21471 14335 21477
rect 14277 21437 14289 21471
rect 14323 21468 14335 21471
rect 14642 21468 14648 21480
rect 14323 21440 14648 21468
rect 14323 21437 14335 21440
rect 14277 21431 14335 21437
rect 10008 21372 13400 21400
rect 13817 21403 13875 21409
rect 10008 21360 10014 21372
rect 13817 21369 13829 21403
rect 13863 21400 13875 21403
rect 13906 21400 13912 21412
rect 13863 21372 13912 21400
rect 13863 21369 13875 21372
rect 13817 21363 13875 21369
rect 13906 21360 13912 21372
rect 13964 21360 13970 21412
rect 3108 21304 3924 21332
rect 3108 21292 3114 21304
rect 5350 21292 5356 21344
rect 5408 21292 5414 21344
rect 5442 21292 5448 21344
rect 5500 21292 5506 21344
rect 6638 21292 6644 21344
rect 6696 21292 6702 21344
rect 7926 21292 7932 21344
rect 7984 21292 7990 21344
rect 8202 21292 8208 21344
rect 8260 21332 8266 21344
rect 10962 21332 10968 21344
rect 8260 21304 10968 21332
rect 8260 21292 8266 21304
rect 10962 21292 10968 21304
rect 11020 21292 11026 21344
rect 11606 21292 11612 21344
rect 11664 21332 11670 21344
rect 14292 21332 14320 21431
rect 14642 21428 14648 21440
rect 14700 21428 14706 21480
rect 11664 21304 14320 21332
rect 15120 21332 15148 21499
rect 15212 21400 15240 21499
rect 15286 21496 15292 21548
rect 15344 21496 15350 21548
rect 15470 21536 15476 21548
rect 15431 21508 15476 21536
rect 15470 21496 15476 21508
rect 15528 21496 15534 21548
rect 15565 21539 15623 21545
rect 15565 21505 15577 21539
rect 15611 21505 15623 21539
rect 15565 21499 15623 21505
rect 15580 21468 15608 21499
rect 15654 21496 15660 21548
rect 15712 21536 15718 21548
rect 16482 21536 16488 21548
rect 15712 21508 16488 21536
rect 15712 21496 15718 21508
rect 16482 21496 16488 21508
rect 16540 21496 16546 21548
rect 17126 21496 17132 21548
rect 17184 21536 17190 21548
rect 17497 21539 17555 21545
rect 17497 21536 17509 21539
rect 17184 21508 17509 21536
rect 17184 21496 17190 21508
rect 17497 21505 17509 21508
rect 17543 21505 17555 21539
rect 17497 21499 17555 21505
rect 17586 21496 17592 21548
rect 17644 21536 17650 21548
rect 17681 21539 17739 21545
rect 17681 21536 17693 21539
rect 17644 21508 17693 21536
rect 17644 21496 17650 21508
rect 17681 21505 17693 21508
rect 17727 21505 17739 21539
rect 17681 21499 17739 21505
rect 17773 21539 17831 21545
rect 17773 21505 17785 21539
rect 17819 21536 17831 21539
rect 17865 21539 17923 21545
rect 17865 21536 17877 21539
rect 17819 21508 17877 21536
rect 17819 21505 17831 21508
rect 17773 21499 17831 21505
rect 17865 21505 17877 21508
rect 17911 21505 17923 21539
rect 17865 21499 17923 21505
rect 16942 21468 16948 21480
rect 15580 21440 16948 21468
rect 16942 21428 16948 21440
rect 17000 21428 17006 21480
rect 17696 21468 17724 21499
rect 17972 21468 18000 21644
rect 18138 21564 18144 21616
rect 18196 21564 18202 21616
rect 18874 21564 18880 21616
rect 18932 21564 18938 21616
rect 19334 21604 19340 21616
rect 19168 21576 19340 21604
rect 18049 21539 18107 21545
rect 18049 21505 18061 21539
rect 18095 21536 18107 21539
rect 18156 21536 18184 21564
rect 19168 21536 19196 21576
rect 19334 21564 19340 21576
rect 19392 21604 19398 21616
rect 19794 21604 19800 21616
rect 19392 21576 19800 21604
rect 19392 21564 19398 21576
rect 19794 21564 19800 21576
rect 19852 21564 19858 21616
rect 20070 21604 20076 21616
rect 19904 21576 20076 21604
rect 18095 21508 19196 21536
rect 18095 21505 18107 21508
rect 18049 21499 18107 21505
rect 19242 21496 19248 21548
rect 19300 21536 19306 21548
rect 19521 21539 19579 21545
rect 19521 21536 19533 21539
rect 19300 21508 19533 21536
rect 19300 21496 19306 21508
rect 19521 21505 19533 21508
rect 19567 21505 19579 21539
rect 19521 21499 19579 21505
rect 17696 21440 18000 21468
rect 18138 21428 18144 21480
rect 18196 21428 18202 21480
rect 18509 21471 18567 21477
rect 18509 21437 18521 21471
rect 18555 21468 18567 21471
rect 18966 21468 18972 21480
rect 18555 21440 18972 21468
rect 18555 21437 18567 21440
rect 18509 21431 18567 21437
rect 18966 21428 18972 21440
rect 19024 21428 19030 21480
rect 19613 21471 19671 21477
rect 19613 21437 19625 21471
rect 19659 21468 19671 21471
rect 19702 21468 19708 21480
rect 19659 21440 19708 21468
rect 19659 21437 19671 21440
rect 19613 21431 19671 21437
rect 19702 21428 19708 21440
rect 19760 21428 19766 21480
rect 19812 21477 19840 21564
rect 19904 21545 19932 21576
rect 20070 21564 20076 21576
rect 20128 21564 20134 21616
rect 20364 21548 20392 21644
rect 22186 21632 22192 21684
rect 22244 21672 22250 21684
rect 22925 21675 22983 21681
rect 22925 21672 22937 21675
rect 22244 21644 22937 21672
rect 22244 21632 22250 21644
rect 22925 21641 22937 21644
rect 22971 21641 22983 21675
rect 25409 21675 25467 21681
rect 22925 21635 22983 21641
rect 23032 21644 23428 21672
rect 19889 21539 19947 21545
rect 19889 21505 19901 21539
rect 19935 21505 19947 21539
rect 19889 21499 19947 21505
rect 19978 21496 19984 21548
rect 20036 21536 20042 21548
rect 20165 21539 20223 21545
rect 20165 21536 20177 21539
rect 20036 21508 20177 21536
rect 20036 21496 20042 21508
rect 20165 21505 20177 21508
rect 20211 21505 20223 21539
rect 20165 21499 20223 21505
rect 20346 21496 20352 21548
rect 20404 21536 20410 21548
rect 20990 21536 20996 21548
rect 20404 21508 20996 21536
rect 20404 21496 20410 21508
rect 20990 21496 20996 21508
rect 21048 21496 21054 21548
rect 22922 21496 22928 21548
rect 22980 21536 22986 21548
rect 23032 21545 23060 21644
rect 23017 21539 23075 21545
rect 23017 21536 23029 21539
rect 22980 21508 23029 21536
rect 22980 21496 22986 21508
rect 23017 21505 23029 21508
rect 23063 21505 23075 21539
rect 23017 21499 23075 21505
rect 23106 21496 23112 21548
rect 23164 21496 23170 21548
rect 23400 21545 23428 21644
rect 25409 21641 25421 21675
rect 25455 21672 25467 21675
rect 25498 21672 25504 21684
rect 25455 21644 25504 21672
rect 25455 21641 25467 21644
rect 25409 21635 25467 21641
rect 25498 21632 25504 21644
rect 25556 21632 25562 21684
rect 25682 21632 25688 21684
rect 25740 21632 25746 21684
rect 25792 21644 27660 21672
rect 23566 21564 23572 21616
rect 23624 21604 23630 21616
rect 24762 21604 24768 21616
rect 23624 21576 24768 21604
rect 23624 21564 23630 21576
rect 24762 21564 24768 21576
rect 24820 21604 24826 21616
rect 25041 21607 25099 21613
rect 24820 21576 24992 21604
rect 24820 21564 24826 21576
rect 23385 21539 23443 21545
rect 23385 21505 23397 21539
rect 23431 21505 23443 21539
rect 23385 21499 23443 21505
rect 24854 21496 24860 21548
rect 24912 21496 24918 21548
rect 24964 21536 24992 21576
rect 25041 21573 25053 21607
rect 25087 21604 25099 21607
rect 25314 21604 25320 21616
rect 25087 21576 25320 21604
rect 25087 21573 25099 21576
rect 25041 21567 25099 21573
rect 25314 21564 25320 21576
rect 25372 21604 25378 21616
rect 25593 21607 25651 21613
rect 25593 21604 25605 21607
rect 25372 21576 25605 21604
rect 25372 21564 25378 21576
rect 25593 21573 25605 21576
rect 25639 21573 25651 21607
rect 25593 21567 25651 21573
rect 25133 21539 25191 21545
rect 25133 21536 25145 21539
rect 24964 21508 25145 21536
rect 25133 21505 25145 21508
rect 25179 21505 25191 21539
rect 25133 21499 25191 21505
rect 25225 21539 25283 21545
rect 25225 21505 25237 21539
rect 25271 21536 25283 21539
rect 25498 21536 25504 21548
rect 25271 21508 25504 21536
rect 25271 21505 25283 21508
rect 25225 21499 25283 21505
rect 25498 21496 25504 21508
rect 25556 21496 25562 21548
rect 25700 21545 25728 21632
rect 25792 21616 25820 21644
rect 25774 21564 25780 21616
rect 25832 21564 25838 21616
rect 27433 21607 27491 21613
rect 27433 21604 27445 21607
rect 26252 21576 27445 21604
rect 25685 21539 25743 21545
rect 25685 21505 25697 21539
rect 25731 21505 25743 21539
rect 25685 21499 25743 21505
rect 19797 21471 19855 21477
rect 19797 21437 19809 21471
rect 19843 21468 19855 21471
rect 20254 21468 20260 21480
rect 19843 21440 20260 21468
rect 19843 21437 19855 21440
rect 19797 21431 19855 21437
rect 20254 21428 20260 21440
rect 20312 21428 20318 21480
rect 22186 21428 22192 21480
rect 22244 21468 22250 21480
rect 22738 21468 22744 21480
rect 22244 21440 22744 21468
rect 22244 21428 22250 21440
rect 22738 21428 22744 21440
rect 22796 21468 22802 21480
rect 23201 21471 23259 21477
rect 23201 21468 23213 21471
rect 22796 21440 23213 21468
rect 22796 21428 22802 21440
rect 23201 21437 23213 21440
rect 23247 21437 23259 21471
rect 26252 21468 26280 21576
rect 27433 21573 27445 21576
rect 27479 21573 27491 21607
rect 27433 21567 27491 21573
rect 27632 21604 27660 21644
rect 28166 21632 28172 21684
rect 28224 21672 28230 21684
rect 32582 21672 32588 21684
rect 28224 21644 32588 21672
rect 28224 21632 28230 21644
rect 32582 21632 32588 21644
rect 32640 21632 32646 21684
rect 34698 21632 34704 21684
rect 34756 21632 34762 21684
rect 35158 21632 35164 21684
rect 35216 21672 35222 21684
rect 35253 21675 35311 21681
rect 35253 21672 35265 21675
rect 35216 21644 35265 21672
rect 35216 21632 35222 21644
rect 35253 21641 35265 21644
rect 35299 21641 35311 21675
rect 35253 21635 35311 21641
rect 35342 21632 35348 21684
rect 35400 21632 35406 21684
rect 35897 21675 35955 21681
rect 35897 21641 35909 21675
rect 35943 21672 35955 21675
rect 36449 21675 36507 21681
rect 36449 21672 36461 21675
rect 35943 21644 36461 21672
rect 35943 21641 35955 21644
rect 35897 21635 35955 21641
rect 36449 21641 36461 21644
rect 36495 21641 36507 21675
rect 36449 21635 36507 21641
rect 28442 21604 28448 21616
rect 27632 21576 28448 21604
rect 23201 21431 23259 21437
rect 23493 21440 26280 21468
rect 27448 21468 27476 21567
rect 27632 21545 27660 21576
rect 28442 21564 28448 21576
rect 28500 21564 28506 21616
rect 29730 21564 29736 21616
rect 29788 21564 29794 21616
rect 29917 21607 29975 21613
rect 29917 21573 29929 21607
rect 29963 21604 29975 21607
rect 30098 21604 30104 21616
rect 29963 21576 30104 21604
rect 29963 21573 29975 21576
rect 29917 21567 29975 21573
rect 30098 21564 30104 21576
rect 30156 21604 30162 21616
rect 30156 21576 30788 21604
rect 30156 21564 30162 21576
rect 27617 21539 27675 21545
rect 27617 21505 27629 21539
rect 27663 21505 27675 21539
rect 27617 21499 27675 21505
rect 27706 21496 27712 21548
rect 27764 21496 27770 21548
rect 30009 21539 30067 21545
rect 30009 21505 30021 21539
rect 30055 21536 30067 21539
rect 30558 21536 30564 21548
rect 30055 21508 30564 21536
rect 30055 21505 30067 21508
rect 30009 21499 30067 21505
rect 30558 21496 30564 21508
rect 30616 21496 30622 21548
rect 30760 21545 30788 21576
rect 33336 21576 33824 21604
rect 33336 21548 33364 21576
rect 30745 21539 30803 21545
rect 30745 21505 30757 21539
rect 30791 21505 30803 21539
rect 30745 21499 30803 21505
rect 30929 21539 30987 21545
rect 30929 21505 30941 21539
rect 30975 21536 30987 21539
rect 31110 21536 31116 21548
rect 30975 21508 31116 21536
rect 30975 21505 30987 21508
rect 30929 21499 30987 21505
rect 31110 21496 31116 21508
rect 31168 21496 31174 21548
rect 32214 21496 32220 21548
rect 32272 21536 32278 21548
rect 32493 21539 32551 21545
rect 32493 21536 32505 21539
rect 32272 21508 32505 21536
rect 32272 21496 32278 21508
rect 32493 21505 32505 21508
rect 32539 21505 32551 21539
rect 32493 21499 32551 21505
rect 32674 21496 32680 21548
rect 32732 21496 32738 21548
rect 33318 21496 33324 21548
rect 33376 21496 33382 21548
rect 33413 21539 33471 21545
rect 33413 21505 33425 21539
rect 33459 21505 33471 21539
rect 33413 21499 33471 21505
rect 33428 21468 33456 21499
rect 33502 21496 33508 21548
rect 33560 21496 33566 21548
rect 33594 21496 33600 21548
rect 33652 21536 33658 21548
rect 33796 21545 33824 21576
rect 33689 21539 33747 21545
rect 33689 21536 33701 21539
rect 33652 21508 33701 21536
rect 33652 21496 33658 21508
rect 33689 21505 33701 21508
rect 33735 21505 33747 21539
rect 33689 21499 33747 21505
rect 33781 21539 33839 21545
rect 33781 21505 33793 21539
rect 33827 21505 33839 21539
rect 33781 21499 33839 21505
rect 33965 21539 34023 21545
rect 33965 21505 33977 21539
rect 34011 21536 34023 21539
rect 34716 21536 34744 21632
rect 35360 21604 35388 21632
rect 35618 21604 35624 21616
rect 35360 21576 35624 21604
rect 34011 21508 34744 21536
rect 35161 21539 35219 21545
rect 34011 21505 34023 21508
rect 33965 21499 34023 21505
rect 35161 21505 35173 21539
rect 35207 21536 35219 21539
rect 35360 21536 35388 21576
rect 35618 21564 35624 21576
rect 35676 21564 35682 21616
rect 35207 21508 35388 21536
rect 35207 21505 35219 21508
rect 35161 21499 35219 21505
rect 33980 21468 34008 21499
rect 35526 21496 35532 21548
rect 35584 21536 35590 21548
rect 35805 21539 35863 21545
rect 35805 21536 35817 21539
rect 35584 21508 35817 21536
rect 35584 21496 35590 21508
rect 35805 21505 35817 21508
rect 35851 21505 35863 21539
rect 35805 21499 35863 21505
rect 36262 21496 36268 21548
rect 36320 21496 36326 21548
rect 36354 21496 36360 21548
rect 36412 21496 36418 21548
rect 36446 21496 36452 21548
rect 36504 21536 36510 21548
rect 36725 21539 36783 21545
rect 36725 21536 36737 21539
rect 36504 21508 36737 21536
rect 36504 21496 36510 21508
rect 36725 21505 36737 21508
rect 36771 21505 36783 21539
rect 36725 21499 36783 21505
rect 27448 21440 33162 21468
rect 33428 21440 34008 21468
rect 15212 21372 16068 21400
rect 16040 21344 16068 21372
rect 16758 21360 16764 21412
rect 16816 21400 16822 21412
rect 23493 21400 23521 21440
rect 16816 21372 23521 21400
rect 23569 21403 23627 21409
rect 16816 21360 16822 21372
rect 23569 21369 23581 21403
rect 23615 21400 23627 21403
rect 27430 21400 27436 21412
rect 23615 21372 27436 21400
rect 23615 21369 23627 21372
rect 23569 21363 23627 21369
rect 27430 21360 27436 21372
rect 27488 21360 27494 21412
rect 28810 21360 28816 21412
rect 28868 21400 28874 21412
rect 33134 21400 33162 21440
rect 35250 21428 35256 21480
rect 35308 21468 35314 21480
rect 35989 21471 36047 21477
rect 35989 21468 36001 21471
rect 35308 21440 36001 21468
rect 35308 21428 35314 21440
rect 35989 21437 36001 21440
rect 36035 21468 36047 21471
rect 36170 21468 36176 21480
rect 36035 21440 36176 21468
rect 36035 21437 36047 21440
rect 35989 21431 36047 21437
rect 36170 21428 36176 21440
rect 36228 21428 36234 21480
rect 37274 21428 37280 21480
rect 37332 21428 37338 21480
rect 37292 21400 37320 21428
rect 28868 21372 31064 21400
rect 33134 21372 37320 21400
rect 28868 21360 28874 21372
rect 15378 21332 15384 21344
rect 15120 21304 15384 21332
rect 11664 21292 11670 21304
rect 15378 21292 15384 21304
rect 15436 21292 15442 21344
rect 15470 21292 15476 21344
rect 15528 21332 15534 21344
rect 15654 21332 15660 21344
rect 15528 21304 15660 21332
rect 15528 21292 15534 21304
rect 15654 21292 15660 21304
rect 15712 21292 15718 21344
rect 16022 21292 16028 21344
rect 16080 21292 16086 21344
rect 16114 21292 16120 21344
rect 16172 21332 16178 21344
rect 19794 21332 19800 21344
rect 16172 21304 19800 21332
rect 16172 21292 16178 21304
rect 19794 21292 19800 21304
rect 19852 21292 19858 21344
rect 20070 21292 20076 21344
rect 20128 21332 20134 21344
rect 20257 21335 20315 21341
rect 20257 21332 20269 21335
rect 20128 21304 20269 21332
rect 20128 21292 20134 21304
rect 20257 21301 20269 21304
rect 20303 21301 20315 21335
rect 20257 21295 20315 21301
rect 23106 21292 23112 21344
rect 23164 21292 23170 21344
rect 24854 21292 24860 21344
rect 24912 21332 24918 21344
rect 25774 21332 25780 21344
rect 24912 21304 25780 21332
rect 24912 21292 24918 21304
rect 25774 21292 25780 21304
rect 25832 21292 25838 21344
rect 27154 21292 27160 21344
rect 27212 21332 27218 21344
rect 27525 21335 27583 21341
rect 27525 21332 27537 21335
rect 27212 21304 27537 21332
rect 27212 21292 27218 21304
rect 27525 21301 27537 21304
rect 27571 21301 27583 21335
rect 27525 21295 27583 21301
rect 29638 21292 29644 21344
rect 29696 21332 29702 21344
rect 29733 21335 29791 21341
rect 29733 21332 29745 21335
rect 29696 21304 29745 21332
rect 29696 21292 29702 21304
rect 29733 21301 29745 21304
rect 29779 21301 29791 21335
rect 29733 21295 29791 21301
rect 30926 21292 30932 21344
rect 30984 21292 30990 21344
rect 31036 21332 31064 21372
rect 33045 21335 33103 21341
rect 33045 21332 33057 21335
rect 31036 21304 33057 21332
rect 33045 21301 33057 21304
rect 33091 21332 33103 21335
rect 33226 21332 33232 21344
rect 33091 21304 33232 21332
rect 33091 21301 33103 21304
rect 33045 21295 33103 21301
rect 33226 21292 33232 21304
rect 33284 21292 33290 21344
rect 33502 21292 33508 21344
rect 33560 21332 33566 21344
rect 33873 21335 33931 21341
rect 33873 21332 33885 21335
rect 33560 21304 33885 21332
rect 33560 21292 33566 21304
rect 33873 21301 33885 21304
rect 33919 21301 33931 21335
rect 33873 21295 33931 21301
rect 35437 21335 35495 21341
rect 35437 21301 35449 21335
rect 35483 21332 35495 21335
rect 35710 21332 35716 21344
rect 35483 21304 35716 21332
rect 35483 21301 35495 21304
rect 35437 21295 35495 21301
rect 35710 21292 35716 21304
rect 35768 21292 35774 21344
rect 1104 21242 38272 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 38272 21242
rect 1104 21168 38272 21190
rect 4341 21131 4399 21137
rect 4341 21097 4353 21131
rect 4387 21128 4399 21131
rect 4614 21128 4620 21140
rect 4387 21100 4620 21128
rect 4387 21097 4399 21100
rect 4341 21091 4399 21097
rect 4614 21088 4620 21100
rect 4672 21088 4678 21140
rect 6822 21088 6828 21140
rect 6880 21128 6886 21140
rect 6917 21131 6975 21137
rect 6917 21128 6929 21131
rect 6880 21100 6929 21128
rect 6880 21088 6886 21100
rect 6917 21097 6929 21100
rect 6963 21097 6975 21131
rect 6917 21091 6975 21097
rect 9493 21131 9551 21137
rect 9493 21097 9505 21131
rect 9539 21128 9551 21131
rect 9766 21128 9772 21140
rect 9539 21100 9772 21128
rect 9539 21097 9551 21100
rect 9493 21091 9551 21097
rect 9766 21088 9772 21100
rect 9824 21088 9830 21140
rect 10134 21088 10140 21140
rect 10192 21088 10198 21140
rect 16758 21128 16764 21140
rect 10980 21100 16764 21128
rect 7193 21063 7251 21069
rect 3712 21032 4200 21060
rect 3712 21004 3740 21032
rect 3694 20952 3700 21004
rect 3752 20952 3758 21004
rect 3786 20952 3792 21004
rect 3844 20992 3850 21004
rect 4172 21001 4200 21032
rect 7193 21029 7205 21063
rect 7239 21029 7251 21063
rect 7193 21023 7251 21029
rect 8588 21032 10180 21060
rect 4065 20995 4123 21001
rect 4065 20992 4077 20995
rect 3844 20964 4077 20992
rect 3844 20952 3850 20964
rect 4065 20961 4077 20964
rect 4111 20961 4123 20995
rect 4065 20955 4123 20961
rect 4157 20995 4215 21001
rect 4157 20961 4169 20995
rect 4203 20961 4215 20995
rect 4157 20955 4215 20961
rect 4890 20952 4896 21004
rect 4948 20992 4954 21004
rect 4948 20964 7052 20992
rect 4948 20952 4954 20964
rect 1765 20927 1823 20933
rect 1765 20893 1777 20927
rect 1811 20924 1823 20927
rect 1854 20924 1860 20936
rect 1811 20896 1860 20924
rect 1811 20893 1823 20896
rect 1765 20887 1823 20893
rect 1854 20884 1860 20896
rect 1912 20884 1918 20936
rect 3602 20884 3608 20936
rect 3660 20924 3666 20936
rect 3881 20927 3939 20933
rect 3881 20924 3893 20927
rect 3660 20896 3893 20924
rect 3660 20884 3666 20896
rect 3881 20893 3893 20896
rect 3927 20893 3939 20927
rect 3881 20887 3939 20893
rect 3896 20856 3924 20887
rect 3970 20884 3976 20936
rect 4028 20884 4034 20936
rect 5445 20927 5503 20933
rect 5445 20924 5457 20927
rect 4264 20896 5457 20924
rect 4264 20856 4292 20896
rect 5445 20893 5457 20896
rect 5491 20893 5503 20927
rect 5445 20887 5503 20893
rect 3896 20828 4292 20856
rect 5258 20816 5264 20868
rect 5316 20816 5322 20868
rect 5626 20816 5632 20868
rect 5684 20816 5690 20868
rect 7024 20856 7052 20964
rect 7101 20927 7159 20933
rect 7101 20893 7113 20927
rect 7147 20924 7159 20927
rect 7208 20924 7236 21023
rect 7742 20952 7748 21004
rect 7800 20952 7806 21004
rect 7147 20896 7236 20924
rect 7561 20927 7619 20933
rect 7147 20893 7159 20896
rect 7101 20887 7159 20893
rect 7561 20893 7573 20927
rect 7607 20924 7619 20927
rect 8588 20924 8616 21032
rect 9324 20964 9996 20992
rect 7607 20896 8616 20924
rect 7607 20893 7619 20896
rect 7561 20887 7619 20893
rect 8662 20884 8668 20936
rect 8720 20924 8726 20936
rect 9324 20933 9352 20964
rect 9968 20936 9996 20964
rect 10152 20936 10180 21032
rect 8941 20927 8999 20933
rect 8941 20924 8953 20927
rect 8720 20896 8953 20924
rect 8720 20884 8726 20896
rect 8941 20893 8953 20896
rect 8987 20893 8999 20927
rect 8941 20887 8999 20893
rect 9309 20927 9367 20933
rect 9309 20893 9321 20927
rect 9355 20893 9367 20927
rect 9309 20887 9367 20893
rect 9582 20884 9588 20936
rect 9640 20884 9646 20936
rect 9861 20927 9919 20933
rect 9861 20924 9873 20927
rect 9692 20896 9873 20924
rect 7653 20859 7711 20865
rect 7653 20856 7665 20859
rect 7024 20828 7665 20856
rect 7653 20825 7665 20828
rect 7699 20856 7711 20859
rect 7926 20856 7932 20868
rect 7699 20828 7932 20856
rect 7699 20825 7711 20828
rect 7653 20819 7711 20825
rect 7926 20816 7932 20828
rect 7984 20816 7990 20868
rect 9125 20859 9183 20865
rect 9125 20825 9137 20859
rect 9171 20825 9183 20859
rect 9125 20819 9183 20825
rect 1486 20748 1492 20800
rect 1544 20748 1550 20800
rect 2866 20748 2872 20800
rect 2924 20788 2930 20800
rect 4062 20788 4068 20800
rect 2924 20760 4068 20788
rect 2924 20748 2930 20760
rect 4062 20748 4068 20760
rect 4120 20788 4126 20800
rect 5276 20788 5304 20816
rect 8202 20788 8208 20800
rect 4120 20760 8208 20788
rect 4120 20748 4126 20760
rect 8202 20748 8208 20760
rect 8260 20748 8266 20800
rect 9140 20788 9168 20819
rect 9214 20816 9220 20868
rect 9272 20816 9278 20868
rect 9490 20816 9496 20868
rect 9548 20856 9554 20868
rect 9692 20856 9720 20896
rect 9861 20893 9873 20896
rect 9907 20893 9919 20927
rect 9861 20887 9919 20893
rect 9950 20884 9956 20936
rect 10008 20884 10014 20936
rect 10134 20884 10140 20936
rect 10192 20884 10198 20936
rect 9548 20828 9720 20856
rect 9769 20859 9827 20865
rect 9548 20816 9554 20828
rect 9769 20825 9781 20859
rect 9815 20825 9827 20859
rect 9769 20819 9827 20825
rect 9674 20788 9680 20800
rect 9140 20760 9680 20788
rect 9674 20748 9680 20760
rect 9732 20788 9738 20800
rect 9784 20788 9812 20819
rect 10042 20816 10048 20868
rect 10100 20856 10106 20868
rect 10226 20856 10232 20868
rect 10100 20828 10232 20856
rect 10100 20816 10106 20828
rect 10226 20816 10232 20828
rect 10284 20816 10290 20868
rect 10060 20788 10088 20816
rect 10980 20800 11008 21100
rect 16758 21088 16764 21100
rect 16816 21088 16822 21140
rect 16945 21131 17003 21137
rect 16945 21097 16957 21131
rect 16991 21128 17003 21131
rect 17034 21128 17040 21140
rect 16991 21100 17040 21128
rect 16991 21097 17003 21100
rect 16945 21091 17003 21097
rect 17034 21088 17040 21100
rect 17092 21088 17098 21140
rect 18322 21128 18328 21140
rect 17512 21100 18328 21128
rect 13998 21020 14004 21072
rect 14056 21060 14062 21072
rect 14458 21060 14464 21072
rect 14056 21032 14464 21060
rect 14056 21020 14062 21032
rect 14458 21020 14464 21032
rect 14516 21060 14522 21072
rect 15473 21063 15531 21069
rect 14516 21032 15332 21060
rect 14516 21020 14522 21032
rect 14366 20952 14372 21004
rect 14424 20952 14430 21004
rect 15102 20992 15108 21004
rect 14476 20964 15108 20992
rect 11514 20884 11520 20936
rect 11572 20924 11578 20936
rect 14476 20924 14504 20964
rect 11572 20896 14504 20924
rect 11572 20884 11578 20896
rect 14550 20884 14556 20936
rect 14608 20884 14614 20936
rect 14734 20884 14740 20936
rect 14792 20884 14798 20936
rect 14844 20933 14872 20964
rect 15102 20952 15108 20964
rect 15160 20952 15166 21004
rect 14829 20927 14887 20933
rect 14829 20893 14841 20927
rect 14875 20893 14887 20927
rect 14829 20887 14887 20893
rect 14918 20884 14924 20936
rect 14976 20884 14982 20936
rect 15304 20933 15332 21032
rect 15473 21029 15485 21063
rect 15519 21060 15531 21063
rect 15562 21060 15568 21072
rect 15519 21032 15568 21060
rect 15519 21029 15531 21032
rect 15473 21023 15531 21029
rect 15562 21020 15568 21032
rect 15620 21020 15626 21072
rect 15746 21020 15752 21072
rect 15804 21060 15810 21072
rect 16301 21063 16359 21069
rect 16301 21060 16313 21063
rect 15804 21032 16313 21060
rect 15804 21020 15810 21032
rect 16301 21029 16313 21032
rect 16347 21029 16359 21063
rect 16301 21023 16359 21029
rect 16666 21020 16672 21072
rect 16724 21060 16730 21072
rect 17512 21060 17540 21100
rect 18322 21088 18328 21100
rect 18380 21088 18386 21140
rect 18414 21088 18420 21140
rect 18472 21088 18478 21140
rect 19978 21128 19984 21140
rect 18524 21100 19984 21128
rect 16724 21032 17540 21060
rect 16724 21020 16730 21032
rect 17862 21020 17868 21072
rect 17920 21060 17926 21072
rect 18524 21060 18552 21100
rect 19978 21088 19984 21100
rect 20036 21128 20042 21140
rect 20530 21128 20536 21140
rect 20036 21100 20536 21128
rect 20036 21088 20042 21100
rect 20530 21088 20536 21100
rect 20588 21128 20594 21140
rect 21082 21128 21088 21140
rect 20588 21100 21088 21128
rect 20588 21088 20594 21100
rect 21082 21088 21088 21100
rect 21140 21088 21146 21140
rect 21177 21131 21235 21137
rect 21177 21097 21189 21131
rect 21223 21128 21235 21131
rect 21910 21128 21916 21140
rect 21223 21100 21916 21128
rect 21223 21097 21235 21100
rect 21177 21091 21235 21097
rect 21910 21088 21916 21100
rect 21968 21088 21974 21140
rect 22002 21088 22008 21140
rect 22060 21088 22066 21140
rect 22830 21088 22836 21140
rect 22888 21088 22894 21140
rect 24946 21088 24952 21140
rect 25004 21128 25010 21140
rect 25041 21131 25099 21137
rect 25041 21128 25053 21131
rect 25004 21100 25053 21128
rect 25004 21088 25010 21100
rect 25041 21097 25053 21100
rect 25087 21097 25099 21131
rect 25041 21091 25099 21097
rect 25314 21088 25320 21140
rect 25372 21088 25378 21140
rect 25682 21088 25688 21140
rect 25740 21088 25746 21140
rect 25866 21088 25872 21140
rect 25924 21128 25930 21140
rect 26510 21128 26516 21140
rect 25924 21100 26516 21128
rect 25924 21088 25930 21100
rect 26510 21088 26516 21100
rect 26568 21088 26574 21140
rect 26789 21131 26847 21137
rect 26789 21097 26801 21131
rect 26835 21128 26847 21131
rect 27338 21128 27344 21140
rect 26835 21100 27344 21128
rect 26835 21097 26847 21100
rect 26789 21091 26847 21097
rect 27338 21088 27344 21100
rect 27396 21088 27402 21140
rect 27522 21088 27528 21140
rect 27580 21088 27586 21140
rect 27614 21088 27620 21140
rect 27672 21088 27678 21140
rect 30561 21131 30619 21137
rect 30561 21097 30573 21131
rect 30607 21128 30619 21131
rect 30926 21128 30932 21140
rect 30607 21100 30932 21128
rect 30607 21097 30619 21100
rect 30561 21091 30619 21097
rect 30926 21088 30932 21100
rect 30984 21088 30990 21140
rect 33594 21088 33600 21140
rect 33652 21128 33658 21140
rect 35250 21128 35256 21140
rect 33652 21100 35256 21128
rect 33652 21088 33658 21100
rect 35250 21088 35256 21100
rect 35308 21088 35314 21140
rect 35618 21088 35624 21140
rect 35676 21088 35682 21140
rect 21818 21060 21824 21072
rect 17920 21032 18552 21060
rect 18616 21032 21824 21060
rect 17920 21020 17926 21032
rect 18616 20992 18644 21032
rect 21818 21020 21824 21032
rect 21876 21020 21882 21072
rect 22370 21060 22376 21072
rect 22204 21032 22376 21060
rect 15396 20964 18644 20992
rect 15197 20927 15255 20933
rect 15197 20893 15209 20927
rect 15243 20893 15255 20927
rect 15197 20887 15255 20893
rect 15294 20927 15352 20933
rect 15294 20893 15306 20927
rect 15340 20893 15352 20927
rect 15294 20887 15352 20893
rect 14182 20816 14188 20868
rect 14240 20856 14246 20868
rect 14936 20856 14964 20884
rect 14240 20828 14964 20856
rect 14240 20816 14246 20828
rect 15102 20816 15108 20868
rect 15160 20816 15166 20868
rect 15212 20856 15240 20887
rect 15396 20856 15424 20964
rect 18690 20952 18696 21004
rect 18748 20992 18754 21004
rect 18969 20995 19027 21001
rect 18969 20992 18981 20995
rect 18748 20964 18981 20992
rect 18748 20952 18754 20964
rect 18969 20961 18981 20964
rect 19015 20961 19027 20995
rect 20257 20995 20315 21001
rect 18969 20955 19027 20961
rect 19444 20964 20208 20992
rect 19444 20936 19472 20964
rect 15562 20884 15568 20936
rect 15620 20924 15626 20936
rect 15930 20924 15936 20936
rect 15620 20896 15936 20924
rect 15620 20884 15626 20896
rect 15930 20884 15936 20896
rect 15988 20884 15994 20936
rect 16114 20884 16120 20936
rect 16172 20884 16178 20936
rect 16209 20927 16267 20933
rect 16209 20893 16221 20927
rect 16255 20893 16267 20927
rect 16209 20887 16267 20893
rect 16393 20927 16451 20933
rect 16393 20893 16405 20927
rect 16439 20893 16451 20927
rect 16393 20887 16451 20893
rect 15212 20828 15424 20856
rect 15746 20816 15752 20868
rect 15804 20816 15810 20868
rect 9732 20760 10088 20788
rect 9732 20748 9738 20760
rect 10962 20748 10968 20800
rect 11020 20748 11026 20800
rect 12158 20748 12164 20800
rect 12216 20788 12222 20800
rect 16132 20788 16160 20884
rect 16224 20800 16252 20887
rect 12216 20760 16160 20788
rect 12216 20748 12222 20760
rect 16206 20748 16212 20800
rect 16264 20748 16270 20800
rect 16298 20748 16304 20800
rect 16356 20788 16362 20800
rect 16408 20788 16436 20887
rect 16942 20884 16948 20936
rect 17000 20884 17006 20936
rect 17126 20933 17132 20936
rect 17124 20924 17132 20933
rect 17087 20896 17132 20924
rect 17124 20887 17132 20896
rect 17126 20884 17132 20887
rect 17184 20884 17190 20936
rect 17497 20927 17555 20933
rect 17497 20893 17509 20927
rect 17543 20924 17555 20927
rect 17954 20924 17960 20936
rect 17543 20896 17960 20924
rect 17543 20893 17555 20896
rect 17497 20887 17555 20893
rect 17954 20884 17960 20896
rect 18012 20924 18018 20936
rect 18542 20927 18600 20933
rect 18542 20924 18554 20927
rect 18012 20896 18554 20924
rect 18012 20884 18018 20896
rect 18542 20893 18554 20896
rect 18588 20893 18600 20927
rect 18542 20887 18600 20893
rect 18782 20884 18788 20936
rect 18840 20924 18846 20936
rect 19061 20927 19119 20933
rect 19061 20924 19073 20927
rect 18840 20896 19073 20924
rect 18840 20884 18846 20896
rect 19061 20893 19073 20896
rect 19107 20893 19119 20927
rect 19061 20887 19119 20893
rect 19337 20927 19395 20933
rect 19337 20893 19349 20927
rect 19383 20893 19395 20927
rect 19337 20887 19395 20893
rect 16960 20856 16988 20884
rect 17221 20859 17279 20865
rect 17221 20856 17233 20859
rect 16960 20828 17233 20856
rect 17221 20825 17233 20828
rect 17267 20825 17279 20859
rect 17221 20819 17279 20825
rect 17313 20859 17371 20865
rect 17313 20825 17325 20859
rect 17359 20856 17371 20859
rect 17402 20856 17408 20868
rect 17359 20828 17408 20856
rect 17359 20825 17371 20828
rect 17313 20819 17371 20825
rect 17034 20788 17040 20800
rect 16356 20760 17040 20788
rect 16356 20748 16362 20760
rect 17034 20748 17040 20760
rect 17092 20748 17098 20800
rect 17236 20788 17264 20819
rect 17402 20816 17408 20828
rect 17460 20856 17466 20868
rect 17460 20828 18552 20856
rect 17460 20816 17466 20828
rect 18524 20800 18552 20828
rect 17862 20788 17868 20800
rect 17236 20760 17868 20788
rect 17862 20748 17868 20760
rect 17920 20748 17926 20800
rect 18506 20748 18512 20800
rect 18564 20788 18570 20800
rect 18601 20791 18659 20797
rect 18601 20788 18613 20791
rect 18564 20760 18613 20788
rect 18564 20748 18570 20760
rect 18601 20757 18613 20760
rect 18647 20788 18659 20791
rect 19352 20788 19380 20887
rect 19426 20884 19432 20936
rect 19484 20884 19490 20936
rect 19518 20884 19524 20936
rect 19576 20884 19582 20936
rect 20180 20933 20208 20964
rect 20257 20961 20269 20995
rect 20303 20992 20315 20995
rect 20898 20992 20904 21004
rect 20303 20964 20904 20992
rect 20303 20961 20315 20964
rect 20257 20955 20315 20961
rect 20898 20952 20904 20964
rect 20956 20992 20962 21004
rect 20956 20964 21036 20992
rect 20956 20952 20962 20964
rect 20165 20927 20223 20933
rect 20165 20893 20177 20927
rect 20211 20893 20223 20927
rect 20165 20887 20223 20893
rect 20346 20884 20352 20936
rect 20404 20884 20410 20936
rect 20530 20884 20536 20936
rect 20588 20884 20594 20936
rect 21008 20933 21036 20964
rect 21174 20952 21180 21004
rect 21232 20992 21238 21004
rect 21232 20964 21772 20992
rect 21232 20952 21238 20964
rect 20681 20927 20739 20933
rect 20681 20893 20693 20927
rect 20727 20924 20739 20927
rect 20998 20927 21056 20933
rect 20727 20893 20760 20924
rect 20681 20887 20760 20893
rect 20998 20893 21010 20927
rect 21044 20893 21056 20927
rect 20998 20887 21056 20893
rect 20364 20856 20392 20884
rect 20732 20856 20760 20887
rect 21358 20884 21364 20936
rect 21416 20884 21422 20936
rect 21450 20884 21456 20936
rect 21508 20884 21514 20936
rect 21744 20933 21772 20964
rect 22204 20936 22232 21032
rect 22370 21020 22376 21032
rect 22428 21060 22434 21072
rect 24578 21060 24584 21072
rect 22428 21032 24584 21060
rect 22428 21020 22434 21032
rect 24578 21020 24584 21032
rect 24636 21020 24642 21072
rect 22646 20992 22652 21004
rect 22480 20964 22652 20992
rect 21729 20927 21787 20933
rect 21729 20893 21741 20927
rect 21775 20893 21787 20927
rect 21729 20887 21787 20893
rect 21826 20927 21884 20933
rect 21826 20893 21838 20927
rect 21872 20893 21884 20927
rect 21826 20887 21884 20893
rect 20364 20828 20760 20856
rect 20806 20816 20812 20868
rect 20864 20816 20870 20868
rect 20901 20859 20959 20865
rect 20901 20825 20913 20859
rect 20947 20856 20959 20859
rect 21082 20856 21088 20868
rect 20947 20828 21088 20856
rect 20947 20825 20959 20828
rect 20901 20819 20959 20825
rect 21082 20816 21088 20828
rect 21140 20816 21146 20868
rect 21266 20816 21272 20868
rect 21324 20856 21330 20868
rect 21637 20859 21695 20865
rect 21637 20856 21649 20859
rect 21324 20828 21649 20856
rect 21324 20816 21330 20828
rect 21637 20825 21649 20828
rect 21683 20825 21695 20859
rect 21637 20819 21695 20825
rect 18647 20760 19380 20788
rect 19429 20791 19487 20797
rect 18647 20757 18659 20760
rect 18601 20751 18659 20757
rect 19429 20757 19441 20791
rect 19475 20788 19487 20791
rect 20346 20788 20352 20800
rect 19475 20760 20352 20788
rect 19475 20757 19487 20760
rect 19429 20751 19487 20757
rect 20346 20748 20352 20760
rect 20404 20788 20410 20800
rect 21841 20788 21869 20887
rect 22186 20884 22192 20936
rect 22244 20884 22250 20936
rect 22370 20884 22376 20936
rect 22428 20884 22434 20936
rect 22480 20933 22508 20964
rect 22646 20952 22652 20964
rect 22704 20992 22710 21004
rect 23290 20992 23296 21004
rect 22704 20964 23296 20992
rect 22704 20952 22710 20964
rect 23290 20952 23296 20964
rect 23348 20952 23354 21004
rect 24670 20952 24676 21004
rect 24728 20992 24734 21004
rect 25133 20995 25191 21001
rect 25133 20992 25145 20995
rect 24728 20964 25145 20992
rect 24728 20952 24734 20964
rect 25133 20961 25145 20964
rect 25179 20961 25191 20995
rect 25133 20955 25191 20961
rect 22465 20927 22523 20933
rect 22465 20893 22477 20927
rect 22511 20893 22523 20927
rect 22465 20887 22523 20893
rect 22557 20927 22615 20933
rect 22557 20893 22569 20927
rect 22603 20924 22615 20927
rect 24394 20924 24400 20936
rect 22603 20896 24400 20924
rect 22603 20893 22615 20896
rect 22557 20887 22615 20893
rect 24394 20884 24400 20896
rect 24452 20884 24458 20936
rect 24854 20884 24860 20936
rect 24912 20924 24918 20936
rect 25332 20933 25360 21088
rect 25700 21060 25728 21088
rect 27246 21060 27252 21072
rect 25700 21032 27252 21060
rect 27246 21020 27252 21032
rect 27304 21020 27310 21072
rect 26694 20952 26700 21004
rect 26752 20992 26758 21004
rect 27540 20992 27568 21088
rect 27632 21060 27660 21088
rect 27632 21032 34836 21060
rect 30466 20992 30472 21004
rect 26752 20964 27108 20992
rect 27540 20964 30472 20992
rect 26752 20952 26758 20964
rect 27080 20936 27108 20964
rect 30466 20952 30472 20964
rect 30524 20952 30530 21004
rect 30650 20952 30656 21004
rect 30708 20952 30714 21004
rect 25041 20927 25099 20933
rect 25041 20924 25053 20927
rect 24912 20896 25053 20924
rect 24912 20884 24918 20896
rect 25041 20893 25053 20896
rect 25087 20893 25099 20927
rect 25041 20887 25099 20893
rect 25317 20927 25375 20933
rect 25317 20893 25329 20927
rect 25363 20893 25375 20927
rect 25317 20887 25375 20893
rect 21910 20816 21916 20868
rect 21968 20816 21974 20868
rect 20404 20760 21869 20788
rect 21928 20788 21956 20816
rect 23106 20788 23112 20800
rect 21928 20760 23112 20788
rect 20404 20748 20410 20760
rect 23106 20748 23112 20760
rect 23164 20748 23170 20800
rect 24854 20748 24860 20800
rect 24912 20748 24918 20800
rect 25056 20788 25084 20887
rect 26878 20884 26884 20936
rect 26936 20924 26942 20936
rect 26973 20927 27031 20933
rect 26973 20924 26985 20927
rect 26936 20896 26985 20924
rect 26936 20884 26942 20896
rect 26973 20893 26985 20896
rect 27019 20893 27031 20927
rect 26973 20887 27031 20893
rect 27062 20884 27068 20936
rect 27120 20884 27126 20936
rect 27338 20884 27344 20936
rect 27396 20926 27402 20936
rect 27396 20924 27476 20926
rect 27522 20924 27528 20936
rect 27396 20898 27528 20924
rect 27396 20884 27402 20898
rect 27448 20896 27528 20898
rect 27522 20884 27528 20896
rect 27580 20884 27586 20936
rect 27617 20927 27675 20933
rect 27617 20893 27629 20927
rect 27663 20893 27675 20927
rect 27617 20887 27675 20893
rect 27801 20927 27859 20933
rect 27801 20893 27813 20927
rect 27847 20924 27859 20927
rect 29362 20924 29368 20936
rect 27847 20896 29368 20924
rect 27847 20893 27859 20896
rect 27801 20887 27859 20893
rect 27157 20859 27215 20865
rect 27157 20825 27169 20859
rect 27203 20856 27215 20859
rect 27433 20859 27491 20865
rect 27433 20856 27445 20859
rect 27203 20828 27445 20856
rect 27203 20825 27215 20828
rect 27157 20819 27215 20825
rect 27433 20825 27445 20828
rect 27479 20825 27491 20859
rect 27632 20856 27660 20887
rect 29362 20884 29368 20896
rect 29420 20884 29426 20936
rect 30374 20884 30380 20936
rect 30432 20884 30438 20936
rect 29822 20856 29828 20868
rect 27632 20828 29828 20856
rect 27433 20819 27491 20825
rect 27172 20788 27200 20819
rect 29822 20816 29828 20828
rect 29880 20856 29886 20868
rect 32398 20856 32404 20868
rect 29880 20828 32404 20856
rect 29880 20816 29886 20828
rect 32398 20816 32404 20828
rect 32456 20816 32462 20868
rect 34514 20816 34520 20868
rect 34572 20856 34578 20868
rect 34701 20859 34759 20865
rect 34701 20856 34713 20859
rect 34572 20828 34713 20856
rect 34572 20816 34578 20828
rect 34701 20825 34713 20828
rect 34747 20825 34759 20859
rect 34701 20819 34759 20825
rect 25056 20760 27200 20788
rect 27246 20748 27252 20800
rect 27304 20788 27310 20800
rect 30098 20788 30104 20800
rect 27304 20760 30104 20788
rect 27304 20748 27310 20760
rect 30098 20748 30104 20760
rect 30156 20748 30162 20800
rect 30193 20791 30251 20797
rect 30193 20757 30205 20791
rect 30239 20788 30251 20791
rect 30282 20788 30288 20800
rect 30239 20760 30288 20788
rect 30239 20757 30251 20760
rect 30193 20751 30251 20757
rect 30282 20748 30288 20760
rect 30340 20748 30346 20800
rect 34808 20788 34836 21032
rect 35636 20992 35664 21088
rect 35710 21020 35716 21072
rect 35768 21020 35774 21072
rect 34991 20964 35664 20992
rect 34991 20933 35019 20964
rect 34976 20927 35034 20933
rect 34976 20893 34988 20927
rect 35022 20893 35034 20927
rect 34976 20887 35034 20893
rect 35066 20884 35072 20936
rect 35124 20884 35130 20936
rect 35161 20927 35219 20933
rect 35161 20893 35173 20927
rect 35207 20893 35219 20927
rect 35161 20887 35219 20893
rect 35176 20856 35204 20887
rect 35250 20884 35256 20936
rect 35308 20924 35314 20936
rect 35452 20933 35480 20964
rect 35345 20927 35403 20933
rect 35345 20924 35357 20927
rect 35308 20896 35357 20924
rect 35308 20884 35314 20896
rect 35345 20893 35357 20896
rect 35391 20893 35403 20927
rect 35345 20887 35403 20893
rect 35437 20927 35495 20933
rect 35437 20893 35449 20927
rect 35483 20893 35495 20927
rect 35437 20887 35495 20893
rect 35621 20927 35679 20933
rect 35621 20893 35633 20927
rect 35667 20924 35679 20927
rect 35728 20924 35756 21020
rect 35667 20896 35756 20924
rect 37185 20927 37243 20933
rect 35667 20893 35679 20896
rect 35621 20887 35679 20893
rect 37185 20893 37197 20927
rect 37231 20893 37243 20927
rect 37185 20887 37243 20893
rect 35529 20859 35587 20865
rect 35529 20856 35541 20859
rect 35176 20828 35541 20856
rect 35529 20825 35541 20828
rect 35575 20825 35587 20859
rect 35529 20819 35587 20825
rect 37200 20788 37228 20887
rect 37553 20859 37611 20865
rect 37553 20856 37565 20859
rect 37384 20828 37565 20856
rect 37384 20797 37412 20828
rect 37553 20825 37565 20828
rect 37599 20825 37611 20859
rect 37553 20819 37611 20825
rect 34808 20760 37228 20788
rect 37369 20791 37427 20797
rect 37369 20757 37381 20791
rect 37415 20757 37427 20791
rect 37369 20751 37427 20757
rect 37829 20791 37887 20797
rect 37829 20757 37841 20791
rect 37875 20788 37887 20791
rect 37875 20760 38424 20788
rect 37875 20757 37887 20760
rect 37829 20751 37887 20757
rect 38396 20732 38424 20760
rect 1104 20698 38272 20720
rect 1104 20646 4874 20698
rect 4926 20646 4938 20698
rect 4990 20646 5002 20698
rect 5054 20646 5066 20698
rect 5118 20646 5130 20698
rect 5182 20646 35594 20698
rect 35646 20646 35658 20698
rect 35710 20646 35722 20698
rect 35774 20646 35786 20698
rect 35838 20646 35850 20698
rect 35902 20646 38272 20698
rect 38378 20680 38384 20732
rect 38436 20680 38442 20732
rect 1104 20624 38272 20646
rect 3697 20587 3755 20593
rect 3697 20553 3709 20587
rect 3743 20584 3755 20587
rect 3878 20584 3884 20596
rect 3743 20556 3884 20584
rect 3743 20553 3755 20556
rect 3697 20547 3755 20553
rect 2777 20451 2835 20457
rect 2777 20417 2789 20451
rect 2823 20448 2835 20451
rect 3142 20448 3148 20460
rect 2823 20420 3148 20448
rect 2823 20417 2835 20420
rect 2777 20411 2835 20417
rect 3142 20408 3148 20420
rect 3200 20448 3206 20460
rect 3513 20451 3571 20457
rect 3200 20420 3372 20448
rect 3200 20408 3206 20420
rect 2866 20340 2872 20392
rect 2924 20340 2930 20392
rect 3050 20340 3056 20392
rect 3108 20340 3114 20392
rect 3344 20389 3372 20420
rect 3513 20417 3525 20451
rect 3559 20448 3571 20451
rect 3602 20448 3608 20460
rect 3559 20420 3608 20448
rect 3559 20417 3571 20420
rect 3513 20411 3571 20417
rect 3602 20408 3608 20420
rect 3660 20408 3666 20460
rect 3804 20457 3832 20556
rect 3878 20544 3884 20556
rect 3936 20544 3942 20596
rect 10410 20544 10416 20596
rect 10468 20584 10474 20596
rect 13630 20584 13636 20596
rect 10468 20556 13636 20584
rect 10468 20544 10474 20556
rect 13630 20544 13636 20556
rect 13688 20544 13694 20596
rect 14274 20544 14280 20596
rect 14332 20544 14338 20596
rect 14550 20544 14556 20596
rect 14608 20544 14614 20596
rect 14829 20587 14887 20593
rect 14829 20553 14841 20587
rect 14875 20584 14887 20587
rect 15194 20584 15200 20596
rect 14875 20556 15200 20584
rect 14875 20553 14887 20556
rect 14829 20547 14887 20553
rect 15194 20544 15200 20556
rect 15252 20544 15258 20596
rect 15841 20587 15899 20593
rect 15841 20553 15853 20587
rect 15887 20584 15899 20587
rect 20165 20587 20223 20593
rect 15887 20556 16068 20584
rect 15887 20553 15899 20556
rect 15841 20547 15899 20553
rect 7561 20519 7619 20525
rect 7561 20485 7573 20519
rect 7607 20516 7619 20519
rect 13170 20516 13176 20528
rect 7607 20488 13176 20516
rect 7607 20485 7619 20488
rect 7561 20479 7619 20485
rect 13170 20476 13176 20488
rect 13228 20476 13234 20528
rect 3789 20451 3847 20457
rect 3789 20417 3801 20451
rect 3835 20417 3847 20451
rect 3789 20411 3847 20417
rect 3970 20408 3976 20460
rect 4028 20408 4034 20460
rect 6546 20408 6552 20460
rect 6604 20448 6610 20460
rect 7653 20451 7711 20457
rect 7653 20448 7665 20451
rect 6604 20420 7665 20448
rect 6604 20408 6610 20420
rect 7653 20417 7665 20420
rect 7699 20448 7711 20451
rect 11701 20451 11759 20457
rect 7699 20420 8432 20448
rect 7699 20417 7711 20420
rect 7653 20411 7711 20417
rect 3329 20383 3387 20389
rect 3329 20349 3341 20383
rect 3375 20380 3387 20383
rect 3988 20380 4016 20408
rect 8404 20392 8432 20420
rect 11701 20417 11713 20451
rect 11747 20448 11759 20451
rect 11974 20448 11980 20460
rect 11747 20420 11980 20448
rect 11747 20417 11759 20420
rect 11701 20411 11759 20417
rect 11974 20408 11980 20420
rect 12032 20448 12038 20460
rect 14292 20448 14320 20544
rect 12032 20420 14320 20448
rect 12032 20408 12038 20420
rect 14366 20408 14372 20460
rect 14424 20448 14430 20460
rect 14568 20448 14596 20544
rect 16040 20528 16068 20556
rect 17880 20556 20116 20584
rect 14642 20476 14648 20528
rect 14700 20476 14706 20528
rect 16022 20476 16028 20528
rect 16080 20476 16086 20528
rect 15764 20448 15884 20452
rect 15933 20451 15991 20457
rect 15933 20448 15945 20451
rect 14424 20424 15945 20448
rect 14424 20420 15792 20424
rect 15856 20420 15945 20424
rect 14424 20408 14430 20420
rect 15933 20417 15945 20420
rect 15979 20417 15991 20451
rect 15933 20411 15991 20417
rect 16574 20408 16580 20460
rect 16632 20448 16638 20460
rect 17310 20448 17316 20460
rect 16632 20420 17316 20448
rect 16632 20408 16638 20420
rect 17310 20408 17316 20420
rect 17368 20448 17374 20460
rect 17880 20448 17908 20556
rect 18322 20476 18328 20528
rect 18380 20516 18386 20528
rect 19797 20519 19855 20525
rect 19797 20516 19809 20519
rect 18380 20488 19809 20516
rect 18380 20476 18386 20488
rect 19797 20485 19809 20488
rect 19843 20485 19855 20519
rect 20088 20516 20116 20556
rect 20165 20553 20177 20587
rect 20211 20584 20223 20587
rect 21082 20584 21088 20596
rect 20211 20556 21088 20584
rect 20211 20553 20223 20556
rect 20165 20547 20223 20553
rect 21082 20544 21088 20556
rect 21140 20544 21146 20596
rect 21269 20587 21327 20593
rect 21269 20553 21281 20587
rect 21315 20584 21327 20587
rect 22922 20584 22928 20596
rect 21315 20556 22928 20584
rect 21315 20553 21327 20556
rect 21269 20547 21327 20553
rect 22922 20544 22928 20556
rect 22980 20544 22986 20596
rect 24394 20544 24400 20596
rect 24452 20584 24458 20596
rect 27801 20587 27859 20593
rect 24452 20556 26004 20584
rect 24452 20544 24458 20556
rect 20533 20519 20591 20525
rect 20088 20488 20484 20516
rect 19797 20479 19855 20485
rect 18049 20451 18107 20457
rect 18049 20448 18061 20451
rect 17368 20420 17632 20448
rect 17880 20420 18061 20448
rect 17368 20408 17374 20420
rect 3375 20352 4016 20380
rect 3375 20349 3387 20352
rect 3329 20343 3387 20349
rect 7742 20340 7748 20392
rect 7800 20340 7806 20392
rect 8386 20340 8392 20392
rect 8444 20340 8450 20392
rect 11606 20340 11612 20392
rect 11664 20340 11670 20392
rect 14277 20383 14335 20389
rect 14277 20349 14289 20383
rect 14323 20380 14335 20383
rect 14826 20380 14832 20392
rect 14323 20352 14832 20380
rect 14323 20349 14335 20352
rect 14277 20343 14335 20349
rect 14826 20340 14832 20352
rect 14884 20340 14890 20392
rect 15470 20340 15476 20392
rect 15528 20340 15534 20392
rect 16298 20340 16304 20392
rect 16356 20340 16362 20392
rect 17604 20389 17632 20420
rect 18049 20417 18061 20420
rect 18095 20417 18107 20451
rect 18049 20411 18107 20417
rect 17589 20383 17647 20389
rect 17589 20349 17601 20383
rect 17635 20349 17647 20383
rect 17589 20343 17647 20349
rect 3786 20272 3792 20324
rect 3844 20312 3850 20324
rect 3844 20284 7328 20312
rect 3844 20272 3850 20284
rect 2406 20204 2412 20256
rect 2464 20204 2470 20256
rect 3881 20247 3939 20253
rect 3881 20213 3893 20247
rect 3927 20244 3939 20247
rect 3970 20244 3976 20256
rect 3927 20216 3976 20244
rect 3927 20213 3939 20216
rect 3881 20207 3939 20213
rect 3970 20204 3976 20216
rect 4028 20204 4034 20256
rect 5074 20204 5080 20256
rect 5132 20244 5138 20256
rect 6362 20244 6368 20256
rect 5132 20216 6368 20244
rect 5132 20204 5138 20216
rect 6362 20204 6368 20216
rect 6420 20204 6426 20256
rect 7190 20204 7196 20256
rect 7248 20204 7254 20256
rect 7300 20244 7328 20284
rect 10042 20272 10048 20324
rect 10100 20312 10106 20324
rect 13906 20312 13912 20324
rect 10100 20284 13912 20312
rect 10100 20272 10106 20284
rect 13906 20272 13912 20284
rect 13964 20272 13970 20324
rect 15657 20315 15715 20321
rect 15657 20281 15669 20315
rect 15703 20312 15715 20315
rect 16316 20312 16344 20340
rect 15703 20284 16344 20312
rect 15703 20281 15715 20284
rect 15657 20275 15715 20281
rect 18064 20256 18092 20411
rect 18138 20408 18144 20460
rect 18196 20408 18202 20460
rect 18506 20408 18512 20460
rect 18564 20408 18570 20460
rect 19245 20451 19303 20457
rect 19245 20417 19257 20451
rect 19291 20448 19303 20451
rect 19334 20448 19340 20460
rect 19291 20420 19340 20448
rect 19291 20417 19303 20420
rect 19245 20411 19303 20417
rect 19334 20408 19340 20420
rect 19392 20408 19398 20460
rect 19981 20451 20039 20457
rect 19981 20417 19993 20451
rect 20027 20448 20039 20451
rect 20070 20448 20076 20460
rect 20027 20420 20076 20448
rect 20027 20417 20039 20420
rect 19981 20411 20039 20417
rect 20070 20408 20076 20420
rect 20128 20408 20134 20460
rect 20346 20408 20352 20460
rect 20404 20408 20410 20460
rect 18156 20312 18184 20408
rect 18598 20340 18604 20392
rect 18656 20380 18662 20392
rect 18782 20380 18788 20392
rect 18656 20352 18788 20380
rect 18656 20340 18662 20352
rect 18782 20340 18788 20352
rect 18840 20340 18846 20392
rect 19153 20383 19211 20389
rect 19153 20349 19165 20383
rect 19199 20349 19211 20383
rect 20456 20380 20484 20488
rect 20533 20485 20545 20519
rect 20579 20516 20591 20519
rect 24486 20516 24492 20528
rect 20579 20488 21128 20516
rect 20579 20485 20591 20488
rect 20533 20479 20591 20485
rect 20622 20408 20628 20460
rect 20680 20408 20686 20460
rect 20718 20451 20776 20457
rect 20718 20417 20730 20451
rect 20764 20417 20776 20451
rect 20718 20411 20776 20417
rect 20732 20380 20760 20411
rect 20898 20408 20904 20460
rect 20956 20408 20962 20460
rect 20990 20408 20996 20460
rect 21048 20408 21054 20460
rect 21100 20457 21128 20488
rect 23768 20488 24492 20516
rect 23768 20460 23796 20488
rect 24486 20476 24492 20488
rect 24544 20516 24550 20528
rect 25866 20516 25872 20528
rect 24544 20488 24624 20516
rect 24544 20476 24550 20488
rect 21090 20451 21148 20457
rect 21090 20417 21102 20451
rect 21136 20417 21148 20451
rect 21090 20411 21148 20417
rect 23750 20408 23756 20460
rect 23808 20408 23814 20460
rect 24305 20451 24363 20457
rect 24305 20417 24317 20451
rect 24351 20417 24363 20451
rect 24305 20411 24363 20417
rect 20456 20352 20760 20380
rect 20916 20380 20944 20408
rect 21266 20380 21272 20392
rect 20916 20352 21272 20380
rect 19153 20343 19211 20349
rect 18414 20312 18420 20324
rect 18156 20284 18420 20312
rect 18414 20272 18420 20284
rect 18472 20312 18478 20324
rect 19168 20312 19196 20343
rect 21266 20340 21272 20352
rect 21324 20340 21330 20392
rect 24320 20380 24348 20411
rect 24394 20408 24400 20460
rect 24452 20408 24458 20460
rect 24596 20457 24624 20488
rect 25148 20488 25872 20516
rect 24581 20451 24639 20457
rect 24581 20417 24593 20451
rect 24627 20417 24639 20451
rect 24581 20411 24639 20417
rect 24854 20408 24860 20460
rect 24912 20408 24918 20460
rect 25148 20457 25176 20488
rect 25866 20476 25872 20488
rect 25924 20476 25930 20528
rect 25976 20516 26004 20556
rect 27801 20553 27813 20587
rect 27847 20584 27859 20587
rect 27982 20584 27988 20596
rect 27847 20556 27988 20584
rect 27847 20553 27859 20556
rect 27801 20547 27859 20553
rect 27982 20544 27988 20556
rect 28040 20544 28046 20596
rect 35434 20544 35440 20596
rect 35492 20544 35498 20596
rect 25976 20488 26280 20516
rect 25133 20451 25191 20457
rect 25133 20417 25145 20451
rect 25179 20417 25191 20451
rect 25133 20411 25191 20417
rect 25222 20408 25228 20460
rect 25280 20408 25286 20460
rect 25314 20408 25320 20460
rect 25372 20448 25378 20460
rect 25777 20451 25835 20457
rect 25777 20448 25789 20451
rect 25372 20420 25789 20448
rect 25372 20408 25378 20420
rect 25777 20417 25789 20420
rect 25823 20417 25835 20451
rect 25777 20411 25835 20417
rect 25958 20408 25964 20460
rect 26016 20408 26022 20460
rect 26053 20451 26111 20457
rect 26053 20417 26065 20451
rect 26099 20417 26111 20451
rect 26053 20411 26111 20417
rect 24489 20383 24547 20389
rect 24320 20352 24440 20380
rect 18472 20284 19196 20312
rect 18472 20272 18478 20284
rect 19610 20272 19616 20324
rect 19668 20312 19674 20324
rect 21450 20312 21456 20324
rect 19668 20284 21456 20312
rect 19668 20272 19674 20284
rect 21450 20272 21456 20284
rect 21508 20272 21514 20324
rect 24412 20312 24440 20352
rect 24489 20349 24501 20383
rect 24535 20380 24547 20383
rect 24872 20380 24900 20408
rect 24535 20352 24900 20380
rect 24535 20349 24547 20352
rect 24489 20343 24547 20349
rect 24670 20312 24676 20324
rect 24412 20284 24676 20312
rect 24670 20272 24676 20284
rect 24728 20312 24734 20324
rect 24728 20284 25084 20312
rect 24728 20272 24734 20284
rect 11422 20244 11428 20256
rect 7300 20216 11428 20244
rect 11422 20204 11428 20216
rect 11480 20204 11486 20256
rect 11882 20204 11888 20256
rect 11940 20244 11946 20256
rect 11977 20247 12035 20253
rect 11977 20244 11989 20247
rect 11940 20216 11989 20244
rect 11940 20204 11946 20216
rect 11977 20213 11989 20216
rect 12023 20213 12035 20247
rect 11977 20207 12035 20213
rect 12158 20204 12164 20256
rect 12216 20244 12222 20256
rect 14274 20244 14280 20256
rect 12216 20216 14280 20244
rect 12216 20204 12222 20216
rect 14274 20204 14280 20216
rect 14332 20204 14338 20256
rect 14645 20247 14703 20253
rect 14645 20213 14657 20247
rect 14691 20244 14703 20247
rect 16298 20244 16304 20256
rect 14691 20216 16304 20244
rect 14691 20213 14703 20216
rect 14645 20207 14703 20213
rect 16298 20204 16304 20216
rect 16356 20204 16362 20256
rect 18046 20204 18052 20256
rect 18104 20204 18110 20256
rect 19426 20204 19432 20256
rect 19484 20204 19490 20256
rect 19518 20204 19524 20256
rect 19576 20244 19582 20256
rect 19705 20247 19763 20253
rect 19705 20244 19717 20247
rect 19576 20216 19717 20244
rect 19576 20204 19582 20216
rect 19705 20213 19717 20216
rect 19751 20213 19763 20247
rect 19705 20207 19763 20213
rect 20162 20204 20168 20256
rect 20220 20244 20226 20256
rect 23290 20244 23296 20256
rect 20220 20216 23296 20244
rect 20220 20204 20226 20216
rect 23290 20204 23296 20216
rect 23348 20204 23354 20256
rect 23934 20204 23940 20256
rect 23992 20244 23998 20256
rect 24121 20247 24179 20253
rect 24121 20244 24133 20247
rect 23992 20216 24133 20244
rect 23992 20204 23998 20216
rect 24121 20213 24133 20216
rect 24167 20213 24179 20247
rect 24121 20207 24179 20213
rect 24854 20204 24860 20256
rect 24912 20244 24918 20256
rect 24949 20247 25007 20253
rect 24949 20244 24961 20247
rect 24912 20216 24961 20244
rect 24912 20204 24918 20216
rect 24949 20213 24961 20216
rect 24995 20213 25007 20247
rect 25056 20244 25084 20284
rect 25314 20272 25320 20324
rect 25372 20312 25378 20324
rect 25976 20312 26004 20408
rect 26068 20324 26096 20411
rect 26142 20408 26148 20460
rect 26200 20408 26206 20460
rect 26252 20380 26280 20488
rect 27062 20476 27068 20528
rect 27120 20516 27126 20528
rect 27525 20519 27583 20525
rect 27525 20516 27537 20519
rect 27120 20488 27537 20516
rect 27120 20476 27126 20488
rect 27525 20485 27537 20488
rect 27571 20516 27583 20519
rect 28258 20516 28264 20528
rect 27571 20488 28264 20516
rect 27571 20485 27583 20488
rect 27525 20479 27583 20485
rect 28258 20476 28264 20488
rect 28316 20476 28322 20528
rect 32030 20516 32036 20528
rect 29196 20488 32036 20516
rect 27249 20451 27307 20457
rect 27249 20417 27261 20451
rect 27295 20448 27307 20451
rect 27338 20448 27344 20460
rect 27295 20420 27344 20448
rect 27295 20417 27307 20420
rect 27249 20411 27307 20417
rect 27338 20408 27344 20420
rect 27396 20408 27402 20460
rect 27433 20451 27491 20457
rect 27433 20417 27445 20451
rect 27479 20417 27491 20451
rect 27433 20411 27491 20417
rect 27448 20380 27476 20411
rect 27614 20408 27620 20460
rect 27672 20408 27678 20460
rect 28534 20408 28540 20460
rect 28592 20448 28598 20460
rect 28905 20451 28963 20457
rect 28905 20448 28917 20451
rect 28592 20420 28917 20448
rect 28592 20408 28598 20420
rect 28905 20417 28917 20420
rect 28951 20417 28963 20451
rect 28905 20411 28963 20417
rect 28994 20408 29000 20460
rect 29052 20448 29058 20460
rect 29089 20451 29147 20457
rect 29089 20448 29101 20451
rect 29052 20420 29101 20448
rect 29052 20408 29058 20420
rect 29089 20417 29101 20420
rect 29135 20417 29147 20451
rect 29089 20411 29147 20417
rect 29196 20380 29224 20488
rect 32030 20476 32036 20488
rect 32088 20516 32094 20528
rect 34422 20516 34428 20528
rect 32088 20488 34428 20516
rect 32088 20476 32094 20488
rect 34422 20476 34428 20488
rect 34480 20476 34486 20528
rect 29733 20451 29791 20457
rect 29733 20417 29745 20451
rect 29779 20448 29791 20451
rect 30285 20451 30343 20457
rect 30285 20448 30297 20451
rect 29779 20420 30297 20448
rect 29779 20417 29791 20420
rect 29733 20411 29791 20417
rect 30285 20417 30297 20420
rect 30331 20448 30343 20451
rect 30374 20448 30380 20460
rect 30331 20420 30380 20448
rect 30331 20417 30343 20420
rect 30285 20411 30343 20417
rect 30374 20408 30380 20420
rect 30432 20408 30438 20460
rect 30561 20451 30619 20457
rect 30561 20417 30573 20451
rect 30607 20448 30619 20451
rect 30650 20448 30656 20460
rect 30607 20420 30656 20448
rect 30607 20417 30619 20420
rect 30561 20411 30619 20417
rect 30650 20408 30656 20420
rect 30708 20408 30714 20460
rect 30745 20451 30803 20457
rect 30745 20417 30757 20451
rect 30791 20448 30803 20451
rect 30926 20448 30932 20460
rect 30791 20420 30932 20448
rect 30791 20417 30803 20420
rect 30745 20411 30803 20417
rect 30926 20408 30932 20420
rect 30984 20408 30990 20460
rect 31021 20451 31079 20457
rect 31021 20417 31033 20451
rect 31067 20448 31079 20451
rect 31110 20448 31116 20460
rect 31067 20420 31116 20448
rect 31067 20417 31079 20420
rect 31021 20411 31079 20417
rect 31110 20408 31116 20420
rect 31168 20408 31174 20460
rect 32582 20408 32588 20460
rect 32640 20448 32646 20460
rect 33137 20451 33195 20457
rect 33137 20448 33149 20451
rect 32640 20420 33149 20448
rect 32640 20408 32646 20420
rect 33137 20417 33149 20420
rect 33183 20417 33195 20451
rect 33137 20411 33195 20417
rect 35894 20408 35900 20460
rect 35952 20408 35958 20460
rect 26252 20352 29224 20380
rect 29638 20340 29644 20392
rect 29696 20340 29702 20392
rect 29748 20352 31754 20380
rect 25372 20284 26004 20312
rect 25372 20272 25378 20284
rect 26050 20272 26056 20324
rect 26108 20272 26114 20324
rect 26234 20272 26240 20324
rect 26292 20312 26298 20324
rect 29748 20312 29776 20352
rect 26292 20284 29776 20312
rect 26292 20272 26298 20284
rect 30650 20272 30656 20324
rect 30708 20272 30714 20324
rect 31726 20312 31754 20352
rect 33226 20340 33232 20392
rect 33284 20340 33290 20392
rect 34422 20340 34428 20392
rect 34480 20380 34486 20392
rect 35621 20383 35679 20389
rect 35621 20380 35633 20383
rect 34480 20352 35633 20380
rect 34480 20340 34486 20352
rect 35621 20349 35633 20352
rect 35667 20349 35679 20383
rect 35621 20343 35679 20349
rect 35713 20383 35771 20389
rect 35713 20349 35725 20383
rect 35759 20349 35771 20383
rect 35713 20343 35771 20349
rect 33134 20312 33140 20324
rect 31726 20284 33140 20312
rect 33134 20272 33140 20284
rect 33192 20272 33198 20324
rect 33505 20315 33563 20321
rect 33505 20281 33517 20315
rect 33551 20312 33563 20315
rect 34514 20312 34520 20324
rect 33551 20284 34520 20312
rect 33551 20281 33563 20284
rect 33505 20275 33563 20281
rect 34514 20272 34520 20284
rect 34572 20272 34578 20324
rect 35728 20312 35756 20343
rect 35802 20340 35808 20392
rect 35860 20340 35866 20392
rect 34808 20284 35756 20312
rect 34808 20256 34836 20284
rect 25958 20244 25964 20256
rect 25056 20216 25964 20244
rect 24949 20207 25007 20213
rect 25958 20204 25964 20216
rect 26016 20204 26022 20256
rect 26329 20247 26387 20253
rect 26329 20213 26341 20247
rect 26375 20244 26387 20247
rect 27154 20244 27160 20256
rect 26375 20216 27160 20244
rect 26375 20213 26387 20216
rect 26329 20207 26387 20213
rect 27154 20204 27160 20216
rect 27212 20204 27218 20256
rect 27430 20204 27436 20256
rect 27488 20244 27494 20256
rect 27614 20244 27620 20256
rect 27488 20216 27620 20244
rect 27488 20204 27494 20216
rect 27614 20204 27620 20216
rect 27672 20204 27678 20256
rect 28905 20247 28963 20253
rect 28905 20213 28917 20247
rect 28951 20244 28963 20247
rect 29546 20244 29552 20256
rect 28951 20216 29552 20244
rect 28951 20213 28963 20216
rect 28905 20207 28963 20213
rect 29546 20204 29552 20216
rect 29604 20204 29610 20256
rect 30009 20247 30067 20253
rect 30009 20213 30021 20247
rect 30055 20244 30067 20247
rect 31202 20244 31208 20256
rect 30055 20216 31208 20244
rect 30055 20213 30067 20216
rect 30009 20207 30067 20213
rect 31202 20204 31208 20216
rect 31260 20204 31266 20256
rect 34790 20204 34796 20256
rect 34848 20204 34854 20256
rect 1104 20154 38272 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 38272 20154
rect 1104 20080 38272 20102
rect 2406 20000 2412 20052
rect 2464 20000 2470 20052
rect 2866 20000 2872 20052
rect 2924 20040 2930 20052
rect 3789 20043 3847 20049
rect 3789 20040 3801 20043
rect 2924 20012 3801 20040
rect 2924 20000 2930 20012
rect 3789 20009 3801 20012
rect 3835 20009 3847 20043
rect 7374 20040 7380 20052
rect 3789 20003 3847 20009
rect 4448 20012 7380 20040
rect 1949 19839 2007 19845
rect 1949 19805 1961 19839
rect 1995 19836 2007 19839
rect 2424 19836 2452 20000
rect 3068 19944 3924 19972
rect 3068 19916 3096 19944
rect 2869 19907 2927 19913
rect 2869 19873 2881 19907
rect 2915 19904 2927 19907
rect 2958 19904 2964 19916
rect 2915 19876 2964 19904
rect 2915 19873 2927 19876
rect 2869 19867 2927 19873
rect 2958 19864 2964 19876
rect 3016 19864 3022 19916
rect 3050 19864 3056 19916
rect 3108 19864 3114 19916
rect 3786 19864 3792 19916
rect 3844 19864 3850 19916
rect 3896 19904 3924 19944
rect 4448 19913 4476 20012
rect 7374 20000 7380 20012
rect 7432 20040 7438 20052
rect 7926 20040 7932 20052
rect 7432 20012 7932 20040
rect 7432 20000 7438 20012
rect 7926 20000 7932 20012
rect 7984 20000 7990 20052
rect 9769 20043 9827 20049
rect 9769 20009 9781 20043
rect 9815 20040 9827 20043
rect 10778 20040 10784 20052
rect 9815 20012 10784 20040
rect 9815 20009 9827 20012
rect 9769 20003 9827 20009
rect 10778 20000 10784 20012
rect 10836 20000 10842 20052
rect 11606 20000 11612 20052
rect 11664 20000 11670 20052
rect 12158 20000 12164 20052
rect 12216 20000 12222 20052
rect 13817 20043 13875 20049
rect 13817 20009 13829 20043
rect 13863 20040 13875 20043
rect 13906 20040 13912 20052
rect 13863 20012 13912 20040
rect 13863 20009 13875 20012
rect 13817 20003 13875 20009
rect 13906 20000 13912 20012
rect 13964 20040 13970 20052
rect 15102 20040 15108 20052
rect 13964 20012 15108 20040
rect 13964 20000 13970 20012
rect 15102 20000 15108 20012
rect 15160 20000 15166 20052
rect 15194 20000 15200 20052
rect 15252 20040 15258 20052
rect 15562 20040 15568 20052
rect 15252 20012 15568 20040
rect 15252 20000 15258 20012
rect 15562 20000 15568 20012
rect 15620 20000 15626 20052
rect 15657 20043 15715 20049
rect 15657 20009 15669 20043
rect 15703 20040 15715 20043
rect 16393 20043 16451 20049
rect 15703 20012 15792 20040
rect 15703 20009 15715 20012
rect 15657 20003 15715 20009
rect 4540 19944 4936 19972
rect 4433 19907 4491 19913
rect 3896 19876 4384 19904
rect 1995 19808 2452 19836
rect 3329 19839 3387 19845
rect 1995 19805 2007 19808
rect 1949 19799 2007 19805
rect 3329 19805 3341 19839
rect 3375 19836 3387 19839
rect 3804 19836 3832 19864
rect 3375 19808 3832 19836
rect 3375 19805 3387 19808
rect 3329 19799 3387 19805
rect 3878 19796 3884 19848
rect 3936 19836 3942 19848
rect 3973 19839 4031 19845
rect 3973 19836 3985 19839
rect 3936 19808 3985 19836
rect 3936 19796 3942 19808
rect 3973 19805 3985 19808
rect 4019 19805 4031 19839
rect 3973 19799 4031 19805
rect 4065 19839 4123 19845
rect 4065 19805 4077 19839
rect 4111 19805 4123 19839
rect 4356 19836 4384 19876
rect 4433 19873 4445 19907
rect 4479 19873 4491 19907
rect 4433 19867 4491 19873
rect 4540 19836 4568 19944
rect 4798 19864 4804 19916
rect 4856 19864 4862 19916
rect 4908 19904 4936 19944
rect 5074 19932 5080 19984
rect 5132 19932 5138 19984
rect 6546 19972 6552 19984
rect 6380 19944 6552 19972
rect 5721 19907 5779 19913
rect 5721 19904 5733 19907
rect 4908 19876 5733 19904
rect 5721 19873 5733 19876
rect 5767 19873 5779 19907
rect 5721 19867 5779 19873
rect 4356 19808 4568 19836
rect 4709 19839 4767 19845
rect 4065 19799 4123 19805
rect 4709 19805 4721 19839
rect 4755 19836 4767 19839
rect 5537 19839 5595 19845
rect 5537 19836 5549 19839
rect 4755 19808 5549 19836
rect 4755 19805 4767 19808
rect 4709 19799 4767 19805
rect 5537 19805 5549 19808
rect 5583 19836 5595 19839
rect 5902 19836 5908 19848
rect 5583 19808 5908 19836
rect 5583 19805 5595 19808
rect 5537 19799 5595 19805
rect 4080 19768 4108 19799
rect 5902 19796 5908 19808
rect 5960 19796 5966 19848
rect 6181 19839 6239 19845
rect 6181 19805 6193 19839
rect 6227 19805 6239 19839
rect 6181 19799 6239 19805
rect 6273 19839 6331 19845
rect 6273 19805 6285 19839
rect 6319 19836 6331 19839
rect 6380 19836 6408 19944
rect 6546 19932 6552 19944
rect 6604 19932 6610 19984
rect 9674 19972 9680 19984
rect 7944 19944 9680 19972
rect 7466 19904 7472 19916
rect 6319 19808 6408 19836
rect 6472 19876 7472 19904
rect 6319 19805 6331 19808
rect 6273 19799 6331 19805
rect 3988 19740 4108 19768
rect 4157 19771 4215 19777
rect 3988 19712 4016 19740
rect 4157 19737 4169 19771
rect 4203 19737 4215 19771
rect 4157 19731 4215 19737
rect 4295 19771 4353 19777
rect 4295 19737 4307 19771
rect 4341 19768 4353 19771
rect 4614 19768 4620 19780
rect 4341 19740 4620 19768
rect 4341 19737 4353 19740
rect 4295 19731 4353 19737
rect 1762 19660 1768 19712
rect 1820 19660 1826 19712
rect 3970 19660 3976 19712
rect 4028 19660 4034 19712
rect 4172 19700 4200 19731
rect 4614 19728 4620 19740
rect 4672 19768 4678 19780
rect 6196 19768 6224 19799
rect 4672 19740 6224 19768
rect 4672 19728 4678 19740
rect 4982 19700 4988 19712
rect 4172 19672 4988 19700
rect 4982 19660 4988 19672
rect 5040 19660 5046 19712
rect 5169 19703 5227 19709
rect 5169 19669 5181 19703
rect 5215 19700 5227 19703
rect 5258 19700 5264 19712
rect 5215 19672 5264 19700
rect 5215 19669 5227 19672
rect 5169 19663 5227 19669
rect 5258 19660 5264 19672
rect 5316 19660 5322 19712
rect 5629 19703 5687 19709
rect 5629 19669 5641 19703
rect 5675 19700 5687 19703
rect 5997 19703 6055 19709
rect 5997 19700 6009 19703
rect 5675 19672 6009 19700
rect 5675 19669 5687 19672
rect 5629 19663 5687 19669
rect 5997 19669 6009 19672
rect 6043 19669 6055 19703
rect 6196 19700 6224 19740
rect 6362 19728 6368 19780
rect 6420 19728 6426 19780
rect 6472 19700 6500 19876
rect 7466 19864 7472 19876
rect 7524 19904 7530 19916
rect 7944 19904 7972 19944
rect 9674 19932 9680 19944
rect 9732 19932 9738 19984
rect 10413 19975 10471 19981
rect 10413 19941 10425 19975
rect 10459 19972 10471 19975
rect 11790 19972 11796 19984
rect 10459 19944 11796 19972
rect 10459 19941 10471 19944
rect 10413 19935 10471 19941
rect 11790 19932 11796 19944
rect 11848 19932 11854 19984
rect 11977 19975 12035 19981
rect 11977 19941 11989 19975
rect 12023 19972 12035 19975
rect 12023 19944 12480 19972
rect 12023 19941 12035 19944
rect 11977 19935 12035 19941
rect 7524 19876 7972 19904
rect 7524 19864 7530 19876
rect 8202 19864 8208 19916
rect 8260 19904 8266 19916
rect 8260 19876 9904 19904
rect 8260 19864 8266 19876
rect 6546 19796 6552 19848
rect 6604 19796 6610 19848
rect 6638 19796 6644 19848
rect 6696 19796 6702 19848
rect 9217 19839 9275 19845
rect 9217 19805 9229 19839
rect 9263 19836 9275 19839
rect 9306 19836 9312 19848
rect 9263 19808 9312 19836
rect 9263 19805 9275 19808
rect 9217 19799 9275 19805
rect 9306 19796 9312 19808
rect 9364 19796 9370 19848
rect 9490 19796 9496 19848
rect 9548 19796 9554 19848
rect 9582 19796 9588 19848
rect 9640 19836 9646 19848
rect 9876 19845 9904 19876
rect 9968 19876 10272 19904
rect 9968 19848 9996 19876
rect 9861 19839 9919 19845
rect 9640 19796 9674 19836
rect 9861 19805 9873 19839
rect 9907 19805 9919 19839
rect 9861 19799 9919 19805
rect 9950 19796 9956 19848
rect 10008 19796 10014 19848
rect 10042 19796 10048 19848
rect 10100 19796 10106 19848
rect 10134 19796 10140 19848
rect 10192 19796 10198 19848
rect 10244 19845 10272 19876
rect 12452 19848 12480 19944
rect 12894 19932 12900 19984
rect 12952 19932 12958 19984
rect 14734 19932 14740 19984
rect 14792 19972 14798 19984
rect 15470 19972 15476 19984
rect 14792 19944 15476 19972
rect 14792 19932 14798 19944
rect 15470 19932 15476 19944
rect 15528 19972 15534 19984
rect 15764 19972 15792 20012
rect 16393 20009 16405 20043
rect 16439 20009 16451 20043
rect 16393 20003 16451 20009
rect 15528 19944 15792 19972
rect 16408 19972 16436 20003
rect 16850 20000 16856 20052
rect 16908 20000 16914 20052
rect 17678 20000 17684 20052
rect 17736 20000 17742 20052
rect 20165 20043 20223 20049
rect 20165 20009 20177 20043
rect 20211 20040 20223 20043
rect 20806 20040 20812 20052
rect 20211 20012 20812 20040
rect 20211 20009 20223 20012
rect 20165 20003 20223 20009
rect 20806 20000 20812 20012
rect 20864 20000 20870 20052
rect 22830 20000 22836 20052
rect 22888 20000 22894 20052
rect 23474 20000 23480 20052
rect 23532 20000 23538 20052
rect 23934 20000 23940 20052
rect 23992 20000 23998 20052
rect 25593 20043 25651 20049
rect 25593 20009 25605 20043
rect 25639 20040 25651 20043
rect 26234 20040 26240 20052
rect 25639 20012 26240 20040
rect 25639 20009 25651 20012
rect 25593 20003 25651 20009
rect 26234 20000 26240 20012
rect 26292 20000 26298 20052
rect 26326 20000 26332 20052
rect 26384 20000 26390 20052
rect 26418 20000 26424 20052
rect 26476 20000 26482 20052
rect 30650 20000 30656 20052
rect 30708 20000 30714 20052
rect 32030 20000 32036 20052
rect 32088 20000 32094 20052
rect 32306 20000 32312 20052
rect 32364 20000 32370 20052
rect 35176 20012 35756 20040
rect 16574 19972 16580 19984
rect 16408 19944 16580 19972
rect 15528 19932 15534 19944
rect 16574 19932 16580 19944
rect 16632 19932 16638 19984
rect 16669 19975 16727 19981
rect 16669 19941 16681 19975
rect 16715 19972 16727 19975
rect 17696 19972 17724 20000
rect 16715 19944 17724 19972
rect 16715 19941 16727 19944
rect 16669 19935 16727 19941
rect 18230 19932 18236 19984
rect 18288 19972 18294 19984
rect 24121 19975 24179 19981
rect 24121 19972 24133 19975
rect 18288 19944 24133 19972
rect 18288 19932 18294 19944
rect 24121 19941 24133 19944
rect 24167 19941 24179 19975
rect 24121 19935 24179 19941
rect 24394 19932 24400 19984
rect 24452 19932 24458 19984
rect 24486 19932 24492 19984
rect 24544 19932 24550 19984
rect 24946 19932 24952 19984
rect 25004 19932 25010 19984
rect 25958 19932 25964 19984
rect 26016 19972 26022 19984
rect 26016 19944 30604 19972
rect 26016 19932 26022 19944
rect 10229 19839 10287 19845
rect 10229 19805 10241 19839
rect 10275 19805 10287 19839
rect 10229 19799 10287 19805
rect 11422 19796 11428 19848
rect 11480 19836 11486 19848
rect 11974 19836 11980 19848
rect 11480 19808 11980 19836
rect 11480 19796 11486 19808
rect 11974 19796 11980 19808
rect 12032 19796 12038 19848
rect 12253 19839 12311 19845
rect 12253 19805 12265 19839
rect 12299 19805 12311 19839
rect 12253 19799 12311 19805
rect 6914 19728 6920 19780
rect 6972 19728 6978 19780
rect 8294 19768 8300 19780
rect 8142 19740 8300 19768
rect 8294 19728 8300 19740
rect 8352 19728 8358 19780
rect 9401 19771 9459 19777
rect 9401 19737 9413 19771
rect 9447 19737 9459 19771
rect 9646 19768 9674 19796
rect 9968 19768 9996 19796
rect 9646 19740 9996 19768
rect 9401 19731 9459 19737
rect 6196 19672 6500 19700
rect 5997 19663 6055 19669
rect 8386 19660 8392 19712
rect 8444 19660 8450 19712
rect 8846 19660 8852 19712
rect 8904 19700 8910 19712
rect 9416 19700 9444 19731
rect 10060 19700 10088 19796
rect 11609 19771 11667 19777
rect 11609 19737 11621 19771
rect 11655 19768 11667 19771
rect 12158 19768 12164 19780
rect 11655 19740 12164 19768
rect 11655 19737 11667 19740
rect 11609 19731 11667 19737
rect 12158 19728 12164 19740
rect 12216 19728 12222 19780
rect 12268 19768 12296 19799
rect 12434 19796 12440 19848
rect 12492 19796 12498 19848
rect 12912 19836 12940 19932
rect 13265 19907 13323 19913
rect 13265 19873 13277 19907
rect 13311 19904 13323 19907
rect 13998 19904 14004 19916
rect 13311 19876 14004 19904
rect 13311 19873 13323 19876
rect 13265 19867 13323 19873
rect 13998 19864 14004 19876
rect 14056 19904 14062 19916
rect 14056 19876 14136 19904
rect 14056 19864 14062 19876
rect 13173 19839 13231 19845
rect 12912 19808 13032 19836
rect 12526 19768 12532 19780
rect 12268 19740 12532 19768
rect 12526 19728 12532 19740
rect 12584 19728 12590 19780
rect 13004 19768 13032 19808
rect 13173 19805 13185 19839
rect 13219 19836 13231 19839
rect 13538 19836 13544 19848
rect 13219 19808 13544 19836
rect 13219 19805 13231 19808
rect 13173 19799 13231 19805
rect 13538 19796 13544 19808
rect 13596 19796 13602 19848
rect 13633 19839 13691 19845
rect 13633 19805 13645 19839
rect 13679 19836 13691 19839
rect 13722 19836 13728 19848
rect 13679 19808 13728 19836
rect 13679 19805 13691 19808
rect 13633 19799 13691 19805
rect 13722 19796 13728 19808
rect 13780 19836 13786 19848
rect 14108 19845 14136 19876
rect 14274 19864 14280 19916
rect 14332 19904 14338 19916
rect 19521 19907 19579 19913
rect 14332 19876 16988 19904
rect 14332 19864 14338 19876
rect 14093 19839 14151 19845
rect 13780 19808 14044 19836
rect 13780 19796 13786 19808
rect 13446 19768 13452 19780
rect 13004 19740 13452 19768
rect 13446 19728 13452 19740
rect 13504 19728 13510 19780
rect 14016 19768 14044 19808
rect 14093 19805 14105 19839
rect 14139 19805 14151 19839
rect 14093 19799 14151 19805
rect 14458 19796 14464 19848
rect 14516 19796 14522 19848
rect 14553 19839 14611 19845
rect 14553 19805 14565 19839
rect 14599 19805 14611 19839
rect 14553 19799 14611 19805
rect 14568 19768 14596 19799
rect 15194 19796 15200 19848
rect 15252 19796 15258 19848
rect 15289 19839 15347 19845
rect 15289 19805 15301 19839
rect 15335 19805 15347 19839
rect 15289 19799 15347 19805
rect 15696 19839 15754 19845
rect 15696 19805 15708 19839
rect 15742 19836 15754 19839
rect 16022 19836 16028 19848
rect 15742 19808 16028 19836
rect 15742 19805 15754 19808
rect 15696 19799 15754 19805
rect 14016 19740 14596 19768
rect 15304 19768 15332 19799
rect 16022 19796 16028 19808
rect 16080 19836 16086 19848
rect 16080 19808 16252 19836
rect 16080 19796 16086 19808
rect 15304 19740 16160 19768
rect 8904 19672 10088 19700
rect 8904 19660 8910 19672
rect 11422 19660 11428 19712
rect 11480 19660 11486 19712
rect 11790 19660 11796 19712
rect 11848 19700 11854 19712
rect 12713 19703 12771 19709
rect 12713 19700 12725 19703
rect 11848 19672 12725 19700
rect 11848 19660 11854 19672
rect 12713 19669 12725 19672
rect 12759 19700 12771 19703
rect 13354 19700 13360 19712
rect 12759 19672 13360 19700
rect 12759 19669 12771 19672
rect 12713 19663 12771 19669
rect 13354 19660 13360 19672
rect 13412 19660 13418 19712
rect 13538 19660 13544 19712
rect 13596 19700 13602 19712
rect 15304 19700 15332 19740
rect 16132 19712 16160 19740
rect 13596 19672 15332 19700
rect 13596 19660 13602 19672
rect 15838 19660 15844 19712
rect 15896 19660 15902 19712
rect 16114 19660 16120 19712
rect 16172 19660 16178 19712
rect 16224 19700 16252 19808
rect 16298 19796 16304 19848
rect 16356 19796 16362 19848
rect 16482 19796 16488 19848
rect 16540 19796 16546 19848
rect 16960 19845 16988 19876
rect 18064 19876 19012 19904
rect 16945 19839 17003 19845
rect 16945 19805 16957 19839
rect 16991 19805 17003 19839
rect 16945 19799 17003 19805
rect 17402 19796 17408 19848
rect 17460 19796 17466 19848
rect 17862 19796 17868 19848
rect 17920 19796 17926 19848
rect 16574 19728 16580 19780
rect 16632 19768 16638 19780
rect 17420 19768 17448 19796
rect 16632 19740 17448 19768
rect 16632 19728 16638 19740
rect 18064 19700 18092 19876
rect 18984 19848 19012 19876
rect 19521 19873 19533 19907
rect 19567 19904 19579 19907
rect 20070 19904 20076 19916
rect 19567 19876 20076 19904
rect 19567 19873 19579 19876
rect 19521 19867 19579 19873
rect 20070 19864 20076 19876
rect 20128 19904 20134 19916
rect 20257 19907 20315 19913
rect 20257 19904 20269 19907
rect 20128 19876 20269 19904
rect 20128 19864 20134 19876
rect 20257 19873 20269 19876
rect 20303 19873 20315 19907
rect 21082 19904 21088 19916
rect 20257 19867 20315 19873
rect 20732 19876 21088 19904
rect 18141 19839 18199 19845
rect 18141 19805 18153 19839
rect 18187 19805 18199 19839
rect 18141 19799 18199 19805
rect 18693 19839 18751 19845
rect 18693 19805 18705 19839
rect 18739 19836 18751 19839
rect 18877 19839 18935 19845
rect 18877 19836 18889 19839
rect 18739 19808 18889 19836
rect 18739 19805 18751 19808
rect 18693 19799 18751 19805
rect 18877 19805 18889 19808
rect 18923 19805 18935 19839
rect 18877 19799 18935 19805
rect 18156 19712 18184 19799
rect 18966 19796 18972 19848
rect 19024 19836 19030 19848
rect 19610 19836 19616 19848
rect 19024 19808 19616 19836
rect 19024 19796 19030 19808
rect 19610 19796 19616 19808
rect 19668 19796 19674 19848
rect 19889 19839 19947 19845
rect 19889 19836 19901 19839
rect 19720 19808 19901 19836
rect 16224 19672 18092 19700
rect 18138 19660 18144 19712
rect 18196 19700 18202 19712
rect 19334 19700 19340 19712
rect 18196 19672 19340 19700
rect 18196 19660 18202 19672
rect 19334 19660 19340 19672
rect 19392 19660 19398 19712
rect 19518 19660 19524 19712
rect 19576 19700 19582 19712
rect 19720 19700 19748 19808
rect 19889 19805 19901 19808
rect 19935 19805 19947 19839
rect 19889 19799 19947 19805
rect 19978 19796 19984 19848
rect 20036 19796 20042 19848
rect 20346 19796 20352 19848
rect 20404 19836 20410 19848
rect 20533 19839 20591 19845
rect 20533 19836 20545 19839
rect 20404 19808 20545 19836
rect 20404 19796 20410 19808
rect 20533 19805 20545 19808
rect 20579 19805 20591 19839
rect 20533 19799 20591 19805
rect 20622 19796 20628 19848
rect 20680 19796 20686 19848
rect 20732 19845 20760 19876
rect 21082 19864 21088 19876
rect 21140 19864 21146 19916
rect 23017 19907 23075 19913
rect 23017 19873 23029 19907
rect 23063 19904 23075 19907
rect 23290 19904 23296 19916
rect 23063 19876 23296 19904
rect 23063 19873 23075 19876
rect 23017 19867 23075 19873
rect 23290 19864 23296 19876
rect 23348 19864 23354 19916
rect 23842 19864 23848 19916
rect 23900 19864 23906 19916
rect 24412 19904 24440 19932
rect 23952 19876 24164 19904
rect 20717 19839 20775 19845
rect 20717 19805 20729 19839
rect 20763 19805 20775 19839
rect 20717 19799 20775 19805
rect 20901 19839 20959 19845
rect 20901 19805 20913 19839
rect 20947 19805 20959 19839
rect 20901 19799 20959 19805
rect 19794 19728 19800 19780
rect 19852 19768 19858 19780
rect 20640 19768 20668 19796
rect 19852 19740 20668 19768
rect 19852 19728 19858 19740
rect 19576 19672 19748 19700
rect 19576 19660 19582 19672
rect 20070 19660 20076 19712
rect 20128 19700 20134 19712
rect 20916 19700 20944 19799
rect 21818 19796 21824 19848
rect 21876 19836 21882 19848
rect 21876 19808 23060 19836
rect 21876 19796 21882 19808
rect 22830 19728 22836 19780
rect 22888 19728 22894 19780
rect 23032 19768 23060 19808
rect 23106 19796 23112 19848
rect 23164 19796 23170 19848
rect 23661 19839 23719 19845
rect 23661 19836 23673 19839
rect 23216 19808 23673 19836
rect 23216 19768 23244 19808
rect 23661 19805 23673 19808
rect 23707 19836 23719 19839
rect 23952 19836 23980 19876
rect 23707 19808 23980 19836
rect 24029 19839 24087 19845
rect 23707 19805 23719 19808
rect 23661 19799 23719 19805
rect 24029 19805 24041 19839
rect 24075 19805 24087 19839
rect 24029 19799 24087 19805
rect 23937 19771 23995 19777
rect 23937 19768 23949 19771
rect 23032 19740 23244 19768
rect 23308 19740 23949 19768
rect 23308 19709 23336 19740
rect 23937 19737 23949 19740
rect 23983 19737 23995 19771
rect 23937 19731 23995 19737
rect 20128 19672 20944 19700
rect 23293 19703 23351 19709
rect 20128 19660 20134 19672
rect 23293 19669 23305 19703
rect 23339 19669 23351 19703
rect 23293 19663 23351 19669
rect 23566 19660 23572 19712
rect 23624 19700 23630 19712
rect 24044 19700 24072 19799
rect 24136 19768 24164 19876
rect 24228 19876 24440 19904
rect 24228 19845 24256 19876
rect 24213 19839 24271 19845
rect 24213 19805 24225 19839
rect 24259 19805 24271 19839
rect 24213 19799 24271 19805
rect 24397 19839 24455 19845
rect 24397 19805 24409 19839
rect 24443 19836 24455 19839
rect 24504 19836 24532 19932
rect 24670 19904 24676 19916
rect 24596 19876 24676 19904
rect 24596 19845 24624 19876
rect 24670 19864 24676 19876
rect 24728 19864 24734 19916
rect 24857 19907 24915 19913
rect 24857 19873 24869 19907
rect 24903 19904 24915 19907
rect 24964 19904 24992 19932
rect 26160 19913 26188 19944
rect 25685 19907 25743 19913
rect 25685 19904 25697 19907
rect 24903 19876 25697 19904
rect 24903 19873 24915 19876
rect 24857 19867 24915 19873
rect 25685 19873 25697 19876
rect 25731 19873 25743 19907
rect 25685 19867 25743 19873
rect 26145 19907 26203 19913
rect 26145 19873 26157 19907
rect 26191 19873 26203 19907
rect 26145 19867 26203 19873
rect 26528 19876 27016 19904
rect 24443 19808 24532 19836
rect 24581 19839 24639 19845
rect 24443 19805 24455 19808
rect 24397 19799 24455 19805
rect 24581 19805 24593 19839
rect 24627 19805 24639 19839
rect 24581 19799 24639 19805
rect 24762 19796 24768 19848
rect 24820 19796 24826 19848
rect 24949 19839 25007 19845
rect 24949 19805 24961 19839
rect 24995 19805 25007 19839
rect 24949 19799 25007 19805
rect 25041 19839 25099 19845
rect 25041 19805 25053 19839
rect 25087 19836 25099 19839
rect 25130 19836 25136 19848
rect 25087 19808 25136 19836
rect 25087 19805 25099 19808
rect 25041 19799 25099 19805
rect 24670 19768 24676 19780
rect 24136 19740 24676 19768
rect 24670 19728 24676 19740
rect 24728 19768 24734 19780
rect 24964 19768 24992 19799
rect 25130 19796 25136 19808
rect 25188 19796 25194 19848
rect 25409 19839 25467 19845
rect 25409 19805 25421 19839
rect 25455 19836 25467 19839
rect 25590 19836 25596 19848
rect 25455 19808 25596 19836
rect 25455 19805 25467 19808
rect 25409 19799 25467 19805
rect 25590 19796 25596 19808
rect 25648 19796 25654 19848
rect 25958 19796 25964 19848
rect 26016 19836 26022 19848
rect 26053 19839 26111 19845
rect 26053 19836 26065 19839
rect 26016 19808 26065 19836
rect 26016 19796 26022 19808
rect 26053 19805 26065 19808
rect 26099 19836 26111 19839
rect 26528 19836 26556 19876
rect 26988 19845 27016 19876
rect 27154 19864 27160 19916
rect 27212 19904 27218 19916
rect 28534 19904 28540 19916
rect 27212 19876 28540 19904
rect 27212 19864 27218 19876
rect 26099 19808 26556 19836
rect 26605 19839 26663 19845
rect 26099 19805 26111 19808
rect 26053 19799 26111 19805
rect 26605 19805 26617 19839
rect 26651 19805 26663 19839
rect 26605 19799 26663 19805
rect 26697 19839 26755 19845
rect 26697 19805 26709 19839
rect 26743 19836 26755 19839
rect 26973 19839 27031 19845
rect 26743 19808 26924 19836
rect 26743 19805 26755 19808
rect 26697 19799 26755 19805
rect 24728 19740 24992 19768
rect 24728 19728 24734 19740
rect 25222 19728 25228 19780
rect 25280 19728 25286 19780
rect 25314 19728 25320 19780
rect 25372 19728 25378 19780
rect 25608 19768 25636 19796
rect 26142 19768 26148 19780
rect 25608 19740 26148 19768
rect 26142 19728 26148 19740
rect 26200 19728 26206 19780
rect 24397 19703 24455 19709
rect 24397 19700 24409 19703
rect 23624 19672 24409 19700
rect 23624 19660 23630 19672
rect 24397 19669 24409 19672
rect 24443 19669 24455 19703
rect 24397 19663 24455 19669
rect 24486 19660 24492 19712
rect 24544 19700 24550 19712
rect 26620 19700 26648 19799
rect 26786 19728 26792 19780
rect 26844 19728 26850 19780
rect 26896 19768 26924 19808
rect 26973 19805 26985 19839
rect 27019 19836 27031 19839
rect 27338 19836 27344 19848
rect 27019 19808 27344 19836
rect 27019 19805 27031 19808
rect 26973 19799 27031 19805
rect 27338 19796 27344 19808
rect 27396 19796 27402 19848
rect 28460 19845 28488 19876
rect 28534 19864 28540 19876
rect 28592 19904 28598 19916
rect 28592 19876 29040 19904
rect 28592 19864 28598 19876
rect 28445 19839 28503 19845
rect 28445 19805 28457 19839
rect 28491 19805 28503 19839
rect 28445 19799 28503 19805
rect 28629 19839 28687 19845
rect 28629 19805 28641 19839
rect 28675 19836 28687 19839
rect 28813 19839 28871 19845
rect 28813 19836 28825 19839
rect 28675 19808 28825 19836
rect 28675 19805 28687 19808
rect 28629 19799 28687 19805
rect 28813 19805 28825 19808
rect 28859 19805 28871 19839
rect 28813 19799 28871 19805
rect 28902 19796 28908 19848
rect 28960 19796 28966 19848
rect 29012 19845 29040 19876
rect 29086 19864 29092 19916
rect 29144 19904 29150 19916
rect 29144 19876 29224 19904
rect 29144 19864 29150 19876
rect 29196 19845 29224 19876
rect 29546 19864 29552 19916
rect 29604 19904 29610 19916
rect 29604 19876 30052 19904
rect 29604 19864 29610 19876
rect 28997 19839 29055 19845
rect 28997 19805 29009 19839
rect 29043 19805 29055 19839
rect 28997 19799 29055 19805
rect 29181 19839 29239 19845
rect 29181 19805 29193 19839
rect 29227 19805 29239 19839
rect 29181 19799 29239 19805
rect 29638 19796 29644 19848
rect 29696 19836 29702 19848
rect 29733 19839 29791 19845
rect 29733 19836 29745 19839
rect 29696 19808 29745 19836
rect 29696 19796 29702 19808
rect 29733 19805 29745 19808
rect 29779 19805 29791 19839
rect 29733 19799 29791 19805
rect 29822 19796 29828 19848
rect 29880 19796 29886 19848
rect 30024 19845 30052 19876
rect 30009 19839 30067 19845
rect 30009 19805 30021 19839
rect 30055 19805 30067 19839
rect 30009 19799 30067 19805
rect 30101 19839 30159 19845
rect 30101 19805 30113 19839
rect 30147 19805 30159 19839
rect 30101 19799 30159 19805
rect 27062 19768 27068 19780
rect 26896 19740 27068 19768
rect 27062 19728 27068 19740
rect 27120 19768 27126 19780
rect 27614 19768 27620 19780
rect 27120 19740 27620 19768
rect 27120 19728 27126 19740
rect 27614 19728 27620 19740
rect 27672 19728 27678 19780
rect 28537 19771 28595 19777
rect 28537 19737 28549 19771
rect 28583 19768 28595 19771
rect 29270 19768 29276 19780
rect 28583 19740 29276 19768
rect 28583 19737 28595 19740
rect 28537 19731 28595 19737
rect 29270 19728 29276 19740
rect 29328 19728 29334 19780
rect 29840 19768 29868 19796
rect 29472 19740 29868 19768
rect 24544 19672 26648 19700
rect 29181 19703 29239 19709
rect 24544 19660 24550 19672
rect 29181 19669 29193 19703
rect 29227 19700 29239 19703
rect 29472 19700 29500 19740
rect 29227 19672 29500 19700
rect 29227 19669 29239 19672
rect 29181 19663 29239 19669
rect 29546 19660 29552 19712
rect 29604 19660 29610 19712
rect 29730 19660 29736 19712
rect 29788 19700 29794 19712
rect 30024 19700 30052 19799
rect 30116 19768 30144 19799
rect 30282 19796 30288 19848
rect 30340 19836 30346 19848
rect 30377 19839 30435 19845
rect 30377 19836 30389 19839
rect 30340 19808 30389 19836
rect 30340 19796 30346 19808
rect 30377 19805 30389 19808
rect 30423 19805 30435 19839
rect 30377 19799 30435 19805
rect 30466 19768 30472 19780
rect 30116 19740 30472 19768
rect 30466 19728 30472 19740
rect 30524 19728 30530 19780
rect 30576 19768 30604 19944
rect 30668 19845 30696 20000
rect 31665 19975 31723 19981
rect 31665 19941 31677 19975
rect 31711 19941 31723 19975
rect 31665 19935 31723 19941
rect 31202 19864 31208 19916
rect 31260 19864 31266 19916
rect 31680 19904 31708 19935
rect 32048 19913 32076 20000
rect 32324 19972 32352 20000
rect 35176 19984 35204 20012
rect 32324 19944 33088 19972
rect 32033 19907 32091 19913
rect 31680 19876 31754 19904
rect 30653 19839 30711 19845
rect 30653 19805 30665 19839
rect 30699 19805 30711 19839
rect 30653 19799 30711 19805
rect 31481 19839 31539 19845
rect 31481 19805 31493 19839
rect 31527 19836 31539 19839
rect 31570 19836 31576 19848
rect 31527 19808 31576 19836
rect 31527 19805 31539 19808
rect 31481 19799 31539 19805
rect 31570 19796 31576 19808
rect 31628 19796 31634 19848
rect 31726 19768 31754 19876
rect 32033 19873 32045 19907
rect 32079 19873 32091 19907
rect 32033 19867 32091 19873
rect 32309 19907 32367 19913
rect 32309 19873 32321 19907
rect 32355 19873 32367 19907
rect 32309 19867 32367 19873
rect 31941 19839 31999 19845
rect 31941 19805 31953 19839
rect 31987 19805 31999 19839
rect 31941 19799 31999 19805
rect 31956 19768 31984 19799
rect 30576 19740 31984 19768
rect 32324 19768 32352 19867
rect 33060 19848 33088 19944
rect 33410 19932 33416 19984
rect 33468 19972 33474 19984
rect 33468 19944 34744 19972
rect 33468 19932 33474 19944
rect 33134 19864 33140 19916
rect 33192 19904 33198 19916
rect 33192 19876 33640 19904
rect 33192 19864 33198 19876
rect 33042 19796 33048 19848
rect 33100 19836 33106 19848
rect 33612 19845 33640 19876
rect 33413 19839 33471 19845
rect 33413 19836 33425 19839
rect 33100 19808 33425 19836
rect 33100 19796 33106 19808
rect 33413 19805 33425 19808
rect 33459 19805 33471 19839
rect 33413 19799 33471 19805
rect 33597 19839 33655 19845
rect 33597 19805 33609 19839
rect 33643 19805 33655 19839
rect 33597 19799 33655 19805
rect 34716 19780 34744 19944
rect 35158 19932 35164 19984
rect 35216 19932 35222 19984
rect 35728 19972 35756 20012
rect 35802 20000 35808 20052
rect 35860 20040 35866 20052
rect 36725 20043 36783 20049
rect 36725 20040 36737 20043
rect 35860 20012 36737 20040
rect 35860 20000 35866 20012
rect 36725 20009 36737 20012
rect 36771 20009 36783 20043
rect 36725 20003 36783 20009
rect 36354 19972 36360 19984
rect 35728 19944 36360 19972
rect 36354 19932 36360 19944
rect 36412 19972 36418 19984
rect 36412 19944 36584 19972
rect 36412 19932 36418 19944
rect 35710 19864 35716 19916
rect 35768 19904 35774 19916
rect 36081 19907 36139 19913
rect 36081 19904 36093 19907
rect 35768 19876 36093 19904
rect 35768 19864 35774 19876
rect 36081 19873 36093 19876
rect 36127 19904 36139 19907
rect 36170 19904 36176 19916
rect 36127 19876 36176 19904
rect 36127 19873 36139 19876
rect 36081 19867 36139 19873
rect 36170 19864 36176 19876
rect 36228 19864 36234 19916
rect 36446 19864 36452 19916
rect 36504 19864 36510 19916
rect 35069 19839 35127 19845
rect 35069 19805 35081 19839
rect 35115 19805 35127 19839
rect 35069 19799 35127 19805
rect 34606 19768 34612 19780
rect 32324 19740 34612 19768
rect 34606 19728 34612 19740
rect 34664 19728 34670 19780
rect 34698 19728 34704 19780
rect 34756 19768 34762 19780
rect 34885 19771 34943 19777
rect 34885 19768 34897 19771
rect 34756 19740 34897 19768
rect 34756 19728 34762 19740
rect 34885 19737 34897 19740
rect 34931 19737 34943 19771
rect 35084 19768 35112 19799
rect 35158 19796 35164 19848
rect 35216 19796 35222 19848
rect 35250 19796 35256 19848
rect 35308 19826 35314 19848
rect 35345 19839 35403 19845
rect 35345 19826 35357 19839
rect 35308 19805 35357 19826
rect 35391 19805 35403 19839
rect 35308 19799 35403 19805
rect 35308 19798 35388 19799
rect 35308 19796 35314 19798
rect 35434 19796 35440 19848
rect 35492 19796 35498 19848
rect 35986 19796 35992 19848
rect 36044 19796 36050 19848
rect 36556 19845 36584 19944
rect 36357 19839 36415 19845
rect 36357 19805 36369 19839
rect 36403 19805 36415 19839
rect 36357 19799 36415 19805
rect 36541 19839 36599 19845
rect 36541 19805 36553 19839
rect 36587 19836 36599 19839
rect 36633 19839 36691 19845
rect 36633 19836 36645 19839
rect 36587 19808 36645 19836
rect 36587 19805 36599 19808
rect 36541 19799 36599 19805
rect 36633 19805 36645 19808
rect 36679 19805 36691 19839
rect 36633 19799 36691 19805
rect 36372 19768 36400 19799
rect 35084 19740 35572 19768
rect 34885 19731 34943 19737
rect 29788 19672 30052 19700
rect 29788 19660 29794 19672
rect 30098 19660 30104 19712
rect 30156 19700 30162 19712
rect 33410 19700 33416 19712
rect 30156 19672 33416 19700
rect 30156 19660 30162 19672
rect 33410 19660 33416 19672
rect 33468 19660 33474 19712
rect 33505 19703 33563 19709
rect 33505 19669 33517 19703
rect 33551 19700 33563 19703
rect 34790 19700 34796 19712
rect 33551 19672 34796 19700
rect 33551 19669 33563 19672
rect 33505 19663 33563 19669
rect 34790 19660 34796 19672
rect 34848 19660 34854 19712
rect 35544 19709 35572 19740
rect 35728 19740 36400 19768
rect 35529 19703 35587 19709
rect 35529 19669 35541 19703
rect 35575 19700 35587 19703
rect 35728 19700 35756 19740
rect 35575 19672 35756 19700
rect 35897 19703 35955 19709
rect 35575 19669 35587 19672
rect 35529 19663 35587 19669
rect 35897 19669 35909 19703
rect 35943 19700 35955 19703
rect 36078 19700 36084 19712
rect 35943 19672 36084 19700
rect 35943 19669 35955 19672
rect 35897 19663 35955 19669
rect 36078 19660 36084 19672
rect 36136 19660 36142 19712
rect 1104 19610 38272 19632
rect 1104 19558 4874 19610
rect 4926 19558 4938 19610
rect 4990 19558 5002 19610
rect 5054 19558 5066 19610
rect 5118 19558 5130 19610
rect 5182 19558 35594 19610
rect 35646 19558 35658 19610
rect 35710 19558 35722 19610
rect 35774 19558 35786 19610
rect 35838 19558 35850 19610
rect 35902 19558 38272 19610
rect 1104 19536 38272 19558
rect 1394 19456 1400 19508
rect 1452 19496 1458 19508
rect 3510 19496 3516 19508
rect 1452 19468 3516 19496
rect 1452 19456 1458 19468
rect 3510 19456 3516 19468
rect 3568 19456 3574 19508
rect 5902 19456 5908 19508
rect 5960 19456 5966 19508
rect 6914 19456 6920 19508
rect 6972 19496 6978 19508
rect 7009 19499 7067 19505
rect 7009 19496 7021 19499
rect 6972 19468 7021 19496
rect 6972 19456 6978 19468
rect 7009 19465 7021 19468
rect 7055 19465 7067 19499
rect 7009 19459 7067 19465
rect 7190 19456 7196 19508
rect 7248 19456 7254 19508
rect 8110 19456 8116 19508
rect 8168 19496 8174 19508
rect 9309 19499 9367 19505
rect 9309 19496 9321 19499
rect 8168 19468 9321 19496
rect 8168 19456 8174 19468
rect 9309 19465 9321 19468
rect 9355 19465 9367 19499
rect 9309 19459 9367 19465
rect 9582 19456 9588 19508
rect 9640 19456 9646 19508
rect 11790 19496 11796 19508
rect 9692 19468 11796 19496
rect 1412 19369 1440 19456
rect 1673 19431 1731 19437
rect 1673 19397 1685 19431
rect 1719 19428 1731 19431
rect 1762 19428 1768 19440
rect 1719 19400 1768 19428
rect 1719 19397 1731 19400
rect 1673 19391 1731 19397
rect 1762 19388 1768 19400
rect 1820 19388 1826 19440
rect 2958 19428 2964 19440
rect 2898 19400 2964 19428
rect 2958 19388 2964 19400
rect 3016 19428 3022 19440
rect 4706 19428 4712 19440
rect 3016 19400 4712 19428
rect 3016 19388 3022 19400
rect 4706 19388 4712 19400
rect 4764 19428 4770 19440
rect 4890 19428 4896 19440
rect 4764 19400 4896 19428
rect 4764 19388 4770 19400
rect 4890 19388 4896 19400
rect 4948 19388 4954 19440
rect 1397 19363 1455 19369
rect 1397 19329 1409 19363
rect 1443 19329 1455 19363
rect 1397 19323 1455 19329
rect 3513 19363 3571 19369
rect 3513 19329 3525 19363
rect 3559 19360 3571 19363
rect 3602 19360 3608 19372
rect 3559 19332 3608 19360
rect 3559 19329 3571 19332
rect 3513 19323 3571 19329
rect 3602 19320 3608 19332
rect 3660 19320 3666 19372
rect 7208 19369 7236 19456
rect 8846 19388 8852 19440
rect 8904 19428 8910 19440
rect 8941 19431 8999 19437
rect 8941 19428 8953 19431
rect 8904 19400 8953 19428
rect 8904 19388 8910 19400
rect 8941 19397 8953 19400
rect 8987 19397 8999 19431
rect 9600 19428 9628 19456
rect 8941 19391 8999 19397
rect 9140 19400 9628 19428
rect 3697 19363 3755 19369
rect 3697 19329 3709 19363
rect 3743 19329 3755 19363
rect 4157 19363 4215 19369
rect 4157 19360 4169 19363
rect 3697 19323 3755 19329
rect 3804 19332 4169 19360
rect 3712 19292 3740 19323
rect 3160 19264 3740 19292
rect 3160 19236 3188 19264
rect 3142 19184 3148 19236
rect 3200 19184 3206 19236
rect 3804 19224 3832 19332
rect 4157 19329 4169 19332
rect 4203 19329 4215 19363
rect 7193 19363 7251 19369
rect 4157 19323 4215 19329
rect 5460 19332 7144 19360
rect 3878 19252 3884 19304
rect 3936 19252 3942 19304
rect 4433 19295 4491 19301
rect 4433 19261 4445 19295
rect 4479 19292 4491 19295
rect 4798 19292 4804 19304
rect 4479 19264 4804 19292
rect 4479 19261 4491 19264
rect 4433 19255 4491 19261
rect 4798 19252 4804 19264
rect 4856 19252 4862 19304
rect 4890 19252 4896 19304
rect 4948 19292 4954 19304
rect 5460 19292 5488 19332
rect 4948 19264 5488 19292
rect 7116 19292 7144 19332
rect 7193 19329 7205 19363
rect 7239 19329 7251 19363
rect 7929 19363 7987 19369
rect 7929 19360 7941 19363
rect 7193 19323 7251 19329
rect 7300 19332 7941 19360
rect 7300 19292 7328 19332
rect 7929 19329 7941 19332
rect 7975 19329 7987 19363
rect 7929 19323 7987 19329
rect 8754 19320 8760 19372
rect 8812 19320 8818 19372
rect 9030 19320 9036 19372
rect 9088 19320 9094 19372
rect 9140 19369 9168 19400
rect 9125 19363 9183 19369
rect 9125 19329 9137 19363
rect 9171 19329 9183 19363
rect 9125 19323 9183 19329
rect 9490 19320 9496 19372
rect 9548 19360 9554 19372
rect 9585 19363 9643 19369
rect 9585 19360 9597 19363
rect 9548 19332 9597 19360
rect 9548 19320 9554 19332
rect 9585 19329 9597 19332
rect 9631 19360 9643 19363
rect 9692 19360 9720 19468
rect 11790 19456 11796 19468
rect 11848 19456 11854 19508
rect 12345 19499 12403 19505
rect 12345 19465 12357 19499
rect 12391 19465 12403 19499
rect 12345 19459 12403 19465
rect 11164 19400 11560 19428
rect 9631 19332 9720 19360
rect 9769 19363 9827 19369
rect 9631 19329 9643 19332
rect 9585 19323 9643 19329
rect 9769 19329 9781 19363
rect 9815 19360 9827 19363
rect 9950 19360 9956 19372
rect 9815 19332 9956 19360
rect 9815 19329 9827 19332
rect 9769 19323 9827 19329
rect 9950 19320 9956 19332
rect 10008 19360 10014 19372
rect 10226 19360 10232 19372
rect 10008 19332 10232 19360
rect 10008 19320 10014 19332
rect 10226 19320 10232 19332
rect 10284 19320 10290 19372
rect 11164 19369 11192 19400
rect 11532 19372 11560 19400
rect 11149 19363 11207 19369
rect 11149 19329 11161 19363
rect 11195 19329 11207 19363
rect 11149 19323 11207 19329
rect 11333 19363 11391 19369
rect 11333 19329 11345 19363
rect 11379 19360 11391 19363
rect 11379 19332 11413 19360
rect 11379 19329 11391 19332
rect 11333 19323 11391 19329
rect 7116 19264 7328 19292
rect 4948 19252 4954 19264
rect 8294 19252 8300 19304
rect 8352 19252 8358 19304
rect 9306 19252 9312 19304
rect 9364 19292 9370 19304
rect 9401 19295 9459 19301
rect 9401 19292 9413 19295
rect 9364 19264 9413 19292
rect 9364 19252 9370 19264
rect 9401 19261 9413 19264
rect 9447 19261 9459 19295
rect 11348 19292 11376 19323
rect 11514 19320 11520 19372
rect 11572 19360 11578 19372
rect 11790 19360 11796 19372
rect 11572 19332 11796 19360
rect 11572 19320 11578 19332
rect 11790 19320 11796 19332
rect 11848 19320 11854 19372
rect 11977 19363 12035 19369
rect 11977 19329 11989 19363
rect 12023 19360 12035 19363
rect 12360 19360 12388 19459
rect 13170 19456 13176 19508
rect 13228 19456 13234 19508
rect 14458 19456 14464 19508
rect 14516 19496 14522 19508
rect 14734 19496 14740 19508
rect 14516 19468 14740 19496
rect 14516 19456 14522 19468
rect 14734 19456 14740 19468
rect 14792 19456 14798 19508
rect 15470 19456 15476 19508
rect 15528 19496 15534 19508
rect 15746 19496 15752 19508
rect 15528 19468 15752 19496
rect 15528 19456 15534 19468
rect 15746 19456 15752 19468
rect 15804 19456 15810 19508
rect 15838 19456 15844 19508
rect 15896 19456 15902 19508
rect 19797 19499 19855 19505
rect 19797 19465 19809 19499
rect 19843 19496 19855 19499
rect 19978 19496 19984 19508
rect 19843 19468 19984 19496
rect 19843 19465 19855 19468
rect 19797 19459 19855 19465
rect 19978 19456 19984 19468
rect 20036 19456 20042 19508
rect 22002 19456 22008 19508
rect 22060 19496 22066 19508
rect 22649 19499 22707 19505
rect 22060 19456 22094 19496
rect 22649 19465 22661 19499
rect 22695 19496 22707 19499
rect 22830 19496 22836 19508
rect 22695 19468 22836 19496
rect 22695 19465 22707 19468
rect 22649 19459 22707 19465
rect 22830 19456 22836 19468
rect 22888 19456 22894 19508
rect 22922 19456 22928 19508
rect 22980 19496 22986 19508
rect 25130 19496 25136 19508
rect 22980 19468 25136 19496
rect 22980 19456 22986 19468
rect 25130 19456 25136 19468
rect 25188 19456 25194 19508
rect 27801 19499 27859 19505
rect 27801 19465 27813 19499
rect 27847 19496 27859 19499
rect 28718 19496 28724 19508
rect 27847 19468 28724 19496
rect 27847 19465 27859 19468
rect 27801 19459 27859 19465
rect 28718 19456 28724 19468
rect 28776 19456 28782 19508
rect 29546 19456 29552 19508
rect 29604 19456 29610 19508
rect 29730 19456 29736 19508
rect 29788 19456 29794 19508
rect 29822 19456 29828 19508
rect 29880 19456 29886 19508
rect 30193 19499 30251 19505
rect 30193 19465 30205 19499
rect 30239 19496 30251 19499
rect 30374 19496 30380 19508
rect 30239 19468 30380 19496
rect 30239 19465 30251 19468
rect 30193 19459 30251 19465
rect 30374 19456 30380 19468
rect 30432 19456 30438 19508
rect 33781 19499 33839 19505
rect 33781 19465 33793 19499
rect 33827 19465 33839 19499
rect 33781 19459 33839 19465
rect 33965 19499 34023 19505
rect 33965 19465 33977 19499
rect 34011 19496 34023 19499
rect 34011 19468 34560 19496
rect 34011 19465 34023 19468
rect 33965 19459 34023 19465
rect 12434 19388 12440 19440
rect 12492 19428 12498 19440
rect 12989 19431 13047 19437
rect 12989 19428 13001 19431
rect 12492 19400 13001 19428
rect 12492 19388 12498 19400
rect 12989 19397 13001 19400
rect 13035 19428 13047 19431
rect 14642 19428 14648 19440
rect 13035 19400 14648 19428
rect 13035 19397 13047 19400
rect 12989 19391 13047 19397
rect 14642 19388 14648 19400
rect 14700 19388 14706 19440
rect 12023 19332 12388 19360
rect 12023 19329 12035 19332
rect 11977 19323 12035 19329
rect 12526 19320 12532 19372
rect 12584 19320 12590 19372
rect 12621 19363 12679 19369
rect 12621 19329 12633 19363
rect 12667 19334 12679 19363
rect 12667 19329 12701 19334
rect 12621 19323 12701 19329
rect 12636 19306 12701 19323
rect 13354 19320 13360 19372
rect 13412 19320 13418 19372
rect 14366 19320 14372 19372
rect 14424 19320 14430 19372
rect 14550 19320 14556 19372
rect 14608 19320 14614 19372
rect 14752 19369 14780 19456
rect 14737 19363 14795 19369
rect 14737 19329 14749 19363
rect 14783 19329 14795 19363
rect 15856 19360 15884 19456
rect 16114 19388 16120 19440
rect 16172 19428 16178 19440
rect 20898 19428 20904 19440
rect 16172 19400 20904 19428
rect 16172 19388 16178 19400
rect 20898 19388 20904 19400
rect 20956 19388 20962 19440
rect 22066 19428 22094 19456
rect 22189 19431 22247 19437
rect 22189 19428 22201 19431
rect 22066 19400 22201 19428
rect 22189 19397 22201 19400
rect 22235 19428 22247 19431
rect 23750 19428 23756 19440
rect 22235 19400 23756 19428
rect 22235 19397 22247 19400
rect 22189 19391 22247 19397
rect 23750 19388 23756 19400
rect 23808 19428 23814 19440
rect 24486 19428 24492 19440
rect 23808 19400 24492 19428
rect 23808 19388 23814 19400
rect 24486 19388 24492 19400
rect 24544 19388 24550 19440
rect 29564 19428 29592 19456
rect 24596 19400 29040 19428
rect 16669 19363 16727 19369
rect 16669 19360 16681 19363
rect 15856 19332 15976 19360
rect 14737 19323 14795 19329
rect 11348 19264 11744 19292
rect 9401 19255 9459 19261
rect 11716 19233 11744 19264
rect 11882 19252 11888 19304
rect 11940 19252 11946 19304
rect 12066 19252 12072 19304
rect 12124 19292 12130 19304
rect 12636 19292 12664 19306
rect 12124 19264 12664 19292
rect 13541 19295 13599 19301
rect 12124 19252 12130 19264
rect 13541 19261 13553 19295
rect 13587 19292 13599 19295
rect 14918 19292 14924 19304
rect 13587 19264 14924 19292
rect 13587 19261 13599 19264
rect 13541 19255 13599 19261
rect 14918 19252 14924 19264
rect 14976 19252 14982 19304
rect 15948 19292 15976 19332
rect 16132 19332 16681 19360
rect 16132 19292 16160 19332
rect 16669 19329 16681 19332
rect 16715 19329 16727 19363
rect 16669 19323 16727 19329
rect 17129 19363 17187 19369
rect 17129 19329 17141 19363
rect 17175 19329 17187 19363
rect 17129 19323 17187 19329
rect 15948 19264 16160 19292
rect 16390 19252 16396 19304
rect 16448 19292 16454 19304
rect 16761 19295 16819 19301
rect 16761 19292 16773 19295
rect 16448 19264 16773 19292
rect 16448 19252 16454 19264
rect 16761 19261 16773 19264
rect 16807 19261 16819 19295
rect 16761 19255 16819 19261
rect 3528 19196 3832 19224
rect 11701 19227 11759 19233
rect 3528 19168 3556 19196
rect 11701 19193 11713 19227
rect 11747 19224 11759 19227
rect 12342 19224 12348 19236
rect 11747 19196 12348 19224
rect 11747 19193 11759 19196
rect 11701 19187 11759 19193
rect 12342 19184 12348 19196
rect 12400 19184 12406 19236
rect 14642 19184 14648 19236
rect 14700 19184 14706 19236
rect 3510 19116 3516 19168
rect 3568 19116 3574 19168
rect 11330 19116 11336 19168
rect 11388 19116 11394 19168
rect 11793 19159 11851 19165
rect 11793 19125 11805 19159
rect 11839 19156 11851 19159
rect 11882 19156 11888 19168
rect 11839 19128 11888 19156
rect 11839 19125 11851 19128
rect 11793 19119 11851 19125
rect 11882 19116 11888 19128
rect 11940 19116 11946 19168
rect 12250 19116 12256 19168
rect 12308 19116 12314 19168
rect 12897 19159 12955 19165
rect 12897 19125 12909 19159
rect 12943 19156 12955 19159
rect 13630 19156 13636 19168
rect 12943 19128 13636 19156
rect 12943 19125 12955 19128
rect 12897 19119 12955 19125
rect 13630 19116 13636 19128
rect 13688 19116 13694 19168
rect 16298 19116 16304 19168
rect 16356 19156 16362 19168
rect 17144 19156 17172 19323
rect 17402 19320 17408 19372
rect 17460 19360 17466 19372
rect 17589 19363 17647 19369
rect 17589 19360 17601 19363
rect 17460 19332 17601 19360
rect 17460 19320 17466 19332
rect 17589 19329 17601 19332
rect 17635 19329 17647 19363
rect 17589 19323 17647 19329
rect 18141 19363 18199 19369
rect 18141 19329 18153 19363
rect 18187 19360 18199 19363
rect 19426 19360 19432 19372
rect 18187 19332 19432 19360
rect 18187 19329 18199 19332
rect 18141 19323 18199 19329
rect 19426 19320 19432 19332
rect 19484 19320 19490 19372
rect 19610 19320 19616 19372
rect 19668 19360 19674 19372
rect 19705 19363 19763 19369
rect 19705 19360 19717 19363
rect 19668 19332 19717 19360
rect 19668 19320 19674 19332
rect 19705 19329 19717 19332
rect 19751 19329 19763 19363
rect 19705 19323 19763 19329
rect 19889 19363 19947 19369
rect 19889 19329 19901 19363
rect 19935 19329 19947 19363
rect 19889 19323 19947 19329
rect 18233 19295 18291 19301
rect 18233 19261 18245 19295
rect 18279 19292 18291 19295
rect 18322 19292 18328 19304
rect 18279 19264 18328 19292
rect 18279 19261 18291 19264
rect 18233 19255 18291 19261
rect 18322 19252 18328 19264
rect 18380 19252 18386 19304
rect 19334 19252 19340 19304
rect 19392 19292 19398 19304
rect 19904 19292 19932 19323
rect 22370 19320 22376 19372
rect 22428 19320 22434 19372
rect 22462 19320 22468 19372
rect 22520 19320 22526 19372
rect 22554 19320 22560 19372
rect 22612 19360 22618 19372
rect 22741 19363 22799 19369
rect 22741 19360 22753 19363
rect 22612 19332 22753 19360
rect 22612 19320 22618 19332
rect 22741 19329 22753 19332
rect 22787 19329 22799 19363
rect 22741 19323 22799 19329
rect 23474 19320 23480 19372
rect 23532 19360 23538 19372
rect 23569 19363 23627 19369
rect 23569 19360 23581 19363
rect 23532 19332 23581 19360
rect 23532 19320 23538 19332
rect 23569 19329 23581 19332
rect 23615 19360 23627 19363
rect 23658 19360 23664 19372
rect 23615 19332 23664 19360
rect 23615 19329 23627 19332
rect 23569 19323 23627 19329
rect 23658 19320 23664 19332
rect 23716 19360 23722 19372
rect 24029 19363 24087 19369
rect 24029 19360 24041 19363
rect 23716 19332 24041 19360
rect 23716 19320 23722 19332
rect 24029 19329 24041 19332
rect 24075 19360 24087 19363
rect 24596 19360 24624 19400
rect 24075 19332 24624 19360
rect 24075 19329 24087 19332
rect 24029 19323 24087 19329
rect 27246 19320 27252 19372
rect 27304 19320 27310 19372
rect 27338 19320 27344 19372
rect 27396 19360 27402 19372
rect 27433 19363 27491 19369
rect 27433 19360 27445 19363
rect 27396 19332 27445 19360
rect 27396 19320 27402 19332
rect 27433 19329 27445 19332
rect 27479 19329 27491 19363
rect 27433 19323 27491 19329
rect 27522 19320 27528 19372
rect 27580 19320 27586 19372
rect 27617 19363 27675 19369
rect 27617 19329 27629 19363
rect 27663 19329 27675 19363
rect 27617 19323 27675 19329
rect 19392 19264 19932 19292
rect 19392 19252 19398 19264
rect 23842 19252 23848 19304
rect 23900 19252 23906 19304
rect 24305 19295 24363 19301
rect 24305 19261 24317 19295
rect 24351 19292 24363 19295
rect 27356 19292 27384 19320
rect 24351 19264 27384 19292
rect 24351 19261 24363 19264
rect 24305 19255 24363 19261
rect 17218 19184 17224 19236
rect 17276 19224 17282 19236
rect 24320 19224 24348 19255
rect 17276 19196 24348 19224
rect 17276 19184 17282 19196
rect 25774 19184 25780 19236
rect 25832 19224 25838 19236
rect 27632 19224 27660 19323
rect 27798 19320 27804 19372
rect 27856 19360 27862 19372
rect 27893 19363 27951 19369
rect 27893 19360 27905 19363
rect 27856 19332 27905 19360
rect 27856 19320 27862 19332
rect 27893 19329 27905 19332
rect 27939 19329 27951 19363
rect 27893 19323 27951 19329
rect 28166 19320 28172 19372
rect 28224 19320 28230 19372
rect 28258 19320 28264 19372
rect 28316 19320 28322 19372
rect 29012 19369 29040 19400
rect 29196 19400 29592 19428
rect 29196 19369 29224 19400
rect 28997 19363 29055 19369
rect 28997 19329 29009 19363
rect 29043 19329 29055 19363
rect 28997 19323 29055 19329
rect 29181 19363 29239 19369
rect 29181 19329 29193 19363
rect 29227 19329 29239 19363
rect 29181 19323 29239 19329
rect 29270 19320 29276 19372
rect 29328 19320 29334 19372
rect 29454 19320 29460 19372
rect 29512 19320 29518 19372
rect 29748 19369 29776 19456
rect 29840 19428 29868 19456
rect 33042 19428 33048 19440
rect 29840 19400 30236 19428
rect 30208 19369 30236 19400
rect 32968 19400 33048 19428
rect 32968 19369 32996 19400
rect 33042 19388 33048 19400
rect 33100 19428 33106 19440
rect 33321 19431 33379 19437
rect 33321 19428 33333 19431
rect 33100 19400 33333 19428
rect 33100 19388 33106 19400
rect 33321 19397 33333 19400
rect 33367 19397 33379 19431
rect 33796 19428 33824 19459
rect 33796 19400 34468 19428
rect 33321 19391 33379 19397
rect 29733 19363 29791 19369
rect 29733 19329 29745 19363
rect 29779 19329 29791 19363
rect 29733 19323 29791 19329
rect 29825 19363 29883 19369
rect 29825 19329 29837 19363
rect 29871 19360 29883 19363
rect 30009 19363 30067 19369
rect 30009 19360 30021 19363
rect 29871 19332 30021 19360
rect 29871 19329 29883 19332
rect 29825 19323 29883 19329
rect 30009 19329 30021 19332
rect 30055 19329 30067 19363
rect 30009 19323 30067 19329
rect 30193 19363 30251 19369
rect 30193 19329 30205 19363
rect 30239 19329 30251 19363
rect 30193 19323 30251 19329
rect 32953 19363 33011 19369
rect 32953 19329 32965 19363
rect 32999 19329 33011 19363
rect 32953 19323 33011 19329
rect 33134 19320 33140 19372
rect 33192 19320 33198 19372
rect 33873 19363 33931 19369
rect 33873 19360 33885 19363
rect 33704 19332 33885 19360
rect 29365 19295 29423 19301
rect 29365 19261 29377 19295
rect 29411 19292 29423 19295
rect 30282 19292 30288 19304
rect 29411 19264 30288 19292
rect 29411 19261 29423 19264
rect 29365 19255 29423 19261
rect 30282 19252 30288 19264
rect 30340 19252 30346 19304
rect 30466 19252 30472 19304
rect 30524 19292 30530 19304
rect 31570 19292 31576 19304
rect 30524 19264 31576 19292
rect 30524 19252 30530 19264
rect 31570 19252 31576 19264
rect 31628 19252 31634 19304
rect 25832 19196 27660 19224
rect 33152 19224 33180 19320
rect 33597 19227 33655 19233
rect 33597 19224 33609 19227
rect 33152 19196 33609 19224
rect 25832 19184 25838 19196
rect 33597 19193 33609 19196
rect 33643 19193 33655 19227
rect 33597 19187 33655 19193
rect 16356 19128 17172 19156
rect 16356 19116 16362 19128
rect 18322 19116 18328 19168
rect 18380 19156 18386 19168
rect 19794 19156 19800 19168
rect 18380 19128 19800 19156
rect 18380 19116 18386 19128
rect 19794 19116 19800 19128
rect 19852 19116 19858 19168
rect 21726 19116 21732 19168
rect 21784 19156 21790 19168
rect 22189 19159 22247 19165
rect 22189 19156 22201 19159
rect 21784 19128 22201 19156
rect 21784 19116 21790 19128
rect 22189 19125 22201 19128
rect 22235 19125 22247 19159
rect 22189 19119 22247 19125
rect 24210 19116 24216 19168
rect 24268 19156 24274 19168
rect 26786 19156 26792 19168
rect 24268 19128 26792 19156
rect 24268 19116 24274 19128
rect 26786 19116 26792 19128
rect 26844 19116 26850 19168
rect 29638 19116 29644 19168
rect 29696 19116 29702 19168
rect 33134 19116 33140 19168
rect 33192 19156 33198 19168
rect 33704 19156 33732 19332
rect 33873 19329 33885 19332
rect 33919 19329 33931 19363
rect 33873 19323 33931 19329
rect 34146 19320 34152 19372
rect 34204 19320 34210 19372
rect 34440 19369 34468 19400
rect 34241 19363 34299 19369
rect 34241 19329 34253 19363
rect 34287 19360 34299 19363
rect 34425 19363 34483 19369
rect 34287 19332 34376 19360
rect 34287 19329 34299 19332
rect 34241 19323 34299 19329
rect 34348 19292 34376 19332
rect 34425 19329 34437 19363
rect 34471 19329 34483 19363
rect 34532 19360 34560 19468
rect 34790 19456 34796 19508
rect 34848 19456 34854 19508
rect 35989 19499 36047 19505
rect 35989 19465 36001 19499
rect 36035 19496 36047 19499
rect 36078 19496 36084 19508
rect 36035 19468 36084 19496
rect 36035 19465 36047 19468
rect 35989 19459 36047 19465
rect 36078 19456 36084 19468
rect 36136 19456 36142 19508
rect 34808 19428 34836 19456
rect 34808 19400 36032 19428
rect 34701 19363 34759 19369
rect 34701 19360 34713 19363
rect 34532 19332 34713 19360
rect 34425 19323 34483 19329
rect 34701 19329 34713 19332
rect 34747 19329 34759 19363
rect 34808 19360 34836 19400
rect 36004 19369 36032 19400
rect 34885 19363 34943 19369
rect 34885 19360 34897 19363
rect 34808 19332 34897 19360
rect 34701 19323 34759 19329
rect 34885 19329 34897 19332
rect 34931 19329 34943 19363
rect 35805 19363 35863 19369
rect 35805 19360 35817 19363
rect 34885 19323 34943 19329
rect 34992 19332 35817 19360
rect 34790 19292 34796 19304
rect 34348 19264 34796 19292
rect 34790 19252 34796 19264
rect 34848 19252 34854 19304
rect 34422 19184 34428 19236
rect 34480 19224 34486 19236
rect 34992 19224 35020 19332
rect 35805 19329 35817 19332
rect 35851 19329 35863 19363
rect 35805 19323 35863 19329
rect 35989 19363 36047 19369
rect 35989 19329 36001 19363
rect 36035 19329 36047 19363
rect 35989 19323 36047 19329
rect 34480 19196 35020 19224
rect 34480 19184 34486 19196
rect 33192 19128 33732 19156
rect 34609 19159 34667 19165
rect 33192 19116 33198 19128
rect 34609 19125 34621 19159
rect 34655 19156 34667 19159
rect 35986 19156 35992 19168
rect 34655 19128 35992 19156
rect 34655 19125 34667 19128
rect 34609 19119 34667 19125
rect 35986 19116 35992 19128
rect 36044 19116 36050 19168
rect 1104 19066 38272 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 38272 19066
rect 1104 18992 38272 19014
rect 4709 18955 4767 18961
rect 4709 18921 4721 18955
rect 4755 18952 4767 18955
rect 4798 18952 4804 18964
rect 4755 18924 4804 18952
rect 4755 18921 4767 18924
rect 4709 18915 4767 18921
rect 4798 18912 4804 18924
rect 4856 18912 4862 18964
rect 17218 18952 17224 18964
rect 5644 18924 17224 18952
rect 3329 18819 3387 18825
rect 3329 18785 3341 18819
rect 3375 18816 3387 18819
rect 4062 18816 4068 18828
rect 3375 18788 4068 18816
rect 3375 18785 3387 18788
rect 3329 18779 3387 18785
rect 4062 18776 4068 18788
rect 4120 18776 4126 18828
rect 3053 18751 3111 18757
rect 3053 18717 3065 18751
rect 3099 18748 3111 18751
rect 3142 18748 3148 18760
rect 3099 18720 3148 18748
rect 3099 18717 3111 18720
rect 3053 18711 3111 18717
rect 3142 18708 3148 18720
rect 3200 18708 3206 18760
rect 4893 18751 4951 18757
rect 4893 18717 4905 18751
rect 4939 18748 4951 18751
rect 5258 18748 5264 18760
rect 4939 18720 5264 18748
rect 4939 18717 4951 18720
rect 4893 18711 4951 18717
rect 5258 18708 5264 18720
rect 5316 18708 5322 18760
rect 5644 18748 5672 18924
rect 17218 18912 17224 18924
rect 17276 18912 17282 18964
rect 18046 18952 18052 18964
rect 17788 18924 18052 18952
rect 11146 18884 11152 18896
rect 9232 18856 11152 18884
rect 9232 18828 9260 18856
rect 11146 18844 11152 18856
rect 11204 18844 11210 18896
rect 13998 18844 14004 18896
rect 14056 18884 14062 18896
rect 17788 18884 17816 18924
rect 18046 18912 18052 18924
rect 18104 18952 18110 18964
rect 18230 18952 18236 18964
rect 18104 18924 18236 18952
rect 18104 18912 18110 18924
rect 18230 18912 18236 18924
rect 18288 18912 18294 18964
rect 18414 18912 18420 18964
rect 18472 18912 18478 18964
rect 19702 18912 19708 18964
rect 19760 18952 19766 18964
rect 19797 18955 19855 18961
rect 19797 18952 19809 18955
rect 19760 18924 19809 18952
rect 19760 18912 19766 18924
rect 19797 18921 19809 18924
rect 19843 18921 19855 18955
rect 19797 18915 19855 18921
rect 20714 18912 20720 18964
rect 20772 18952 20778 18964
rect 20809 18955 20867 18961
rect 20809 18952 20821 18955
rect 20772 18924 20821 18952
rect 20772 18912 20778 18924
rect 20809 18921 20821 18924
rect 20855 18921 20867 18955
rect 20809 18915 20867 18921
rect 20993 18955 21051 18961
rect 20993 18921 21005 18955
rect 21039 18952 21051 18955
rect 21082 18952 21088 18964
rect 21039 18924 21088 18952
rect 21039 18921 21051 18924
rect 20993 18915 21051 18921
rect 21082 18912 21088 18924
rect 21140 18912 21146 18964
rect 22094 18912 22100 18964
rect 22152 18952 22158 18964
rect 22462 18952 22468 18964
rect 22152 18924 22468 18952
rect 22152 18912 22158 18924
rect 22462 18912 22468 18924
rect 22520 18952 22526 18964
rect 22557 18955 22615 18961
rect 22557 18952 22569 18955
rect 22520 18924 22569 18952
rect 22520 18912 22526 18924
rect 22557 18921 22569 18924
rect 22603 18921 22615 18955
rect 22557 18915 22615 18921
rect 26786 18912 26792 18964
rect 26844 18952 26850 18964
rect 32858 18952 32864 18964
rect 26844 18924 32864 18952
rect 26844 18912 26850 18924
rect 32858 18912 32864 18924
rect 32916 18912 32922 18964
rect 32953 18955 33011 18961
rect 32953 18921 32965 18955
rect 32999 18952 33011 18955
rect 34422 18952 34428 18964
rect 32999 18924 34428 18952
rect 32999 18921 33011 18924
rect 32953 18915 33011 18921
rect 34422 18912 34428 18924
rect 34480 18912 34486 18964
rect 14056 18856 17816 18884
rect 17865 18887 17923 18893
rect 14056 18844 14062 18856
rect 17865 18853 17877 18887
rect 17911 18884 17923 18887
rect 18325 18887 18383 18893
rect 18325 18884 18337 18887
rect 17911 18856 18337 18884
rect 17911 18853 17923 18856
rect 17865 18847 17923 18853
rect 18325 18853 18337 18856
rect 18371 18853 18383 18887
rect 18325 18847 18383 18853
rect 5721 18819 5779 18825
rect 5721 18785 5733 18819
rect 5767 18816 5779 18819
rect 5902 18816 5908 18828
rect 5767 18788 5908 18816
rect 5767 18785 5779 18788
rect 5721 18779 5779 18785
rect 5902 18776 5908 18788
rect 5960 18776 5966 18828
rect 9214 18776 9220 18828
rect 9272 18776 9278 18828
rect 9858 18776 9864 18828
rect 9916 18816 9922 18828
rect 10870 18816 10876 18828
rect 9916 18788 10876 18816
rect 9916 18776 9922 18788
rect 10870 18776 10876 18788
rect 10928 18776 10934 18828
rect 11330 18776 11336 18828
rect 11388 18816 11394 18828
rect 15930 18816 15936 18828
rect 11388 18788 12204 18816
rect 11388 18776 11394 18788
rect 5552 18720 5672 18748
rect 934 18640 940 18692
rect 992 18680 998 18692
rect 1397 18683 1455 18689
rect 1397 18680 1409 18683
rect 992 18652 1409 18680
rect 992 18640 998 18652
rect 1397 18649 1409 18652
rect 1443 18649 1455 18683
rect 1397 18643 1455 18649
rect 1762 18640 1768 18692
rect 1820 18640 1826 18692
rect 5552 18680 5580 18720
rect 5994 18708 6000 18760
rect 6052 18708 6058 18760
rect 6089 18751 6147 18757
rect 6089 18717 6101 18751
rect 6135 18747 6147 18751
rect 10781 18751 10839 18757
rect 6196 18747 9076 18748
rect 6135 18720 9076 18747
rect 6135 18719 6224 18720
rect 6135 18717 6147 18719
rect 6089 18711 6147 18717
rect 3160 18652 5580 18680
rect 1946 18572 1952 18624
rect 2004 18612 2010 18624
rect 3160 18621 3188 18652
rect 5626 18640 5632 18692
rect 5684 18680 5690 18692
rect 5810 18680 5816 18692
rect 5684 18652 5816 18680
rect 5684 18640 5690 18652
rect 5810 18640 5816 18652
rect 5868 18680 5874 18692
rect 8846 18680 8852 18692
rect 5868 18652 8852 18680
rect 5868 18640 5874 18652
rect 8846 18640 8852 18652
rect 8904 18640 8910 18692
rect 9048 18680 9076 18720
rect 10781 18717 10793 18751
rect 10827 18748 10839 18751
rect 11422 18748 11428 18760
rect 10827 18720 11428 18748
rect 10827 18717 10839 18720
rect 10781 18711 10839 18717
rect 11422 18708 11428 18720
rect 11480 18708 11486 18760
rect 11790 18708 11796 18760
rect 11848 18708 11854 18760
rect 11882 18708 11888 18760
rect 11940 18708 11946 18760
rect 11977 18751 12035 18757
rect 11977 18717 11989 18751
rect 12023 18748 12035 18751
rect 12066 18748 12072 18760
rect 12023 18720 12072 18748
rect 12023 18717 12035 18720
rect 11977 18711 12035 18717
rect 12066 18708 12072 18720
rect 12124 18708 12130 18760
rect 12176 18757 12204 18788
rect 15672 18788 15936 18816
rect 15672 18760 15700 18788
rect 15930 18776 15936 18788
rect 15988 18816 15994 18828
rect 18432 18816 18460 18912
rect 18506 18844 18512 18896
rect 18564 18884 18570 18896
rect 21726 18884 21732 18896
rect 18564 18856 21732 18884
rect 18564 18844 18570 18856
rect 21726 18844 21732 18856
rect 21784 18844 21790 18896
rect 22005 18887 22063 18893
rect 22005 18853 22017 18887
rect 22051 18884 22063 18887
rect 25958 18884 25964 18896
rect 22051 18856 25964 18884
rect 22051 18853 22063 18856
rect 22005 18847 22063 18853
rect 25958 18844 25964 18856
rect 26016 18844 26022 18896
rect 33597 18887 33655 18893
rect 33597 18884 33609 18887
rect 30944 18856 33609 18884
rect 15988 18788 18460 18816
rect 15988 18776 15994 18788
rect 12161 18751 12219 18757
rect 12161 18717 12173 18751
rect 12207 18717 12219 18751
rect 12161 18711 12219 18717
rect 15654 18708 15660 18760
rect 15712 18708 15718 18760
rect 17126 18708 17132 18760
rect 17184 18748 17190 18760
rect 17184 18720 17632 18748
rect 17184 18708 17190 18720
rect 10689 18683 10747 18689
rect 9048 18652 10456 18680
rect 2685 18615 2743 18621
rect 2685 18612 2697 18615
rect 2004 18584 2697 18612
rect 2004 18572 2010 18584
rect 2685 18581 2697 18584
rect 2731 18581 2743 18615
rect 2685 18575 2743 18581
rect 3145 18615 3203 18621
rect 3145 18581 3157 18615
rect 3191 18581 3203 18615
rect 3145 18575 3203 18581
rect 4246 18572 4252 18624
rect 4304 18612 4310 18624
rect 6273 18615 6331 18621
rect 6273 18612 6285 18615
rect 4304 18584 6285 18612
rect 4304 18572 4310 18584
rect 6273 18581 6285 18584
rect 6319 18581 6331 18615
rect 6273 18575 6331 18581
rect 6546 18572 6552 18624
rect 6604 18612 6610 18624
rect 10042 18612 10048 18624
rect 6604 18584 10048 18612
rect 6604 18572 6610 18584
rect 10042 18572 10048 18584
rect 10100 18572 10106 18624
rect 10318 18572 10324 18624
rect 10376 18572 10382 18624
rect 10428 18612 10456 18652
rect 10689 18649 10701 18683
rect 10735 18680 10747 18683
rect 11517 18683 11575 18689
rect 11517 18680 11529 18683
rect 10735 18652 11529 18680
rect 10735 18649 10747 18652
rect 10689 18643 10747 18649
rect 11517 18649 11529 18652
rect 11563 18649 11575 18683
rect 14369 18683 14427 18689
rect 14369 18680 14381 18683
rect 11517 18643 11575 18649
rect 14108 18652 14381 18680
rect 13906 18612 13912 18624
rect 10428 18584 13912 18612
rect 13906 18572 13912 18584
rect 13964 18612 13970 18624
rect 14108 18612 14136 18652
rect 14369 18649 14381 18652
rect 14415 18649 14427 18683
rect 14369 18643 14427 18649
rect 14553 18683 14611 18689
rect 14553 18649 14565 18683
rect 14599 18680 14611 18683
rect 17034 18680 17040 18692
rect 14599 18652 17040 18680
rect 14599 18649 14611 18652
rect 14553 18643 14611 18649
rect 17034 18640 17040 18652
rect 17092 18640 17098 18692
rect 17604 18680 17632 18720
rect 17678 18708 17684 18760
rect 17736 18708 17742 18760
rect 18064 18757 18092 18788
rect 17957 18751 18015 18757
rect 17957 18717 17969 18751
rect 18003 18717 18015 18751
rect 17957 18711 18015 18717
rect 18049 18751 18107 18757
rect 18049 18717 18061 18751
rect 18095 18748 18107 18751
rect 18233 18751 18291 18757
rect 18095 18720 18129 18748
rect 18095 18717 18107 18720
rect 18049 18711 18107 18717
rect 18233 18717 18245 18751
rect 18279 18748 18291 18751
rect 18432 18748 18460 18788
rect 19334 18776 19340 18828
rect 19392 18776 19398 18828
rect 20165 18819 20223 18825
rect 20165 18816 20177 18819
rect 19536 18788 20177 18816
rect 18506 18748 18512 18760
rect 18279 18720 18368 18748
rect 18432 18720 18512 18748
rect 18279 18717 18291 18720
rect 18233 18711 18291 18717
rect 17972 18680 18000 18711
rect 18340 18689 18368 18720
rect 18506 18708 18512 18720
rect 18564 18708 18570 18760
rect 18601 18751 18659 18757
rect 18601 18717 18613 18751
rect 18647 18748 18659 18751
rect 18647 18720 18828 18748
rect 18647 18717 18659 18720
rect 18601 18711 18659 18717
rect 17604 18652 18000 18680
rect 18325 18683 18383 18689
rect 18325 18649 18337 18683
rect 18371 18680 18383 18683
rect 18690 18680 18696 18692
rect 18371 18652 18696 18680
rect 18371 18649 18383 18652
rect 18325 18643 18383 18649
rect 18690 18640 18696 18652
rect 18748 18640 18754 18692
rect 18800 18680 18828 18720
rect 18966 18708 18972 18760
rect 19024 18748 19030 18760
rect 19245 18751 19303 18757
rect 19245 18748 19257 18751
rect 19024 18720 19257 18748
rect 19024 18708 19030 18720
rect 19245 18717 19257 18720
rect 19291 18717 19303 18751
rect 19245 18711 19303 18717
rect 19426 18708 19432 18760
rect 19484 18748 19490 18760
rect 19536 18757 19564 18788
rect 20165 18785 20177 18788
rect 20211 18785 20223 18819
rect 20165 18779 20223 18785
rect 20441 18819 20499 18825
rect 20441 18785 20453 18819
rect 20487 18785 20499 18819
rect 20441 18779 20499 18785
rect 19521 18751 19579 18757
rect 19521 18748 19533 18751
rect 19484 18720 19533 18748
rect 19484 18708 19490 18720
rect 19521 18717 19533 18720
rect 19567 18717 19579 18751
rect 19521 18711 19579 18717
rect 19613 18751 19671 18757
rect 19613 18717 19625 18751
rect 19659 18748 19671 18751
rect 19702 18748 19708 18760
rect 19659 18720 19708 18748
rect 19659 18717 19671 18720
rect 19613 18711 19671 18717
rect 19628 18680 19656 18711
rect 19702 18708 19708 18720
rect 19760 18708 19766 18760
rect 19978 18748 19984 18760
rect 20036 18757 20042 18760
rect 19944 18720 19984 18748
rect 19978 18708 19984 18720
rect 20036 18711 20044 18757
rect 20456 18748 20484 18779
rect 20622 18776 20628 18828
rect 20680 18776 20686 18828
rect 20088 18720 20484 18748
rect 20533 18751 20591 18757
rect 20036 18708 20042 18711
rect 20088 18692 20116 18720
rect 20533 18717 20545 18751
rect 20579 18717 20591 18751
rect 20640 18748 20668 18776
rect 21545 18751 21603 18757
rect 21545 18748 21557 18751
rect 20640 18720 21557 18748
rect 20533 18711 20591 18717
rect 21545 18717 21557 18720
rect 21591 18717 21603 18751
rect 21545 18711 21603 18717
rect 18800 18652 19656 18680
rect 18800 18624 18828 18652
rect 20070 18640 20076 18692
rect 20128 18640 20134 18692
rect 20548 18680 20576 18711
rect 21634 18708 21640 18760
rect 21692 18708 21698 18760
rect 20364 18652 20576 18680
rect 20364 18624 20392 18652
rect 21174 18640 21180 18692
rect 21232 18640 21238 18692
rect 21744 18680 21772 18844
rect 21821 18819 21879 18825
rect 21821 18785 21833 18819
rect 21867 18816 21879 18819
rect 22649 18819 22707 18825
rect 22649 18816 22661 18819
rect 21867 18788 22661 18816
rect 21867 18785 21879 18788
rect 21821 18779 21879 18785
rect 22649 18785 22661 18788
rect 22695 18816 22707 18819
rect 23474 18816 23480 18828
rect 22695 18788 23480 18816
rect 22695 18785 22707 18788
rect 22649 18779 22707 18785
rect 23474 18776 23480 18788
rect 23532 18776 23538 18828
rect 22370 18708 22376 18760
rect 22428 18708 22434 18760
rect 27338 18708 27344 18760
rect 27396 18748 27402 18760
rect 30944 18748 30972 18856
rect 33597 18853 33609 18856
rect 33643 18853 33655 18887
rect 33597 18847 33655 18853
rect 33134 18816 33140 18828
rect 31036 18788 31616 18816
rect 31036 18757 31064 18788
rect 27396 18720 30972 18748
rect 31021 18751 31079 18757
rect 27396 18708 27402 18720
rect 31021 18717 31033 18751
rect 31067 18717 31079 18751
rect 31021 18711 31079 18717
rect 24670 18680 24676 18692
rect 21744 18652 24676 18680
rect 24670 18640 24676 18652
rect 24728 18680 24734 18692
rect 25682 18680 25688 18692
rect 24728 18652 25688 18680
rect 24728 18640 24734 18652
rect 25682 18640 25688 18652
rect 25740 18640 25746 18692
rect 30742 18640 30748 18692
rect 30800 18680 30806 18692
rect 31036 18680 31064 18711
rect 31202 18708 31208 18760
rect 31260 18708 31266 18760
rect 31386 18708 31392 18760
rect 31444 18708 31450 18760
rect 31588 18757 31616 18788
rect 32508 18788 33140 18816
rect 32508 18757 32536 18788
rect 33134 18776 33140 18788
rect 33192 18776 33198 18828
rect 35342 18816 35348 18828
rect 34716 18788 35348 18816
rect 31573 18751 31631 18757
rect 31573 18717 31585 18751
rect 31619 18717 31631 18751
rect 31573 18711 31631 18717
rect 32401 18751 32459 18757
rect 32401 18717 32413 18751
rect 32447 18717 32459 18751
rect 32401 18711 32459 18717
rect 32493 18751 32551 18757
rect 32493 18717 32505 18751
rect 32539 18717 32551 18751
rect 32493 18711 32551 18717
rect 30800 18652 31064 18680
rect 31481 18683 31539 18689
rect 30800 18640 30806 18652
rect 31481 18649 31493 18683
rect 31527 18680 31539 18683
rect 32416 18680 32444 18711
rect 32674 18708 32680 18760
rect 32732 18708 32738 18760
rect 32766 18708 32772 18760
rect 32824 18708 32830 18760
rect 33042 18708 33048 18760
rect 33100 18748 33106 18760
rect 33689 18751 33747 18757
rect 33100 18720 33272 18748
rect 33100 18708 33106 18720
rect 33244 18680 33272 18720
rect 33689 18717 33701 18751
rect 33735 18748 33747 18751
rect 33962 18748 33968 18760
rect 33735 18720 33968 18748
rect 33735 18717 33747 18720
rect 33689 18711 33747 18717
rect 33962 18708 33968 18720
rect 34020 18708 34026 18760
rect 34716 18689 34744 18788
rect 35342 18776 35348 18788
rect 35400 18776 35406 18828
rect 36722 18776 36728 18828
rect 36780 18776 36786 18828
rect 34977 18751 35035 18757
rect 34977 18717 34989 18751
rect 35023 18748 35035 18751
rect 36909 18751 36967 18757
rect 36909 18748 36921 18751
rect 35023 18720 35204 18748
rect 35023 18717 35035 18720
rect 34977 18711 35035 18717
rect 34701 18683 34759 18689
rect 34701 18680 34713 18683
rect 31527 18652 33180 18680
rect 33244 18652 34713 18680
rect 31527 18649 31539 18652
rect 31481 18643 31539 18649
rect 33152 18624 33180 18652
rect 34701 18649 34713 18652
rect 34747 18649 34759 18683
rect 34701 18643 34759 18649
rect 35176 18624 35204 18720
rect 36832 18720 36921 18748
rect 36832 18692 36860 18720
rect 36909 18717 36921 18720
rect 36955 18717 36967 18751
rect 36909 18711 36967 18717
rect 36814 18640 36820 18692
rect 36872 18640 36878 18692
rect 13964 18584 14136 18612
rect 13964 18572 13970 18584
rect 14182 18572 14188 18624
rect 14240 18572 14246 18624
rect 16206 18572 16212 18624
rect 16264 18612 16270 18624
rect 17497 18615 17555 18621
rect 17497 18612 17509 18615
rect 16264 18584 17509 18612
rect 16264 18572 16270 18584
rect 17497 18581 17509 18584
rect 17543 18581 17555 18615
rect 17497 18575 17555 18581
rect 18046 18572 18052 18624
rect 18104 18572 18110 18624
rect 18782 18572 18788 18624
rect 18840 18572 18846 18624
rect 20346 18572 20352 18624
rect 20404 18572 20410 18624
rect 20622 18572 20628 18624
rect 20680 18612 20686 18624
rect 20967 18615 21025 18621
rect 20967 18612 20979 18615
rect 20680 18584 20979 18612
rect 20680 18572 20686 18584
rect 20967 18581 20979 18584
rect 21013 18581 21025 18615
rect 20967 18575 21025 18581
rect 22186 18572 22192 18624
rect 22244 18572 22250 18624
rect 25130 18572 25136 18624
rect 25188 18612 25194 18624
rect 25958 18612 25964 18624
rect 25188 18584 25964 18612
rect 25188 18572 25194 18584
rect 25958 18572 25964 18584
rect 26016 18612 26022 18624
rect 28350 18612 28356 18624
rect 26016 18584 28356 18612
rect 26016 18572 26022 18584
rect 28350 18572 28356 18584
rect 28408 18612 28414 18624
rect 30926 18612 30932 18624
rect 28408 18584 30932 18612
rect 28408 18572 28414 18584
rect 30926 18572 30932 18584
rect 30984 18572 30990 18624
rect 31202 18572 31208 18624
rect 31260 18572 31266 18624
rect 32306 18572 32312 18624
rect 32364 18612 32370 18624
rect 33042 18612 33048 18624
rect 32364 18584 33048 18612
rect 32364 18572 32370 18584
rect 33042 18572 33048 18584
rect 33100 18572 33106 18624
rect 33134 18572 33140 18624
rect 33192 18572 33198 18624
rect 34790 18572 34796 18624
rect 34848 18621 34854 18624
rect 34848 18575 34857 18621
rect 34885 18615 34943 18621
rect 34885 18581 34897 18615
rect 34931 18612 34943 18615
rect 34974 18612 34980 18624
rect 34931 18584 34980 18612
rect 34931 18581 34943 18584
rect 34885 18575 34943 18581
rect 34848 18572 34854 18575
rect 34974 18572 34980 18584
rect 35032 18572 35038 18624
rect 35158 18572 35164 18624
rect 35216 18572 35222 18624
rect 37090 18572 37096 18624
rect 37148 18572 37154 18624
rect 1104 18522 38272 18544
rect 1104 18470 4874 18522
rect 4926 18470 4938 18522
rect 4990 18470 5002 18522
rect 5054 18470 5066 18522
rect 5118 18470 5130 18522
rect 5182 18470 35594 18522
rect 35646 18470 35658 18522
rect 35710 18470 35722 18522
rect 35774 18470 35786 18522
rect 35838 18470 35850 18522
rect 35902 18470 38272 18522
rect 1104 18448 38272 18470
rect 4246 18408 4252 18420
rect 2332 18380 4252 18408
rect 2332 18281 2360 18380
rect 4246 18368 4252 18380
rect 4304 18368 4310 18420
rect 13814 18408 13820 18420
rect 4356 18380 9536 18408
rect 4356 18349 4384 18380
rect 4341 18343 4399 18349
rect 4341 18309 4353 18343
rect 4387 18309 4399 18343
rect 4341 18303 4399 18309
rect 8294 18300 8300 18352
rect 8352 18300 8358 18352
rect 9508 18349 9536 18380
rect 10796 18380 13820 18408
rect 9493 18343 9551 18349
rect 9493 18309 9505 18343
rect 9539 18340 9551 18343
rect 10226 18340 10232 18352
rect 9539 18312 10232 18340
rect 9539 18309 9551 18312
rect 9493 18303 9551 18309
rect 10226 18300 10232 18312
rect 10284 18300 10290 18352
rect 1857 18275 1915 18281
rect 1857 18241 1869 18275
rect 1903 18272 1915 18275
rect 2317 18275 2375 18281
rect 1903 18244 2268 18272
rect 1903 18241 1915 18244
rect 1857 18235 1915 18241
rect 1670 18164 1676 18216
rect 1728 18204 1734 18216
rect 2133 18207 2191 18213
rect 2133 18204 2145 18207
rect 1728 18176 2145 18204
rect 1728 18164 1734 18176
rect 2133 18173 2145 18176
rect 2179 18173 2191 18207
rect 2240 18204 2268 18244
rect 2317 18241 2329 18275
rect 2363 18241 2375 18275
rect 2317 18235 2375 18241
rect 6181 18275 6239 18281
rect 6181 18241 6193 18275
rect 6227 18272 6239 18275
rect 6546 18272 6552 18284
rect 6227 18244 6552 18272
rect 6227 18241 6239 18244
rect 6181 18235 6239 18241
rect 6546 18232 6552 18244
rect 6604 18232 6610 18284
rect 4062 18204 4068 18216
rect 2240 18176 4068 18204
rect 2133 18167 2191 18173
rect 2148 18136 2176 18167
rect 4062 18164 4068 18176
rect 4120 18164 4126 18216
rect 5902 18164 5908 18216
rect 5960 18164 5966 18216
rect 6638 18204 6644 18216
rect 6196 18176 6644 18204
rect 3418 18136 3424 18148
rect 2148 18108 3424 18136
rect 3418 18096 3424 18108
rect 3476 18136 3482 18148
rect 3694 18136 3700 18148
rect 3476 18108 3700 18136
rect 3476 18096 3482 18108
rect 3694 18096 3700 18108
rect 3752 18096 3758 18148
rect 6196 18080 6224 18176
rect 6638 18164 6644 18176
rect 6696 18204 6702 18216
rect 7561 18207 7619 18213
rect 7561 18204 7573 18207
rect 6696 18176 7573 18204
rect 6696 18164 6702 18176
rect 7561 18173 7573 18176
rect 7607 18173 7619 18207
rect 7561 18167 7619 18173
rect 7837 18207 7895 18213
rect 7837 18173 7849 18207
rect 7883 18204 7895 18207
rect 7926 18204 7932 18216
rect 7883 18176 7932 18204
rect 7883 18173 7895 18176
rect 7837 18167 7895 18173
rect 2038 18028 2044 18080
rect 2096 18028 2102 18080
rect 2498 18028 2504 18080
rect 2556 18028 2562 18080
rect 2958 18028 2964 18080
rect 3016 18068 3022 18080
rect 3053 18071 3111 18077
rect 3053 18068 3065 18071
rect 3016 18040 3065 18068
rect 3016 18028 3022 18040
rect 3053 18037 3065 18040
rect 3099 18068 3111 18071
rect 3510 18068 3516 18080
rect 3099 18040 3516 18068
rect 3099 18037 3111 18040
rect 3053 18031 3111 18037
rect 3510 18028 3516 18040
rect 3568 18028 3574 18080
rect 6178 18028 6184 18080
rect 6236 18028 6242 18080
rect 7576 18068 7604 18167
rect 7926 18164 7932 18176
rect 7984 18164 7990 18216
rect 9030 18164 9036 18216
rect 9088 18204 9094 18216
rect 9309 18207 9367 18213
rect 9309 18204 9321 18207
rect 9088 18176 9321 18204
rect 9088 18164 9094 18176
rect 9309 18173 9321 18176
rect 9355 18173 9367 18207
rect 9309 18167 9367 18173
rect 10796 18145 10824 18380
rect 13814 18368 13820 18380
rect 13872 18368 13878 18420
rect 13906 18368 13912 18420
rect 13964 18368 13970 18420
rect 14182 18368 14188 18420
rect 14240 18368 14246 18420
rect 15378 18368 15384 18420
rect 15436 18368 15442 18420
rect 18506 18368 18512 18420
rect 18564 18408 18570 18420
rect 18564 18380 18920 18408
rect 18564 18368 18570 18380
rect 12069 18343 12127 18349
rect 12069 18309 12081 18343
rect 12115 18340 12127 18343
rect 12250 18340 12256 18352
rect 12115 18312 12256 18340
rect 12115 18309 12127 18312
rect 12069 18303 12127 18309
rect 12250 18300 12256 18312
rect 12308 18300 12314 18352
rect 14200 18340 14228 18368
rect 15013 18343 15071 18349
rect 14200 18312 14504 18340
rect 11330 18232 11336 18284
rect 11388 18272 11394 18284
rect 11517 18275 11575 18281
rect 11517 18272 11529 18275
rect 11388 18244 11529 18272
rect 11388 18232 11394 18244
rect 11517 18241 11529 18244
rect 11563 18241 11575 18275
rect 11517 18235 11575 18241
rect 11701 18275 11759 18281
rect 11701 18241 11713 18275
rect 11747 18241 11759 18275
rect 11701 18235 11759 18241
rect 12345 18275 12403 18281
rect 12345 18241 12357 18275
rect 12391 18241 12403 18275
rect 12345 18235 12403 18241
rect 11422 18164 11428 18216
rect 11480 18204 11486 18216
rect 11716 18204 11744 18235
rect 11480 18176 11744 18204
rect 11480 18164 11486 18176
rect 12066 18164 12072 18216
rect 12124 18204 12130 18216
rect 12161 18207 12219 18213
rect 12161 18204 12173 18207
rect 12124 18176 12173 18204
rect 12124 18164 12130 18176
rect 12161 18173 12173 18176
rect 12207 18173 12219 18207
rect 12161 18167 12219 18173
rect 10781 18139 10839 18145
rect 10781 18136 10793 18139
rect 8864 18108 10793 18136
rect 8864 18068 8892 18108
rect 10781 18105 10793 18108
rect 10827 18105 10839 18139
rect 10781 18099 10839 18105
rect 11146 18096 11152 18148
rect 11204 18136 11210 18148
rect 11701 18139 11759 18145
rect 11701 18136 11713 18139
rect 11204 18108 11713 18136
rect 11204 18096 11210 18108
rect 11701 18105 11713 18108
rect 11747 18105 11759 18139
rect 12360 18136 12388 18235
rect 12526 18232 12532 18284
rect 12584 18232 12590 18284
rect 13814 18232 13820 18284
rect 13872 18272 13878 18284
rect 14093 18275 14151 18281
rect 14093 18272 14105 18275
rect 13872 18244 14105 18272
rect 13872 18232 13878 18244
rect 14093 18241 14105 18244
rect 14139 18241 14151 18275
rect 14093 18235 14151 18241
rect 14274 18232 14280 18284
rect 14332 18232 14338 18284
rect 14476 18281 14504 18312
rect 15013 18309 15025 18343
rect 15059 18340 15071 18343
rect 15102 18340 15108 18352
rect 15059 18312 15108 18340
rect 15059 18309 15071 18312
rect 15013 18303 15071 18309
rect 15102 18300 15108 18312
rect 15160 18300 15166 18352
rect 18892 18284 18920 18380
rect 19702 18368 19708 18420
rect 19760 18408 19766 18420
rect 19889 18411 19947 18417
rect 19889 18408 19901 18411
rect 19760 18380 19901 18408
rect 19760 18368 19766 18380
rect 19889 18377 19901 18380
rect 19935 18377 19947 18411
rect 19889 18371 19947 18377
rect 20162 18368 20168 18420
rect 20220 18408 20226 18420
rect 25593 18411 25651 18417
rect 20220 18380 22232 18408
rect 20220 18368 20226 18380
rect 22204 18340 22232 18380
rect 25593 18377 25605 18411
rect 25639 18408 25651 18411
rect 30742 18408 30748 18420
rect 25639 18380 30748 18408
rect 25639 18377 25651 18380
rect 25593 18371 25651 18377
rect 30742 18368 30748 18380
rect 30800 18408 30806 18420
rect 30800 18380 30972 18408
rect 30800 18368 30806 18380
rect 22646 18340 22652 18352
rect 19168 18312 20024 18340
rect 22204 18312 22652 18340
rect 14461 18275 14519 18281
rect 14461 18241 14473 18275
rect 14507 18241 14519 18275
rect 15657 18275 15715 18281
rect 15657 18272 15669 18275
rect 14461 18235 14519 18241
rect 15396 18244 15669 18272
rect 15396 18216 15424 18244
rect 15657 18241 15669 18244
rect 15703 18272 15715 18275
rect 16114 18272 16120 18284
rect 15703 18244 16120 18272
rect 15703 18241 15715 18244
rect 15657 18235 15715 18241
rect 16114 18232 16120 18244
rect 16172 18232 16178 18284
rect 16482 18232 16488 18284
rect 16540 18272 16546 18284
rect 16758 18272 16764 18284
rect 16540 18244 16764 18272
rect 16540 18232 16546 18244
rect 16758 18232 16764 18244
rect 16816 18232 16822 18284
rect 16942 18232 16948 18284
rect 17000 18272 17006 18284
rect 17129 18275 17187 18281
rect 17129 18272 17141 18275
rect 17000 18244 17141 18272
rect 17000 18232 17006 18244
rect 17129 18241 17141 18244
rect 17175 18241 17187 18275
rect 17129 18235 17187 18241
rect 18230 18232 18236 18284
rect 18288 18272 18294 18284
rect 18785 18275 18843 18281
rect 18785 18272 18797 18275
rect 18288 18244 18797 18272
rect 18288 18232 18294 18244
rect 18785 18241 18797 18244
rect 18831 18241 18843 18275
rect 18785 18235 18843 18241
rect 18874 18232 18880 18284
rect 18932 18232 18938 18284
rect 19168 18281 19196 18312
rect 19996 18284 20024 18312
rect 22646 18300 22652 18312
rect 22704 18300 22710 18352
rect 25222 18340 25228 18352
rect 24964 18312 25228 18340
rect 24964 18284 24992 18312
rect 25222 18300 25228 18312
rect 25280 18300 25286 18352
rect 27614 18300 27620 18352
rect 27672 18340 27678 18352
rect 27672 18312 28212 18340
rect 27672 18300 27678 18312
rect 19168 18275 19245 18281
rect 19168 18244 19199 18275
rect 19187 18241 19199 18244
rect 19233 18241 19245 18275
rect 19187 18235 19245 18241
rect 19521 18275 19579 18281
rect 19521 18241 19533 18275
rect 19567 18241 19579 18275
rect 19521 18235 19579 18241
rect 19675 18275 19733 18281
rect 19675 18241 19687 18275
rect 19721 18272 19733 18275
rect 19794 18272 19800 18284
rect 19721 18244 19800 18272
rect 19721 18241 19733 18244
rect 19675 18235 19733 18241
rect 15378 18164 15384 18216
rect 15436 18164 15442 18216
rect 15565 18207 15623 18213
rect 15565 18173 15577 18207
rect 15611 18204 15623 18207
rect 15746 18204 15752 18216
rect 15611 18176 15752 18204
rect 15611 18173 15623 18176
rect 15565 18167 15623 18173
rect 15746 18164 15752 18176
rect 15804 18164 15810 18216
rect 15930 18164 15936 18216
rect 15988 18204 15994 18216
rect 16025 18207 16083 18213
rect 16025 18204 16037 18207
rect 15988 18176 16037 18204
rect 15988 18164 15994 18176
rect 16025 18173 16037 18176
rect 16071 18173 16083 18207
rect 19536 18204 19564 18235
rect 19794 18232 19800 18244
rect 19852 18232 19858 18284
rect 19978 18232 19984 18284
rect 20036 18232 20042 18284
rect 20530 18232 20536 18284
rect 20588 18232 20594 18284
rect 22370 18232 22376 18284
rect 22428 18232 22434 18284
rect 22462 18232 22468 18284
rect 22520 18232 22526 18284
rect 22554 18232 22560 18284
rect 22612 18272 22618 18284
rect 22741 18275 22799 18281
rect 22741 18272 22753 18275
rect 22612 18244 22753 18272
rect 22612 18232 22618 18244
rect 22741 18241 22753 18244
rect 22787 18241 22799 18275
rect 22741 18235 22799 18241
rect 23293 18275 23351 18281
rect 23293 18241 23305 18275
rect 23339 18272 23351 18275
rect 23566 18272 23572 18284
rect 23339 18244 23572 18272
rect 23339 18241 23351 18244
rect 23293 18235 23351 18241
rect 23566 18232 23572 18244
rect 23624 18232 23630 18284
rect 24946 18232 24952 18284
rect 25004 18232 25010 18284
rect 25038 18232 25044 18284
rect 25096 18232 25102 18284
rect 25317 18275 25375 18281
rect 25317 18241 25329 18275
rect 25363 18241 25375 18275
rect 25317 18235 25375 18241
rect 25409 18275 25467 18281
rect 25409 18241 25421 18275
rect 25455 18272 25467 18275
rect 25590 18272 25596 18284
rect 25455 18244 25596 18272
rect 25455 18241 25467 18244
rect 25409 18235 25467 18241
rect 20548 18204 20576 18232
rect 19536 18176 20576 18204
rect 22388 18204 22416 18232
rect 22925 18207 22983 18213
rect 22925 18204 22937 18207
rect 22388 18176 22937 18204
rect 16025 18167 16083 18173
rect 22925 18173 22937 18176
rect 22971 18173 22983 18207
rect 22925 18167 22983 18173
rect 23658 18164 23664 18216
rect 23716 18204 23722 18216
rect 25332 18204 25360 18235
rect 23716 18176 25360 18204
rect 23716 18164 23722 18176
rect 11701 18099 11759 18105
rect 12084 18108 12388 18136
rect 12084 18080 12112 18108
rect 19426 18096 19432 18148
rect 19484 18096 19490 18148
rect 23569 18139 23627 18145
rect 19536 18108 20392 18136
rect 7576 18040 8892 18068
rect 8938 18028 8944 18080
rect 8996 18068 9002 18080
rect 10502 18068 10508 18080
rect 8996 18040 10508 18068
rect 8996 18028 9002 18040
rect 10502 18028 10508 18040
rect 10560 18028 10566 18080
rect 11054 18028 11060 18080
rect 11112 18068 11118 18080
rect 11514 18068 11520 18080
rect 11112 18040 11520 18068
rect 11112 18028 11118 18040
rect 11514 18028 11520 18040
rect 11572 18068 11578 18080
rect 12066 18068 12072 18080
rect 11572 18040 12072 18068
rect 11572 18028 11578 18040
rect 12066 18028 12072 18040
rect 12124 18028 12130 18080
rect 12710 18028 12716 18080
rect 12768 18068 12774 18080
rect 14182 18068 14188 18080
rect 12768 18040 14188 18068
rect 12768 18028 12774 18040
rect 14182 18028 14188 18040
rect 14240 18028 14246 18080
rect 17954 18028 17960 18080
rect 18012 18068 18018 18080
rect 18417 18071 18475 18077
rect 18417 18068 18429 18071
rect 18012 18040 18429 18068
rect 18012 18028 18018 18040
rect 18417 18037 18429 18040
rect 18463 18068 18475 18071
rect 18506 18068 18512 18080
rect 18463 18040 18512 18068
rect 18463 18037 18475 18040
rect 18417 18031 18475 18037
rect 18506 18028 18512 18040
rect 18564 18028 18570 18080
rect 18598 18028 18604 18080
rect 18656 18068 18662 18080
rect 19245 18071 19303 18077
rect 19245 18068 19257 18071
rect 18656 18040 19257 18068
rect 18656 18028 18662 18040
rect 19245 18037 19257 18040
rect 19291 18068 19303 18071
rect 19536 18068 19564 18108
rect 20364 18080 20392 18108
rect 23569 18105 23581 18139
rect 23615 18105 23627 18139
rect 23569 18099 23627 18105
rect 19291 18040 19564 18068
rect 19291 18037 19303 18040
rect 19245 18031 19303 18037
rect 19978 18028 19984 18080
rect 20036 18068 20042 18080
rect 20254 18068 20260 18080
rect 20036 18040 20260 18068
rect 20036 18028 20042 18040
rect 20254 18028 20260 18040
rect 20312 18028 20318 18080
rect 20346 18028 20352 18080
rect 20404 18028 20410 18080
rect 20438 18028 20444 18080
rect 20496 18068 20502 18080
rect 21542 18068 21548 18080
rect 20496 18040 21548 18068
rect 20496 18028 20502 18040
rect 21542 18028 21548 18040
rect 21600 18028 21606 18080
rect 23584 18068 23612 18099
rect 23842 18096 23848 18148
rect 23900 18136 23906 18148
rect 25424 18136 25452 18235
rect 25590 18232 25596 18244
rect 25648 18232 25654 18284
rect 25869 18275 25927 18281
rect 25869 18241 25881 18275
rect 25915 18272 25927 18275
rect 25958 18272 25964 18284
rect 25915 18244 25964 18272
rect 25915 18241 25927 18244
rect 25869 18235 25927 18241
rect 25958 18232 25964 18244
rect 26016 18232 26022 18284
rect 27982 18232 27988 18284
rect 28040 18232 28046 18284
rect 28184 18281 28212 18312
rect 30300 18312 30696 18340
rect 30300 18284 30328 18312
rect 28169 18275 28227 18281
rect 28169 18241 28181 18275
rect 28215 18272 28227 18275
rect 28626 18272 28632 18284
rect 28215 18244 28632 18272
rect 28215 18241 28227 18244
rect 28169 18235 28227 18241
rect 28626 18232 28632 18244
rect 28684 18232 28690 18284
rect 29362 18232 29368 18284
rect 29420 18272 29426 18284
rect 29546 18272 29552 18284
rect 29420 18244 29552 18272
rect 29420 18232 29426 18244
rect 29546 18232 29552 18244
rect 29604 18232 29610 18284
rect 29733 18275 29791 18281
rect 29733 18241 29745 18275
rect 29779 18272 29791 18275
rect 29779 18244 29868 18272
rect 29779 18241 29791 18244
rect 29733 18235 29791 18241
rect 25774 18164 25780 18216
rect 25832 18164 25838 18216
rect 23900 18108 25452 18136
rect 23900 18096 23906 18108
rect 26234 18096 26240 18148
rect 26292 18096 26298 18148
rect 28442 18096 28448 18148
rect 28500 18136 28506 18148
rect 29840 18136 29868 18244
rect 30282 18232 30288 18284
rect 30340 18232 30346 18284
rect 30374 18232 30380 18284
rect 30432 18232 30438 18284
rect 30668 18281 30696 18312
rect 30834 18300 30840 18352
rect 30892 18300 30898 18352
rect 30944 18340 30972 18380
rect 31202 18368 31208 18420
rect 31260 18408 31266 18420
rect 32769 18411 32827 18417
rect 31260 18380 31754 18408
rect 31260 18368 31266 18380
rect 31021 18343 31079 18349
rect 31021 18340 31033 18343
rect 30944 18312 31033 18340
rect 31021 18309 31033 18312
rect 31067 18309 31079 18343
rect 31726 18340 31754 18380
rect 32769 18377 32781 18411
rect 32815 18408 32827 18411
rect 34146 18408 34152 18420
rect 32815 18380 34152 18408
rect 32815 18377 32827 18380
rect 32769 18371 32827 18377
rect 34146 18368 34152 18380
rect 34204 18408 34210 18420
rect 34241 18411 34299 18417
rect 34241 18408 34253 18411
rect 34204 18380 34253 18408
rect 34204 18368 34210 18380
rect 34241 18377 34253 18380
rect 34287 18377 34299 18411
rect 34241 18371 34299 18377
rect 34790 18368 34796 18420
rect 34848 18368 34854 18420
rect 37090 18368 37096 18420
rect 37148 18368 37154 18420
rect 32125 18343 32183 18349
rect 32125 18340 32137 18343
rect 31021 18303 31079 18309
rect 31680 18312 32137 18340
rect 30653 18275 30711 18281
rect 30653 18241 30665 18275
rect 30699 18241 30711 18275
rect 30852 18272 30880 18300
rect 31205 18275 31263 18281
rect 31205 18272 31217 18275
rect 30852 18244 31217 18272
rect 30653 18235 30711 18241
rect 31205 18241 31217 18244
rect 31251 18272 31263 18275
rect 31294 18272 31300 18284
rect 31251 18244 31300 18272
rect 31251 18241 31263 18244
rect 31205 18235 31263 18241
rect 31294 18232 31300 18244
rect 31352 18232 31358 18284
rect 31680 18281 31708 18312
rect 32125 18309 32137 18312
rect 32171 18309 32183 18343
rect 32674 18340 32680 18352
rect 32125 18303 32183 18309
rect 32324 18312 32680 18340
rect 31389 18275 31447 18281
rect 31389 18241 31401 18275
rect 31435 18272 31447 18275
rect 31481 18275 31539 18281
rect 31481 18272 31493 18275
rect 31435 18244 31493 18272
rect 31435 18241 31447 18244
rect 31389 18235 31447 18241
rect 31481 18241 31493 18244
rect 31527 18241 31539 18275
rect 31481 18235 31539 18241
rect 31665 18275 31723 18281
rect 31665 18241 31677 18275
rect 31711 18241 31723 18275
rect 32324 18272 32352 18312
rect 32674 18300 32680 18312
rect 32732 18340 32738 18352
rect 32953 18343 33011 18349
rect 32953 18340 32965 18343
rect 32732 18312 32965 18340
rect 32732 18300 32738 18312
rect 32953 18309 32965 18312
rect 32999 18309 33011 18343
rect 32953 18303 33011 18309
rect 33134 18300 33140 18352
rect 33192 18300 33198 18352
rect 34072 18312 34744 18340
rect 31665 18235 31723 18241
rect 31956 18244 32352 18272
rect 28500 18108 29868 18136
rect 30300 18136 30328 18232
rect 31956 18216 31984 18244
rect 32766 18232 32772 18284
rect 32824 18272 32830 18284
rect 32861 18275 32919 18281
rect 32861 18272 32873 18275
rect 32824 18244 32873 18272
rect 32824 18232 32830 18244
rect 32861 18241 32873 18244
rect 32907 18241 32919 18275
rect 32861 18235 32919 18241
rect 30466 18164 30472 18216
rect 30524 18204 30530 18216
rect 31110 18204 31116 18216
rect 30524 18176 31116 18204
rect 30524 18164 30530 18176
rect 31110 18164 31116 18176
rect 31168 18164 31174 18216
rect 31849 18207 31907 18213
rect 31849 18173 31861 18207
rect 31895 18204 31907 18207
rect 31938 18204 31944 18216
rect 31895 18176 31944 18204
rect 31895 18173 31907 18176
rect 31849 18167 31907 18173
rect 31938 18164 31944 18176
rect 31996 18164 32002 18216
rect 32490 18164 32496 18216
rect 32548 18164 32554 18216
rect 32582 18164 32588 18216
rect 32640 18164 32646 18216
rect 34072 18213 34100 18312
rect 34333 18275 34391 18281
rect 34333 18241 34345 18275
rect 34379 18241 34391 18275
rect 34333 18235 34391 18241
rect 34057 18207 34115 18213
rect 34057 18204 34069 18207
rect 33060 18176 34069 18204
rect 31478 18136 31484 18148
rect 30300 18108 31484 18136
rect 28500 18096 28506 18108
rect 26510 18068 26516 18080
rect 23584 18040 26516 18068
rect 26510 18028 26516 18040
rect 26568 18028 26574 18080
rect 27890 18028 27896 18080
rect 27948 18068 27954 18080
rect 28077 18071 28135 18077
rect 28077 18068 28089 18071
rect 27948 18040 28089 18068
rect 27948 18028 27954 18040
rect 28077 18037 28089 18040
rect 28123 18037 28135 18071
rect 28077 18031 28135 18037
rect 29454 18028 29460 18080
rect 29512 18068 29518 18080
rect 29549 18071 29607 18077
rect 29549 18068 29561 18071
rect 29512 18040 29561 18068
rect 29512 18028 29518 18040
rect 29549 18037 29561 18040
rect 29595 18037 29607 18071
rect 29840 18068 29868 18108
rect 31478 18096 31484 18108
rect 31536 18136 31542 18148
rect 33060 18136 33088 18176
rect 34057 18173 34069 18176
rect 34103 18173 34115 18207
rect 34057 18167 34115 18173
rect 31536 18108 33088 18136
rect 33137 18139 33195 18145
rect 31536 18096 31542 18108
rect 33137 18105 33149 18139
rect 33183 18136 33195 18139
rect 34348 18136 34376 18235
rect 34716 18204 34744 18312
rect 34808 18281 34836 18368
rect 35434 18340 35440 18352
rect 35084 18312 35440 18340
rect 34793 18275 34851 18281
rect 34793 18241 34805 18275
rect 34839 18241 34851 18275
rect 34793 18235 34851 18241
rect 34974 18232 34980 18284
rect 35032 18232 35038 18284
rect 35084 18204 35112 18312
rect 35434 18300 35440 18312
rect 35492 18300 35498 18352
rect 35158 18232 35164 18284
rect 35216 18232 35222 18284
rect 36909 18275 36967 18281
rect 36909 18241 36921 18275
rect 36955 18272 36967 18275
rect 37108 18272 37136 18368
rect 37274 18300 37280 18352
rect 37332 18340 37338 18352
rect 37553 18343 37611 18349
rect 37553 18340 37565 18343
rect 37332 18312 37565 18340
rect 37332 18300 37338 18312
rect 37553 18309 37565 18312
rect 37599 18309 37611 18343
rect 37553 18303 37611 18309
rect 36955 18244 37136 18272
rect 36955 18241 36967 18244
rect 36909 18235 36967 18241
rect 34716 18176 35112 18204
rect 33183 18108 34376 18136
rect 34701 18139 34759 18145
rect 33183 18105 33195 18108
rect 33137 18099 33195 18105
rect 34701 18105 34713 18139
rect 34747 18136 34759 18139
rect 35176 18136 35204 18232
rect 34747 18108 35204 18136
rect 34747 18105 34759 18108
rect 34701 18099 34759 18105
rect 32030 18068 32036 18080
rect 29840 18040 32036 18068
rect 29549 18031 29607 18037
rect 32030 18028 32036 18040
rect 32088 18028 32094 18080
rect 33962 18028 33968 18080
rect 34020 18068 34026 18080
rect 34885 18071 34943 18077
rect 34885 18068 34897 18071
rect 34020 18040 34897 18068
rect 34020 18028 34026 18040
rect 34885 18037 34897 18040
rect 34931 18037 34943 18071
rect 34885 18031 34943 18037
rect 37093 18071 37151 18077
rect 37093 18037 37105 18071
rect 37139 18068 37151 18071
rect 37550 18068 37556 18080
rect 37139 18040 37556 18068
rect 37139 18037 37151 18040
rect 37093 18031 37151 18037
rect 37550 18028 37556 18040
rect 37608 18028 37614 18080
rect 37829 18071 37887 18077
rect 37829 18037 37841 18071
rect 37875 18068 37887 18071
rect 37875 18040 38424 18068
rect 37875 18037 37887 18040
rect 37829 18031 37887 18037
rect 38396 18012 38424 18040
rect 1104 17978 38272 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 38272 17978
rect 38378 17960 38384 18012
rect 38436 17960 38442 18012
rect 1104 17904 38272 17926
rect 1762 17824 1768 17876
rect 1820 17864 1826 17876
rect 2041 17867 2099 17873
rect 2041 17864 2053 17867
rect 1820 17836 2053 17864
rect 1820 17824 1826 17836
rect 2041 17833 2053 17836
rect 2087 17833 2099 17867
rect 2041 17827 2099 17833
rect 2130 17824 2136 17876
rect 2188 17864 2194 17876
rect 2961 17867 3019 17873
rect 2961 17864 2973 17867
rect 2188 17836 2973 17864
rect 2188 17824 2194 17836
rect 2961 17833 2973 17836
rect 3007 17833 3019 17867
rect 5626 17864 5632 17876
rect 2961 17827 3019 17833
rect 3344 17836 5632 17864
rect 1581 17731 1639 17737
rect 1581 17697 1593 17731
rect 1627 17728 1639 17731
rect 1670 17728 1676 17740
rect 1627 17700 1676 17728
rect 1627 17697 1639 17700
rect 1581 17691 1639 17697
rect 1670 17688 1676 17700
rect 1728 17688 1734 17740
rect 1765 17663 1823 17669
rect 1765 17629 1777 17663
rect 1811 17660 1823 17663
rect 1946 17660 1952 17672
rect 1811 17632 1952 17660
rect 1811 17629 1823 17632
rect 1765 17623 1823 17629
rect 1946 17620 1952 17632
rect 2004 17620 2010 17672
rect 2038 17620 2044 17672
rect 2096 17660 2102 17672
rect 3344 17669 3372 17836
rect 5626 17824 5632 17836
rect 5684 17824 5690 17876
rect 6914 17824 6920 17876
rect 6972 17864 6978 17876
rect 6972 17836 7604 17864
rect 6972 17824 6978 17836
rect 7576 17796 7604 17836
rect 7650 17824 7656 17876
rect 7708 17864 7714 17876
rect 7837 17867 7895 17873
rect 7837 17864 7849 17867
rect 7708 17836 7849 17864
rect 7708 17824 7714 17836
rect 7837 17833 7849 17836
rect 7883 17833 7895 17867
rect 7837 17827 7895 17833
rect 7926 17824 7932 17876
rect 7984 17864 7990 17876
rect 8021 17867 8079 17873
rect 8021 17864 8033 17867
rect 7984 17836 8033 17864
rect 7984 17824 7990 17836
rect 8021 17833 8033 17836
rect 8067 17833 8079 17867
rect 9766 17864 9772 17876
rect 8021 17827 8079 17833
rect 8864 17836 9772 17864
rect 8294 17796 8300 17808
rect 7576 17768 8300 17796
rect 8294 17756 8300 17768
rect 8352 17756 8358 17808
rect 3510 17688 3516 17740
rect 3568 17728 3574 17740
rect 3973 17731 4031 17737
rect 3973 17728 3985 17731
rect 3568 17700 3985 17728
rect 3568 17688 3574 17700
rect 3973 17697 3985 17700
rect 4019 17697 4031 17731
rect 8864 17728 8892 17836
rect 9766 17824 9772 17836
rect 9824 17824 9830 17876
rect 11333 17867 11391 17873
rect 11333 17833 11345 17867
rect 11379 17864 11391 17867
rect 11422 17864 11428 17876
rect 11379 17836 11428 17864
rect 11379 17833 11391 17836
rect 11333 17827 11391 17833
rect 11422 17824 11428 17836
rect 11480 17824 11486 17876
rect 12434 17864 12440 17876
rect 11716 17836 12440 17864
rect 8941 17799 8999 17805
rect 8941 17765 8953 17799
rect 8987 17765 8999 17799
rect 8941 17759 8999 17765
rect 11241 17799 11299 17805
rect 11241 17765 11253 17799
rect 11287 17796 11299 17799
rect 11716 17796 11744 17836
rect 12434 17824 12440 17836
rect 12492 17824 12498 17876
rect 12526 17824 12532 17876
rect 12584 17864 12590 17876
rect 12805 17867 12863 17873
rect 12805 17864 12817 17867
rect 12584 17836 12817 17864
rect 12584 17824 12590 17836
rect 12805 17833 12817 17836
rect 12851 17833 12863 17867
rect 12805 17827 12863 17833
rect 13081 17867 13139 17873
rect 13081 17833 13093 17867
rect 13127 17864 13139 17867
rect 13354 17864 13360 17876
rect 13127 17836 13360 17864
rect 13127 17833 13139 17836
rect 13081 17827 13139 17833
rect 13354 17824 13360 17836
rect 13412 17824 13418 17876
rect 15286 17824 15292 17876
rect 15344 17824 15350 17876
rect 17678 17824 17684 17876
rect 17736 17824 17742 17876
rect 20625 17867 20683 17873
rect 20625 17864 20637 17867
rect 17788 17836 20637 17864
rect 11287 17768 11744 17796
rect 11287 17765 11299 17768
rect 11241 17759 11299 17765
rect 3973 17691 4031 17697
rect 5644 17700 8892 17728
rect 2225 17663 2283 17669
rect 2225 17660 2237 17663
rect 2096 17632 2237 17660
rect 2096 17620 2102 17632
rect 2225 17629 2237 17632
rect 2271 17629 2283 17663
rect 2225 17623 2283 17629
rect 3237 17663 3295 17669
rect 3237 17629 3249 17663
rect 3283 17629 3295 17663
rect 3237 17623 3295 17629
rect 3329 17663 3387 17669
rect 3329 17629 3341 17663
rect 3375 17629 3387 17663
rect 3329 17623 3387 17629
rect 1946 17484 1952 17536
rect 2004 17484 2010 17536
rect 3252 17524 3280 17623
rect 3418 17620 3424 17672
rect 3476 17620 3482 17672
rect 3605 17663 3663 17669
rect 3605 17629 3617 17663
rect 3651 17660 3663 17663
rect 3694 17660 3700 17672
rect 3651 17632 3700 17660
rect 3651 17629 3663 17632
rect 3605 17623 3663 17629
rect 3694 17620 3700 17632
rect 3752 17620 3758 17672
rect 4246 17552 4252 17604
rect 4304 17552 4310 17604
rect 4706 17552 4712 17604
rect 4764 17552 4770 17604
rect 5644 17524 5672 17700
rect 6089 17663 6147 17669
rect 6089 17629 6101 17663
rect 6135 17629 6147 17663
rect 6089 17623 6147 17629
rect 8205 17663 8263 17669
rect 8205 17629 8217 17663
rect 8251 17660 8263 17663
rect 8956 17660 8984 17759
rect 12710 17756 12716 17808
rect 12768 17756 12774 17808
rect 12894 17756 12900 17808
rect 12952 17756 12958 17808
rect 14182 17756 14188 17808
rect 14240 17796 14246 17808
rect 16025 17799 16083 17805
rect 16025 17796 16037 17799
rect 14240 17768 16037 17796
rect 14240 17756 14246 17768
rect 16025 17765 16037 17768
rect 16071 17765 16083 17799
rect 16025 17759 16083 17765
rect 9030 17688 9036 17740
rect 9088 17728 9094 17740
rect 9401 17731 9459 17737
rect 9401 17728 9413 17731
rect 9088 17700 9413 17728
rect 9088 17688 9094 17700
rect 9401 17697 9413 17700
rect 9447 17697 9459 17731
rect 9401 17691 9459 17697
rect 9493 17731 9551 17737
rect 9493 17697 9505 17731
rect 9539 17697 9551 17731
rect 9493 17691 9551 17697
rect 8251 17632 8984 17660
rect 8251 17629 8263 17632
rect 8205 17623 8263 17629
rect 6104 17592 6132 17623
rect 6104 17564 6224 17592
rect 6196 17536 6224 17564
rect 6362 17552 6368 17604
rect 6420 17552 6426 17604
rect 6914 17552 6920 17604
rect 6972 17552 6978 17604
rect 9508 17592 9536 17691
rect 10042 17688 10048 17740
rect 10100 17728 10106 17740
rect 10873 17731 10931 17737
rect 10100 17700 10548 17728
rect 10100 17688 10106 17700
rect 10520 17672 10548 17700
rect 10873 17697 10885 17731
rect 10919 17728 10931 17731
rect 11146 17728 11152 17740
rect 10919 17700 11152 17728
rect 10919 17697 10931 17700
rect 10873 17691 10931 17697
rect 11146 17688 11152 17700
rect 11204 17688 11210 17740
rect 11698 17728 11704 17740
rect 11256 17700 11704 17728
rect 10137 17663 10195 17669
rect 10137 17629 10149 17663
rect 10183 17629 10195 17663
rect 10137 17623 10195 17629
rect 7760 17564 9536 17592
rect 10152 17592 10180 17623
rect 10318 17620 10324 17672
rect 10376 17660 10382 17672
rect 10413 17663 10471 17669
rect 10413 17660 10425 17663
rect 10376 17632 10425 17660
rect 10376 17620 10382 17632
rect 10413 17629 10425 17632
rect 10459 17629 10471 17663
rect 10413 17623 10471 17629
rect 10502 17620 10508 17672
rect 10560 17620 10566 17672
rect 11054 17620 11060 17672
rect 11112 17620 11118 17672
rect 11256 17669 11284 17700
rect 11698 17688 11704 17700
rect 11756 17688 11762 17740
rect 11977 17731 12035 17737
rect 11977 17697 11989 17731
rect 12023 17697 12035 17731
rect 11977 17691 12035 17697
rect 11241 17663 11299 17669
rect 11241 17629 11253 17663
rect 11287 17629 11299 17663
rect 11241 17623 11299 17629
rect 11606 17620 11612 17672
rect 11664 17660 11670 17672
rect 11793 17663 11851 17669
rect 11793 17660 11805 17663
rect 11664 17632 11805 17660
rect 11664 17620 11670 17632
rect 11793 17629 11805 17632
rect 11839 17629 11851 17663
rect 11793 17623 11851 17629
rect 11992 17604 12020 17691
rect 12250 17688 12256 17740
rect 12308 17688 12314 17740
rect 12728 17728 12756 17756
rect 12636 17700 12756 17728
rect 12912 17728 12940 17756
rect 14090 17728 14096 17740
rect 12912 17700 13032 17728
rect 10870 17592 10876 17604
rect 10152 17564 10876 17592
rect 7760 17536 7788 17564
rect 10870 17552 10876 17564
rect 10928 17552 10934 17604
rect 11698 17552 11704 17604
rect 11756 17552 11762 17604
rect 11974 17552 11980 17604
rect 12032 17552 12038 17604
rect 3252 17496 5672 17524
rect 5718 17484 5724 17536
rect 5776 17484 5782 17536
rect 6178 17484 6184 17536
rect 6236 17484 6242 17536
rect 7742 17484 7748 17536
rect 7800 17484 7806 17536
rect 9309 17527 9367 17533
rect 9309 17493 9321 17527
rect 9355 17524 9367 17527
rect 9582 17524 9588 17536
rect 9355 17496 9588 17524
rect 9355 17493 9367 17496
rect 9309 17487 9367 17493
rect 9582 17484 9588 17496
rect 9640 17484 9646 17536
rect 12268 17533 12296 17688
rect 12342 17620 12348 17672
rect 12400 17660 12406 17672
rect 12636 17669 12664 17700
rect 12437 17663 12495 17669
rect 12437 17660 12449 17663
rect 12400 17632 12449 17660
rect 12400 17620 12406 17632
rect 12437 17629 12449 17632
rect 12483 17629 12495 17663
rect 12437 17623 12495 17629
rect 12621 17663 12679 17669
rect 12621 17629 12633 17663
rect 12667 17629 12679 17663
rect 12621 17623 12679 17629
rect 12710 17620 12716 17672
rect 12768 17620 12774 17672
rect 13004 17671 13032 17700
rect 13740 17700 14096 17728
rect 12890 17663 12948 17669
rect 12890 17660 12902 17663
rect 12820 17632 12902 17660
rect 12820 17592 12848 17632
rect 12890 17629 12902 17632
rect 12936 17629 12948 17663
rect 12890 17623 12948 17629
rect 12989 17665 13047 17671
rect 13740 17669 13768 17700
rect 14090 17688 14096 17700
rect 14148 17688 14154 17740
rect 14826 17688 14832 17740
rect 14884 17688 14890 17740
rect 15473 17731 15531 17737
rect 15473 17697 15485 17731
rect 15519 17728 15531 17731
rect 16206 17728 16212 17740
rect 15519 17700 16212 17728
rect 15519 17697 15531 17700
rect 15473 17691 15531 17697
rect 16206 17688 16212 17700
rect 16264 17688 16270 17740
rect 17788 17728 17816 17836
rect 20625 17833 20637 17836
rect 20671 17864 20683 17867
rect 20806 17864 20812 17876
rect 20671 17836 20812 17864
rect 20671 17833 20683 17836
rect 20625 17827 20683 17833
rect 20806 17824 20812 17836
rect 20864 17864 20870 17876
rect 21634 17864 21640 17876
rect 20864 17836 21640 17864
rect 20864 17824 20870 17836
rect 21634 17824 21640 17836
rect 21692 17824 21698 17876
rect 22094 17824 22100 17876
rect 22152 17864 22158 17876
rect 22152 17836 22324 17864
rect 22152 17824 22158 17836
rect 18598 17796 18604 17808
rect 16408 17700 17816 17728
rect 18248 17768 18604 17796
rect 12989 17631 13001 17665
rect 13035 17631 13047 17665
rect 12989 17625 13047 17631
rect 13173 17663 13231 17669
rect 13173 17629 13185 17663
rect 13219 17629 13231 17663
rect 13173 17623 13231 17629
rect 13725 17663 13783 17669
rect 13725 17629 13737 17663
rect 13771 17629 13783 17663
rect 13725 17623 13783 17629
rect 13909 17663 13967 17669
rect 13909 17629 13921 17663
rect 13955 17660 13967 17663
rect 13955 17632 14136 17660
rect 13955 17629 13967 17632
rect 13909 17623 13967 17629
rect 13188 17592 13216 17623
rect 12820 17564 14044 17592
rect 14016 17536 14044 17564
rect 12253 17527 12311 17533
rect 12253 17493 12265 17527
rect 12299 17493 12311 17527
rect 12253 17487 12311 17493
rect 13633 17527 13691 17533
rect 13633 17493 13645 17527
rect 13679 17524 13691 17527
rect 13722 17524 13728 17536
rect 13679 17496 13728 17524
rect 13679 17493 13691 17496
rect 13633 17487 13691 17493
rect 13722 17484 13728 17496
rect 13780 17484 13786 17536
rect 13998 17484 14004 17536
rect 14056 17484 14062 17536
rect 14108 17524 14136 17632
rect 14182 17620 14188 17672
rect 14240 17660 14246 17672
rect 14277 17663 14335 17669
rect 14277 17660 14289 17663
rect 14240 17632 14289 17660
rect 14240 17620 14246 17632
rect 14277 17629 14289 17632
rect 14323 17629 14335 17663
rect 14844 17660 14872 17688
rect 16408 17672 16436 17700
rect 15565 17663 15623 17669
rect 15565 17660 15577 17663
rect 14844 17632 15577 17660
rect 14277 17623 14335 17629
rect 15565 17629 15577 17632
rect 15611 17629 15623 17663
rect 15565 17623 15623 17629
rect 15838 17620 15844 17672
rect 15896 17620 15902 17672
rect 16022 17620 16028 17672
rect 16080 17660 16086 17672
rect 16301 17663 16359 17669
rect 16301 17660 16313 17663
rect 16080 17632 16313 17660
rect 16080 17620 16086 17632
rect 16301 17629 16313 17632
rect 16347 17629 16359 17663
rect 16301 17623 16359 17629
rect 16390 17620 16396 17672
rect 16448 17620 16454 17672
rect 16482 17620 16488 17672
rect 16540 17620 16546 17672
rect 16574 17620 16580 17672
rect 16632 17660 16638 17672
rect 16669 17663 16727 17669
rect 16669 17660 16681 17663
rect 16632 17632 16681 17660
rect 16632 17620 16638 17632
rect 16669 17629 16681 17632
rect 16715 17660 16727 17663
rect 17218 17660 17224 17672
rect 16715 17632 17224 17660
rect 16715 17629 16727 17632
rect 16669 17623 16727 17629
rect 17218 17620 17224 17632
rect 17276 17620 17282 17672
rect 17310 17620 17316 17672
rect 17368 17660 17374 17672
rect 17405 17663 17463 17669
rect 17405 17660 17417 17663
rect 17368 17632 17417 17660
rect 17368 17620 17374 17632
rect 17405 17629 17417 17632
rect 17451 17629 17463 17663
rect 17405 17623 17463 17629
rect 17497 17663 17555 17669
rect 17497 17629 17509 17663
rect 17543 17660 17555 17663
rect 17865 17663 17923 17669
rect 17543 17632 17816 17660
rect 17543 17629 17555 17632
rect 17497 17623 17555 17629
rect 14366 17552 14372 17604
rect 14424 17592 14430 17604
rect 14645 17595 14703 17601
rect 14645 17592 14657 17595
rect 14424 17564 14657 17592
rect 14424 17552 14430 17564
rect 14645 17561 14657 17564
rect 14691 17561 14703 17595
rect 14645 17555 14703 17561
rect 15933 17595 15991 17601
rect 15933 17561 15945 17595
rect 15979 17592 15991 17595
rect 16206 17592 16212 17604
rect 15979 17564 16212 17592
rect 15979 17561 15991 17564
rect 15933 17555 15991 17561
rect 16206 17552 16212 17564
rect 16264 17552 16270 17604
rect 17034 17552 17040 17604
rect 17092 17592 17098 17604
rect 17788 17592 17816 17632
rect 17865 17629 17877 17663
rect 17911 17657 17923 17663
rect 17954 17657 17960 17672
rect 17911 17629 17960 17657
rect 17865 17623 17923 17629
rect 17954 17620 17960 17629
rect 18012 17620 18018 17672
rect 18046 17620 18052 17672
rect 18104 17620 18110 17672
rect 18138 17620 18144 17672
rect 18196 17620 18202 17672
rect 18248 17669 18276 17768
rect 18598 17756 18604 17768
rect 18656 17756 18662 17808
rect 19150 17756 19156 17808
rect 19208 17796 19214 17808
rect 19208 17768 22094 17796
rect 19208 17756 19214 17768
rect 18690 17728 18696 17740
rect 18340 17700 18696 17728
rect 18233 17663 18291 17669
rect 18233 17629 18245 17663
rect 18279 17629 18291 17663
rect 18233 17623 18291 17629
rect 18340 17592 18368 17700
rect 18690 17688 18696 17700
rect 18748 17728 18754 17740
rect 18748 17700 20208 17728
rect 18748 17688 18754 17700
rect 20180 17672 20208 17700
rect 20254 17688 20260 17740
rect 20312 17728 20318 17740
rect 20622 17728 20628 17740
rect 20312 17700 20628 17728
rect 20312 17688 20318 17700
rect 20622 17688 20628 17700
rect 20680 17688 20686 17740
rect 18417 17663 18475 17669
rect 18417 17629 18429 17663
rect 18463 17629 18475 17663
rect 18417 17623 18475 17629
rect 17092 17564 17632 17592
rect 17788 17564 18368 17592
rect 18432 17592 18460 17623
rect 18782 17620 18788 17672
rect 18840 17620 18846 17672
rect 18969 17663 19027 17669
rect 18969 17629 18981 17663
rect 19015 17660 19027 17663
rect 19518 17660 19524 17672
rect 19015 17632 19524 17660
rect 19015 17629 19027 17632
rect 18969 17623 19027 17629
rect 19518 17620 19524 17632
rect 19576 17620 19582 17672
rect 20070 17620 20076 17672
rect 20128 17620 20134 17672
rect 20162 17620 20168 17672
rect 20220 17660 20226 17672
rect 20349 17663 20407 17669
rect 20349 17660 20361 17663
rect 20220 17632 20361 17660
rect 20220 17620 20226 17632
rect 20349 17629 20361 17632
rect 20395 17660 20407 17663
rect 21174 17660 21180 17672
rect 20395 17632 21180 17660
rect 20395 17629 20407 17632
rect 20349 17623 20407 17629
rect 21174 17620 21180 17632
rect 21232 17620 21238 17672
rect 19242 17592 19248 17604
rect 18432 17564 19248 17592
rect 17092 17552 17098 17564
rect 14274 17524 14280 17536
rect 14108 17496 14280 17524
rect 14274 17484 14280 17496
rect 14332 17524 14338 17536
rect 16390 17524 16396 17536
rect 14332 17496 16396 17524
rect 14332 17484 14338 17496
rect 16390 17484 16396 17496
rect 16448 17484 16454 17536
rect 16482 17484 16488 17536
rect 16540 17524 16546 17536
rect 17494 17524 17500 17536
rect 16540 17496 17500 17524
rect 16540 17484 16546 17496
rect 17494 17484 17500 17496
rect 17552 17484 17558 17536
rect 17604 17524 17632 17564
rect 18432 17524 18460 17564
rect 19242 17552 19248 17564
rect 19300 17552 19306 17604
rect 19794 17552 19800 17604
rect 19852 17592 19858 17604
rect 20088 17592 20116 17620
rect 20533 17595 20591 17601
rect 20533 17592 20545 17595
rect 19852 17564 20545 17592
rect 19852 17552 19858 17564
rect 20533 17561 20545 17564
rect 20579 17561 20591 17595
rect 22066 17592 22094 17768
rect 22296 17669 22324 17836
rect 22646 17824 22652 17876
rect 22704 17824 22710 17876
rect 22925 17867 22983 17873
rect 22925 17833 22937 17867
rect 22971 17864 22983 17867
rect 23198 17864 23204 17876
rect 22971 17836 23204 17864
rect 22971 17833 22983 17836
rect 22925 17827 22983 17833
rect 23198 17824 23204 17836
rect 23256 17824 23262 17876
rect 26234 17824 26240 17876
rect 26292 17824 26298 17876
rect 26878 17824 26884 17876
rect 26936 17864 26942 17876
rect 27341 17867 27399 17873
rect 26936 17836 27108 17864
rect 26936 17824 26942 17836
rect 22664 17728 22692 17824
rect 23937 17799 23995 17805
rect 22572 17700 22692 17728
rect 23400 17768 23612 17796
rect 22281 17663 22339 17669
rect 22281 17629 22293 17663
rect 22327 17629 22339 17663
rect 22281 17623 22339 17629
rect 22462 17620 22468 17672
rect 22520 17620 22526 17672
rect 22572 17669 22600 17700
rect 22557 17663 22615 17669
rect 22557 17629 22569 17663
rect 22603 17629 22615 17663
rect 22557 17623 22615 17629
rect 22649 17663 22707 17669
rect 22649 17629 22661 17663
rect 22695 17660 22707 17663
rect 23400 17660 23428 17768
rect 23474 17688 23480 17740
rect 23532 17688 23538 17740
rect 23584 17728 23612 17768
rect 23937 17765 23949 17799
rect 23983 17796 23995 17799
rect 25593 17799 25651 17805
rect 23983 17768 25268 17796
rect 23983 17765 23995 17768
rect 23937 17759 23995 17765
rect 23584 17700 24624 17728
rect 22695 17632 23428 17660
rect 23569 17663 23627 17669
rect 22695 17629 22707 17632
rect 22649 17623 22707 17629
rect 23569 17629 23581 17663
rect 23615 17660 23627 17663
rect 23750 17660 23756 17672
rect 23615 17632 23756 17660
rect 23615 17629 23627 17632
rect 23569 17623 23627 17629
rect 23750 17620 23756 17632
rect 23808 17620 23814 17672
rect 24596 17669 24624 17700
rect 24670 17688 24676 17740
rect 24728 17688 24734 17740
rect 24949 17731 25007 17737
rect 24949 17697 24961 17731
rect 24995 17728 25007 17731
rect 25133 17731 25191 17737
rect 25133 17728 25145 17731
rect 24995 17700 25145 17728
rect 24995 17697 25007 17700
rect 24949 17691 25007 17697
rect 25133 17697 25145 17700
rect 25179 17697 25191 17731
rect 25133 17691 25191 17697
rect 24581 17663 24639 17669
rect 24581 17629 24593 17663
rect 24627 17660 24639 17663
rect 24762 17660 24768 17672
rect 24627 17632 24768 17660
rect 24627 17629 24639 17632
rect 24581 17623 24639 17629
rect 24762 17620 24768 17632
rect 24820 17620 24826 17672
rect 25240 17669 25268 17768
rect 25593 17765 25605 17799
rect 25639 17765 25651 17799
rect 25593 17759 25651 17765
rect 25225 17663 25283 17669
rect 25225 17629 25237 17663
rect 25271 17629 25283 17663
rect 25608 17660 25636 17759
rect 26252 17728 26280 17824
rect 26605 17799 26663 17805
rect 26605 17765 26617 17799
rect 26651 17796 26663 17799
rect 27080 17796 27108 17836
rect 27341 17833 27353 17867
rect 27387 17864 27399 17867
rect 27982 17864 27988 17876
rect 27387 17836 27988 17864
rect 27387 17833 27399 17836
rect 27341 17827 27399 17833
rect 27982 17824 27988 17836
rect 28040 17824 28046 17876
rect 31202 17864 31208 17876
rect 28092 17836 31208 17864
rect 28092 17796 28120 17836
rect 31202 17824 31208 17836
rect 31260 17824 31266 17876
rect 31297 17867 31355 17873
rect 31297 17833 31309 17867
rect 31343 17864 31355 17867
rect 31386 17864 31392 17876
rect 31343 17836 31392 17864
rect 31343 17833 31355 17836
rect 31297 17827 31355 17833
rect 31386 17824 31392 17836
rect 31444 17824 31450 17876
rect 32125 17867 32183 17873
rect 32125 17833 32137 17867
rect 32171 17864 32183 17867
rect 32490 17864 32496 17876
rect 32171 17836 32496 17864
rect 32171 17833 32183 17836
rect 32125 17827 32183 17833
rect 32490 17824 32496 17836
rect 32548 17824 32554 17876
rect 32306 17796 32312 17808
rect 26651 17768 27016 17796
rect 27080 17768 28120 17796
rect 29932 17768 32312 17796
rect 26651 17765 26663 17768
rect 26605 17759 26663 17765
rect 26988 17737 27016 17768
rect 26329 17731 26387 17737
rect 26329 17728 26341 17731
rect 26252 17700 26341 17728
rect 26329 17697 26341 17700
rect 26375 17697 26387 17731
rect 26329 17691 26387 17697
rect 26973 17731 27031 17737
rect 26973 17697 26985 17731
rect 27019 17697 27031 17731
rect 26973 17691 27031 17697
rect 27706 17688 27712 17740
rect 27764 17688 27770 17740
rect 29932 17728 29960 17768
rect 32306 17756 32312 17768
rect 32364 17756 32370 17808
rect 32398 17756 32404 17808
rect 32456 17796 32462 17808
rect 32456 17768 32812 17796
rect 32456 17756 32462 17768
rect 28184 17700 29960 17728
rect 28184 17672 28212 17700
rect 26237 17663 26295 17669
rect 26237 17660 26249 17663
rect 25608 17632 26249 17660
rect 25225 17623 25283 17629
rect 26237 17629 26249 17632
rect 26283 17629 26295 17663
rect 26237 17623 26295 17629
rect 27065 17663 27123 17669
rect 27065 17629 27077 17663
rect 27111 17660 27123 17663
rect 27430 17660 27436 17672
rect 27111 17632 27436 17660
rect 27111 17629 27123 17632
rect 27065 17623 27123 17629
rect 27430 17620 27436 17632
rect 27488 17620 27494 17672
rect 27890 17620 27896 17672
rect 27948 17620 27954 17672
rect 28166 17620 28172 17672
rect 28224 17620 28230 17672
rect 28350 17620 28356 17672
rect 28408 17620 28414 17672
rect 28537 17663 28595 17669
rect 28537 17629 28549 17663
rect 28583 17629 28595 17663
rect 28537 17623 28595 17629
rect 22066 17564 28212 17592
rect 20533 17555 20591 17561
rect 17604 17496 18460 17524
rect 18598 17484 18604 17536
rect 18656 17484 18662 17536
rect 18874 17484 18880 17536
rect 18932 17484 18938 17536
rect 18966 17484 18972 17536
rect 19024 17524 19030 17536
rect 23658 17524 23664 17536
rect 19024 17496 23664 17524
rect 19024 17484 19030 17496
rect 23658 17484 23664 17496
rect 23716 17484 23722 17536
rect 28184 17524 28212 17564
rect 28258 17552 28264 17604
rect 28316 17592 28322 17604
rect 28552 17592 28580 17623
rect 28626 17620 28632 17672
rect 28684 17660 28690 17672
rect 28997 17663 29055 17669
rect 28997 17660 29009 17663
rect 28684 17632 29009 17660
rect 28684 17620 28690 17632
rect 28997 17629 29009 17632
rect 29043 17660 29055 17663
rect 29549 17663 29607 17669
rect 29549 17660 29561 17663
rect 29043 17632 29561 17660
rect 29043 17629 29055 17632
rect 28997 17623 29055 17629
rect 29549 17629 29561 17632
rect 29595 17629 29607 17663
rect 29549 17623 29607 17629
rect 29730 17620 29736 17672
rect 29788 17620 29794 17672
rect 29932 17669 29960 17700
rect 30006 17688 30012 17740
rect 30064 17728 30070 17740
rect 32582 17728 32588 17740
rect 30064 17700 32588 17728
rect 30064 17688 30070 17700
rect 29825 17663 29883 17669
rect 29825 17629 29837 17663
rect 29871 17629 29883 17663
rect 29825 17623 29883 17629
rect 29917 17663 29975 17669
rect 29917 17629 29929 17663
rect 29963 17629 29975 17663
rect 29917 17623 29975 17629
rect 28316 17564 28580 17592
rect 29840 17592 29868 17623
rect 30282 17620 30288 17672
rect 30340 17620 30346 17672
rect 30484 17669 30512 17700
rect 32582 17688 32588 17700
rect 32640 17688 32646 17740
rect 30469 17663 30527 17669
rect 30469 17629 30481 17663
rect 30515 17629 30527 17663
rect 30469 17623 30527 17629
rect 31205 17663 31263 17669
rect 31205 17629 31217 17663
rect 31251 17660 31263 17663
rect 31294 17660 31300 17672
rect 31251 17632 31300 17660
rect 31251 17629 31263 17632
rect 31205 17623 31263 17629
rect 31294 17620 31300 17632
rect 31352 17620 31358 17672
rect 32033 17663 32091 17669
rect 32033 17660 32045 17663
rect 31956 17632 32045 17660
rect 31956 17604 31984 17632
rect 32033 17629 32045 17632
rect 32079 17629 32091 17663
rect 32784 17660 32812 17768
rect 34054 17756 34060 17808
rect 34112 17756 34118 17808
rect 32950 17660 32956 17672
rect 32784 17632 32956 17660
rect 32033 17623 32091 17629
rect 32950 17620 32956 17632
rect 33008 17660 33014 17672
rect 33781 17663 33839 17669
rect 33781 17660 33793 17663
rect 33008 17632 33793 17660
rect 33008 17620 33014 17632
rect 33781 17629 33793 17632
rect 33827 17629 33839 17663
rect 33781 17623 33839 17629
rect 33962 17620 33968 17672
rect 34020 17660 34026 17672
rect 34057 17663 34115 17669
rect 34057 17660 34069 17663
rect 34020 17632 34069 17660
rect 34020 17620 34026 17632
rect 34057 17629 34069 17632
rect 34103 17629 34115 17663
rect 34057 17623 34115 17629
rect 29840 17564 30420 17592
rect 28316 17552 28322 17564
rect 29178 17524 29184 17536
rect 28184 17496 29184 17524
rect 29178 17484 29184 17496
rect 29236 17484 29242 17536
rect 30190 17484 30196 17536
rect 30248 17484 30254 17536
rect 30392 17533 30420 17564
rect 31938 17552 31944 17604
rect 31996 17552 32002 17604
rect 30377 17527 30435 17533
rect 30377 17493 30389 17527
rect 30423 17524 30435 17527
rect 32490 17524 32496 17536
rect 30423 17496 32496 17524
rect 30423 17493 30435 17496
rect 30377 17487 30435 17493
rect 32490 17484 32496 17496
rect 32548 17484 32554 17536
rect 33778 17484 33784 17536
rect 33836 17524 33842 17536
rect 33873 17527 33931 17533
rect 33873 17524 33885 17527
rect 33836 17496 33885 17524
rect 33836 17484 33842 17496
rect 33873 17493 33885 17496
rect 33919 17493 33931 17527
rect 33873 17487 33931 17493
rect 1104 17434 38272 17456
rect 1104 17382 4874 17434
rect 4926 17382 4938 17434
rect 4990 17382 5002 17434
rect 5054 17382 5066 17434
rect 5118 17382 5130 17434
rect 5182 17382 35594 17434
rect 35646 17382 35658 17434
rect 35710 17382 35722 17434
rect 35774 17382 35786 17434
rect 35838 17382 35850 17434
rect 35902 17382 38272 17434
rect 1104 17360 38272 17382
rect 3418 17280 3424 17332
rect 3476 17280 3482 17332
rect 4246 17280 4252 17332
rect 4304 17280 4310 17332
rect 4525 17323 4583 17329
rect 4525 17289 4537 17323
rect 4571 17289 4583 17323
rect 4525 17283 4583 17289
rect 3053 17255 3111 17261
rect 3053 17221 3065 17255
rect 3099 17252 3111 17255
rect 3099 17224 3832 17252
rect 3099 17221 3111 17224
rect 3053 17215 3111 17221
rect 3804 17196 3832 17224
rect 3234 17144 3240 17196
rect 3292 17144 3298 17196
rect 3786 17144 3792 17196
rect 3844 17144 3850 17196
rect 4433 17187 4491 17193
rect 4433 17153 4445 17187
rect 4479 17184 4491 17187
rect 4540 17184 4568 17283
rect 5718 17280 5724 17332
rect 5776 17280 5782 17332
rect 6362 17280 6368 17332
rect 6420 17320 6426 17332
rect 6549 17323 6607 17329
rect 6549 17320 6561 17323
rect 6420 17292 6561 17320
rect 6420 17280 6426 17292
rect 6549 17289 6561 17292
rect 6595 17289 6607 17323
rect 6549 17283 6607 17289
rect 6917 17323 6975 17329
rect 6917 17289 6929 17323
rect 6963 17289 6975 17323
rect 6917 17283 6975 17289
rect 7377 17323 7435 17329
rect 7377 17289 7389 17323
rect 7423 17320 7435 17323
rect 7650 17320 7656 17332
rect 7423 17292 7656 17320
rect 7423 17289 7435 17292
rect 7377 17283 7435 17289
rect 4798 17212 4804 17264
rect 4856 17252 4862 17264
rect 4893 17255 4951 17261
rect 4893 17252 4905 17255
rect 4856 17224 4905 17252
rect 4856 17212 4862 17224
rect 4893 17221 4905 17224
rect 4939 17252 4951 17255
rect 5736 17252 5764 17280
rect 5905 17255 5963 17261
rect 5905 17252 5917 17255
rect 4939 17224 5917 17252
rect 4939 17221 4951 17224
rect 4893 17215 4951 17221
rect 5905 17221 5917 17224
rect 5951 17221 5963 17255
rect 5905 17215 5963 17221
rect 4479 17156 4568 17184
rect 4985 17187 5043 17193
rect 4479 17153 4491 17156
rect 4433 17147 4491 17153
rect 4985 17153 4997 17187
rect 5031 17184 5043 17187
rect 5258 17184 5264 17196
rect 5031 17156 5264 17184
rect 5031 17153 5043 17156
rect 4985 17147 5043 17153
rect 5258 17144 5264 17156
rect 5316 17144 5322 17196
rect 5721 17187 5779 17193
rect 5721 17184 5733 17187
rect 5644 17156 5733 17184
rect 3050 17076 3056 17128
rect 3108 17116 3114 17128
rect 5077 17119 5135 17125
rect 5077 17116 5089 17119
rect 3108 17088 5089 17116
rect 3108 17076 3114 17088
rect 5077 17085 5089 17088
rect 5123 17085 5135 17119
rect 5077 17079 5135 17085
rect 3786 16940 3792 16992
rect 3844 16980 3850 16992
rect 4062 16980 4068 16992
rect 3844 16952 4068 16980
rect 3844 16940 3850 16952
rect 4062 16940 4068 16952
rect 4120 16980 4126 16992
rect 5644 16980 5672 17156
rect 5721 17153 5733 17156
rect 5767 17153 5779 17187
rect 5721 17147 5779 17153
rect 6733 17187 6791 17193
rect 6733 17153 6745 17187
rect 6779 17184 6791 17187
rect 6932 17184 6960 17283
rect 7650 17280 7656 17292
rect 7708 17280 7714 17332
rect 9214 17320 9220 17332
rect 8956 17292 9220 17320
rect 6779 17156 6960 17184
rect 7285 17187 7343 17193
rect 6779 17153 6791 17156
rect 6733 17147 6791 17153
rect 7285 17153 7297 17187
rect 7331 17184 7343 17187
rect 8478 17184 8484 17196
rect 7331 17156 8484 17184
rect 7331 17153 7343 17156
rect 7285 17147 7343 17153
rect 8478 17144 8484 17156
rect 8536 17144 8542 17196
rect 8956 17193 8984 17292
rect 9214 17280 9220 17292
rect 9272 17320 9278 17332
rect 10134 17320 10140 17332
rect 9272 17292 10140 17320
rect 9272 17280 9278 17292
rect 10134 17280 10140 17292
rect 10192 17280 10198 17332
rect 10870 17280 10876 17332
rect 10928 17280 10934 17332
rect 11606 17280 11612 17332
rect 11664 17280 11670 17332
rect 11974 17280 11980 17332
rect 12032 17280 12038 17332
rect 12342 17320 12348 17332
rect 12084 17292 12348 17320
rect 9490 17212 9496 17264
rect 9548 17212 9554 17264
rect 9674 17212 9680 17264
rect 9732 17252 9738 17264
rect 9953 17255 10011 17261
rect 9953 17252 9965 17255
rect 9732 17224 9965 17252
rect 9732 17212 9738 17224
rect 9953 17221 9965 17224
rect 9999 17221 10011 17255
rect 9953 17215 10011 17221
rect 8941 17187 8999 17193
rect 8941 17153 8953 17187
rect 8987 17153 8999 17187
rect 8941 17147 8999 17153
rect 9030 17144 9036 17196
rect 9088 17184 9094 17196
rect 9125 17187 9183 17193
rect 9125 17184 9137 17187
rect 9088 17156 9137 17184
rect 9088 17144 9094 17156
rect 9125 17153 9137 17156
rect 9171 17184 9183 17187
rect 9508 17184 9536 17212
rect 9171 17156 9536 17184
rect 10228 17187 10286 17193
rect 9171 17153 9183 17156
rect 9125 17147 9183 17153
rect 10228 17153 10240 17187
rect 10274 17153 10286 17187
rect 10228 17147 10286 17153
rect 7561 17119 7619 17125
rect 7561 17085 7573 17119
rect 7607 17116 7619 17119
rect 7650 17116 7656 17128
rect 7607 17088 7656 17116
rect 7607 17085 7619 17088
rect 7561 17079 7619 17085
rect 7650 17076 7656 17088
rect 7708 17076 7714 17128
rect 10243 17116 10271 17147
rect 10318 17144 10324 17196
rect 10376 17144 10382 17196
rect 10410 17144 10416 17196
rect 10468 17144 10474 17196
rect 10597 17187 10655 17193
rect 10597 17153 10609 17187
rect 10643 17184 10655 17187
rect 10888 17184 10916 17280
rect 11624 17252 11652 17280
rect 12084 17252 12112 17292
rect 12342 17280 12348 17292
rect 12400 17280 12406 17332
rect 12434 17280 12440 17332
rect 12492 17280 12498 17332
rect 12710 17280 12716 17332
rect 12768 17320 12774 17332
rect 13814 17320 13820 17332
rect 12768 17292 13820 17320
rect 12768 17280 12774 17292
rect 13814 17280 13820 17292
rect 13872 17280 13878 17332
rect 13998 17280 14004 17332
rect 14056 17320 14062 17332
rect 15746 17320 15752 17332
rect 14056 17292 15752 17320
rect 14056 17280 14062 17292
rect 15746 17280 15752 17292
rect 15804 17280 15810 17332
rect 16206 17280 16212 17332
rect 16264 17320 16270 17332
rect 16574 17320 16580 17332
rect 16264 17292 16580 17320
rect 16264 17280 16270 17292
rect 16574 17280 16580 17292
rect 16632 17320 16638 17332
rect 21082 17320 21088 17332
rect 16632 17292 21088 17320
rect 16632 17280 16638 17292
rect 12452 17252 12480 17280
rect 18966 17252 18972 17264
rect 11624 17224 12112 17252
rect 12176 17224 12480 17252
rect 14108 17224 18972 17252
rect 10643 17156 10916 17184
rect 10643 17153 10655 17156
rect 10597 17147 10655 17153
rect 11790 17144 11796 17196
rect 11848 17184 11854 17196
rect 12176 17193 12204 17224
rect 11977 17187 12035 17193
rect 11977 17184 11989 17187
rect 11848 17156 11989 17184
rect 11848 17144 11854 17156
rect 11977 17153 11989 17156
rect 12023 17153 12035 17187
rect 11977 17147 12035 17153
rect 12161 17187 12219 17193
rect 12161 17153 12173 17187
rect 12207 17153 12219 17187
rect 12161 17147 12219 17153
rect 12253 17187 12311 17193
rect 12253 17153 12265 17187
rect 12299 17153 12311 17187
rect 12253 17147 12311 17153
rect 12437 17187 12495 17193
rect 12437 17153 12449 17187
rect 12483 17184 12495 17187
rect 12526 17184 12532 17196
rect 12483 17156 12532 17184
rect 12483 17153 12495 17156
rect 12437 17147 12495 17153
rect 11146 17116 11152 17128
rect 10243 17088 11152 17116
rect 11146 17076 11152 17088
rect 11204 17076 11210 17128
rect 12066 17076 12072 17128
rect 12124 17116 12130 17128
rect 12268 17116 12296 17147
rect 12526 17144 12532 17156
rect 12584 17144 12590 17196
rect 13538 17144 13544 17196
rect 13596 17144 13602 17196
rect 13556 17116 13584 17144
rect 12124 17088 13584 17116
rect 12124 17076 12130 17088
rect 7926 17008 7932 17060
rect 7984 17048 7990 17060
rect 14108 17048 14136 17224
rect 18966 17212 18972 17224
rect 19024 17212 19030 17264
rect 19150 17212 19156 17264
rect 19208 17212 19214 17264
rect 19306 17224 19748 17252
rect 15746 17144 15752 17196
rect 15804 17184 15810 17196
rect 16669 17187 16727 17193
rect 16669 17184 16681 17187
rect 15804 17156 16681 17184
rect 15804 17144 15810 17156
rect 16669 17153 16681 17156
rect 16715 17153 16727 17187
rect 16669 17147 16727 17153
rect 16850 17144 16856 17196
rect 16908 17144 16914 17196
rect 17310 17144 17316 17196
rect 17368 17144 17374 17196
rect 18046 17144 18052 17196
rect 18104 17184 18110 17196
rect 18414 17184 18420 17196
rect 18104 17156 18420 17184
rect 18104 17144 18110 17156
rect 18414 17144 18420 17156
rect 18472 17144 18478 17196
rect 14458 17076 14464 17128
rect 14516 17076 14522 17128
rect 17328 17116 17356 17144
rect 14568 17088 17356 17116
rect 7984 17020 14136 17048
rect 7984 17008 7990 17020
rect 14182 17008 14188 17060
rect 14240 17048 14246 17060
rect 14568 17048 14596 17088
rect 17494 17076 17500 17128
rect 17552 17116 17558 17128
rect 18782 17116 18788 17128
rect 17552 17088 18788 17116
rect 17552 17076 17558 17088
rect 18782 17076 18788 17088
rect 18840 17076 18846 17128
rect 14240 17020 14596 17048
rect 14240 17008 14246 17020
rect 15838 17008 15844 17060
rect 15896 17048 15902 17060
rect 16390 17048 16396 17060
rect 15896 17020 16396 17048
rect 15896 17008 15902 17020
rect 16390 17008 16396 17020
rect 16448 17008 16454 17060
rect 19168 17048 19196 17212
rect 16592 17020 19196 17048
rect 4120 16952 5672 16980
rect 4120 16940 4126 16952
rect 6086 16940 6092 16992
rect 6144 16940 6150 16992
rect 9309 16983 9367 16989
rect 9309 16949 9321 16983
rect 9355 16980 9367 16983
rect 9582 16980 9588 16992
rect 9355 16952 9588 16980
rect 9355 16949 9367 16952
rect 9309 16943 9367 16949
rect 9582 16940 9588 16952
rect 9640 16940 9646 16992
rect 11790 16940 11796 16992
rect 11848 16980 11854 16992
rect 16592 16980 16620 17020
rect 11848 16952 16620 16980
rect 11848 16940 11854 16952
rect 16666 16940 16672 16992
rect 16724 16940 16730 16992
rect 17037 16983 17095 16989
rect 17037 16949 17049 16983
rect 17083 16980 17095 16983
rect 17678 16980 17684 16992
rect 17083 16952 17684 16980
rect 17083 16949 17095 16952
rect 17037 16943 17095 16949
rect 17678 16940 17684 16952
rect 17736 16940 17742 16992
rect 18322 16940 18328 16992
rect 18380 16980 18386 16992
rect 19306 16980 19334 17224
rect 19720 17196 19748 17224
rect 19794 17212 19800 17264
rect 19852 17212 19858 17264
rect 19904 17261 19932 17292
rect 21082 17280 21088 17292
rect 21140 17280 21146 17332
rect 23106 17320 23112 17332
rect 22388 17292 23112 17320
rect 19889 17255 19947 17261
rect 19889 17221 19901 17255
rect 19935 17221 19947 17255
rect 19889 17215 19947 17221
rect 20162 17212 20168 17264
rect 20220 17212 20226 17264
rect 19613 17187 19671 17193
rect 19613 17153 19625 17187
rect 19659 17153 19671 17187
rect 19613 17147 19671 17153
rect 19628 17048 19656 17147
rect 19702 17144 19708 17196
rect 19760 17144 19766 17196
rect 19812 17184 19840 17212
rect 19981 17187 20039 17193
rect 19981 17184 19993 17187
rect 19812 17156 19993 17184
rect 19981 17153 19993 17156
rect 20027 17153 20039 17187
rect 19981 17147 20039 17153
rect 20078 17187 20136 17193
rect 20078 17153 20090 17187
rect 20124 17184 20136 17187
rect 20180 17184 20208 17212
rect 20625 17187 20683 17193
rect 20625 17184 20637 17187
rect 20124 17156 20208 17184
rect 20272 17156 20637 17184
rect 20124 17153 20136 17156
rect 20078 17147 20136 17153
rect 20162 17076 20168 17128
rect 20220 17116 20226 17128
rect 20272 17116 20300 17156
rect 20625 17153 20637 17156
rect 20671 17153 20683 17187
rect 20625 17147 20683 17153
rect 20717 17187 20775 17193
rect 20717 17153 20729 17187
rect 20763 17153 20775 17187
rect 20717 17147 20775 17153
rect 20220 17088 20300 17116
rect 20220 17076 20226 17088
rect 20346 17076 20352 17128
rect 20404 17076 20410 17128
rect 20438 17076 20444 17128
rect 20496 17116 20502 17128
rect 20732 17116 20760 17147
rect 20806 17144 20812 17196
rect 20864 17144 20870 17196
rect 22388 17193 22416 17292
rect 23106 17280 23112 17292
rect 23164 17280 23170 17332
rect 28162 17323 28220 17329
rect 28162 17289 28174 17323
rect 28208 17320 28220 17323
rect 28258 17320 28264 17332
rect 28208 17292 28264 17320
rect 28208 17289 28220 17292
rect 28162 17283 28220 17289
rect 28258 17280 28264 17292
rect 28316 17280 28322 17332
rect 28350 17280 28356 17332
rect 28408 17280 28414 17332
rect 28521 17323 28579 17329
rect 28521 17289 28533 17323
rect 28567 17320 28579 17323
rect 28567 17292 28856 17320
rect 28567 17289 28579 17292
rect 28521 17283 28579 17289
rect 28536 17252 28564 17283
rect 22572 17224 22968 17252
rect 22572 17196 22600 17224
rect 20993 17187 21051 17193
rect 20993 17153 21005 17187
rect 21039 17153 21051 17187
rect 20993 17147 21051 17153
rect 22373 17187 22431 17193
rect 22373 17153 22385 17187
rect 22419 17153 22431 17187
rect 22373 17147 22431 17153
rect 20496 17088 20760 17116
rect 20496 17076 20502 17088
rect 20714 17048 20720 17060
rect 19628 17020 20720 17048
rect 20714 17008 20720 17020
rect 20772 17008 20778 17060
rect 18380 16952 19334 16980
rect 20257 16983 20315 16989
rect 18380 16940 18386 16952
rect 20257 16949 20269 16983
rect 20303 16980 20315 16983
rect 21008 16980 21036 17147
rect 22554 17144 22560 17196
rect 22612 17144 22618 17196
rect 22940 17193 22968 17224
rect 28000 17224 28564 17252
rect 22925 17187 22983 17193
rect 22925 17153 22937 17187
rect 22971 17153 22983 17187
rect 22925 17147 22983 17153
rect 23477 17187 23535 17193
rect 23477 17153 23489 17187
rect 23523 17184 23535 17187
rect 27798 17184 27804 17196
rect 23523 17156 27804 17184
rect 23523 17153 23535 17156
rect 23477 17147 23535 17153
rect 27798 17144 27804 17156
rect 27856 17144 27862 17196
rect 28000 17193 28028 17224
rect 28626 17212 28632 17264
rect 28684 17252 28690 17264
rect 28721 17255 28779 17261
rect 28721 17252 28733 17255
rect 28684 17224 28733 17252
rect 28684 17212 28690 17224
rect 28721 17221 28733 17224
rect 28767 17221 28779 17255
rect 28721 17215 28779 17221
rect 27985 17187 28043 17193
rect 27985 17153 27997 17187
rect 28031 17153 28043 17187
rect 27985 17147 28043 17153
rect 28077 17187 28135 17193
rect 28077 17153 28089 17187
rect 28123 17153 28135 17187
rect 28077 17147 28135 17153
rect 28261 17187 28319 17193
rect 28261 17153 28273 17187
rect 28307 17184 28319 17187
rect 28644 17184 28672 17212
rect 28307 17156 28672 17184
rect 28307 17153 28319 17156
rect 28261 17147 28319 17153
rect 22465 17119 22523 17125
rect 22465 17085 22477 17119
rect 22511 17085 22523 17119
rect 22465 17079 22523 17085
rect 22480 17048 22508 17079
rect 23290 17076 23296 17128
rect 23348 17076 23354 17128
rect 28092 17116 28120 17147
rect 28828 17116 28856 17292
rect 29178 17280 29184 17332
rect 29236 17280 29242 17332
rect 30190 17280 30196 17332
rect 30248 17280 30254 17332
rect 31938 17320 31944 17332
rect 31680 17292 31944 17320
rect 30208 17252 30236 17280
rect 31680 17261 31708 17292
rect 31938 17280 31944 17292
rect 31996 17320 32002 17332
rect 32398 17320 32404 17332
rect 31996 17292 32404 17320
rect 31996 17280 32002 17292
rect 32398 17280 32404 17292
rect 32456 17280 32462 17332
rect 32858 17280 32864 17332
rect 32916 17320 32922 17332
rect 33042 17320 33048 17332
rect 32916 17292 33048 17320
rect 32916 17280 32922 17292
rect 33042 17280 33048 17292
rect 33100 17320 33106 17332
rect 33137 17323 33195 17329
rect 33137 17320 33149 17323
rect 33100 17292 33149 17320
rect 33100 17280 33106 17292
rect 33137 17289 33149 17292
rect 33183 17289 33195 17323
rect 33137 17283 33195 17289
rect 33962 17280 33968 17332
rect 34020 17329 34026 17332
rect 34020 17323 34039 17329
rect 34027 17289 34039 17323
rect 34020 17283 34039 17289
rect 34149 17323 34207 17329
rect 34149 17289 34161 17323
rect 34195 17289 34207 17323
rect 34149 17283 34207 17289
rect 34020 17280 34026 17283
rect 29012 17224 30236 17252
rect 31665 17255 31723 17261
rect 29012 17193 29040 17224
rect 31665 17221 31677 17255
rect 31711 17221 31723 17255
rect 31665 17215 31723 17221
rect 31849 17255 31907 17261
rect 31849 17221 31861 17255
rect 31895 17252 31907 17255
rect 32490 17252 32496 17264
rect 31895 17224 32496 17252
rect 31895 17221 31907 17224
rect 31849 17215 31907 17221
rect 32490 17212 32496 17224
rect 32548 17212 32554 17264
rect 33778 17212 33784 17264
rect 33836 17212 33842 17264
rect 28997 17187 29055 17193
rect 28997 17153 29009 17187
rect 29043 17153 29055 17187
rect 28997 17147 29055 17153
rect 29178 17144 29184 17196
rect 29236 17144 29242 17196
rect 29549 17187 29607 17193
rect 29549 17153 29561 17187
rect 29595 17184 29607 17187
rect 29638 17184 29644 17196
rect 29595 17156 29644 17184
rect 29595 17153 29607 17156
rect 29549 17147 29607 17153
rect 29638 17144 29644 17156
rect 29696 17144 29702 17196
rect 31941 17187 31999 17193
rect 31941 17153 31953 17187
rect 31987 17184 31999 17187
rect 32122 17184 32128 17196
rect 31987 17156 32128 17184
rect 31987 17153 31999 17156
rect 31941 17147 31999 17153
rect 32122 17144 32128 17156
rect 32180 17184 32186 17196
rect 32861 17187 32919 17193
rect 32861 17184 32873 17187
rect 32180 17156 32628 17184
rect 32180 17144 32186 17156
rect 28092 17088 28580 17116
rect 28828 17088 29500 17116
rect 23308 17048 23336 17076
rect 22480 17020 23336 17048
rect 23474 17008 23480 17060
rect 23532 17008 23538 17060
rect 28552 17048 28580 17088
rect 29362 17048 29368 17060
rect 28552 17020 29368 17048
rect 20303 16952 21036 16980
rect 22741 16983 22799 16989
rect 20303 16949 20315 16952
rect 20257 16943 20315 16949
rect 22741 16949 22753 16983
rect 22787 16980 22799 16983
rect 23492 16980 23520 17008
rect 28552 16989 28580 17020
rect 29362 17008 29368 17020
rect 29420 17008 29426 17060
rect 22787 16952 23520 16980
rect 28537 16983 28595 16989
rect 22787 16949 22799 16952
rect 22741 16943 22799 16949
rect 28537 16949 28549 16983
rect 28583 16949 28595 16983
rect 29472 16980 29500 17088
rect 32306 17076 32312 17128
rect 32364 17076 32370 17128
rect 32398 17076 32404 17128
rect 32456 17076 32462 17128
rect 32490 17076 32496 17128
rect 32548 17076 32554 17128
rect 32600 17125 32628 17156
rect 32692 17156 32873 17184
rect 32585 17119 32643 17125
rect 32585 17085 32597 17119
rect 32631 17085 32643 17119
rect 32585 17079 32643 17085
rect 31665 17051 31723 17057
rect 31665 17017 31677 17051
rect 31711 17048 31723 17051
rect 32692 17048 32720 17156
rect 32861 17153 32873 17156
rect 32907 17153 32919 17187
rect 32861 17147 32919 17153
rect 33045 17187 33103 17193
rect 33045 17153 33057 17187
rect 33091 17153 33103 17187
rect 34164 17184 34192 17283
rect 34514 17212 34520 17264
rect 34572 17252 34578 17264
rect 34572 17224 35204 17252
rect 34572 17212 34578 17224
rect 34425 17187 34483 17193
rect 34425 17184 34437 17187
rect 34164 17156 34437 17184
rect 33045 17147 33103 17153
rect 34425 17153 34437 17156
rect 34471 17184 34483 17187
rect 34885 17187 34943 17193
rect 34471 17156 34652 17184
rect 34471 17153 34483 17156
rect 34425 17147 34483 17153
rect 32769 17119 32827 17125
rect 32769 17085 32781 17119
rect 32815 17116 32827 17119
rect 33060 17116 33088 17147
rect 32815 17088 33088 17116
rect 32815 17085 32827 17088
rect 32769 17079 32827 17085
rect 34054 17076 34060 17128
rect 34112 17076 34118 17128
rect 34514 17076 34520 17128
rect 34572 17076 34578 17128
rect 34624 17116 34652 17156
rect 34885 17153 34897 17187
rect 34931 17184 34943 17187
rect 34931 17156 35112 17184
rect 34931 17153 34943 17156
rect 34885 17147 34943 17153
rect 34977 17119 35035 17125
rect 34977 17116 34989 17119
rect 34624 17088 34989 17116
rect 34977 17085 34989 17088
rect 35023 17085 35035 17119
rect 34977 17079 35035 17085
rect 31711 17020 32720 17048
rect 31711 17017 31723 17020
rect 31665 17011 31723 17017
rect 31846 16980 31852 16992
rect 29472 16952 31852 16980
rect 28537 16943 28595 16949
rect 31846 16940 31852 16952
rect 31904 16940 31910 16992
rect 32950 16940 32956 16992
rect 33008 16980 33014 16992
rect 33965 16983 34023 16989
rect 33965 16980 33977 16983
rect 33008 16952 33977 16980
rect 33008 16940 33014 16952
rect 33965 16949 33977 16952
rect 34011 16949 34023 16983
rect 34072 16980 34100 17076
rect 35084 17048 35112 17156
rect 35176 17125 35204 17224
rect 35161 17119 35219 17125
rect 35161 17085 35173 17119
rect 35207 17085 35219 17119
rect 35161 17079 35219 17085
rect 34440 17020 35112 17048
rect 34440 16989 34468 17020
rect 34425 16983 34483 16989
rect 34425 16980 34437 16983
rect 34072 16952 34437 16980
rect 33965 16943 34023 16949
rect 34425 16949 34437 16952
rect 34471 16949 34483 16983
rect 34425 16943 34483 16949
rect 34514 16940 34520 16992
rect 34572 16980 34578 16992
rect 34698 16980 34704 16992
rect 34572 16952 34704 16980
rect 34572 16940 34578 16952
rect 34698 16940 34704 16952
rect 34756 16940 34762 16992
rect 34790 16940 34796 16992
rect 34848 16940 34854 16992
rect 35069 16983 35127 16989
rect 35069 16949 35081 16983
rect 35115 16980 35127 16983
rect 35342 16980 35348 16992
rect 35115 16952 35348 16980
rect 35115 16949 35127 16952
rect 35069 16943 35127 16949
rect 35342 16940 35348 16952
rect 35400 16940 35406 16992
rect 1104 16890 38272 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 38272 16890
rect 1104 16816 38272 16838
rect 3602 16736 3608 16788
rect 3660 16776 3666 16788
rect 3660 16748 4660 16776
rect 3660 16736 3666 16748
rect 3789 16711 3847 16717
rect 3789 16708 3801 16711
rect 2792 16680 3801 16708
rect 2792 16649 2820 16680
rect 3789 16677 3801 16680
rect 3835 16677 3847 16711
rect 3789 16671 3847 16677
rect 2777 16643 2835 16649
rect 2777 16609 2789 16643
rect 2823 16609 2835 16643
rect 2777 16603 2835 16609
rect 2961 16643 3019 16649
rect 2961 16609 2973 16643
rect 3007 16640 3019 16643
rect 3050 16640 3056 16652
rect 3007 16612 3056 16640
rect 3007 16609 3019 16612
rect 2961 16603 3019 16609
rect 3050 16600 3056 16612
rect 3108 16600 3114 16652
rect 4430 16600 4436 16652
rect 4488 16600 4494 16652
rect 1949 16575 2007 16581
rect 1949 16541 1961 16575
rect 1995 16572 2007 16575
rect 2130 16572 2136 16584
rect 1995 16544 2136 16572
rect 1995 16541 2007 16544
rect 1949 16535 2007 16541
rect 2130 16532 2136 16544
rect 2188 16532 2194 16584
rect 2225 16575 2283 16581
rect 2225 16541 2237 16575
rect 2271 16572 2283 16575
rect 2271 16544 2360 16572
rect 2271 16541 2283 16544
rect 2225 16535 2283 16541
rect 1762 16396 1768 16448
rect 1820 16396 1826 16448
rect 1946 16396 1952 16448
rect 2004 16436 2010 16448
rect 2332 16445 2360 16544
rect 3970 16532 3976 16584
rect 4028 16532 4034 16584
rect 4154 16532 4160 16584
rect 4212 16574 4218 16584
rect 4525 16575 4583 16581
rect 4212 16572 4384 16574
rect 4212 16546 4476 16572
rect 4212 16532 4218 16546
rect 4356 16544 4476 16546
rect 4065 16507 4123 16513
rect 4065 16473 4077 16507
rect 4111 16473 4123 16507
rect 4065 16467 4123 16473
rect 2041 16439 2099 16445
rect 2041 16436 2053 16439
rect 2004 16408 2053 16436
rect 2004 16396 2010 16408
rect 2041 16405 2053 16408
rect 2087 16405 2099 16439
rect 2041 16399 2099 16405
rect 2317 16439 2375 16445
rect 2317 16405 2329 16439
rect 2363 16405 2375 16439
rect 2317 16399 2375 16405
rect 2685 16439 2743 16445
rect 2685 16405 2697 16439
rect 2731 16436 2743 16439
rect 3142 16436 3148 16448
rect 2731 16408 3148 16436
rect 2731 16405 2743 16408
rect 2685 16399 2743 16405
rect 3142 16396 3148 16408
rect 3200 16396 3206 16448
rect 4080 16436 4108 16467
rect 4246 16464 4252 16516
rect 4304 16513 4310 16516
rect 4304 16507 4353 16513
rect 4304 16473 4307 16507
rect 4341 16473 4353 16507
rect 4448 16504 4476 16544
rect 4525 16541 4537 16575
rect 4571 16572 4583 16575
rect 4632 16572 4660 16748
rect 6086 16736 6092 16788
rect 6144 16776 6150 16788
rect 6144 16748 12434 16776
rect 6144 16736 6150 16748
rect 8389 16711 8447 16717
rect 8389 16677 8401 16711
rect 8435 16708 8447 16711
rect 8478 16708 8484 16720
rect 8435 16680 8484 16708
rect 8435 16677 8447 16680
rect 8389 16671 8447 16677
rect 8478 16668 8484 16680
rect 8536 16668 8542 16720
rect 9030 16708 9036 16720
rect 8585 16680 9036 16708
rect 6178 16600 6184 16652
rect 6236 16640 6242 16652
rect 6236 16612 8524 16640
rect 6236 16600 6242 16612
rect 4571 16544 4660 16572
rect 4571 16541 4583 16544
rect 4525 16535 4583 16541
rect 5902 16504 5908 16516
rect 4448 16476 5908 16504
rect 4304 16467 4353 16473
rect 4304 16464 4310 16467
rect 5902 16464 5908 16476
rect 5960 16464 5966 16516
rect 8496 16504 8524 16612
rect 8585 16584 8613 16680
rect 9030 16668 9036 16680
rect 9088 16668 9094 16720
rect 12406 16708 12434 16748
rect 12986 16736 12992 16788
rect 13044 16776 13050 16788
rect 16022 16776 16028 16788
rect 13044 16748 16028 16776
rect 13044 16736 13050 16748
rect 16022 16736 16028 16748
rect 16080 16736 16086 16788
rect 16485 16779 16543 16785
rect 16485 16745 16497 16779
rect 16531 16776 16543 16779
rect 16574 16776 16580 16788
rect 16531 16748 16580 16776
rect 16531 16745 16543 16748
rect 16485 16739 16543 16745
rect 16574 16736 16580 16748
rect 16632 16736 16638 16788
rect 16666 16736 16672 16788
rect 16724 16736 16730 16788
rect 22462 16776 22468 16788
rect 17236 16748 22468 16776
rect 17236 16708 17264 16748
rect 22462 16736 22468 16748
rect 22520 16736 22526 16788
rect 27798 16736 27804 16788
rect 27856 16736 27862 16788
rect 29178 16736 29184 16788
rect 29236 16776 29242 16788
rect 30101 16779 30159 16785
rect 30101 16776 30113 16779
rect 29236 16748 30113 16776
rect 29236 16736 29242 16748
rect 30101 16745 30113 16748
rect 30147 16745 30159 16779
rect 30101 16739 30159 16745
rect 31202 16736 31208 16788
rect 31260 16736 31266 16788
rect 31846 16736 31852 16788
rect 31904 16776 31910 16788
rect 31904 16748 32076 16776
rect 31904 16736 31910 16748
rect 12406 16680 17264 16708
rect 18156 16680 20668 16708
rect 9125 16643 9183 16649
rect 9125 16640 9137 16643
rect 8680 16612 9137 16640
rect 8570 16532 8576 16584
rect 8628 16532 8634 16584
rect 8680 16504 8708 16612
rect 9125 16609 9137 16612
rect 9171 16609 9183 16643
rect 9125 16603 9183 16609
rect 15654 16600 15660 16652
rect 15712 16640 15718 16652
rect 16117 16643 16175 16649
rect 16117 16640 16129 16643
rect 15712 16612 16129 16640
rect 15712 16600 15718 16612
rect 16117 16609 16129 16612
rect 16163 16609 16175 16643
rect 16117 16603 16175 16609
rect 16390 16600 16396 16652
rect 16448 16640 16454 16652
rect 16761 16643 16819 16649
rect 16761 16640 16773 16643
rect 16448 16612 16773 16640
rect 16448 16600 16454 16612
rect 16761 16609 16773 16612
rect 16807 16609 16819 16643
rect 17681 16643 17739 16649
rect 17681 16640 17693 16643
rect 16761 16603 16819 16609
rect 17052 16612 17693 16640
rect 8757 16575 8815 16581
rect 8757 16541 8769 16575
rect 8803 16572 8815 16575
rect 8938 16572 8944 16584
rect 8803 16544 8944 16572
rect 8803 16541 8815 16544
rect 8757 16535 8815 16541
rect 8938 16532 8944 16544
rect 8996 16532 9002 16584
rect 14182 16532 14188 16584
rect 14240 16532 14246 16584
rect 15013 16575 15071 16581
rect 15013 16572 15025 16575
rect 14476 16544 15025 16572
rect 8496 16476 8708 16504
rect 9398 16464 9404 16516
rect 9456 16464 9462 16516
rect 9674 16464 9680 16516
rect 9732 16504 9738 16516
rect 9732 16476 9890 16504
rect 9732 16464 9738 16476
rect 11238 16464 11244 16516
rect 11296 16504 11302 16516
rect 13078 16504 13084 16516
rect 11296 16476 13084 16504
rect 11296 16464 11302 16476
rect 13078 16464 13084 16476
rect 13136 16464 13142 16516
rect 14476 16448 14504 16544
rect 15013 16541 15025 16544
rect 15059 16572 15071 16575
rect 15059 16544 16436 16572
rect 15059 16541 15071 16544
rect 15013 16535 15071 16541
rect 15686 16476 15792 16504
rect 4617 16439 4675 16445
rect 4617 16436 4629 16439
rect 4080 16408 4629 16436
rect 4617 16405 4629 16408
rect 4663 16405 4675 16439
rect 4617 16399 4675 16405
rect 10873 16439 10931 16445
rect 10873 16405 10885 16439
rect 10919 16436 10931 16439
rect 11054 16436 11060 16448
rect 10919 16408 11060 16436
rect 10919 16405 10931 16408
rect 10873 16399 10931 16405
rect 11054 16396 11060 16408
rect 11112 16436 11118 16448
rect 12250 16436 12256 16448
rect 11112 16408 12256 16436
rect 11112 16396 11118 16408
rect 12250 16396 12256 16408
rect 12308 16396 12314 16448
rect 14458 16396 14464 16448
rect 14516 16396 14522 16448
rect 15764 16436 15792 16476
rect 16298 16436 16304 16448
rect 15764 16408 16304 16436
rect 16298 16396 16304 16408
rect 16356 16396 16362 16448
rect 16408 16436 16436 16544
rect 16666 16532 16672 16584
rect 16724 16572 16730 16584
rect 16945 16575 17003 16581
rect 16945 16572 16957 16575
rect 16724 16544 16957 16572
rect 16724 16532 16730 16544
rect 16945 16541 16957 16544
rect 16991 16541 17003 16575
rect 16945 16535 17003 16541
rect 16574 16464 16580 16516
rect 16632 16504 16638 16516
rect 17052 16504 17080 16612
rect 17681 16609 17693 16612
rect 17727 16609 17739 16643
rect 17681 16603 17739 16609
rect 17221 16575 17279 16581
rect 17221 16541 17233 16575
rect 17267 16572 17279 16575
rect 17586 16572 17592 16584
rect 17267 16544 17592 16572
rect 17267 16541 17279 16544
rect 17221 16535 17279 16541
rect 17420 16516 17448 16544
rect 17586 16532 17592 16544
rect 17644 16532 17650 16584
rect 18156 16581 18184 16680
rect 20640 16652 20668 16680
rect 20714 16668 20720 16720
rect 20772 16668 20778 16720
rect 22278 16668 22284 16720
rect 22336 16708 22342 16720
rect 23106 16708 23112 16720
rect 22336 16680 23112 16708
rect 22336 16668 22342 16680
rect 23106 16668 23112 16680
rect 23164 16668 23170 16720
rect 27816 16708 27844 16736
rect 30282 16708 30288 16720
rect 27816 16680 30288 16708
rect 30282 16668 30288 16680
rect 30340 16708 30346 16720
rect 32048 16708 32076 16748
rect 32122 16736 32128 16788
rect 32180 16736 32186 16788
rect 35161 16779 35219 16785
rect 35161 16745 35173 16779
rect 35207 16776 35219 16779
rect 35250 16776 35256 16788
rect 35207 16748 35256 16776
rect 35207 16745 35219 16748
rect 35161 16739 35219 16745
rect 35250 16736 35256 16748
rect 35308 16736 35314 16788
rect 35434 16736 35440 16788
rect 35492 16736 35498 16788
rect 34333 16711 34391 16717
rect 34333 16708 34345 16711
rect 30340 16680 31892 16708
rect 32048 16680 34345 16708
rect 30340 16668 30346 16680
rect 18230 16600 18236 16652
rect 18288 16640 18294 16652
rect 18288 16612 18368 16640
rect 18288 16600 18294 16612
rect 18340 16581 18368 16612
rect 20162 16600 20168 16652
rect 20220 16640 20226 16652
rect 20530 16640 20536 16652
rect 20220 16612 20536 16640
rect 20220 16600 20226 16612
rect 20530 16600 20536 16612
rect 20588 16600 20594 16652
rect 20622 16600 20628 16652
rect 20680 16600 20686 16652
rect 20732 16640 20760 16668
rect 20732 16612 21404 16640
rect 17957 16575 18015 16581
rect 17957 16541 17969 16575
rect 18003 16541 18015 16575
rect 17957 16535 18015 16541
rect 18141 16575 18199 16581
rect 18141 16541 18153 16575
rect 18187 16541 18199 16575
rect 18141 16535 18199 16541
rect 18325 16575 18383 16581
rect 18325 16541 18337 16575
rect 18371 16541 18383 16575
rect 18325 16535 18383 16541
rect 16632 16476 17080 16504
rect 16632 16464 16638 16476
rect 17402 16464 17408 16516
rect 17460 16464 17466 16516
rect 17972 16504 18000 16535
rect 18598 16532 18604 16584
rect 18656 16532 18662 16584
rect 18782 16532 18788 16584
rect 18840 16572 18846 16584
rect 20070 16572 20076 16584
rect 18840 16544 20076 16572
rect 18840 16532 18846 16544
rect 20070 16532 20076 16544
rect 20128 16572 20134 16584
rect 20257 16575 20315 16581
rect 20257 16572 20269 16575
rect 20128 16544 20269 16572
rect 20128 16532 20134 16544
rect 20257 16541 20269 16544
rect 20303 16541 20315 16575
rect 20257 16535 20315 16541
rect 20346 16532 20352 16584
rect 20404 16572 20410 16584
rect 20548 16572 20576 16600
rect 20806 16581 20812 16584
rect 20763 16575 20812 16581
rect 20404 16544 20449 16572
rect 20548 16544 20668 16572
rect 20404 16532 20410 16544
rect 18690 16504 18696 16516
rect 17972 16476 18696 16504
rect 18690 16464 18696 16476
rect 18748 16464 18754 16516
rect 19058 16464 19064 16516
rect 19116 16464 19122 16516
rect 20640 16513 20668 16544
rect 20763 16541 20775 16575
rect 20809 16541 20812 16575
rect 20763 16535 20812 16541
rect 20806 16532 20812 16535
rect 20864 16532 20870 16584
rect 20990 16532 20996 16584
rect 21048 16532 21054 16584
rect 21376 16581 21404 16612
rect 23198 16600 23204 16652
rect 23256 16600 23262 16652
rect 23493 16643 23551 16649
rect 23493 16640 23505 16643
rect 23308 16612 23505 16640
rect 23308 16584 23336 16612
rect 23493 16609 23505 16612
rect 23539 16640 23551 16643
rect 23842 16640 23848 16652
rect 23539 16612 23848 16640
rect 23539 16609 23551 16612
rect 23493 16603 23551 16609
rect 23842 16600 23848 16612
rect 23900 16600 23906 16652
rect 23937 16643 23995 16649
rect 23937 16609 23949 16643
rect 23983 16640 23995 16643
rect 24854 16640 24860 16652
rect 23983 16612 24860 16640
rect 23983 16609 23995 16612
rect 23937 16603 23995 16609
rect 24854 16600 24860 16612
rect 24912 16640 24918 16652
rect 25593 16643 25651 16649
rect 24912 16612 25544 16640
rect 24912 16600 24918 16612
rect 21361 16575 21419 16581
rect 21361 16541 21373 16575
rect 21407 16541 21419 16575
rect 21361 16535 21419 16541
rect 21821 16575 21879 16581
rect 21821 16541 21833 16575
rect 21867 16541 21879 16575
rect 21821 16535 21879 16541
rect 20533 16507 20591 16513
rect 20533 16473 20545 16507
rect 20579 16473 20591 16507
rect 20533 16467 20591 16473
rect 20625 16507 20683 16513
rect 20625 16473 20637 16507
rect 20671 16473 20683 16507
rect 21836 16504 21864 16535
rect 22278 16532 22284 16584
rect 22336 16532 22342 16584
rect 23290 16532 23296 16584
rect 23348 16532 23354 16584
rect 23382 16532 23388 16584
rect 23440 16581 23446 16584
rect 23440 16575 23467 16581
rect 23455 16541 23467 16575
rect 23440 16535 23467 16541
rect 23440 16532 23446 16535
rect 25222 16532 25228 16584
rect 25280 16532 25286 16584
rect 25409 16575 25467 16581
rect 25409 16541 25421 16575
rect 25455 16541 25467 16575
rect 25516 16572 25544 16612
rect 25593 16609 25605 16643
rect 25639 16640 25651 16643
rect 26234 16640 26240 16652
rect 25639 16612 26240 16640
rect 25639 16609 25651 16612
rect 25593 16603 25651 16609
rect 26234 16600 26240 16612
rect 26292 16600 26298 16652
rect 31754 16640 31760 16652
rect 30024 16612 31760 16640
rect 26050 16572 26056 16584
rect 25516 16544 26056 16572
rect 25409 16535 25467 16541
rect 20625 16467 20683 16473
rect 20916 16476 21864 16504
rect 22097 16507 22155 16513
rect 16485 16439 16543 16445
rect 16485 16436 16497 16439
rect 16408 16408 16497 16436
rect 16485 16405 16497 16408
rect 16531 16405 16543 16439
rect 16485 16399 16543 16405
rect 16942 16396 16948 16448
rect 17000 16436 17006 16448
rect 17129 16439 17187 16445
rect 17129 16436 17141 16439
rect 17000 16408 17141 16436
rect 17000 16396 17006 16408
rect 17129 16405 17141 16408
rect 17175 16405 17187 16439
rect 17129 16399 17187 16405
rect 17678 16396 17684 16448
rect 17736 16436 17742 16448
rect 18046 16436 18052 16448
rect 17736 16408 18052 16436
rect 17736 16396 17742 16408
rect 18046 16396 18052 16408
rect 18104 16396 18110 16448
rect 18138 16396 18144 16448
rect 18196 16436 18202 16448
rect 18506 16436 18512 16448
rect 18196 16408 18512 16436
rect 18196 16396 18202 16408
rect 18506 16396 18512 16408
rect 18564 16436 18570 16448
rect 20548 16436 20576 16467
rect 20916 16448 20944 16476
rect 22097 16473 22109 16507
rect 22143 16504 22155 16507
rect 22462 16504 22468 16516
rect 22143 16476 22468 16504
rect 22143 16473 22155 16476
rect 22097 16467 22155 16473
rect 22462 16464 22468 16476
rect 22520 16464 22526 16516
rect 22833 16507 22891 16513
rect 22833 16473 22845 16507
rect 22879 16504 22891 16507
rect 23198 16504 23204 16516
rect 22879 16476 23204 16504
rect 22879 16473 22891 16476
rect 22833 16467 22891 16473
rect 23198 16464 23204 16476
rect 23256 16464 23262 16516
rect 23750 16464 23756 16516
rect 23808 16464 23814 16516
rect 25424 16504 25452 16535
rect 26050 16532 26056 16544
rect 26108 16532 26114 16584
rect 30024 16581 30052 16612
rect 31754 16600 31760 16612
rect 31812 16600 31818 16652
rect 30009 16575 30067 16581
rect 30009 16541 30021 16575
rect 30055 16541 30067 16575
rect 30009 16535 30067 16541
rect 30190 16532 30196 16584
rect 30248 16532 30254 16584
rect 30282 16532 30288 16584
rect 30340 16572 30346 16584
rect 30561 16575 30619 16581
rect 30561 16572 30573 16575
rect 30340 16544 30573 16572
rect 30340 16532 30346 16544
rect 30561 16541 30573 16544
rect 30607 16541 30619 16575
rect 30561 16535 30619 16541
rect 30650 16532 30656 16584
rect 30708 16572 30714 16584
rect 30745 16575 30803 16581
rect 30745 16572 30757 16575
rect 30708 16544 30757 16572
rect 30708 16532 30714 16544
rect 30745 16541 30757 16544
rect 30791 16572 30803 16575
rect 31110 16572 31116 16584
rect 30791 16544 31116 16572
rect 30791 16541 30803 16544
rect 30745 16535 30803 16541
rect 31110 16532 31116 16544
rect 31168 16532 31174 16584
rect 31389 16575 31447 16581
rect 31389 16541 31401 16575
rect 31435 16572 31447 16575
rect 31478 16572 31484 16584
rect 31435 16544 31484 16572
rect 31435 16541 31447 16544
rect 31389 16535 31447 16541
rect 31478 16532 31484 16544
rect 31536 16532 31542 16584
rect 31864 16572 31892 16680
rect 34333 16677 34345 16680
rect 34379 16677 34391 16711
rect 34333 16671 34391 16677
rect 34425 16711 34483 16717
rect 34425 16677 34437 16711
rect 34471 16708 34483 16711
rect 35345 16711 35403 16717
rect 35345 16708 35357 16711
rect 34471 16680 35357 16708
rect 34471 16677 34483 16680
rect 34425 16671 34483 16677
rect 35345 16677 35357 16680
rect 35391 16708 35403 16711
rect 35391 16680 35664 16708
rect 35391 16677 35403 16680
rect 35345 16671 35403 16677
rect 34241 16643 34299 16649
rect 34241 16609 34253 16643
rect 34287 16640 34299 16643
rect 34698 16640 34704 16652
rect 34287 16612 34704 16640
rect 34287 16609 34299 16612
rect 34241 16603 34299 16609
rect 34698 16600 34704 16612
rect 34756 16640 34762 16652
rect 35529 16643 35587 16649
rect 35529 16640 35541 16643
rect 34756 16612 35541 16640
rect 34756 16600 34762 16612
rect 35529 16609 35541 16612
rect 35575 16609 35587 16643
rect 35529 16603 35587 16609
rect 32309 16575 32367 16581
rect 32309 16572 32321 16575
rect 31864 16544 32321 16572
rect 32309 16541 32321 16544
rect 32355 16541 32367 16575
rect 34517 16575 34575 16581
rect 32309 16535 32367 16541
rect 32416 16544 34376 16572
rect 25148 16476 25452 16504
rect 25148 16448 25176 16476
rect 25958 16464 25964 16516
rect 26016 16504 26022 16516
rect 26237 16507 26295 16513
rect 26237 16504 26249 16507
rect 26016 16476 26249 16504
rect 26016 16464 26022 16476
rect 26237 16473 26249 16476
rect 26283 16473 26295 16507
rect 26237 16467 26295 16473
rect 29362 16464 29368 16516
rect 29420 16504 29426 16516
rect 32416 16504 32444 16544
rect 29420 16476 32444 16504
rect 32493 16507 32551 16513
rect 29420 16464 29426 16476
rect 32493 16473 32505 16507
rect 32539 16504 32551 16507
rect 32766 16504 32772 16516
rect 32539 16476 32772 16504
rect 32539 16473 32551 16476
rect 32493 16467 32551 16473
rect 32766 16464 32772 16476
rect 32824 16464 32830 16516
rect 18564 16408 20576 16436
rect 18564 16396 18570 16408
rect 20898 16396 20904 16448
rect 20956 16396 20962 16448
rect 22646 16396 22652 16448
rect 22704 16436 22710 16448
rect 23293 16439 23351 16445
rect 23293 16436 23305 16439
rect 22704 16408 23305 16436
rect 22704 16396 22710 16408
rect 23293 16405 23305 16408
rect 23339 16436 23351 16439
rect 24946 16436 24952 16448
rect 23339 16408 24952 16436
rect 23339 16405 23351 16408
rect 23293 16399 23351 16405
rect 24946 16396 24952 16408
rect 25004 16396 25010 16448
rect 25130 16396 25136 16448
rect 25188 16396 25194 16448
rect 26418 16396 26424 16448
rect 26476 16396 26482 16448
rect 27154 16396 27160 16448
rect 27212 16436 27218 16448
rect 30650 16436 30656 16448
rect 27212 16408 30656 16436
rect 27212 16396 27218 16408
rect 30650 16396 30656 16408
rect 30708 16396 30714 16448
rect 30742 16396 30748 16448
rect 30800 16396 30806 16448
rect 34348 16436 34376 16544
rect 34517 16541 34529 16575
rect 34563 16572 34575 16575
rect 35066 16572 35072 16584
rect 34563 16544 35072 16572
rect 34563 16541 34575 16544
rect 34517 16535 34575 16541
rect 35066 16532 35072 16544
rect 35124 16532 35130 16584
rect 35437 16575 35495 16581
rect 35437 16541 35449 16575
rect 35483 16572 35495 16575
rect 35636 16572 35664 16680
rect 35483 16544 35664 16572
rect 35483 16541 35495 16544
rect 35437 16535 35495 16541
rect 34790 16464 34796 16516
rect 34848 16504 34854 16516
rect 34977 16507 35035 16513
rect 34977 16504 34989 16507
rect 34848 16476 34989 16504
rect 34848 16464 34854 16476
rect 34977 16473 34989 16476
rect 35023 16473 35035 16507
rect 34977 16467 35035 16473
rect 35084 16476 35848 16504
rect 35084 16436 35112 16476
rect 34348 16408 35112 16436
rect 35158 16396 35164 16448
rect 35216 16445 35222 16448
rect 35820 16445 35848 16476
rect 35216 16439 35235 16445
rect 35223 16405 35235 16439
rect 35216 16399 35235 16405
rect 35805 16439 35863 16445
rect 35805 16405 35817 16439
rect 35851 16405 35863 16439
rect 35805 16399 35863 16405
rect 35216 16396 35222 16399
rect 1104 16346 38272 16368
rect 1104 16294 4874 16346
rect 4926 16294 4938 16346
rect 4990 16294 5002 16346
rect 5054 16294 5066 16346
rect 5118 16294 5130 16346
rect 5182 16294 35594 16346
rect 35646 16294 35658 16346
rect 35710 16294 35722 16346
rect 35774 16294 35786 16346
rect 35838 16294 35850 16346
rect 35902 16294 38272 16346
rect 1104 16272 38272 16294
rect 1394 16192 1400 16244
rect 1452 16232 1458 16244
rect 2958 16232 2964 16244
rect 1452 16204 2964 16232
rect 1452 16192 1458 16204
rect 2958 16192 2964 16204
rect 3016 16192 3022 16244
rect 3602 16192 3608 16244
rect 3660 16232 3666 16244
rect 3881 16235 3939 16241
rect 3881 16232 3893 16235
rect 3660 16204 3893 16232
rect 3660 16192 3666 16204
rect 3881 16201 3893 16204
rect 3927 16201 3939 16235
rect 3881 16195 3939 16201
rect 4049 16235 4107 16241
rect 4049 16201 4061 16235
rect 4095 16232 4107 16235
rect 4614 16232 4620 16244
rect 4095 16204 4620 16232
rect 4095 16201 4107 16204
rect 4049 16195 4107 16201
rect 4614 16192 4620 16204
rect 4672 16192 4678 16244
rect 5169 16235 5227 16241
rect 5169 16201 5181 16235
rect 5215 16232 5227 16235
rect 5258 16232 5264 16244
rect 5215 16204 5264 16232
rect 5215 16201 5227 16204
rect 5169 16195 5227 16201
rect 5258 16192 5264 16204
rect 5316 16192 5322 16244
rect 9398 16192 9404 16244
rect 9456 16232 9462 16244
rect 9493 16235 9551 16241
rect 9493 16232 9505 16235
rect 9456 16204 9505 16232
rect 9456 16192 9462 16204
rect 9493 16201 9505 16204
rect 9539 16201 9551 16235
rect 9493 16195 9551 16201
rect 9769 16235 9827 16241
rect 9769 16201 9781 16235
rect 9815 16201 9827 16235
rect 9769 16195 9827 16201
rect 10137 16235 10195 16241
rect 10137 16201 10149 16235
rect 10183 16232 10195 16235
rect 11238 16232 11244 16244
rect 10183 16204 11244 16232
rect 10183 16201 10195 16204
rect 10137 16195 10195 16201
rect 1673 16167 1731 16173
rect 1673 16133 1685 16167
rect 1719 16164 1731 16167
rect 1946 16164 1952 16176
rect 1719 16136 1952 16164
rect 1719 16133 1731 16136
rect 1673 16127 1731 16133
rect 1946 16124 1952 16136
rect 2004 16124 2010 16176
rect 4249 16167 4307 16173
rect 4249 16133 4261 16167
rect 4295 16164 4307 16167
rect 4798 16164 4804 16176
rect 4295 16136 4804 16164
rect 4295 16133 4307 16136
rect 4249 16127 4307 16133
rect 4798 16124 4804 16136
rect 4856 16124 4862 16176
rect 5460 16136 6040 16164
rect 4706 16096 4712 16108
rect 2806 16068 4712 16096
rect 4706 16056 4712 16068
rect 4764 16056 4770 16108
rect 1394 15988 1400 16040
rect 1452 15988 1458 16040
rect 2130 15988 2136 16040
rect 2188 16028 2194 16040
rect 5460 16028 5488 16136
rect 5537 16099 5595 16105
rect 5537 16065 5549 16099
rect 5583 16065 5595 16099
rect 5537 16059 5595 16065
rect 2188 16000 5488 16028
rect 2188 15988 2194 16000
rect 5552 15960 5580 16059
rect 5626 15988 5632 16040
rect 5684 15988 5690 16040
rect 5813 16031 5871 16037
rect 5813 15997 5825 16031
rect 5859 16028 5871 16031
rect 5902 16028 5908 16040
rect 5859 16000 5908 16028
rect 5859 15997 5871 16000
rect 5813 15991 5871 15997
rect 5902 15988 5908 16000
rect 5960 15988 5966 16040
rect 6012 16028 6040 16136
rect 9677 16099 9735 16105
rect 9677 16065 9689 16099
rect 9723 16096 9735 16099
rect 9784 16096 9812 16195
rect 11238 16192 11244 16204
rect 11296 16192 11302 16244
rect 14090 16192 14096 16244
rect 14148 16232 14154 16244
rect 14277 16235 14335 16241
rect 14277 16232 14289 16235
rect 14148 16204 14289 16232
rect 14148 16192 14154 16204
rect 14277 16201 14289 16204
rect 14323 16201 14335 16235
rect 14277 16195 14335 16201
rect 16666 16192 16672 16244
rect 16724 16232 16730 16244
rect 16853 16235 16911 16241
rect 16853 16232 16865 16235
rect 16724 16204 16865 16232
rect 16724 16192 16730 16204
rect 16853 16201 16865 16204
rect 16899 16201 16911 16235
rect 16853 16195 16911 16201
rect 17037 16235 17095 16241
rect 17037 16201 17049 16235
rect 17083 16232 17095 16235
rect 18230 16232 18236 16244
rect 17083 16204 18236 16232
rect 17083 16201 17095 16204
rect 17037 16195 17095 16201
rect 18230 16192 18236 16204
rect 18288 16232 18294 16244
rect 18288 16204 19012 16232
rect 18288 16192 18294 16204
rect 10229 16167 10287 16173
rect 10229 16133 10241 16167
rect 10275 16164 10287 16167
rect 11054 16164 11060 16176
rect 10275 16136 11060 16164
rect 10275 16133 10287 16136
rect 10229 16127 10287 16133
rect 11054 16124 11060 16136
rect 11112 16124 11118 16176
rect 12618 16124 12624 16176
rect 12676 16164 12682 16176
rect 12676 16136 16344 16164
rect 12676 16124 12682 16136
rect 9723 16068 9812 16096
rect 9876 16068 12204 16096
rect 9723 16065 9735 16068
rect 9677 16059 9735 16065
rect 9876 16028 9904 16068
rect 12176 16040 12204 16068
rect 12250 16056 12256 16108
rect 12308 16056 12314 16108
rect 12342 16056 12348 16108
rect 12400 16056 12406 16108
rect 14458 16056 14464 16108
rect 14516 16056 14522 16108
rect 14734 16056 14740 16108
rect 14792 16056 14798 16108
rect 14826 16056 14832 16108
rect 14884 16056 14890 16108
rect 6012 16000 9904 16028
rect 10318 15988 10324 16040
rect 10376 15988 10382 16040
rect 12158 15988 12164 16040
rect 12216 15988 12222 16040
rect 12526 15988 12532 16040
rect 12584 15988 12590 16040
rect 14645 16031 14703 16037
rect 14645 15997 14657 16031
rect 14691 16028 14703 16031
rect 14844 16028 14872 16056
rect 14691 16000 14872 16028
rect 16316 16028 16344 16136
rect 16758 16124 16764 16176
rect 16816 16164 16822 16176
rect 17221 16167 17279 16173
rect 17221 16164 17233 16167
rect 16816 16136 17233 16164
rect 16816 16124 16822 16136
rect 17221 16133 17233 16136
rect 17267 16164 17279 16167
rect 17310 16164 17316 16176
rect 17267 16136 17316 16164
rect 17267 16133 17279 16136
rect 17221 16127 17279 16133
rect 17310 16124 17316 16136
rect 17368 16124 17374 16176
rect 17497 16167 17555 16173
rect 17497 16164 17509 16167
rect 17420 16136 17509 16164
rect 16390 16056 16396 16108
rect 16448 16096 16454 16108
rect 16945 16099 17003 16105
rect 16945 16096 16957 16099
rect 16448 16068 16957 16096
rect 16448 16056 16454 16068
rect 16945 16065 16957 16068
rect 16991 16065 17003 16099
rect 16945 16059 17003 16065
rect 17420 16028 17448 16136
rect 17497 16133 17509 16136
rect 17543 16133 17555 16167
rect 17697 16167 17755 16173
rect 17697 16164 17709 16167
rect 17497 16127 17555 16133
rect 17696 16133 17709 16164
rect 17743 16133 17755 16167
rect 17696 16127 17755 16133
rect 16316 16000 17448 16028
rect 14691 15997 14703 16000
rect 14645 15991 14703 15997
rect 11885 15963 11943 15969
rect 11885 15960 11897 15963
rect 5552 15932 11897 15960
rect 11885 15929 11897 15932
rect 11931 15929 11943 15963
rect 16758 15960 16764 15972
rect 11885 15923 11943 15929
rect 12406 15932 16764 15960
rect 3142 15852 3148 15904
rect 3200 15892 3206 15904
rect 3878 15892 3884 15904
rect 3200 15864 3884 15892
rect 3200 15852 3206 15864
rect 3878 15852 3884 15864
rect 3936 15892 3942 15904
rect 4065 15895 4123 15901
rect 4065 15892 4077 15895
rect 3936 15864 4077 15892
rect 3936 15852 3942 15864
rect 4065 15861 4077 15864
rect 4111 15892 4123 15895
rect 12406 15892 12434 15932
rect 16758 15920 16764 15932
rect 16816 15920 16822 15972
rect 17420 15960 17448 16000
rect 17494 15988 17500 16040
rect 17552 16028 17558 16040
rect 17696 16028 17724 16127
rect 17862 16124 17868 16176
rect 17920 16164 17926 16176
rect 18785 16167 18843 16173
rect 18785 16164 18797 16167
rect 17920 16136 18797 16164
rect 17920 16124 17926 16136
rect 18785 16133 18797 16136
rect 18831 16133 18843 16167
rect 18984 16164 19012 16204
rect 19058 16192 19064 16244
rect 19116 16232 19122 16244
rect 19116 16204 20684 16232
rect 19116 16192 19122 16204
rect 20165 16167 20223 16173
rect 20165 16164 20177 16167
rect 18984 16136 20177 16164
rect 18785 16127 18843 16133
rect 20165 16133 20177 16136
rect 20211 16133 20223 16167
rect 20165 16127 20223 16133
rect 20346 16124 20352 16176
rect 20404 16124 20410 16176
rect 20549 16167 20607 16173
rect 20549 16164 20561 16167
rect 20548 16133 20561 16164
rect 20595 16133 20607 16167
rect 20656 16164 20684 16204
rect 20714 16192 20720 16244
rect 20772 16192 20778 16244
rect 21453 16235 21511 16241
rect 21453 16201 21465 16235
rect 21499 16232 21511 16235
rect 22278 16232 22284 16244
rect 21499 16204 22284 16232
rect 21499 16201 21511 16204
rect 21453 16195 21511 16201
rect 22278 16192 22284 16204
rect 22336 16192 22342 16244
rect 29273 16235 29331 16241
rect 22940 16204 27108 16232
rect 22940 16164 22968 16204
rect 20656 16136 22968 16164
rect 20548 16127 20607 16133
rect 17957 16099 18015 16105
rect 17957 16096 17969 16099
rect 17552 16000 17724 16028
rect 17756 16068 17969 16096
rect 17552 15988 17558 16000
rect 17586 15960 17592 15972
rect 17420 15932 17592 15960
rect 17586 15920 17592 15932
rect 17644 15960 17650 15972
rect 17756 15960 17784 16068
rect 17957 16065 17969 16068
rect 18003 16065 18015 16099
rect 17957 16059 18015 16065
rect 18046 16056 18052 16108
rect 18104 16056 18110 16108
rect 18138 16056 18144 16108
rect 18196 16056 18202 16108
rect 18233 16099 18291 16105
rect 18233 16065 18245 16099
rect 18279 16065 18291 16099
rect 18233 16059 18291 16065
rect 18325 16099 18383 16105
rect 18325 16065 18337 16099
rect 18371 16096 18383 16099
rect 18874 16096 18880 16108
rect 18371 16068 18880 16096
rect 18371 16065 18383 16068
rect 18325 16059 18383 16065
rect 18064 16028 18092 16056
rect 18248 16028 18276 16059
rect 18064 16000 18276 16028
rect 17644 15932 17784 15960
rect 17644 15920 17650 15932
rect 17862 15920 17868 15972
rect 17920 15920 17926 15972
rect 4111 15864 12434 15892
rect 4111 15861 4123 15864
rect 4065 15855 4123 15861
rect 14182 15852 14188 15904
rect 14240 15892 14246 15904
rect 14734 15892 14740 15904
rect 14240 15864 14740 15892
rect 14240 15852 14246 15864
rect 14734 15852 14740 15864
rect 14792 15852 14798 15904
rect 16666 15852 16672 15904
rect 16724 15852 16730 15904
rect 17681 15895 17739 15901
rect 17681 15861 17693 15895
rect 17727 15892 17739 15895
rect 18340 15892 18368 16059
rect 18874 16056 18880 16068
rect 18932 16056 18938 16108
rect 19702 16056 19708 16108
rect 19760 16096 19766 16108
rect 20257 16099 20315 16105
rect 20257 16096 20269 16099
rect 19760 16068 20269 16096
rect 19760 16056 19766 16068
rect 20257 16065 20269 16068
rect 20303 16096 20315 16099
rect 20438 16096 20444 16108
rect 20303 16068 20444 16096
rect 20303 16065 20315 16068
rect 20257 16059 20315 16065
rect 20438 16056 20444 16068
rect 20496 16056 20502 16108
rect 20548 16040 20576 16127
rect 23014 16124 23020 16176
rect 23072 16124 23078 16176
rect 25130 16124 25136 16176
rect 25188 16164 25194 16176
rect 27080 16164 27108 16204
rect 29273 16201 29285 16235
rect 29319 16232 29331 16235
rect 29319 16204 30144 16232
rect 29319 16201 29331 16204
rect 29273 16195 29331 16201
rect 27246 16164 27252 16176
rect 25188 16136 26280 16164
rect 27080 16136 27252 16164
rect 25188 16124 25194 16136
rect 20898 16056 20904 16108
rect 20956 16096 20962 16108
rect 21269 16099 21327 16105
rect 21269 16096 21281 16099
rect 20956 16068 21281 16096
rect 20956 16056 20962 16068
rect 21269 16065 21281 16068
rect 21315 16065 21327 16099
rect 21269 16059 21327 16065
rect 21542 16056 21548 16108
rect 21600 16096 21606 16108
rect 22002 16096 22008 16108
rect 21600 16068 22008 16096
rect 21600 16056 21606 16068
rect 22002 16056 22008 16068
rect 22060 16096 22066 16108
rect 22833 16099 22891 16105
rect 22833 16096 22845 16099
rect 22060 16068 22845 16096
rect 22060 16056 22066 16068
rect 22833 16065 22845 16068
rect 22879 16065 22891 16099
rect 22833 16059 22891 16065
rect 23109 16099 23167 16105
rect 23109 16065 23121 16099
rect 23155 16065 23167 16099
rect 23109 16059 23167 16065
rect 23201 16099 23259 16105
rect 23201 16065 23213 16099
rect 23247 16096 23259 16099
rect 23290 16096 23296 16108
rect 23247 16068 23296 16096
rect 23247 16065 23259 16068
rect 23201 16059 23259 16065
rect 20530 15988 20536 16040
rect 20588 15988 20594 16040
rect 20990 15988 20996 16040
rect 21048 15988 21054 16040
rect 20346 15920 20352 15972
rect 20404 15960 20410 15972
rect 23124 15960 23152 16059
rect 20404 15932 23152 15960
rect 20404 15920 20410 15932
rect 17727 15864 18368 15892
rect 17727 15861 17739 15864
rect 17681 15855 17739 15861
rect 18598 15852 18604 15904
rect 18656 15852 18662 15904
rect 18874 15852 18880 15904
rect 18932 15852 18938 15904
rect 20162 15852 20168 15904
rect 20220 15892 20226 15904
rect 20533 15895 20591 15901
rect 20533 15892 20545 15895
rect 20220 15864 20545 15892
rect 20220 15852 20226 15864
rect 20533 15861 20545 15864
rect 20579 15861 20591 15895
rect 20533 15855 20591 15861
rect 20714 15852 20720 15904
rect 20772 15892 20778 15904
rect 21085 15895 21143 15901
rect 21085 15892 21097 15895
rect 20772 15864 21097 15892
rect 20772 15852 20778 15864
rect 21085 15861 21097 15864
rect 21131 15861 21143 15895
rect 21085 15855 21143 15861
rect 22922 15852 22928 15904
rect 22980 15892 22986 15904
rect 23216 15892 23244 16059
rect 23290 16056 23296 16068
rect 23348 16056 23354 16108
rect 24670 16056 24676 16108
rect 24728 16056 24734 16108
rect 24854 16056 24860 16108
rect 24912 16096 24918 16108
rect 26252 16105 26280 16136
rect 25225 16099 25283 16105
rect 25225 16096 25237 16099
rect 24912 16068 25237 16096
rect 24912 16056 24918 16068
rect 25225 16065 25237 16068
rect 25271 16065 25283 16099
rect 25225 16059 25283 16065
rect 26237 16099 26295 16105
rect 26237 16065 26249 16099
rect 26283 16065 26295 16099
rect 26237 16059 26295 16065
rect 26329 16099 26387 16105
rect 26329 16065 26341 16099
rect 26375 16065 26387 16099
rect 26329 16059 26387 16065
rect 25222 15920 25228 15972
rect 25280 15960 25286 15972
rect 26344 15960 26372 16059
rect 26418 16056 26424 16108
rect 26476 16096 26482 16108
rect 27172 16105 27200 16136
rect 27246 16124 27252 16136
rect 27304 16164 27310 16176
rect 29365 16167 29423 16173
rect 29365 16164 29377 16167
rect 27304 16136 29377 16164
rect 27304 16124 27310 16136
rect 27065 16099 27123 16105
rect 27065 16096 27077 16099
rect 26476 16068 27077 16096
rect 26476 16056 26482 16068
rect 27065 16065 27077 16068
rect 27111 16065 27123 16099
rect 27065 16059 27123 16065
rect 27157 16099 27215 16105
rect 27157 16065 27169 16099
rect 27203 16065 27215 16099
rect 27157 16059 27215 16065
rect 27338 16056 27344 16108
rect 27396 16056 27402 16108
rect 29104 16105 29132 16136
rect 29365 16133 29377 16136
rect 29411 16164 29423 16167
rect 30116 16164 30144 16204
rect 30190 16192 30196 16244
rect 30248 16232 30254 16244
rect 30469 16235 30527 16241
rect 30469 16232 30481 16235
rect 30248 16204 30481 16232
rect 30248 16192 30254 16204
rect 30469 16201 30481 16204
rect 30515 16201 30527 16235
rect 30469 16195 30527 16201
rect 30742 16192 30748 16244
rect 30800 16232 30806 16244
rect 30837 16235 30895 16241
rect 30837 16232 30849 16235
rect 30800 16204 30849 16232
rect 30800 16192 30806 16204
rect 30837 16201 30849 16204
rect 30883 16201 30895 16235
rect 30837 16195 30895 16201
rect 34790 16192 34796 16244
rect 34848 16232 34854 16244
rect 34977 16235 35035 16241
rect 34977 16232 34989 16235
rect 34848 16204 34989 16232
rect 34848 16192 34854 16204
rect 34977 16201 34989 16204
rect 35023 16201 35035 16235
rect 34977 16195 35035 16201
rect 35066 16192 35072 16244
rect 35124 16232 35130 16244
rect 35434 16232 35440 16244
rect 35124 16204 35440 16232
rect 35124 16192 35130 16204
rect 35434 16192 35440 16204
rect 35492 16192 35498 16244
rect 30282 16164 30288 16176
rect 29411 16136 29684 16164
rect 29411 16133 29423 16136
rect 29365 16127 29423 16133
rect 29656 16108 29684 16136
rect 30116 16136 30288 16164
rect 29089 16099 29147 16105
rect 29089 16065 29101 16099
rect 29135 16065 29147 16099
rect 29089 16059 29147 16065
rect 29273 16099 29331 16105
rect 29273 16065 29285 16099
rect 29319 16096 29331 16099
rect 29546 16096 29552 16108
rect 29319 16094 29408 16096
rect 29472 16094 29552 16096
rect 29319 16068 29552 16094
rect 29319 16065 29331 16068
rect 29380 16066 29500 16068
rect 29273 16059 29331 16065
rect 29546 16056 29552 16068
rect 29604 16056 29610 16108
rect 29638 16056 29644 16108
rect 29696 16056 29702 16108
rect 30116 16105 30144 16136
rect 30282 16124 30288 16136
rect 30340 16164 30346 16176
rect 31021 16167 31079 16173
rect 31021 16164 31033 16167
rect 30340 16136 31033 16164
rect 30340 16124 30346 16136
rect 31021 16133 31033 16136
rect 31067 16133 31079 16167
rect 31021 16127 31079 16133
rect 31110 16124 31116 16176
rect 31168 16164 31174 16176
rect 31205 16167 31263 16173
rect 31205 16164 31217 16167
rect 31168 16136 31217 16164
rect 31168 16124 31174 16136
rect 31205 16133 31217 16136
rect 31251 16133 31263 16167
rect 31205 16127 31263 16133
rect 34716 16136 37688 16164
rect 30101 16099 30159 16105
rect 30101 16065 30113 16099
rect 30147 16065 30159 16099
rect 30101 16059 30159 16065
rect 30653 16099 30711 16105
rect 30653 16065 30665 16099
rect 30699 16065 30711 16099
rect 30653 16059 30711 16065
rect 30929 16099 30987 16105
rect 30929 16065 30941 16099
rect 30975 16065 30987 16099
rect 30929 16059 30987 16065
rect 26513 16031 26571 16037
rect 26513 15997 26525 16031
rect 26559 16028 26571 16031
rect 27249 16031 27307 16037
rect 27249 16028 27261 16031
rect 26559 16000 27261 16028
rect 26559 15997 26571 16000
rect 26513 15991 26571 15997
rect 27249 15997 27261 16000
rect 27295 16028 27307 16031
rect 29178 16028 29184 16040
rect 27295 16000 29184 16028
rect 27295 15997 27307 16000
rect 27249 15991 27307 15997
rect 29178 15988 29184 16000
rect 29236 15988 29242 16040
rect 29733 16031 29791 16037
rect 29733 15997 29745 16031
rect 29779 16028 29791 16031
rect 29917 16031 29975 16037
rect 29917 16028 29929 16031
rect 29779 16000 29929 16028
rect 29779 15997 29791 16000
rect 29733 15991 29791 15997
rect 29917 15997 29929 16000
rect 29963 15997 29975 16031
rect 29917 15991 29975 15997
rect 25280 15932 26372 15960
rect 25280 15920 25286 15932
rect 27338 15920 27344 15972
rect 27396 15960 27402 15972
rect 30668 15960 30696 16059
rect 30944 16028 30972 16059
rect 32214 16028 32220 16040
rect 30944 16000 32220 16028
rect 32214 15988 32220 16000
rect 32272 15988 32278 16040
rect 34716 15960 34744 16136
rect 34885 16099 34943 16105
rect 34885 16065 34897 16099
rect 34931 16065 34943 16099
rect 34885 16059 34943 16065
rect 34900 16028 34928 16059
rect 35158 16056 35164 16108
rect 35216 16096 35222 16108
rect 37660 16105 37688 16136
rect 37645 16099 37703 16105
rect 35216 16068 35388 16096
rect 35216 16056 35222 16068
rect 35250 16028 35256 16040
rect 34900 16000 35256 16028
rect 35250 15988 35256 16000
rect 35308 15988 35314 16040
rect 27396 15932 30696 15960
rect 30760 15932 34744 15960
rect 27396 15920 27402 15932
rect 22980 15864 23244 15892
rect 23385 15895 23443 15901
rect 22980 15852 22986 15864
rect 23385 15861 23397 15895
rect 23431 15892 23443 15895
rect 24026 15892 24032 15904
rect 23431 15864 24032 15892
rect 23431 15861 23443 15864
rect 23385 15855 23443 15861
rect 24026 15852 24032 15864
rect 24084 15852 24090 15904
rect 25038 15852 25044 15904
rect 25096 15892 25102 15904
rect 26053 15895 26111 15901
rect 26053 15892 26065 15895
rect 25096 15864 26065 15892
rect 25096 15852 25102 15864
rect 26053 15861 26065 15864
rect 26099 15892 26111 15895
rect 27154 15892 27160 15904
rect 26099 15864 27160 15892
rect 26099 15861 26111 15864
rect 26053 15855 26111 15861
rect 27154 15852 27160 15864
rect 27212 15852 27218 15904
rect 27525 15895 27583 15901
rect 27525 15861 27537 15895
rect 27571 15892 27583 15895
rect 30006 15892 30012 15904
rect 27571 15864 30012 15892
rect 27571 15861 27583 15864
rect 27525 15855 27583 15861
rect 30006 15852 30012 15864
rect 30064 15852 30070 15904
rect 30190 15852 30196 15904
rect 30248 15892 30254 15904
rect 30285 15895 30343 15901
rect 30285 15892 30297 15895
rect 30248 15864 30297 15892
rect 30248 15852 30254 15864
rect 30285 15861 30297 15864
rect 30331 15861 30343 15895
rect 30285 15855 30343 15861
rect 30374 15852 30380 15904
rect 30432 15892 30438 15904
rect 30760 15892 30788 15932
rect 35066 15920 35072 15972
rect 35124 15960 35130 15972
rect 35161 15963 35219 15969
rect 35161 15960 35173 15963
rect 35124 15932 35173 15960
rect 35124 15920 35130 15932
rect 35161 15929 35173 15932
rect 35207 15929 35219 15963
rect 35161 15923 35219 15929
rect 35360 15904 35388 16068
rect 37645 16065 37657 16099
rect 37691 16065 37703 16099
rect 37645 16059 37703 16065
rect 30432 15864 30788 15892
rect 30432 15852 30438 15864
rect 31386 15852 31392 15904
rect 31444 15852 31450 15904
rect 31754 15852 31760 15904
rect 31812 15892 31818 15904
rect 32490 15892 32496 15904
rect 31812 15864 32496 15892
rect 31812 15852 31818 15864
rect 32490 15852 32496 15864
rect 32548 15852 32554 15904
rect 35342 15852 35348 15904
rect 35400 15852 35406 15904
rect 37826 15852 37832 15904
rect 37884 15852 37890 15904
rect 1104 15802 38272 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 38272 15802
rect 1104 15728 38272 15750
rect 934 15648 940 15700
rect 992 15688 998 15700
rect 1489 15691 1547 15697
rect 1489 15688 1501 15691
rect 992 15660 1501 15688
rect 992 15648 998 15660
rect 1489 15657 1501 15660
rect 1535 15657 1547 15691
rect 1489 15651 1547 15657
rect 3789 15691 3847 15697
rect 3789 15657 3801 15691
rect 3835 15688 3847 15691
rect 3970 15688 3976 15700
rect 3835 15660 3976 15688
rect 3835 15657 3847 15660
rect 3789 15651 3847 15657
rect 3970 15648 3976 15660
rect 4028 15648 4034 15700
rect 4706 15648 4712 15700
rect 4764 15648 4770 15700
rect 4985 15691 5043 15697
rect 4985 15657 4997 15691
rect 5031 15688 5043 15691
rect 5626 15688 5632 15700
rect 5031 15660 5632 15688
rect 5031 15657 5043 15660
rect 4985 15651 5043 15657
rect 5626 15648 5632 15660
rect 5684 15648 5690 15700
rect 7926 15648 7932 15700
rect 7984 15648 7990 15700
rect 9490 15648 9496 15700
rect 9548 15688 9554 15700
rect 10226 15688 10232 15700
rect 9548 15660 10232 15688
rect 9548 15648 9554 15660
rect 10226 15648 10232 15660
rect 10284 15648 10290 15700
rect 12526 15688 12532 15700
rect 11532 15660 12532 15688
rect 4614 15620 4620 15632
rect 4540 15592 4620 15620
rect 4540 15561 4568 15592
rect 4614 15580 4620 15592
rect 4672 15580 4678 15632
rect 4724 15620 4752 15648
rect 4724 15592 6316 15620
rect 4065 15555 4123 15561
rect 4065 15521 4077 15555
rect 4111 15552 4123 15555
rect 4525 15555 4583 15561
rect 4111 15524 4476 15552
rect 4111 15521 4123 15524
rect 4065 15515 4123 15521
rect 1762 15444 1768 15496
rect 1820 15444 1826 15496
rect 3878 15444 3884 15496
rect 3936 15444 3942 15496
rect 3970 15444 3976 15496
rect 4028 15444 4034 15496
rect 4154 15444 4160 15496
rect 4212 15444 4218 15496
rect 4249 15487 4307 15493
rect 4249 15453 4261 15487
rect 4295 15453 4307 15487
rect 4448 15484 4476 15524
rect 4525 15521 4537 15555
rect 4571 15521 4583 15555
rect 4525 15515 4583 15521
rect 6178 15512 6184 15564
rect 6236 15512 6242 15564
rect 6288 15552 6316 15592
rect 6288 15524 10640 15552
rect 4617 15487 4675 15493
rect 4617 15484 4629 15487
rect 4448 15456 4629 15484
rect 4249 15447 4307 15453
rect 4617 15453 4629 15456
rect 4663 15484 4675 15487
rect 4798 15484 4804 15496
rect 4663 15456 4804 15484
rect 4663 15453 4675 15456
rect 4617 15447 4675 15453
rect 3896 15416 3924 15444
rect 4264 15416 4292 15447
rect 4798 15444 4804 15456
rect 4856 15444 4862 15496
rect 3896 15388 4292 15416
rect 6196 15416 6224 15512
rect 7834 15444 7840 15496
rect 7892 15484 7898 15496
rect 8941 15487 8999 15493
rect 8941 15484 8953 15487
rect 7892 15456 8953 15484
rect 7892 15444 7898 15456
rect 8941 15453 8953 15456
rect 8987 15453 8999 15487
rect 10612 15484 10640 15524
rect 11238 15512 11244 15564
rect 11296 15552 11302 15564
rect 11532 15561 11560 15660
rect 12526 15648 12532 15660
rect 12584 15648 12590 15700
rect 14182 15648 14188 15700
rect 14240 15688 14246 15700
rect 14277 15691 14335 15697
rect 14277 15688 14289 15691
rect 14240 15660 14289 15688
rect 14240 15648 14246 15660
rect 14277 15657 14289 15660
rect 14323 15657 14335 15691
rect 14277 15651 14335 15657
rect 14737 15691 14795 15697
rect 14737 15657 14749 15691
rect 14783 15688 14795 15691
rect 15470 15688 15476 15700
rect 14783 15660 15476 15688
rect 14783 15657 14795 15660
rect 14737 15651 14795 15657
rect 15470 15648 15476 15660
rect 15528 15648 15534 15700
rect 17770 15648 17776 15700
rect 17828 15688 17834 15700
rect 18141 15691 18199 15697
rect 18141 15688 18153 15691
rect 17828 15660 18153 15688
rect 17828 15648 17834 15660
rect 18141 15657 18153 15660
rect 18187 15657 18199 15691
rect 20809 15691 20867 15697
rect 18141 15651 18199 15657
rect 18248 15660 19196 15688
rect 14108 15592 16528 15620
rect 11517 15555 11575 15561
rect 11517 15552 11529 15555
rect 11296 15524 11529 15552
rect 11296 15512 11302 15524
rect 11517 15521 11529 15524
rect 11563 15521 11575 15555
rect 14108 15552 14136 15592
rect 16500 15564 16528 15592
rect 15473 15555 15531 15561
rect 15473 15552 15485 15555
rect 11517 15515 11575 15521
rect 11624 15524 14136 15552
rect 14200 15524 15485 15552
rect 11146 15484 11152 15496
rect 10612 15456 11152 15484
rect 8941 15447 8999 15453
rect 11146 15444 11152 15456
rect 11204 15444 11210 15496
rect 11422 15444 11428 15496
rect 11480 15444 11486 15496
rect 6362 15416 6368 15428
rect 6196 15388 6368 15416
rect 6362 15376 6368 15388
rect 6420 15376 6426 15428
rect 6454 15376 6460 15428
rect 6512 15376 6518 15428
rect 6914 15376 6920 15428
rect 6972 15376 6978 15428
rect 7760 15388 11008 15416
rect 5350 15308 5356 15360
rect 5408 15348 5414 15360
rect 7760 15348 7788 15388
rect 10980 15357 11008 15388
rect 5408 15320 7788 15348
rect 10965 15351 11023 15357
rect 5408 15308 5414 15320
rect 10965 15317 10977 15351
rect 11011 15317 11023 15351
rect 11164 15348 11192 15444
rect 11624 15428 11652 15524
rect 11882 15444 11888 15496
rect 11940 15444 11946 15496
rect 13909 15487 13967 15493
rect 13909 15453 13921 15487
rect 13955 15484 13967 15487
rect 14090 15484 14096 15496
rect 13955 15456 14096 15484
rect 13955 15453 13967 15456
rect 13909 15447 13967 15453
rect 14090 15444 14096 15456
rect 14148 15444 14154 15496
rect 14200 15493 14228 15524
rect 15473 15521 15485 15524
rect 15519 15521 15531 15555
rect 15473 15515 15531 15521
rect 15657 15555 15715 15561
rect 15657 15521 15669 15555
rect 15703 15552 15715 15555
rect 16209 15555 16267 15561
rect 16209 15552 16221 15555
rect 15703 15524 16221 15552
rect 15703 15521 15715 15524
rect 15657 15515 15715 15521
rect 16209 15521 16221 15524
rect 16255 15521 16267 15555
rect 16390 15552 16396 15564
rect 16209 15515 16267 15521
rect 16316 15524 16396 15552
rect 14185 15487 14243 15493
rect 14185 15453 14197 15487
rect 14231 15453 14243 15487
rect 14185 15447 14243 15453
rect 14553 15487 14611 15493
rect 14553 15453 14565 15487
rect 14599 15484 14611 15487
rect 14642 15484 14648 15496
rect 14599 15456 14648 15484
rect 14599 15453 14611 15456
rect 14553 15447 14611 15453
rect 14642 15444 14648 15456
rect 14700 15444 14706 15496
rect 15746 15444 15752 15496
rect 15804 15444 15810 15496
rect 15838 15444 15844 15496
rect 15896 15444 15902 15496
rect 15930 15444 15936 15496
rect 15988 15444 15994 15496
rect 16316 15493 16344 15524
rect 16390 15512 16396 15524
rect 16448 15512 16454 15564
rect 16482 15512 16488 15564
rect 16540 15512 16546 15564
rect 18248 15496 18276 15660
rect 18969 15623 19027 15629
rect 18969 15589 18981 15623
rect 19015 15620 19027 15623
rect 19058 15620 19064 15632
rect 19015 15592 19064 15620
rect 19015 15589 19027 15592
rect 18969 15583 19027 15589
rect 19058 15580 19064 15592
rect 19116 15580 19122 15632
rect 18598 15512 18604 15564
rect 18656 15552 18662 15564
rect 18785 15555 18843 15561
rect 18785 15552 18797 15555
rect 18656 15524 18797 15552
rect 18656 15512 18662 15524
rect 18785 15521 18797 15524
rect 18831 15521 18843 15555
rect 19168 15552 19196 15660
rect 20809 15657 20821 15691
rect 20855 15688 20867 15691
rect 21082 15688 21088 15700
rect 20855 15660 21088 15688
rect 20855 15657 20867 15660
rect 20809 15651 20867 15657
rect 21082 15648 21088 15660
rect 21140 15648 21146 15700
rect 24486 15648 24492 15700
rect 24544 15688 24550 15700
rect 26329 15691 26387 15697
rect 24544 15660 25452 15688
rect 24544 15648 24550 15660
rect 19242 15580 19248 15632
rect 19300 15620 19306 15632
rect 19300 15592 19656 15620
rect 19300 15580 19306 15592
rect 19168 15524 19380 15552
rect 18785 15515 18843 15521
rect 16117 15487 16175 15493
rect 16117 15486 16129 15487
rect 16040 15458 16129 15486
rect 11333 15419 11391 15425
rect 11333 15385 11345 15419
rect 11379 15416 11391 15419
rect 11606 15416 11612 15428
rect 11379 15388 11612 15416
rect 11379 15385 11391 15388
rect 11333 15379 11391 15385
rect 11606 15376 11612 15388
rect 11664 15376 11670 15428
rect 12161 15419 12219 15425
rect 12161 15385 12173 15419
rect 12207 15416 12219 15419
rect 12434 15416 12440 15428
rect 12207 15388 12440 15416
rect 12207 15385 12219 15388
rect 12161 15379 12219 15385
rect 12434 15376 12440 15388
rect 12492 15376 12498 15428
rect 12544 15388 12650 15416
rect 12544 15348 12572 15388
rect 13814 15376 13820 15428
rect 13872 15416 13878 15428
rect 14734 15416 14740 15428
rect 13872 15388 14740 15416
rect 13872 15376 13878 15388
rect 14734 15376 14740 15388
rect 14792 15376 14798 15428
rect 15654 15376 15660 15428
rect 15712 15416 15718 15428
rect 15856 15416 15884 15444
rect 15712 15388 15884 15416
rect 15712 15376 15718 15388
rect 11164 15320 12572 15348
rect 14752 15348 14780 15376
rect 16040 15348 16068 15458
rect 16117 15453 16129 15458
rect 16163 15453 16175 15487
rect 16117 15447 16175 15453
rect 16301 15487 16359 15493
rect 16301 15453 16313 15487
rect 16347 15453 16359 15487
rect 16301 15447 16359 15453
rect 18230 15444 18236 15496
rect 18288 15444 18294 15496
rect 19352 15493 19380 15524
rect 19062 15487 19120 15493
rect 19062 15453 19074 15487
rect 19108 15453 19120 15487
rect 19062 15447 19120 15453
rect 19337 15487 19395 15493
rect 19337 15453 19349 15487
rect 19383 15453 19395 15487
rect 19628 15484 19656 15592
rect 23768 15592 24992 15620
rect 20622 15512 20628 15564
rect 20680 15552 20686 15564
rect 22646 15552 22652 15564
rect 20680 15524 22652 15552
rect 20680 15512 20686 15524
rect 22646 15512 22652 15524
rect 22704 15512 22710 15564
rect 22738 15512 22744 15564
rect 22796 15552 22802 15564
rect 23768 15552 23796 15592
rect 22796 15524 23428 15552
rect 22796 15512 22802 15524
rect 19981 15487 20039 15493
rect 19981 15484 19993 15487
rect 19628 15456 19993 15484
rect 19337 15447 19395 15453
rect 19981 15453 19993 15456
rect 20027 15453 20039 15487
rect 19981 15447 20039 15453
rect 20717 15487 20775 15493
rect 20717 15453 20729 15487
rect 20763 15453 20775 15487
rect 20717 15447 20775 15453
rect 18417 15419 18475 15425
rect 18417 15385 18429 15419
rect 18463 15385 18475 15419
rect 18417 15379 18475 15385
rect 14752 15320 16068 15348
rect 18432 15348 18460 15379
rect 18690 15376 18696 15428
rect 18748 15416 18754 15428
rect 19077 15416 19105 15447
rect 19610 15416 19616 15428
rect 18748 15388 19012 15416
rect 19077 15388 19616 15416
rect 18748 15376 18754 15388
rect 18601 15351 18659 15357
rect 18601 15348 18613 15351
rect 18432 15320 18613 15348
rect 10965 15311 11023 15317
rect 18601 15317 18613 15320
rect 18647 15348 18659 15351
rect 18782 15348 18788 15360
rect 18647 15320 18788 15348
rect 18647 15317 18659 15320
rect 18601 15311 18659 15317
rect 18782 15308 18788 15320
rect 18840 15308 18846 15360
rect 18984 15348 19012 15388
rect 19610 15376 19616 15388
rect 19668 15376 19674 15428
rect 20070 15376 20076 15428
rect 20128 15416 20134 15428
rect 20530 15416 20536 15428
rect 20128 15388 20536 15416
rect 20128 15376 20134 15388
rect 20530 15376 20536 15388
rect 20588 15416 20594 15428
rect 20732 15416 20760 15447
rect 22002 15444 22008 15496
rect 22060 15484 22066 15496
rect 22925 15487 22983 15493
rect 22925 15484 22937 15487
rect 22060 15456 22937 15484
rect 22060 15444 22066 15456
rect 22925 15453 22937 15456
rect 22971 15453 22983 15487
rect 22925 15447 22983 15453
rect 23014 15444 23020 15496
rect 23072 15484 23078 15496
rect 23400 15493 23428 15524
rect 23584 15524 23796 15552
rect 23109 15487 23167 15493
rect 23109 15484 23121 15487
rect 23072 15456 23121 15484
rect 23072 15444 23078 15456
rect 23109 15453 23121 15456
rect 23155 15453 23167 15487
rect 23109 15447 23167 15453
rect 23385 15487 23443 15493
rect 23385 15453 23397 15487
rect 23431 15453 23443 15487
rect 23385 15447 23443 15453
rect 23584 15428 23612 15524
rect 23768 15493 23796 15524
rect 23661 15487 23719 15493
rect 23661 15453 23673 15487
rect 23707 15453 23719 15487
rect 23661 15447 23719 15453
rect 23753 15487 23811 15493
rect 23753 15453 23765 15487
rect 23799 15453 23811 15487
rect 23753 15447 23811 15453
rect 20588 15388 20760 15416
rect 20588 15376 20594 15388
rect 23566 15376 23572 15428
rect 23624 15376 23630 15428
rect 23676 15416 23704 15447
rect 24486 15444 24492 15496
rect 24544 15444 24550 15496
rect 24670 15444 24676 15496
rect 24728 15484 24734 15496
rect 24964 15493 24992 15592
rect 24765 15487 24823 15493
rect 24765 15484 24777 15487
rect 24728 15456 24777 15484
rect 24728 15444 24734 15456
rect 24765 15453 24777 15456
rect 24811 15453 24823 15487
rect 24765 15447 24823 15453
rect 24949 15487 25007 15493
rect 24949 15453 24961 15487
rect 24995 15484 25007 15487
rect 25222 15484 25228 15496
rect 24995 15456 25228 15484
rect 24995 15453 25007 15456
rect 24949 15447 25007 15453
rect 25222 15444 25228 15456
rect 25280 15444 25286 15496
rect 25424 15493 25452 15660
rect 26329 15657 26341 15691
rect 26375 15688 26387 15691
rect 27338 15688 27344 15700
rect 26375 15660 27344 15688
rect 26375 15657 26387 15660
rect 26329 15651 26387 15657
rect 27338 15648 27344 15660
rect 27396 15648 27402 15700
rect 30742 15648 30748 15700
rect 30800 15648 30806 15700
rect 31386 15648 31392 15700
rect 31444 15648 31450 15700
rect 32214 15648 32220 15700
rect 32272 15688 32278 15700
rect 32309 15691 32367 15697
rect 32309 15688 32321 15691
rect 32272 15660 32321 15688
rect 32272 15648 32278 15660
rect 32309 15657 32321 15660
rect 32355 15657 32367 15691
rect 32309 15651 32367 15657
rect 32490 15648 32496 15700
rect 32548 15688 32554 15700
rect 32769 15691 32827 15697
rect 32769 15688 32781 15691
rect 32548 15660 32781 15688
rect 32548 15648 32554 15660
rect 32769 15657 32781 15660
rect 32815 15657 32827 15691
rect 32769 15651 32827 15657
rect 32858 15648 32864 15700
rect 32916 15688 32922 15700
rect 33229 15691 33287 15697
rect 33229 15688 33241 15691
rect 32916 15660 33241 15688
rect 32916 15648 32922 15660
rect 33229 15657 33241 15660
rect 33275 15657 33287 15691
rect 33229 15651 33287 15657
rect 34698 15648 34704 15700
rect 34756 15648 34762 15700
rect 35161 15691 35219 15697
rect 35161 15657 35173 15691
rect 35207 15688 35219 15691
rect 35342 15688 35348 15700
rect 35207 15660 35348 15688
rect 35207 15657 35219 15660
rect 35161 15651 35219 15657
rect 35342 15648 35348 15660
rect 35400 15648 35406 15700
rect 35437 15691 35495 15697
rect 35437 15657 35449 15691
rect 35483 15657 35495 15691
rect 35437 15651 35495 15657
rect 27709 15555 27767 15561
rect 27709 15521 27721 15555
rect 27755 15552 27767 15555
rect 27985 15555 28043 15561
rect 27985 15552 27997 15555
rect 27755 15524 27997 15552
rect 27755 15521 27767 15524
rect 27709 15515 27767 15521
rect 27985 15521 27997 15524
rect 28031 15521 28043 15555
rect 27985 15515 28043 15521
rect 29178 15512 29184 15564
rect 29236 15552 29242 15564
rect 29546 15552 29552 15564
rect 29236 15524 29552 15552
rect 29236 15512 29242 15524
rect 29546 15512 29552 15524
rect 29604 15552 29610 15564
rect 29604 15524 29868 15552
rect 29604 15512 29610 15524
rect 25409 15487 25467 15493
rect 25409 15453 25421 15487
rect 25455 15453 25467 15487
rect 25409 15447 25467 15453
rect 25498 15444 25504 15496
rect 25556 15484 25562 15496
rect 25958 15484 25964 15496
rect 25556 15456 25964 15484
rect 25556 15444 25562 15456
rect 25958 15444 25964 15456
rect 26016 15444 26022 15496
rect 26050 15444 26056 15496
rect 26108 15484 26114 15496
rect 26145 15487 26203 15493
rect 26145 15484 26157 15487
rect 26108 15456 26157 15484
rect 26108 15444 26114 15456
rect 26145 15453 26157 15456
rect 26191 15453 26203 15487
rect 26145 15447 26203 15453
rect 26234 15444 26240 15496
rect 26292 15484 26298 15496
rect 26421 15487 26479 15493
rect 26421 15484 26433 15487
rect 26292 15456 26433 15484
rect 26292 15444 26298 15456
rect 26421 15453 26433 15456
rect 26467 15453 26479 15487
rect 26421 15447 26479 15453
rect 27154 15444 27160 15496
rect 27212 15484 27218 15496
rect 27614 15484 27620 15496
rect 27212 15456 27620 15484
rect 27212 15444 27218 15456
rect 27614 15444 27620 15456
rect 27672 15444 27678 15496
rect 28169 15487 28227 15493
rect 28169 15453 28181 15487
rect 28215 15453 28227 15487
rect 28169 15447 28227 15453
rect 28445 15487 28503 15493
rect 28445 15453 28457 15487
rect 28491 15484 28503 15487
rect 28629 15487 28687 15493
rect 28629 15484 28641 15487
rect 28491 15456 28641 15484
rect 28491 15453 28503 15456
rect 28445 15447 28503 15453
rect 28629 15453 28641 15456
rect 28675 15453 28687 15487
rect 28629 15447 28687 15453
rect 28721 15487 28779 15493
rect 28721 15453 28733 15487
rect 28767 15484 28779 15487
rect 29638 15484 29644 15496
rect 28767 15456 29644 15484
rect 28767 15453 28779 15456
rect 28721 15447 28779 15453
rect 25314 15416 25320 15428
rect 23676 15388 25320 15416
rect 25314 15376 25320 15388
rect 25372 15376 25378 15428
rect 28184 15416 28212 15447
rect 29638 15444 29644 15456
rect 29696 15444 29702 15496
rect 29840 15493 29868 15524
rect 29825 15487 29883 15493
rect 29825 15453 29837 15487
rect 29871 15453 29883 15487
rect 30760 15484 30788 15648
rect 31404 15552 31432 15648
rect 32401 15623 32459 15629
rect 32401 15589 32413 15623
rect 32447 15620 32459 15623
rect 34716 15620 34744 15648
rect 35452 15620 35480 15651
rect 32447 15592 33456 15620
rect 34716 15592 35480 15620
rect 32447 15589 32459 15592
rect 32401 15583 32459 15589
rect 31849 15555 31907 15561
rect 31404 15524 31708 15552
rect 31680 15493 31708 15524
rect 31849 15521 31861 15555
rect 31895 15552 31907 15555
rect 32217 15555 32275 15561
rect 32217 15552 32229 15555
rect 31895 15524 32229 15552
rect 31895 15521 31907 15524
rect 31849 15515 31907 15521
rect 32217 15521 32229 15524
rect 32263 15552 32275 15555
rect 33321 15555 33379 15561
rect 33321 15552 33333 15555
rect 32263 15524 33333 15552
rect 32263 15521 32275 15524
rect 32217 15515 32275 15521
rect 33321 15521 33333 15524
rect 33367 15521 33379 15555
rect 33321 15515 33379 15521
rect 33428 15496 33456 15592
rect 34514 15512 34520 15564
rect 34572 15552 34578 15564
rect 34572 15524 34744 15552
rect 34572 15512 34578 15524
rect 31481 15487 31539 15493
rect 31481 15484 31493 15487
rect 30760 15456 31493 15484
rect 29825 15447 29883 15453
rect 31481 15453 31493 15456
rect 31527 15453 31539 15487
rect 31481 15447 31539 15453
rect 31665 15487 31723 15493
rect 31665 15453 31677 15487
rect 31711 15453 31723 15487
rect 31665 15447 31723 15453
rect 32493 15487 32551 15493
rect 32493 15453 32505 15487
rect 32539 15484 32551 15487
rect 32858 15484 32864 15496
rect 32539 15456 32864 15484
rect 32539 15453 32551 15456
rect 32493 15447 32551 15453
rect 32858 15444 32864 15456
rect 32916 15444 32922 15496
rect 33410 15444 33416 15496
rect 33468 15444 33474 15496
rect 34606 15444 34612 15496
rect 34664 15444 34670 15496
rect 34716 15484 34744 15524
rect 34790 15512 34796 15564
rect 34848 15512 34854 15564
rect 35342 15512 35348 15564
rect 35400 15552 35406 15564
rect 35621 15555 35679 15561
rect 35621 15552 35633 15555
rect 35400 15524 35633 15552
rect 35400 15512 35406 15524
rect 35621 15521 35633 15524
rect 35667 15521 35679 15555
rect 35621 15515 35679 15521
rect 34885 15487 34943 15493
rect 34885 15484 34897 15487
rect 34716 15456 34897 15484
rect 34885 15453 34897 15456
rect 34931 15453 34943 15487
rect 34885 15447 34943 15453
rect 35713 15487 35771 15493
rect 35713 15453 35725 15487
rect 35759 15453 35771 15487
rect 35713 15447 35771 15453
rect 30742 15416 30748 15428
rect 26712 15388 27476 15416
rect 28184 15388 30748 15416
rect 26712 15360 26740 15388
rect 19150 15348 19156 15360
rect 18984 15320 19156 15348
rect 19150 15308 19156 15320
rect 19208 15348 19214 15360
rect 22922 15348 22928 15360
rect 19208 15320 22928 15348
rect 19208 15308 19214 15320
rect 22922 15308 22928 15320
rect 22980 15308 22986 15360
rect 24670 15308 24676 15360
rect 24728 15348 24734 15360
rect 25498 15348 25504 15360
rect 24728 15320 25504 15348
rect 24728 15308 24734 15320
rect 25498 15308 25504 15320
rect 25556 15308 25562 15360
rect 25593 15351 25651 15357
rect 25593 15317 25605 15351
rect 25639 15348 25651 15351
rect 25682 15348 25688 15360
rect 25639 15320 25688 15348
rect 25639 15317 25651 15320
rect 25593 15311 25651 15317
rect 25682 15308 25688 15320
rect 25740 15308 25746 15360
rect 26605 15351 26663 15357
rect 26605 15317 26617 15351
rect 26651 15348 26663 15351
rect 26694 15348 26700 15360
rect 26651 15320 26700 15348
rect 26651 15317 26663 15320
rect 26605 15311 26663 15317
rect 26694 15308 26700 15320
rect 26752 15308 26758 15360
rect 27249 15351 27307 15357
rect 27249 15317 27261 15351
rect 27295 15348 27307 15351
rect 27338 15348 27344 15360
rect 27295 15320 27344 15348
rect 27295 15317 27307 15320
rect 27249 15311 27307 15317
rect 27338 15308 27344 15320
rect 27396 15308 27402 15360
rect 27448 15348 27476 15388
rect 30742 15376 30748 15388
rect 30800 15376 30806 15428
rect 32214 15376 32220 15428
rect 32272 15416 32278 15428
rect 32737 15419 32795 15425
rect 32737 15416 32749 15419
rect 32272 15388 32749 15416
rect 32272 15376 32278 15388
rect 32737 15385 32749 15388
rect 32783 15385 32795 15419
rect 32737 15379 32795 15385
rect 32953 15419 33011 15425
rect 32953 15385 32965 15419
rect 32999 15416 33011 15419
rect 34624 15416 34652 15444
rect 35728 15416 35756 15447
rect 32999 15388 33088 15416
rect 34624 15388 35756 15416
rect 32999 15385 33011 15388
rect 32953 15379 33011 15385
rect 28350 15348 28356 15360
rect 27448 15320 28356 15348
rect 28350 15308 28356 15320
rect 28408 15308 28414 15360
rect 30466 15308 30472 15360
rect 30524 15348 30530 15360
rect 30653 15351 30711 15357
rect 30653 15348 30665 15351
rect 30524 15320 30665 15348
rect 30524 15308 30530 15320
rect 30653 15317 30665 15320
rect 30699 15317 30711 15351
rect 30653 15311 30711 15317
rect 32582 15308 32588 15360
rect 32640 15308 32646 15360
rect 33060 15357 33088 15388
rect 33045 15351 33103 15357
rect 33045 15317 33057 15351
rect 33091 15317 33103 15351
rect 33045 15311 33103 15317
rect 1104 15258 38272 15280
rect 1104 15206 4874 15258
rect 4926 15206 4938 15258
rect 4990 15206 5002 15258
rect 5054 15206 5066 15258
rect 5118 15206 5130 15258
rect 5182 15206 35594 15258
rect 35646 15206 35658 15258
rect 35710 15206 35722 15258
rect 35774 15206 35786 15258
rect 35838 15206 35850 15258
rect 35902 15206 38272 15258
rect 1104 15184 38272 15206
rect 2961 15147 3019 15153
rect 2961 15113 2973 15147
rect 3007 15144 3019 15147
rect 3697 15147 3755 15153
rect 3697 15144 3709 15147
rect 3007 15116 3709 15144
rect 3007 15113 3019 15116
rect 2961 15107 3019 15113
rect 3697 15113 3709 15116
rect 3743 15113 3755 15147
rect 3697 15107 3755 15113
rect 4065 15147 4123 15153
rect 4065 15113 4077 15147
rect 4111 15144 4123 15147
rect 5350 15144 5356 15156
rect 4111 15116 5356 15144
rect 4111 15113 4123 15116
rect 4065 15107 4123 15113
rect 5350 15104 5356 15116
rect 5408 15104 5414 15156
rect 6454 15104 6460 15156
rect 6512 15144 6518 15156
rect 6641 15147 6699 15153
rect 6641 15144 6653 15147
rect 6512 15116 6653 15144
rect 6512 15104 6518 15116
rect 6641 15113 6653 15116
rect 6687 15113 6699 15147
rect 6641 15107 6699 15113
rect 7561 15147 7619 15153
rect 7561 15113 7573 15147
rect 7607 15144 7619 15147
rect 7926 15144 7932 15156
rect 7607 15116 7932 15144
rect 7607 15113 7619 15116
rect 7561 15107 7619 15113
rect 7926 15104 7932 15116
rect 7984 15104 7990 15156
rect 8202 15144 8208 15156
rect 8036 15116 8208 15144
rect 4154 15076 4160 15088
rect 3436 15048 4160 15076
rect 2869 15011 2927 15017
rect 2869 14977 2881 15011
rect 2915 15008 2927 15011
rect 3234 15008 3240 15020
rect 2915 14980 3240 15008
rect 2915 14977 2927 14980
rect 2869 14971 2927 14977
rect 3234 14968 3240 14980
rect 3292 15008 3298 15020
rect 3436 15017 3464 15048
rect 4154 15036 4160 15048
rect 4212 15076 4218 15088
rect 4212 15048 4568 15076
rect 4212 15036 4218 15048
rect 3421 15011 3479 15017
rect 3421 15008 3433 15011
rect 3292 14980 3433 15008
rect 3292 14968 3298 14980
rect 3421 14977 3433 14980
rect 3467 14977 3479 15011
rect 3421 14971 3479 14977
rect 3605 15011 3663 15017
rect 3605 14977 3617 15011
rect 3651 15008 3663 15011
rect 3970 15008 3976 15020
rect 3651 14980 3976 15008
rect 3651 14977 3663 14980
rect 3605 14971 3663 14977
rect 3970 14968 3976 14980
rect 4028 15008 4034 15020
rect 4028 14980 4384 15008
rect 4028 14968 4034 14980
rect 3142 14900 3148 14952
rect 3200 14900 3206 14952
rect 4157 14943 4215 14949
rect 4157 14940 4169 14943
rect 4080 14912 4169 14940
rect 4080 14884 4108 14912
rect 4157 14909 4169 14912
rect 4203 14909 4215 14943
rect 4157 14903 4215 14909
rect 4246 14900 4252 14952
rect 4304 14900 4310 14952
rect 4062 14832 4068 14884
rect 4120 14832 4126 14884
rect 2498 14764 2504 14816
rect 2556 14764 2562 14816
rect 3602 14764 3608 14816
rect 3660 14764 3666 14816
rect 3878 14764 3884 14816
rect 3936 14804 3942 14816
rect 4264 14804 4292 14900
rect 4356 14872 4384 14980
rect 4540 14949 4568 15048
rect 4614 15036 4620 15088
rect 4672 15076 4678 15088
rect 4893 15079 4951 15085
rect 4893 15076 4905 15079
rect 4672 15048 4905 15076
rect 4672 15036 4678 15048
rect 4893 15045 4905 15048
rect 4939 15045 4951 15079
rect 4893 15039 4951 15045
rect 4706 14968 4712 15020
rect 4764 14968 4770 15020
rect 8036 15017 8064 15116
rect 8202 15104 8208 15116
rect 8260 15104 8266 15156
rect 8570 15104 8576 15156
rect 8628 15104 8634 15156
rect 8754 15104 8760 15156
rect 8812 15104 8818 15156
rect 9214 15104 9220 15156
rect 9272 15104 9278 15156
rect 12434 15104 12440 15156
rect 12492 15144 12498 15156
rect 13909 15147 13967 15153
rect 13909 15144 13921 15147
rect 12492 15116 13921 15144
rect 12492 15104 12498 15116
rect 13909 15113 13921 15116
rect 13955 15113 13967 15147
rect 15562 15144 15568 15156
rect 13909 15107 13967 15113
rect 14200 15116 15568 15144
rect 8588 15076 8616 15104
rect 8128 15048 8616 15076
rect 8128 15017 8156 15048
rect 6825 15011 6883 15017
rect 6825 14977 6837 15011
rect 6871 15008 6883 15011
rect 7469 15011 7527 15017
rect 6871 14980 7144 15008
rect 6871 14977 6883 14980
rect 6825 14971 6883 14977
rect 4525 14943 4583 14949
rect 4525 14909 4537 14943
rect 4571 14909 4583 14943
rect 4525 14903 4583 14909
rect 4724 14872 4752 14968
rect 7116 14881 7144 14980
rect 7469 14977 7481 15011
rect 7515 14977 7527 15011
rect 7469 14971 7527 14977
rect 8021 15011 8079 15017
rect 8021 14977 8033 15011
rect 8067 14977 8079 15011
rect 8021 14971 8079 14977
rect 8113 15011 8171 15017
rect 8113 14977 8125 15011
rect 8159 14977 8171 15011
rect 8113 14971 8171 14977
rect 4356 14844 4752 14872
rect 7101 14875 7159 14881
rect 7101 14841 7113 14875
rect 7147 14841 7159 14875
rect 7101 14835 7159 14841
rect 3936 14776 4292 14804
rect 7484 14804 7512 14971
rect 8386 14968 8392 15020
rect 8444 15008 8450 15020
rect 8772 15008 8800 15104
rect 9033 15079 9091 15085
rect 9033 15076 9045 15079
rect 8956 15048 9045 15076
rect 8956 15020 8984 15048
rect 9033 15045 9045 15048
rect 9079 15045 9091 15079
rect 9033 15039 9091 15045
rect 8444 14980 8800 15008
rect 8444 14968 8450 14980
rect 8938 14968 8944 15020
rect 8996 14968 9002 15020
rect 9232 15008 9260 15104
rect 9582 15036 9588 15088
rect 9640 15076 9646 15088
rect 11054 15076 11060 15088
rect 9640 15048 11060 15076
rect 9640 15036 9646 15048
rect 11054 15036 11060 15048
rect 11112 15076 11118 15088
rect 11885 15079 11943 15085
rect 11885 15076 11897 15079
rect 11112 15048 11897 15076
rect 11112 15036 11118 15048
rect 11885 15045 11897 15048
rect 11931 15045 11943 15079
rect 11885 15039 11943 15045
rect 11977 15079 12035 15085
rect 11977 15045 11989 15079
rect 12023 15076 12035 15079
rect 12066 15076 12072 15088
rect 12023 15048 12072 15076
rect 12023 15045 12035 15048
rect 11977 15039 12035 15045
rect 12066 15036 12072 15048
rect 12124 15076 12130 15088
rect 12894 15076 12900 15088
rect 12124 15048 12900 15076
rect 12124 15036 12130 15048
rect 12894 15036 12900 15048
rect 12952 15036 12958 15088
rect 10505 15011 10563 15017
rect 9232 14980 9628 15008
rect 7650 14900 7656 14952
rect 7708 14900 7714 14952
rect 9398 14940 9404 14952
rect 8312 14912 9404 14940
rect 8312 14813 8340 14912
rect 9398 14900 9404 14912
rect 9456 14940 9462 14952
rect 9600 14949 9628 14980
rect 10505 14977 10517 15011
rect 10551 15008 10563 15011
rect 10551 14980 11560 15008
rect 10551 14977 10563 14980
rect 10505 14971 10563 14977
rect 9493 14943 9551 14949
rect 9493 14940 9505 14943
rect 9456 14912 9505 14940
rect 9456 14900 9462 14912
rect 9493 14909 9505 14912
rect 9539 14909 9551 14943
rect 9493 14903 9551 14909
rect 9585 14943 9643 14949
rect 9585 14909 9597 14943
rect 9631 14909 9643 14943
rect 9585 14903 9643 14909
rect 9030 14832 9036 14884
rect 9088 14832 9094 14884
rect 11532 14881 11560 14980
rect 12986 14968 12992 15020
rect 13044 14968 13050 15020
rect 13354 14968 13360 15020
rect 13412 14968 13418 15020
rect 14090 14968 14096 15020
rect 14148 14968 14154 15020
rect 14200 15017 14228 15116
rect 15562 15104 15568 15116
rect 15620 15104 15626 15156
rect 15749 15147 15807 15153
rect 15749 15113 15761 15147
rect 15795 15144 15807 15147
rect 16390 15144 16396 15156
rect 15795 15116 16396 15144
rect 15795 15113 15807 15116
rect 15749 15107 15807 15113
rect 16390 15104 16396 15116
rect 16448 15104 16454 15156
rect 16482 15104 16488 15156
rect 16540 15104 16546 15156
rect 19058 15144 19064 15156
rect 16776 15116 19064 15144
rect 14737 15079 14795 15085
rect 14737 15045 14749 15079
rect 14783 15076 14795 15079
rect 15013 15079 15071 15085
rect 15013 15076 15025 15079
rect 14783 15048 15025 15076
rect 14783 15045 14795 15048
rect 14737 15039 14795 15045
rect 15013 15045 15025 15048
rect 15059 15045 15071 15079
rect 16114 15076 16120 15088
rect 15013 15039 15071 15045
rect 15580 15048 16120 15076
rect 14185 15011 14243 15017
rect 14185 14977 14197 15011
rect 14231 14977 14243 15011
rect 14185 14971 14243 14977
rect 14277 15011 14335 15017
rect 14277 14977 14289 15011
rect 14323 14977 14335 15011
rect 14277 14971 14335 14977
rect 12161 14943 12219 14949
rect 12161 14909 12173 14943
rect 12207 14940 12219 14943
rect 12526 14940 12532 14952
rect 12207 14912 12532 14940
rect 12207 14909 12219 14912
rect 12161 14903 12219 14909
rect 12526 14900 12532 14912
rect 12584 14900 12590 14952
rect 11517 14875 11575 14881
rect 11517 14841 11529 14875
rect 11563 14841 11575 14875
rect 11517 14835 11575 14841
rect 12250 14832 12256 14884
rect 12308 14872 12314 14884
rect 14200 14872 14228 14971
rect 14292 14940 14320 14971
rect 14366 14968 14372 15020
rect 14424 15008 14430 15020
rect 14461 15011 14519 15017
rect 14461 15008 14473 15011
rect 14424 14980 14473 15008
rect 14424 14968 14430 14980
rect 14461 14977 14473 14980
rect 14507 14977 14519 15011
rect 14461 14971 14519 14977
rect 14553 15011 14611 15017
rect 14553 14977 14565 15011
rect 14599 14977 14611 15011
rect 14553 14971 14611 14977
rect 14292 14912 14504 14940
rect 14476 14884 14504 14912
rect 12308 14844 14228 14872
rect 12308 14832 12314 14844
rect 14458 14832 14464 14884
rect 14516 14832 14522 14884
rect 14568 14872 14596 14971
rect 14826 14968 14832 15020
rect 14884 14968 14890 15020
rect 15105 15011 15163 15017
rect 15105 14977 15117 15011
rect 15151 14977 15163 15011
rect 15105 14971 15163 14977
rect 14642 14900 14648 14952
rect 14700 14940 14706 14952
rect 14700 14912 14872 14940
rect 14700 14900 14706 14912
rect 14734 14872 14740 14884
rect 14568 14844 14740 14872
rect 14734 14832 14740 14844
rect 14792 14832 14798 14884
rect 14844 14881 14872 14912
rect 14829 14875 14887 14881
rect 14829 14841 14841 14875
rect 14875 14841 14887 14875
rect 15120 14872 15148 14971
rect 15378 14968 15384 15020
rect 15436 14968 15442 15020
rect 15580 15017 15608 15048
rect 16114 15036 16120 15048
rect 16172 15036 16178 15088
rect 15565 15011 15623 15017
rect 15565 14977 15577 15011
rect 15611 14977 15623 15011
rect 15565 14971 15623 14977
rect 16206 14968 16212 15020
rect 16264 14968 16270 15020
rect 16408 15008 16436 15104
rect 16500 15076 16528 15104
rect 16776 15076 16804 15116
rect 19058 15104 19064 15116
rect 19116 15104 19122 15156
rect 20162 15104 20168 15156
rect 20220 15104 20226 15156
rect 26050 15104 26056 15156
rect 26108 15104 26114 15156
rect 27065 15147 27123 15153
rect 27065 15113 27077 15147
rect 27111 15144 27123 15147
rect 27338 15144 27344 15156
rect 27111 15116 27344 15144
rect 27111 15113 27123 15116
rect 27065 15107 27123 15113
rect 27338 15104 27344 15116
rect 27396 15144 27402 15156
rect 27706 15144 27712 15156
rect 27396 15116 27712 15144
rect 27396 15104 27402 15116
rect 27706 15104 27712 15116
rect 27764 15104 27770 15156
rect 32582 15144 32588 15156
rect 27816 15116 32588 15144
rect 16500 15048 16804 15076
rect 16776 15017 16804 15048
rect 17862 15036 17868 15088
rect 17920 15076 17926 15088
rect 24210 15076 24216 15088
rect 17920 15048 24216 15076
rect 17920 15036 17926 15048
rect 24210 15036 24216 15048
rect 24268 15036 24274 15088
rect 26068 15076 26096 15104
rect 25516 15048 26096 15076
rect 16485 15011 16543 15017
rect 16485 15008 16497 15011
rect 16408 14980 16497 15008
rect 16485 14977 16497 14980
rect 16531 14977 16543 15011
rect 16485 14971 16543 14977
rect 16761 15011 16819 15017
rect 16761 14977 16773 15011
rect 16807 14977 16819 15011
rect 16761 14971 16819 14977
rect 17034 14968 17040 15020
rect 17092 14968 17098 15020
rect 17129 15011 17187 15017
rect 17129 14977 17141 15011
rect 17175 14977 17187 15011
rect 17129 14971 17187 14977
rect 16298 14900 16304 14952
rect 16356 14940 16362 14952
rect 17144 14940 17172 14971
rect 17586 14968 17592 15020
rect 17644 14968 17650 15020
rect 17678 14968 17684 15020
rect 17736 14968 17742 15020
rect 18230 14968 18236 15020
rect 18288 14968 18294 15020
rect 18598 14968 18604 15020
rect 18656 15008 18662 15020
rect 18785 15011 18843 15017
rect 18785 15008 18797 15011
rect 18656 14980 18797 15008
rect 18656 14968 18662 14980
rect 18785 14977 18797 14980
rect 18831 14977 18843 15011
rect 18785 14971 18843 14977
rect 19058 14968 19064 15020
rect 19116 15008 19122 15020
rect 19153 15011 19211 15017
rect 19153 15008 19165 15011
rect 19116 14980 19165 15008
rect 19116 14968 19122 14980
rect 19153 14977 19165 14980
rect 19199 14977 19211 15011
rect 19153 14971 19211 14977
rect 19610 14968 19616 15020
rect 19668 14968 19674 15020
rect 20070 14968 20076 15020
rect 20128 14968 20134 15020
rect 20349 15011 20407 15017
rect 20349 14977 20361 15011
rect 20395 15008 20407 15011
rect 20990 15008 20996 15020
rect 20395 14980 20996 15008
rect 20395 14977 20407 14980
rect 20349 14971 20407 14977
rect 16356 14912 17172 14940
rect 16356 14900 16362 14912
rect 18690 14900 18696 14952
rect 18748 14900 18754 14952
rect 19426 14900 19432 14952
rect 19484 14940 19490 14952
rect 20088 14940 20116 14968
rect 19484 14912 20116 14940
rect 19484 14900 19490 14912
rect 15933 14875 15991 14881
rect 15933 14872 15945 14875
rect 15120 14844 15945 14872
rect 14829 14835 14887 14841
rect 15933 14841 15945 14844
rect 15979 14841 15991 14875
rect 20364 14872 20392 14971
rect 20990 14968 20996 14980
rect 21048 14968 21054 15020
rect 21910 14968 21916 15020
rect 21968 15008 21974 15020
rect 25516 15017 25544 15048
rect 22005 15011 22063 15017
rect 22005 15008 22017 15011
rect 21968 14980 22017 15008
rect 21968 14968 21974 14980
rect 22005 14977 22017 14980
rect 22051 14977 22063 15011
rect 22005 14971 22063 14977
rect 22189 15011 22247 15017
rect 22189 14977 22201 15011
rect 22235 15008 22247 15011
rect 22649 15011 22707 15017
rect 22649 15008 22661 15011
rect 22235 14980 22661 15008
rect 22235 14977 22247 14980
rect 22189 14971 22247 14977
rect 22649 14977 22661 14980
rect 22695 14977 22707 15011
rect 22649 14971 22707 14977
rect 25501 15011 25559 15017
rect 25501 14977 25513 15011
rect 25547 14977 25559 15011
rect 25501 14971 25559 14977
rect 25682 14968 25688 15020
rect 25740 15008 25746 15020
rect 25777 15011 25835 15017
rect 25777 15008 25789 15011
rect 25740 14980 25789 15008
rect 25740 14968 25746 14980
rect 25777 14977 25789 14980
rect 25823 14977 25835 15011
rect 25777 14971 25835 14977
rect 25961 15011 26019 15017
rect 25961 14977 25973 15011
rect 26007 15008 26019 15011
rect 26068 15008 26096 15048
rect 26007 14980 26096 15008
rect 26007 14977 26019 14980
rect 25961 14971 26019 14977
rect 21818 14900 21824 14952
rect 21876 14900 21882 14952
rect 23201 14943 23259 14949
rect 23201 14909 23213 14943
rect 23247 14940 23259 14943
rect 23290 14940 23296 14952
rect 23247 14912 23296 14940
rect 23247 14909 23259 14912
rect 23201 14903 23259 14909
rect 23290 14900 23296 14912
rect 23348 14940 23354 14952
rect 25590 14940 25596 14952
rect 23348 14912 25596 14940
rect 23348 14900 23354 14912
rect 25590 14900 25596 14912
rect 25648 14900 25654 14952
rect 25792 14940 25820 14971
rect 26418 14968 26424 15020
rect 26476 15008 26482 15020
rect 26973 15011 27031 15017
rect 26973 15008 26985 15011
rect 26476 14980 26985 15008
rect 26476 14968 26482 14980
rect 26973 14977 26985 14980
rect 27019 14977 27031 15011
rect 26973 14971 27031 14977
rect 27154 14968 27160 15020
rect 27212 15008 27218 15020
rect 27816 15017 27844 15116
rect 32582 15104 32588 15116
rect 32640 15104 32646 15156
rect 34333 15147 34391 15153
rect 34333 15113 34345 15147
rect 34379 15144 34391 15147
rect 34790 15144 34796 15156
rect 34379 15116 34796 15144
rect 34379 15113 34391 15116
rect 34333 15107 34391 15113
rect 34790 15104 34796 15116
rect 34848 15104 34854 15156
rect 27982 15036 27988 15088
rect 28040 15076 28046 15088
rect 28997 15079 29055 15085
rect 28040 15048 28488 15076
rect 28040 15036 28046 15048
rect 27249 15011 27307 15017
rect 27249 15008 27261 15011
rect 27212 14980 27261 15008
rect 27212 14968 27218 14980
rect 27249 14977 27261 14980
rect 27295 14977 27307 15011
rect 27249 14971 27307 14977
rect 27801 15011 27859 15017
rect 27801 14977 27813 15011
rect 27847 14977 27859 15011
rect 27801 14971 27859 14977
rect 27890 14968 27896 15020
rect 27948 14968 27954 15020
rect 28460 15017 28488 15048
rect 28552 15048 28948 15076
rect 28552 15017 28580 15048
rect 28077 15011 28135 15017
rect 28077 14977 28089 15011
rect 28123 15008 28135 15011
rect 28261 15011 28319 15017
rect 28261 15008 28273 15011
rect 28123 14980 28273 15008
rect 28123 14977 28135 14980
rect 28077 14971 28135 14977
rect 28261 14977 28273 14980
rect 28307 14977 28319 15011
rect 28261 14971 28319 14977
rect 28445 15011 28503 15017
rect 28445 14977 28457 15011
rect 28491 14977 28503 15011
rect 28445 14971 28503 14977
rect 28537 15011 28595 15017
rect 28537 14977 28549 15011
rect 28583 14977 28595 15011
rect 28537 14971 28595 14977
rect 26142 14940 26148 14952
rect 25792 14912 26148 14940
rect 26142 14900 26148 14912
rect 26200 14940 26206 14952
rect 28276 14940 28304 14971
rect 28810 14968 28816 15020
rect 28868 14968 28874 15020
rect 28920 15008 28948 15048
rect 28997 15045 29009 15079
rect 29043 15076 29055 15079
rect 29043 15048 34008 15076
rect 29043 15045 29055 15048
rect 28997 15039 29055 15045
rect 28920 14980 29500 15008
rect 29472 14952 29500 14980
rect 30466 14968 30472 15020
rect 30524 15008 30530 15020
rect 30653 15011 30711 15017
rect 30653 15008 30665 15011
rect 30524 14980 30665 15008
rect 30524 14968 30530 14980
rect 30653 14977 30665 14980
rect 30699 14977 30711 15011
rect 30653 14971 30711 14977
rect 30742 14968 30748 15020
rect 30800 14968 30806 15020
rect 30834 14968 30840 15020
rect 30892 14968 30898 15020
rect 30929 15011 30987 15017
rect 30929 14977 30941 15011
rect 30975 14977 30987 15011
rect 30929 14971 30987 14977
rect 28629 14943 28687 14949
rect 26200 14912 28120 14940
rect 28276 14912 28580 14940
rect 26200 14900 26206 14912
rect 15933 14835 15991 14841
rect 16040 14844 20392 14872
rect 8297 14807 8355 14813
rect 8297 14804 8309 14807
rect 7484 14776 8309 14804
rect 3936 14764 3942 14776
rect 8297 14773 8309 14776
rect 8343 14773 8355 14807
rect 8297 14767 8355 14773
rect 8662 14764 8668 14816
rect 8720 14764 8726 14816
rect 8849 14807 8907 14813
rect 8849 14773 8861 14807
rect 8895 14804 8907 14807
rect 8938 14804 8944 14816
rect 8895 14776 8944 14804
rect 8895 14773 8907 14776
rect 8849 14767 8907 14773
rect 8938 14764 8944 14776
rect 8996 14764 9002 14816
rect 9766 14764 9772 14816
rect 9824 14764 9830 14816
rect 10226 14764 10232 14816
rect 10284 14804 10290 14816
rect 10321 14807 10379 14813
rect 10321 14804 10333 14807
rect 10284 14776 10333 14804
rect 10284 14764 10290 14776
rect 10321 14773 10333 14776
rect 10367 14773 10379 14807
rect 10321 14767 10379 14773
rect 13538 14764 13544 14816
rect 13596 14804 13602 14816
rect 16040 14804 16068 14844
rect 21266 14832 21272 14884
rect 21324 14872 21330 14884
rect 23658 14872 23664 14884
rect 21324 14844 23664 14872
rect 21324 14832 21330 14844
rect 23658 14832 23664 14844
rect 23716 14832 23722 14884
rect 24762 14832 24768 14884
rect 24820 14872 24826 14884
rect 27433 14875 27491 14881
rect 24820 14844 26464 14872
rect 24820 14832 24826 14844
rect 13596 14776 16068 14804
rect 13596 14764 13602 14776
rect 16390 14764 16396 14816
rect 16448 14764 16454 14816
rect 16574 14764 16580 14816
rect 16632 14804 16638 14816
rect 17678 14804 17684 14816
rect 16632 14776 17684 14804
rect 16632 14764 16638 14776
rect 17678 14764 17684 14776
rect 17736 14764 17742 14816
rect 18782 14764 18788 14816
rect 18840 14804 18846 14816
rect 19242 14804 19248 14816
rect 18840 14776 19248 14804
rect 18840 14764 18846 14776
rect 19242 14764 19248 14776
rect 19300 14764 19306 14816
rect 20530 14764 20536 14816
rect 20588 14764 20594 14816
rect 20806 14764 20812 14816
rect 20864 14804 20870 14816
rect 22186 14804 22192 14816
rect 20864 14776 22192 14804
rect 20864 14764 20870 14776
rect 22186 14764 22192 14776
rect 22244 14764 22250 14816
rect 25590 14764 25596 14816
rect 25648 14764 25654 14816
rect 25961 14807 26019 14813
rect 25961 14773 25973 14807
rect 26007 14804 26019 14807
rect 26326 14804 26332 14816
rect 26007 14776 26332 14804
rect 26007 14773 26019 14776
rect 25961 14767 26019 14773
rect 26326 14764 26332 14776
rect 26384 14764 26390 14816
rect 26436 14804 26464 14844
rect 27433 14841 27445 14875
rect 27479 14872 27491 14875
rect 27985 14875 28043 14881
rect 27985 14872 27997 14875
rect 27479 14844 27997 14872
rect 27479 14841 27491 14844
rect 27433 14835 27491 14841
rect 27985 14841 27997 14844
rect 28031 14841 28043 14875
rect 27985 14835 28043 14841
rect 27617 14807 27675 14813
rect 27617 14804 27629 14807
rect 26436 14776 27629 14804
rect 27617 14773 27629 14776
rect 27663 14773 27675 14807
rect 28092 14804 28120 14912
rect 28552 14884 28580 14912
rect 28629 14909 28641 14943
rect 28675 14940 28687 14943
rect 28718 14940 28724 14952
rect 28675 14912 28724 14940
rect 28675 14909 28687 14912
rect 28629 14903 28687 14909
rect 28718 14900 28724 14912
rect 28776 14940 28782 14952
rect 28776 14912 28994 14940
rect 28776 14900 28782 14912
rect 28534 14832 28540 14884
rect 28592 14832 28598 14884
rect 28810 14832 28816 14884
rect 28868 14832 28874 14884
rect 28966 14872 28994 14912
rect 29454 14900 29460 14952
rect 29512 14900 29518 14952
rect 30374 14900 30380 14952
rect 30432 14940 30438 14952
rect 30944 14940 30972 14971
rect 31110 14968 31116 15020
rect 31168 14968 31174 15020
rect 33042 14968 33048 15020
rect 33100 14968 33106 15020
rect 33980 15017 34008 15048
rect 33965 15011 34023 15017
rect 33965 14977 33977 15011
rect 34011 14977 34023 15011
rect 33965 14971 34023 14977
rect 30432 14912 30972 14940
rect 30432 14900 30438 14912
rect 31662 14900 31668 14952
rect 31720 14900 31726 14952
rect 32950 14900 32956 14952
rect 33008 14900 33014 14952
rect 33873 14943 33931 14949
rect 33873 14940 33885 14943
rect 33428 14912 33885 14940
rect 31680 14872 31708 14900
rect 33428 14881 33456 14912
rect 33873 14909 33885 14912
rect 33919 14909 33931 14943
rect 33873 14903 33931 14909
rect 28966 14844 31708 14872
rect 33413 14875 33471 14881
rect 33413 14841 33425 14875
rect 33459 14841 33471 14875
rect 33413 14835 33471 14841
rect 28828 14804 28856 14832
rect 28092 14776 28856 14804
rect 31021 14807 31079 14813
rect 27617 14767 27675 14773
rect 31021 14773 31033 14807
rect 31067 14804 31079 14807
rect 31202 14804 31208 14816
rect 31067 14776 31208 14804
rect 31067 14773 31079 14776
rect 31021 14767 31079 14773
rect 31202 14764 31208 14776
rect 31260 14764 31266 14816
rect 1104 14714 38272 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 38272 14714
rect 1104 14640 38272 14662
rect 3145 14603 3203 14609
rect 3145 14569 3157 14603
rect 3191 14600 3203 14603
rect 3234 14600 3240 14612
rect 3191 14572 3240 14600
rect 3191 14569 3203 14572
rect 3145 14563 3203 14569
rect 3234 14560 3240 14572
rect 3292 14560 3298 14612
rect 3602 14560 3608 14612
rect 3660 14560 3666 14612
rect 4062 14560 4068 14612
rect 4120 14560 4126 14612
rect 7374 14560 7380 14612
rect 7432 14560 7438 14612
rect 8662 14560 8668 14612
rect 8720 14600 8726 14612
rect 8846 14600 8852 14612
rect 8720 14572 8852 14600
rect 8720 14560 8726 14572
rect 8846 14560 8852 14572
rect 8904 14560 8910 14612
rect 13449 14603 13507 14609
rect 13449 14569 13461 14603
rect 13495 14600 13507 14603
rect 14090 14600 14096 14612
rect 13495 14572 14096 14600
rect 13495 14569 13507 14572
rect 13449 14563 13507 14569
rect 14090 14560 14096 14572
rect 14148 14560 14154 14612
rect 14826 14560 14832 14612
rect 14884 14560 14890 14612
rect 15562 14560 15568 14612
rect 15620 14560 15626 14612
rect 15930 14560 15936 14612
rect 15988 14600 15994 14612
rect 16574 14600 16580 14612
rect 15988 14572 16580 14600
rect 15988 14560 15994 14572
rect 16574 14560 16580 14572
rect 16632 14560 16638 14612
rect 17034 14560 17040 14612
rect 17092 14560 17098 14612
rect 17402 14560 17408 14612
rect 17460 14600 17466 14612
rect 19613 14603 19671 14609
rect 19613 14600 19625 14603
rect 17460 14572 19625 14600
rect 17460 14560 17466 14572
rect 19613 14569 19625 14572
rect 19659 14569 19671 14603
rect 19613 14563 19671 14569
rect 22922 14560 22928 14612
rect 22980 14600 22986 14612
rect 22980 14572 27614 14600
rect 22980 14560 22986 14572
rect 1394 14356 1400 14408
rect 1452 14356 1458 14408
rect 2774 14356 2780 14408
rect 2832 14356 2838 14408
rect 3620 14396 3648 14560
rect 9122 14492 9128 14544
rect 9180 14532 9186 14544
rect 9180 14504 9352 14532
rect 9180 14492 9186 14504
rect 3694 14424 3700 14476
rect 3752 14464 3758 14476
rect 3752 14436 8984 14464
rect 3752 14424 3758 14436
rect 4065 14399 4123 14405
rect 4065 14396 4077 14399
rect 3620 14368 4077 14396
rect 4065 14365 4077 14368
rect 4111 14365 4123 14399
rect 4065 14359 4123 14365
rect 4249 14399 4307 14405
rect 4249 14365 4261 14399
rect 4295 14396 4307 14399
rect 4614 14396 4620 14408
rect 4295 14368 4620 14396
rect 4295 14365 4307 14368
rect 4249 14359 4307 14365
rect 4614 14356 4620 14368
rect 4672 14356 4678 14408
rect 5626 14356 5632 14408
rect 5684 14356 5690 14408
rect 8956 14405 8984 14436
rect 8941 14399 8999 14405
rect 8941 14365 8953 14399
rect 8987 14365 8999 14399
rect 8941 14359 8999 14365
rect 9030 14356 9036 14408
rect 9088 14396 9094 14408
rect 9324 14405 9352 14504
rect 10137 14467 10195 14473
rect 10137 14433 10149 14467
rect 10183 14464 10195 14467
rect 10226 14464 10232 14476
rect 10183 14436 10232 14464
rect 10183 14433 10195 14436
rect 10137 14427 10195 14433
rect 10226 14424 10232 14436
rect 10284 14424 10290 14476
rect 11885 14467 11943 14473
rect 11885 14433 11897 14467
rect 11931 14464 11943 14467
rect 12066 14464 12072 14476
rect 11931 14436 12072 14464
rect 11931 14433 11943 14436
rect 11885 14427 11943 14433
rect 12066 14424 12072 14436
rect 12124 14424 12130 14476
rect 12526 14424 12532 14476
rect 12584 14464 12590 14476
rect 12805 14467 12863 14473
rect 12805 14464 12817 14467
rect 12584 14436 12817 14464
rect 12584 14424 12590 14436
rect 12805 14433 12817 14436
rect 12851 14433 12863 14467
rect 12805 14427 12863 14433
rect 12989 14467 13047 14473
rect 12989 14433 13001 14467
rect 13035 14464 13047 14467
rect 14366 14464 14372 14476
rect 13035 14436 14372 14464
rect 13035 14433 13047 14436
rect 12989 14427 13047 14433
rect 14366 14424 14372 14436
rect 14424 14424 14430 14476
rect 14844 14464 14872 14560
rect 15580 14532 15608 14560
rect 15580 14504 18000 14532
rect 15473 14467 15531 14473
rect 15473 14464 15485 14467
rect 14844 14436 15485 14464
rect 15473 14433 15485 14436
rect 15519 14433 15531 14467
rect 15473 14427 15531 14433
rect 9125 14399 9183 14405
rect 9125 14396 9137 14399
rect 9088 14368 9137 14396
rect 9088 14356 9094 14368
rect 9125 14365 9137 14368
rect 9171 14365 9183 14399
rect 9125 14359 9183 14365
rect 9217 14399 9275 14405
rect 9217 14365 9229 14399
rect 9263 14365 9275 14399
rect 9217 14359 9275 14365
rect 9309 14399 9367 14405
rect 9309 14365 9321 14399
rect 9355 14365 9367 14399
rect 9309 14359 9367 14365
rect 1670 14288 1676 14340
rect 1728 14288 1734 14340
rect 5902 14288 5908 14340
rect 5960 14288 5966 14340
rect 6914 14288 6920 14340
rect 6972 14288 6978 14340
rect 8754 14288 8760 14340
rect 8812 14328 8818 14340
rect 9232 14328 9260 14359
rect 9858 14356 9864 14408
rect 9916 14356 9922 14408
rect 11146 14356 11152 14408
rect 11204 14396 11210 14408
rect 11698 14396 11704 14408
rect 11204 14368 11704 14396
rect 11204 14356 11210 14368
rect 11698 14356 11704 14368
rect 11756 14356 11762 14408
rect 14458 14356 14464 14408
rect 14516 14396 14522 14408
rect 14826 14396 14832 14408
rect 14516 14368 14832 14396
rect 14516 14356 14522 14368
rect 14826 14356 14832 14368
rect 14884 14356 14890 14408
rect 15286 14356 15292 14408
rect 15344 14356 15350 14408
rect 15488 14396 15516 14427
rect 16390 14424 16396 14476
rect 16448 14464 16454 14476
rect 16448 14436 17632 14464
rect 16448 14424 16454 14436
rect 16482 14396 16488 14408
rect 15488 14368 16488 14396
rect 16482 14356 16488 14368
rect 16540 14356 16546 14408
rect 16577 14399 16635 14405
rect 16577 14365 16589 14399
rect 16623 14396 16635 14399
rect 16666 14396 16672 14408
rect 16623 14368 16672 14396
rect 16623 14365 16635 14368
rect 16577 14359 16635 14365
rect 16666 14356 16672 14368
rect 16724 14356 16730 14408
rect 17052 14405 17080 14436
rect 16761 14399 16819 14405
rect 16761 14365 16773 14399
rect 16807 14365 16819 14399
rect 16761 14359 16819 14365
rect 17037 14399 17095 14405
rect 17037 14365 17049 14399
rect 17083 14365 17095 14399
rect 17037 14359 17095 14365
rect 17221 14399 17279 14405
rect 17221 14365 17233 14399
rect 17267 14365 17279 14399
rect 17221 14359 17279 14365
rect 8812 14300 9260 14328
rect 8812 14288 8818 14300
rect 9582 14288 9588 14340
rect 9640 14288 9646 14340
rect 12406 14300 13124 14328
rect 8662 14220 8668 14272
rect 8720 14260 8726 14272
rect 12406 14260 12434 14300
rect 13096 14269 13124 14300
rect 15562 14288 15568 14340
rect 15620 14328 15626 14340
rect 16776 14328 16804 14359
rect 16942 14328 16948 14340
rect 15620 14300 16948 14328
rect 15620 14288 15626 14300
rect 16942 14288 16948 14300
rect 17000 14288 17006 14340
rect 8720 14232 12434 14260
rect 13081 14263 13139 14269
rect 8720 14220 8726 14232
rect 13081 14229 13093 14263
rect 13127 14260 13139 14263
rect 13998 14260 14004 14272
rect 13127 14232 14004 14260
rect 13127 14229 13139 14232
rect 13081 14223 13139 14229
rect 13998 14220 14004 14232
rect 14056 14220 14062 14272
rect 16114 14220 16120 14272
rect 16172 14260 16178 14272
rect 17236 14260 17264 14359
rect 17310 14356 17316 14408
rect 17368 14356 17374 14408
rect 17604 14328 17632 14436
rect 17972 14405 18000 14504
rect 20530 14492 20536 14544
rect 20588 14492 20594 14544
rect 20622 14492 20628 14544
rect 20680 14532 20686 14544
rect 23109 14535 23167 14541
rect 20680 14504 21312 14532
rect 20680 14492 20686 14504
rect 18046 14424 18052 14476
rect 18104 14464 18110 14476
rect 20548 14464 20576 14492
rect 20993 14467 21051 14473
rect 20993 14464 21005 14467
rect 18104 14436 18184 14464
rect 20548 14436 21005 14464
rect 18104 14424 18110 14436
rect 18156 14405 18184 14436
rect 20993 14433 21005 14436
rect 21039 14433 21051 14467
rect 20993 14427 21051 14433
rect 17957 14399 18015 14405
rect 17957 14365 17969 14399
rect 18003 14365 18015 14399
rect 17957 14359 18015 14365
rect 18141 14399 18199 14405
rect 18141 14365 18153 14399
rect 18187 14365 18199 14399
rect 19245 14399 19303 14405
rect 19245 14396 19257 14399
rect 18141 14359 18199 14365
rect 18248 14368 19257 14396
rect 18049 14331 18107 14337
rect 18049 14328 18061 14331
rect 17604 14300 18061 14328
rect 18049 14297 18061 14300
rect 18095 14328 18107 14331
rect 18248 14328 18276 14368
rect 19245 14365 19257 14368
rect 19291 14365 19303 14399
rect 19245 14359 19303 14365
rect 19889 14399 19947 14405
rect 19889 14365 19901 14399
rect 19935 14365 19947 14399
rect 19889 14359 19947 14365
rect 20533 14399 20591 14405
rect 20533 14365 20545 14399
rect 20579 14365 20591 14399
rect 20533 14359 20591 14365
rect 20809 14399 20867 14405
rect 20809 14365 20821 14399
rect 20855 14396 20867 14399
rect 20898 14396 20904 14408
rect 20855 14368 20904 14396
rect 20855 14365 20867 14368
rect 20809 14359 20867 14365
rect 19518 14328 19524 14340
rect 18095 14300 18276 14328
rect 19306 14300 19524 14328
rect 18095 14297 18107 14300
rect 18049 14291 18107 14297
rect 19306 14260 19334 14300
rect 19518 14288 19524 14300
rect 19576 14288 19582 14340
rect 19904 14328 19932 14359
rect 20438 14328 20444 14340
rect 19904 14300 20444 14328
rect 20438 14288 20444 14300
rect 20496 14328 20502 14340
rect 20548 14328 20576 14359
rect 20898 14356 20904 14368
rect 20956 14356 20962 14408
rect 21082 14356 21088 14408
rect 21140 14356 21146 14408
rect 21284 14405 21312 14504
rect 23109 14501 23121 14535
rect 23155 14532 23167 14535
rect 23934 14532 23940 14544
rect 23155 14504 23940 14532
rect 23155 14501 23167 14504
rect 23109 14495 23167 14501
rect 23934 14492 23940 14504
rect 23992 14492 23998 14544
rect 27586 14532 27614 14572
rect 28350 14560 28356 14612
rect 28408 14600 28414 14612
rect 31754 14600 31760 14612
rect 28408 14572 31760 14600
rect 28408 14560 28414 14572
rect 31754 14560 31760 14572
rect 31812 14560 31818 14612
rect 31941 14603 31999 14609
rect 31941 14569 31953 14603
rect 31987 14600 31999 14603
rect 32950 14600 32956 14612
rect 31987 14572 32956 14600
rect 31987 14569 31999 14572
rect 31941 14563 31999 14569
rect 32950 14560 32956 14572
rect 33008 14560 33014 14612
rect 29178 14532 29184 14544
rect 27586 14504 29184 14532
rect 29178 14492 29184 14504
rect 29236 14492 29242 14544
rect 31294 14492 31300 14544
rect 31352 14532 31358 14544
rect 31352 14504 31524 14532
rect 31352 14492 31358 14504
rect 21637 14467 21695 14473
rect 21637 14433 21649 14467
rect 21683 14464 21695 14467
rect 21910 14464 21916 14476
rect 21683 14436 21916 14464
rect 21683 14433 21695 14436
rect 21637 14427 21695 14433
rect 21910 14424 21916 14436
rect 21968 14464 21974 14476
rect 21968 14436 22692 14464
rect 21968 14424 21974 14436
rect 22664 14405 22692 14436
rect 23290 14424 23296 14476
rect 23348 14424 23354 14476
rect 23385 14467 23443 14473
rect 23385 14433 23397 14467
rect 23431 14464 23443 14467
rect 23431 14436 23704 14464
rect 23431 14433 23443 14436
rect 23385 14427 23443 14433
rect 21269 14399 21327 14405
rect 21269 14365 21281 14399
rect 21315 14365 21327 14399
rect 21269 14359 21327 14365
rect 22005 14399 22063 14405
rect 22005 14365 22017 14399
rect 22051 14365 22063 14399
rect 22005 14359 22063 14365
rect 22649 14399 22707 14405
rect 22649 14365 22661 14399
rect 22695 14365 22707 14399
rect 22649 14359 22707 14365
rect 23569 14399 23627 14405
rect 23569 14365 23581 14399
rect 23615 14365 23627 14399
rect 23676 14396 23704 14436
rect 30834 14424 30840 14476
rect 30892 14424 30898 14476
rect 24118 14396 24124 14408
rect 23676 14368 24124 14396
rect 23569 14359 23627 14365
rect 20496 14300 20576 14328
rect 21100 14328 21128 14356
rect 21818 14328 21824 14340
rect 21100 14300 21824 14328
rect 20496 14288 20502 14300
rect 21818 14288 21824 14300
rect 21876 14328 21882 14340
rect 22020 14328 22048 14359
rect 21876 14300 22048 14328
rect 21876 14288 21882 14300
rect 23198 14288 23204 14340
rect 23256 14328 23262 14340
rect 23584 14328 23612 14359
rect 24118 14356 24124 14368
rect 24176 14356 24182 14408
rect 24486 14356 24492 14408
rect 24544 14356 24550 14408
rect 30285 14399 30343 14405
rect 30285 14365 30297 14399
rect 30331 14365 30343 14399
rect 30285 14359 30343 14365
rect 30377 14399 30435 14405
rect 30377 14365 30389 14399
rect 30423 14396 30435 14399
rect 30852 14396 30880 14424
rect 30423 14368 30972 14396
rect 30423 14365 30435 14368
rect 30377 14359 30435 14365
rect 24504 14328 24532 14356
rect 23256 14300 24532 14328
rect 23256 14288 23262 14300
rect 26234 14288 26240 14340
rect 26292 14328 26298 14340
rect 27154 14328 27160 14340
rect 26292 14300 27160 14328
rect 26292 14288 26298 14300
rect 27154 14288 27160 14300
rect 27212 14288 27218 14340
rect 30300 14328 30328 14359
rect 30466 14328 30472 14340
rect 30300 14300 30472 14328
rect 30300 14272 30328 14300
rect 30466 14288 30472 14300
rect 30524 14288 30530 14340
rect 30561 14331 30619 14337
rect 30561 14297 30573 14331
rect 30607 14328 30619 14331
rect 30653 14331 30711 14337
rect 30653 14328 30665 14331
rect 30607 14300 30665 14328
rect 30607 14297 30619 14300
rect 30561 14291 30619 14297
rect 30653 14297 30665 14300
rect 30699 14297 30711 14331
rect 30653 14291 30711 14297
rect 30742 14288 30748 14340
rect 30800 14328 30806 14340
rect 30837 14331 30895 14337
rect 30837 14328 30849 14331
rect 30800 14300 30849 14328
rect 30800 14288 30806 14300
rect 30837 14297 30849 14300
rect 30883 14297 30895 14331
rect 30944 14328 30972 14368
rect 31202 14356 31208 14408
rect 31260 14356 31266 14408
rect 31386 14356 31392 14408
rect 31444 14356 31450 14408
rect 31496 14405 31524 14504
rect 31573 14467 31631 14473
rect 31573 14433 31585 14467
rect 31619 14464 31631 14467
rect 31662 14464 31668 14476
rect 31619 14436 31668 14464
rect 31619 14433 31631 14436
rect 31573 14427 31631 14433
rect 31662 14424 31668 14436
rect 31720 14464 31726 14476
rect 33778 14464 33784 14476
rect 31720 14436 33784 14464
rect 31720 14424 31726 14436
rect 33778 14424 33784 14436
rect 33836 14464 33842 14476
rect 33836 14436 34100 14464
rect 33836 14424 33842 14436
rect 34072 14408 34100 14436
rect 31481 14399 31539 14405
rect 31481 14365 31493 14399
rect 31527 14365 31539 14399
rect 31481 14359 31539 14365
rect 31754 14356 31760 14408
rect 31812 14356 31818 14408
rect 34054 14356 34060 14408
rect 34112 14356 34118 14408
rect 30944 14300 31156 14328
rect 30837 14291 30895 14297
rect 16172 14232 19334 14260
rect 16172 14220 16178 14232
rect 19426 14220 19432 14272
rect 19484 14260 19490 14272
rect 19622 14263 19680 14269
rect 19622 14260 19634 14263
rect 19484 14232 19634 14260
rect 19484 14220 19490 14232
rect 19622 14229 19634 14232
rect 19668 14229 19680 14263
rect 19622 14223 19680 14229
rect 23753 14263 23811 14269
rect 23753 14229 23765 14263
rect 23799 14260 23811 14263
rect 23842 14260 23848 14272
rect 23799 14232 23848 14260
rect 23799 14229 23811 14232
rect 23753 14223 23811 14229
rect 23842 14220 23848 14232
rect 23900 14260 23906 14272
rect 26418 14260 26424 14272
rect 23900 14232 26424 14260
rect 23900 14220 23906 14232
rect 26418 14220 26424 14232
rect 26476 14220 26482 14272
rect 30282 14220 30288 14272
rect 30340 14220 30346 14272
rect 30374 14220 30380 14272
rect 30432 14260 30438 14272
rect 31021 14263 31079 14269
rect 31021 14260 31033 14263
rect 30432 14232 31033 14260
rect 30432 14220 30438 14232
rect 31021 14229 31033 14232
rect 31067 14229 31079 14263
rect 31128 14260 31156 14300
rect 32122 14260 32128 14272
rect 31128 14232 32128 14260
rect 31021 14223 31079 14229
rect 32122 14220 32128 14232
rect 32180 14220 32186 14272
rect 1104 14170 38272 14192
rect 1104 14118 4874 14170
rect 4926 14118 4938 14170
rect 4990 14118 5002 14170
rect 5054 14118 5066 14170
rect 5118 14118 5130 14170
rect 5182 14118 35594 14170
rect 35646 14118 35658 14170
rect 35710 14118 35722 14170
rect 35774 14118 35786 14170
rect 35838 14118 35850 14170
rect 35902 14118 38272 14170
rect 1104 14096 38272 14118
rect 1670 14016 1676 14068
rect 1728 14056 1734 14068
rect 1949 14059 2007 14065
rect 1949 14056 1961 14059
rect 1728 14028 1961 14056
rect 1728 14016 1734 14028
rect 1949 14025 1961 14028
rect 1995 14025 2007 14059
rect 1949 14019 2007 14025
rect 2498 14016 2504 14068
rect 2556 14016 2562 14068
rect 5902 14016 5908 14068
rect 5960 14056 5966 14068
rect 6365 14059 6423 14065
rect 6365 14056 6377 14059
rect 5960 14028 6377 14056
rect 5960 14016 5966 14028
rect 6365 14025 6377 14028
rect 6411 14025 6423 14059
rect 6365 14019 6423 14025
rect 6641 14059 6699 14065
rect 6641 14025 6653 14059
rect 6687 14025 6699 14059
rect 6641 14019 6699 14025
rect 7009 14059 7067 14065
rect 7009 14025 7021 14059
rect 7055 14056 7067 14059
rect 8662 14056 8668 14068
rect 7055 14028 8668 14056
rect 7055 14025 7067 14028
rect 7009 14019 7067 14025
rect 1765 13923 1823 13929
rect 1765 13889 1777 13923
rect 1811 13889 1823 13923
rect 1765 13883 1823 13889
rect 2133 13923 2191 13929
rect 2133 13889 2145 13923
rect 2179 13920 2191 13923
rect 2516 13920 2544 14016
rect 2179 13892 2544 13920
rect 6549 13923 6607 13929
rect 2179 13889 2191 13892
rect 2133 13883 2191 13889
rect 6549 13889 6561 13923
rect 6595 13920 6607 13923
rect 6656 13920 6684 14019
rect 8662 14016 8668 14028
rect 8720 14016 8726 14068
rect 16758 14016 16764 14068
rect 16816 14056 16822 14068
rect 17773 14059 17831 14065
rect 17773 14056 17785 14059
rect 16816 14028 17785 14056
rect 16816 14016 16822 14028
rect 17773 14025 17785 14028
rect 17819 14025 17831 14059
rect 17773 14019 17831 14025
rect 17862 14016 17868 14068
rect 17920 14016 17926 14068
rect 19797 14059 19855 14065
rect 19797 14025 19809 14059
rect 19843 14056 19855 14059
rect 21082 14056 21088 14068
rect 19843 14028 21088 14056
rect 19843 14025 19855 14028
rect 19797 14019 19855 14025
rect 21082 14016 21088 14028
rect 21140 14016 21146 14068
rect 23477 14059 23535 14065
rect 23477 14025 23489 14059
rect 23523 14056 23535 14059
rect 23523 14028 25912 14056
rect 23523 14025 23535 14028
rect 23477 14019 23535 14025
rect 7101 13991 7159 13997
rect 7101 13957 7113 13991
rect 7147 13988 7159 13991
rect 7374 13988 7380 14000
rect 7147 13960 7380 13988
rect 7147 13957 7159 13960
rect 7101 13951 7159 13957
rect 7374 13948 7380 13960
rect 7432 13948 7438 14000
rect 8570 13988 8576 14000
rect 8496 13960 8576 13988
rect 6595 13892 6684 13920
rect 6595 13889 6607 13892
rect 6549 13883 6607 13889
rect 1486 13812 1492 13864
rect 1544 13812 1550 13864
rect 1780 13852 1808 13883
rect 8386 13880 8392 13932
rect 8444 13880 8450 13932
rect 8496 13929 8524 13960
rect 8570 13948 8576 13960
rect 8628 13988 8634 14000
rect 10134 13988 10140 14000
rect 8628 13960 10140 13988
rect 8628 13948 8634 13960
rect 10134 13948 10140 13960
rect 10192 13948 10198 14000
rect 12986 13948 12992 14000
rect 13044 13988 13050 14000
rect 13262 13988 13268 14000
rect 13044 13960 13268 13988
rect 13044 13948 13050 13960
rect 13262 13948 13268 13960
rect 13320 13988 13326 14000
rect 15102 13988 15108 14000
rect 13320 13960 15108 13988
rect 13320 13948 13326 13960
rect 8481 13923 8539 13929
rect 8481 13889 8493 13923
rect 8527 13889 8539 13923
rect 8481 13883 8539 13889
rect 9950 13880 9956 13932
rect 10008 13920 10014 13932
rect 12434 13920 12440 13932
rect 10008 13892 12440 13920
rect 10008 13880 10014 13892
rect 12434 13880 12440 13892
rect 12492 13880 12498 13932
rect 13354 13880 13360 13932
rect 13412 13880 13418 13932
rect 14660 13929 14688 13960
rect 15102 13948 15108 13960
rect 15160 13988 15166 14000
rect 17221 13991 17279 13997
rect 15160 13960 16804 13988
rect 15160 13948 15166 13960
rect 14645 13923 14703 13929
rect 14645 13889 14657 13923
rect 14691 13889 14703 13923
rect 14645 13883 14703 13889
rect 15194 13880 15200 13932
rect 15252 13920 15258 13932
rect 16776 13929 16804 13960
rect 17221 13957 17233 13991
rect 17267 13988 17279 13991
rect 17494 13988 17500 14000
rect 17267 13960 17500 13988
rect 17267 13957 17279 13960
rect 17221 13951 17279 13957
rect 17494 13948 17500 13960
rect 17552 13948 17558 14000
rect 20530 13948 20536 14000
rect 20588 13988 20594 14000
rect 20588 13960 21128 13988
rect 20588 13948 20594 13960
rect 15289 13923 15347 13929
rect 15289 13920 15301 13923
rect 15252 13892 15301 13920
rect 15252 13880 15258 13892
rect 15289 13889 15301 13892
rect 15335 13920 15347 13923
rect 16209 13923 16267 13929
rect 16209 13920 16221 13923
rect 15335 13892 16221 13920
rect 15335 13889 15347 13892
rect 15289 13883 15347 13889
rect 16209 13889 16221 13892
rect 16255 13920 16267 13923
rect 16669 13923 16727 13929
rect 16669 13920 16681 13923
rect 16255 13892 16681 13920
rect 16255 13889 16267 13892
rect 16209 13883 16267 13889
rect 16669 13889 16681 13892
rect 16715 13889 16727 13923
rect 16669 13883 16727 13889
rect 16761 13923 16819 13929
rect 16761 13889 16773 13923
rect 16807 13920 16819 13923
rect 17310 13920 17316 13932
rect 16807 13892 17316 13920
rect 16807 13889 16819 13892
rect 16761 13883 16819 13889
rect 17310 13880 17316 13892
rect 17368 13880 17374 13932
rect 19702 13880 19708 13932
rect 19760 13880 19766 13932
rect 20257 13923 20315 13929
rect 20257 13920 20269 13923
rect 19812 13892 20269 13920
rect 5994 13852 6000 13864
rect 1780 13824 6000 13852
rect 5994 13812 6000 13824
rect 6052 13812 6058 13864
rect 7193 13855 7251 13861
rect 7193 13821 7205 13855
rect 7239 13852 7251 13855
rect 7650 13852 7656 13864
rect 7239 13824 7656 13852
rect 7239 13821 7251 13824
rect 7193 13815 7251 13821
rect 7208 13784 7236 13815
rect 7650 13812 7656 13824
rect 7708 13812 7714 13864
rect 13372 13852 13400 13880
rect 15562 13852 15568 13864
rect 13372 13824 15568 13852
rect 15562 13812 15568 13824
rect 15620 13812 15626 13864
rect 17957 13855 18015 13861
rect 17957 13821 17969 13855
rect 18003 13821 18015 13855
rect 17957 13815 18015 13821
rect 7116 13756 7236 13784
rect 7116 13728 7144 13756
rect 10962 13744 10968 13796
rect 11020 13784 11026 13796
rect 17972 13784 18000 13815
rect 11020 13756 18000 13784
rect 11020 13744 11026 13756
rect 18414 13744 18420 13796
rect 18472 13784 18478 13796
rect 18966 13784 18972 13796
rect 18472 13756 18972 13784
rect 18472 13744 18478 13756
rect 18966 13744 18972 13756
rect 19024 13744 19030 13796
rect 7098 13676 7104 13728
rect 7156 13676 7162 13728
rect 15013 13719 15071 13725
rect 15013 13685 15025 13719
rect 15059 13716 15071 13719
rect 15654 13716 15660 13728
rect 15059 13688 15660 13716
rect 15059 13685 15071 13688
rect 15013 13679 15071 13685
rect 15654 13676 15660 13688
rect 15712 13676 15718 13728
rect 17402 13676 17408 13728
rect 17460 13676 17466 13728
rect 17862 13676 17868 13728
rect 17920 13716 17926 13728
rect 19610 13716 19616 13728
rect 17920 13688 19616 13716
rect 17920 13676 17926 13688
rect 19610 13676 19616 13688
rect 19668 13716 19674 13728
rect 19812 13716 19840 13892
rect 20257 13889 20269 13892
rect 20303 13889 20315 13923
rect 20257 13883 20315 13889
rect 20438 13880 20444 13932
rect 20496 13920 20502 13932
rect 20625 13923 20683 13929
rect 20625 13920 20637 13923
rect 20496 13892 20637 13920
rect 20496 13880 20502 13892
rect 20625 13889 20637 13892
rect 20671 13889 20683 13923
rect 20625 13883 20683 13889
rect 20640 13852 20668 13883
rect 20714 13880 20720 13932
rect 20772 13920 20778 13932
rect 21100 13929 21128 13960
rect 22554 13948 22560 14000
rect 22612 13988 22618 14000
rect 22833 13991 22891 13997
rect 22833 13988 22845 13991
rect 22612 13960 22845 13988
rect 22612 13948 22618 13960
rect 22833 13957 22845 13960
rect 22879 13988 22891 13991
rect 25409 13991 25467 13997
rect 25409 13988 25421 13991
rect 22879 13960 24624 13988
rect 22879 13957 22891 13960
rect 22833 13951 22891 13957
rect 20901 13923 20959 13929
rect 20901 13920 20913 13923
rect 20772 13892 20913 13920
rect 20772 13880 20778 13892
rect 20901 13889 20913 13892
rect 20947 13889 20959 13923
rect 20901 13883 20959 13889
rect 21085 13923 21143 13929
rect 21085 13889 21097 13923
rect 21131 13889 21143 13923
rect 21085 13883 21143 13889
rect 21177 13923 21235 13929
rect 21177 13889 21189 13923
rect 21223 13889 21235 13923
rect 21177 13883 21235 13889
rect 21270 13913 21328 13919
rect 21192 13852 21220 13883
rect 21270 13879 21282 13913
rect 21316 13879 21328 13913
rect 22094 13880 22100 13932
rect 22152 13880 22158 13932
rect 22281 13923 22339 13929
rect 22281 13889 22293 13923
rect 22327 13920 22339 13923
rect 22649 13923 22707 13929
rect 22649 13920 22661 13923
rect 22327 13892 22661 13920
rect 22327 13889 22339 13892
rect 22281 13883 22339 13889
rect 22649 13889 22661 13892
rect 22695 13920 22707 13923
rect 24118 13920 24124 13932
rect 22695 13892 24124 13920
rect 22695 13889 22707 13892
rect 22649 13883 22707 13889
rect 24118 13880 24124 13892
rect 24176 13880 24182 13932
rect 24486 13880 24492 13932
rect 24544 13880 24550 13932
rect 21270 13873 21328 13879
rect 20640 13824 21220 13852
rect 20898 13744 20904 13796
rect 20956 13784 20962 13796
rect 21285 13784 21313 13873
rect 21913 13855 21971 13861
rect 21913 13852 21925 13855
rect 21560 13824 21925 13852
rect 20956 13756 21313 13784
rect 20956 13744 20962 13756
rect 21358 13744 21364 13796
rect 21416 13784 21422 13796
rect 21560 13793 21588 13824
rect 21913 13821 21925 13824
rect 21959 13821 21971 13855
rect 21913 13815 21971 13821
rect 22462 13812 22468 13864
rect 22520 13812 22526 13864
rect 22922 13812 22928 13864
rect 22980 13852 22986 13864
rect 23017 13855 23075 13861
rect 23017 13852 23029 13855
rect 22980 13824 23029 13852
rect 22980 13812 22986 13824
rect 23017 13821 23029 13824
rect 23063 13821 23075 13855
rect 23017 13815 23075 13821
rect 23106 13812 23112 13864
rect 23164 13812 23170 13864
rect 23198 13812 23204 13864
rect 23256 13812 23262 13864
rect 23293 13855 23351 13861
rect 23293 13821 23305 13855
rect 23339 13821 23351 13855
rect 23293 13815 23351 13821
rect 21545 13787 21603 13793
rect 21545 13784 21557 13787
rect 21416 13756 21557 13784
rect 21416 13744 21422 13756
rect 21545 13753 21557 13756
rect 21591 13753 21603 13787
rect 21545 13747 21603 13753
rect 22738 13744 22744 13796
rect 22796 13784 22802 13796
rect 23308 13784 23336 13815
rect 23382 13812 23388 13864
rect 23440 13852 23446 13864
rect 23658 13852 23664 13864
rect 23440 13824 23664 13852
rect 23440 13812 23446 13824
rect 23658 13812 23664 13824
rect 23716 13812 23722 13864
rect 24302 13852 24308 13864
rect 23768 13824 24308 13852
rect 23768 13784 23796 13824
rect 24302 13812 24308 13824
rect 24360 13812 24366 13864
rect 22796 13756 23796 13784
rect 22796 13744 22802 13756
rect 24210 13744 24216 13796
rect 24268 13784 24274 13796
rect 24397 13787 24455 13793
rect 24397 13784 24409 13787
rect 24268 13756 24409 13784
rect 24268 13744 24274 13756
rect 24397 13753 24409 13756
rect 24443 13753 24455 13787
rect 24504 13784 24532 13880
rect 24596 13852 24624 13960
rect 24872 13960 25421 13988
rect 24762 13880 24768 13932
rect 24820 13880 24826 13932
rect 24872 13929 24900 13960
rect 25409 13957 25421 13960
rect 25455 13957 25467 13991
rect 25409 13951 25467 13957
rect 24857 13923 24915 13929
rect 24857 13889 24869 13923
rect 24903 13889 24915 13923
rect 24857 13883 24915 13889
rect 25038 13880 25044 13932
rect 25096 13880 25102 13932
rect 25133 13923 25191 13929
rect 25133 13889 25145 13923
rect 25179 13889 25191 13923
rect 25133 13883 25191 13889
rect 25593 13923 25651 13929
rect 25593 13889 25605 13923
rect 25639 13889 25651 13923
rect 25593 13883 25651 13889
rect 25685 13923 25743 13929
rect 25685 13889 25697 13923
rect 25731 13920 25743 13923
rect 25774 13920 25780 13932
rect 25731 13892 25780 13920
rect 25731 13889 25743 13892
rect 25685 13883 25743 13889
rect 25148 13852 25176 13883
rect 25608 13852 25636 13883
rect 25774 13880 25780 13892
rect 25832 13880 25838 13932
rect 25884 13929 25912 14028
rect 26326 14016 26332 14068
rect 26384 14056 26390 14068
rect 26384 14028 26556 14056
rect 26384 14016 26390 14028
rect 26421 13991 26479 13997
rect 26421 13988 26433 13991
rect 25976 13960 26433 13988
rect 25976 13929 26004 13960
rect 26421 13957 26433 13960
rect 26467 13957 26479 13991
rect 26421 13951 26479 13957
rect 25869 13923 25927 13929
rect 25869 13889 25881 13923
rect 25915 13889 25927 13923
rect 25869 13883 25927 13889
rect 25961 13923 26019 13929
rect 25961 13889 25973 13923
rect 26007 13889 26019 13923
rect 25961 13883 26019 13889
rect 26050 13880 26056 13932
rect 26108 13880 26114 13932
rect 26142 13880 26148 13932
rect 26200 13920 26206 13932
rect 26528 13929 26556 14028
rect 27246 14016 27252 14068
rect 27304 14016 27310 14068
rect 28534 14016 28540 14068
rect 28592 14056 28598 14068
rect 29089 14059 29147 14065
rect 29089 14056 29101 14059
rect 28592 14028 29101 14056
rect 28592 14016 28598 14028
rect 29089 14025 29101 14028
rect 29135 14025 29147 14059
rect 29089 14019 29147 14025
rect 29270 14016 29276 14068
rect 29328 14056 29334 14068
rect 30190 14056 30196 14068
rect 29328 14028 30196 14056
rect 29328 14016 29334 14028
rect 30190 14016 30196 14028
rect 30248 14056 30254 14068
rect 31389 14059 31447 14065
rect 30248 14028 30788 14056
rect 30248 14016 30254 14028
rect 27264 13988 27292 14016
rect 26804 13960 27292 13988
rect 26237 13923 26295 13929
rect 26237 13920 26249 13923
rect 26200 13892 26249 13920
rect 26200 13880 26206 13892
rect 26237 13889 26249 13892
rect 26283 13889 26295 13923
rect 26237 13883 26295 13889
rect 26329 13923 26387 13929
rect 26329 13889 26341 13923
rect 26375 13920 26387 13923
rect 26513 13923 26571 13929
rect 26375 13892 26464 13920
rect 26375 13889 26387 13892
rect 26329 13883 26387 13889
rect 24596 13824 25176 13852
rect 25240 13824 25636 13852
rect 25792 13852 25820 13880
rect 26436 13864 26464 13892
rect 26513 13889 26525 13923
rect 26559 13889 26571 13923
rect 26513 13883 26571 13889
rect 26605 13923 26663 13929
rect 26605 13889 26617 13923
rect 26651 13920 26663 13923
rect 26694 13920 26700 13932
rect 26651 13892 26700 13920
rect 26651 13889 26663 13892
rect 26605 13883 26663 13889
rect 25792 13824 26192 13852
rect 25038 13784 25044 13796
rect 24504 13756 25044 13784
rect 24397 13747 24455 13753
rect 25038 13744 25044 13756
rect 25096 13744 25102 13796
rect 19668 13688 19840 13716
rect 19668 13676 19674 13688
rect 23106 13676 23112 13728
rect 23164 13716 23170 13728
rect 25240 13716 25268 13824
rect 25317 13787 25375 13793
rect 25317 13753 25329 13787
rect 25363 13784 25375 13787
rect 25958 13784 25964 13796
rect 25363 13756 25964 13784
rect 25363 13753 25375 13756
rect 25317 13747 25375 13753
rect 25958 13744 25964 13756
rect 26016 13744 26022 13796
rect 26164 13784 26192 13824
rect 26418 13812 26424 13864
rect 26476 13812 26482 13864
rect 26620 13784 26648 13883
rect 26694 13880 26700 13892
rect 26752 13880 26758 13932
rect 26804 13929 26832 13960
rect 27264 13929 27292 13960
rect 27798 13948 27804 14000
rect 27856 13988 27862 14000
rect 30760 13988 30788 14028
rect 31389 14025 31401 14059
rect 31435 14056 31447 14059
rect 31478 14056 31484 14068
rect 31435 14028 31484 14056
rect 31435 14025 31447 14028
rect 31389 14019 31447 14025
rect 31478 14016 31484 14028
rect 31536 14016 31542 14068
rect 32858 14016 32864 14068
rect 32916 14016 32922 14068
rect 32876 13988 32904 14016
rect 27856 13960 30236 13988
rect 27856 13948 27862 13960
rect 26789 13923 26847 13929
rect 26789 13889 26801 13923
rect 26835 13889 26847 13923
rect 27249 13923 27307 13929
rect 26789 13883 26847 13889
rect 27065 13913 27123 13919
rect 27065 13879 27077 13913
rect 27111 13879 27123 13913
rect 27249 13889 27261 13923
rect 27295 13889 27307 13923
rect 27249 13883 27307 13889
rect 27614 13880 27620 13932
rect 27672 13920 27678 13932
rect 28810 13920 28816 13932
rect 27672 13892 28816 13920
rect 27672 13880 27678 13892
rect 28810 13880 28816 13892
rect 28868 13880 28874 13932
rect 29089 13923 29147 13929
rect 29089 13889 29101 13923
rect 29135 13889 29147 13923
rect 29089 13883 29147 13889
rect 27065 13873 27123 13879
rect 27080 13784 27108 13873
rect 28905 13855 28963 13861
rect 28905 13821 28917 13855
rect 28951 13852 28963 13855
rect 28994 13852 29000 13864
rect 28951 13824 29000 13852
rect 28951 13821 28963 13824
rect 28905 13815 28963 13821
rect 28994 13812 29000 13824
rect 29052 13812 29058 13864
rect 29104 13784 29132 13883
rect 29178 13880 29184 13932
rect 29236 13920 29242 13932
rect 30208 13929 30236 13960
rect 30760 13960 32812 13988
rect 32876 13960 33088 13988
rect 29273 13923 29331 13929
rect 29273 13920 29285 13923
rect 29236 13892 29285 13920
rect 29236 13880 29242 13892
rect 29273 13889 29285 13892
rect 29319 13889 29331 13923
rect 29273 13883 29331 13889
rect 30193 13923 30251 13929
rect 30193 13889 30205 13923
rect 30239 13889 30251 13923
rect 30193 13883 30251 13889
rect 29288 13852 29316 13883
rect 30374 13880 30380 13932
rect 30432 13880 30438 13932
rect 30466 13880 30472 13932
rect 30524 13880 30530 13932
rect 30760 13929 30788 13960
rect 32784 13929 32812 13960
rect 30745 13923 30803 13929
rect 30745 13889 30757 13923
rect 30791 13889 30803 13923
rect 30745 13883 30803 13889
rect 30929 13923 30987 13929
rect 30929 13889 30941 13923
rect 30975 13920 30987 13923
rect 31941 13923 31999 13929
rect 31941 13920 31953 13923
rect 30975 13892 31953 13920
rect 30975 13889 30987 13892
rect 30929 13883 30987 13889
rect 31941 13889 31953 13892
rect 31987 13889 31999 13923
rect 31941 13883 31999 13889
rect 32769 13923 32827 13929
rect 32769 13889 32781 13923
rect 32815 13920 32827 13923
rect 32815 13892 32904 13920
rect 32815 13889 32827 13892
rect 32769 13883 32827 13889
rect 29288 13824 30420 13852
rect 26164 13756 27108 13784
rect 28552 13756 29132 13784
rect 30392 13784 30420 13824
rect 30558 13812 30564 13864
rect 30616 13812 30622 13864
rect 31665 13855 31723 13861
rect 30668 13824 31616 13852
rect 30668 13784 30696 13824
rect 30392 13756 30696 13784
rect 31588 13784 31616 13824
rect 31665 13821 31677 13855
rect 31711 13852 31723 13855
rect 32398 13852 32404 13864
rect 31711 13824 32404 13852
rect 31711 13821 31723 13824
rect 31665 13815 31723 13821
rect 32398 13812 32404 13824
rect 32456 13812 32462 13864
rect 32582 13784 32588 13796
rect 31588 13756 32588 13784
rect 28552 13728 28580 13756
rect 23164 13688 25268 13716
rect 23164 13676 23170 13688
rect 26050 13676 26056 13728
rect 26108 13716 26114 13728
rect 26145 13719 26203 13725
rect 26145 13716 26157 13719
rect 26108 13688 26157 13716
rect 26108 13676 26114 13688
rect 26145 13685 26157 13688
rect 26191 13685 26203 13719
rect 26145 13679 26203 13685
rect 26234 13676 26240 13728
rect 26292 13716 26298 13728
rect 26789 13719 26847 13725
rect 26789 13716 26801 13719
rect 26292 13688 26801 13716
rect 26292 13676 26298 13688
rect 26789 13685 26801 13688
rect 26835 13716 26847 13719
rect 26970 13716 26976 13728
rect 26835 13688 26976 13716
rect 26835 13685 26847 13688
rect 26789 13679 26847 13685
rect 26970 13676 26976 13688
rect 27028 13676 27034 13728
rect 27157 13719 27215 13725
rect 27157 13685 27169 13719
rect 27203 13716 27215 13719
rect 27338 13716 27344 13728
rect 27203 13688 27344 13716
rect 27203 13685 27215 13688
rect 27157 13679 27215 13685
rect 27338 13676 27344 13688
rect 27396 13676 27402 13728
rect 28534 13676 28540 13728
rect 28592 13676 28598 13728
rect 29104 13716 29132 13756
rect 32582 13744 32588 13756
rect 32640 13744 32646 13796
rect 32876 13784 32904 13892
rect 32950 13880 32956 13932
rect 33008 13880 33014 13932
rect 33060 13929 33088 13960
rect 33045 13923 33103 13929
rect 33045 13889 33057 13923
rect 33091 13889 33103 13923
rect 33045 13883 33103 13889
rect 33226 13880 33232 13932
rect 33284 13880 33290 13932
rect 32876 13756 33548 13784
rect 33520 13728 33548 13756
rect 29362 13716 29368 13728
rect 29104 13688 29368 13716
rect 29362 13676 29368 13688
rect 29420 13676 29426 13728
rect 30190 13676 30196 13728
rect 30248 13716 30254 13728
rect 30466 13716 30472 13728
rect 30248 13688 30472 13716
rect 30248 13676 30254 13688
rect 30466 13676 30472 13688
rect 30524 13676 30530 13728
rect 31846 13676 31852 13728
rect 31904 13676 31910 13728
rect 33134 13676 33140 13728
rect 33192 13716 33198 13728
rect 33229 13719 33287 13725
rect 33229 13716 33241 13719
rect 33192 13688 33241 13716
rect 33192 13676 33198 13688
rect 33229 13685 33241 13688
rect 33275 13685 33287 13719
rect 33229 13679 33287 13685
rect 33502 13676 33508 13728
rect 33560 13676 33566 13728
rect 1104 13626 38272 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 38272 13626
rect 1104 13552 38272 13574
rect 4249 13515 4307 13521
rect 4249 13481 4261 13515
rect 4295 13512 4307 13515
rect 9030 13512 9036 13524
rect 4295 13484 9036 13512
rect 4295 13481 4307 13484
rect 4249 13475 4307 13481
rect 9030 13472 9036 13484
rect 9088 13472 9094 13524
rect 10318 13472 10324 13524
rect 10376 13472 10382 13524
rect 10410 13472 10416 13524
rect 10468 13512 10474 13524
rect 10505 13515 10563 13521
rect 10505 13512 10517 13515
rect 10468 13484 10517 13512
rect 10468 13472 10474 13484
rect 10505 13481 10517 13484
rect 10551 13481 10563 13515
rect 11238 13512 11244 13524
rect 10505 13475 10563 13481
rect 10612 13484 11244 13512
rect 9125 13447 9183 13453
rect 9125 13413 9137 13447
rect 9171 13413 9183 13447
rect 9125 13407 9183 13413
rect 1394 13336 1400 13388
rect 1452 13376 1458 13388
rect 4341 13379 4399 13385
rect 4341 13376 4353 13379
rect 1452 13348 4353 13376
rect 1452 13336 1458 13348
rect 4341 13345 4353 13348
rect 4387 13376 4399 13379
rect 5626 13376 5632 13388
rect 4387 13348 5632 13376
rect 4387 13345 4399 13348
rect 4341 13339 4399 13345
rect 5626 13336 5632 13348
rect 5684 13336 5690 13388
rect 6270 13336 6276 13388
rect 6328 13376 6334 13388
rect 6365 13379 6423 13385
rect 6365 13376 6377 13379
rect 6328 13348 6377 13376
rect 6328 13336 6334 13348
rect 6365 13345 6377 13348
rect 6411 13345 6423 13379
rect 6914 13376 6920 13388
rect 6365 13339 6423 13345
rect 6472 13348 6920 13376
rect 2958 13268 2964 13320
rect 3016 13308 3022 13320
rect 3786 13308 3792 13320
rect 3016 13280 3792 13308
rect 3016 13268 3022 13280
rect 3786 13268 3792 13280
rect 3844 13308 3850 13320
rect 3881 13311 3939 13317
rect 3881 13308 3893 13311
rect 3844 13280 3893 13308
rect 3844 13268 3850 13280
rect 3881 13277 3893 13280
rect 3927 13277 3939 13311
rect 3881 13271 3939 13277
rect 3970 13200 3976 13252
rect 4028 13240 4034 13252
rect 4065 13243 4123 13249
rect 4065 13240 4077 13243
rect 4028 13212 4077 13240
rect 4028 13200 4034 13212
rect 4065 13209 4077 13212
rect 4111 13209 4123 13243
rect 4065 13203 4123 13209
rect 4614 13200 4620 13252
rect 4672 13200 4678 13252
rect 5000 13212 5106 13240
rect 2774 13132 2780 13184
rect 2832 13172 2838 13184
rect 5000 13172 5028 13212
rect 6472 13172 6500 13348
rect 6914 13336 6920 13348
rect 6972 13336 6978 13388
rect 7098 13336 7104 13388
rect 7156 13336 7162 13388
rect 8757 13311 8815 13317
rect 8757 13277 8769 13311
rect 8803 13308 8815 13311
rect 9140 13308 9168 13407
rect 9582 13336 9588 13388
rect 9640 13336 9646 13388
rect 9769 13379 9827 13385
rect 9769 13345 9781 13379
rect 9815 13376 9827 13379
rect 10336 13376 10364 13472
rect 9815 13348 10364 13376
rect 9815 13345 9827 13348
rect 9769 13339 9827 13345
rect 8803 13280 9168 13308
rect 8803 13277 8815 13280
rect 8757 13271 8815 13277
rect 9214 13268 9220 13320
rect 9272 13308 9278 13320
rect 9600 13308 9628 13336
rect 9272 13280 10088 13308
rect 9272 13268 9278 13280
rect 6917 13243 6975 13249
rect 6917 13209 6929 13243
rect 6963 13240 6975 13243
rect 9950 13240 9956 13252
rect 6963 13212 9956 13240
rect 6963 13209 6975 13212
rect 6917 13203 6975 13209
rect 9950 13200 9956 13212
rect 10008 13200 10014 13252
rect 10060 13240 10088 13280
rect 10134 13268 10140 13320
rect 10192 13268 10198 13320
rect 10612 13317 10640 13484
rect 11238 13472 11244 13484
rect 11296 13472 11302 13524
rect 15286 13472 15292 13524
rect 15344 13512 15350 13524
rect 15381 13515 15439 13521
rect 15381 13512 15393 13515
rect 15344 13484 15393 13512
rect 15344 13472 15350 13484
rect 15381 13481 15393 13484
rect 15427 13481 15439 13515
rect 15381 13475 15439 13481
rect 16669 13515 16727 13521
rect 16669 13481 16681 13515
rect 16715 13481 16727 13515
rect 16669 13475 16727 13481
rect 13541 13447 13599 13453
rect 13541 13413 13553 13447
rect 13587 13413 13599 13447
rect 16684 13444 16712 13475
rect 16850 13472 16856 13524
rect 16908 13512 16914 13524
rect 17862 13512 17868 13524
rect 16908 13484 17868 13512
rect 16908 13472 16914 13484
rect 17862 13472 17868 13484
rect 17920 13472 17926 13524
rect 18414 13472 18420 13524
rect 18472 13472 18478 13524
rect 18877 13515 18935 13521
rect 18877 13512 18889 13515
rect 18524 13484 18889 13512
rect 16758 13444 16764 13456
rect 16684 13416 16764 13444
rect 13541 13407 13599 13413
rect 10965 13379 11023 13385
rect 10965 13345 10977 13379
rect 11011 13376 11023 13379
rect 11882 13376 11888 13388
rect 11011 13348 11888 13376
rect 11011 13345 11023 13348
rect 10965 13339 11023 13345
rect 11882 13336 11888 13348
rect 11940 13336 11946 13388
rect 12526 13336 12532 13388
rect 12584 13376 12590 13388
rect 12897 13379 12955 13385
rect 12897 13376 12909 13379
rect 12584 13348 12909 13376
rect 12584 13336 12590 13348
rect 12897 13345 12909 13348
rect 12943 13345 12955 13379
rect 12897 13339 12955 13345
rect 10229 13311 10287 13317
rect 10229 13277 10241 13311
rect 10275 13277 10287 13311
rect 10229 13271 10287 13277
rect 10597 13311 10655 13317
rect 10597 13277 10609 13311
rect 10643 13277 10655 13311
rect 10597 13271 10655 13277
rect 10689 13311 10747 13317
rect 10689 13277 10701 13311
rect 10735 13277 10747 13311
rect 10689 13271 10747 13277
rect 10244 13240 10272 13271
rect 10060 13212 10272 13240
rect 10704 13240 10732 13271
rect 13078 13268 13084 13320
rect 13136 13308 13142 13320
rect 13173 13311 13231 13317
rect 13173 13308 13185 13311
rect 13136 13280 13185 13308
rect 13136 13268 13142 13280
rect 13173 13277 13185 13280
rect 13219 13277 13231 13311
rect 13556 13308 13584 13407
rect 16758 13404 16764 13416
rect 16816 13444 16822 13456
rect 17586 13444 17592 13456
rect 16816 13416 17592 13444
rect 16816 13404 16822 13416
rect 17586 13404 17592 13416
rect 17644 13404 17650 13456
rect 18524 13444 18552 13484
rect 18877 13481 18889 13484
rect 18923 13481 18935 13515
rect 18877 13475 18935 13481
rect 19702 13472 19708 13524
rect 19760 13472 19766 13524
rect 20625 13515 20683 13521
rect 20625 13512 20637 13515
rect 19996 13484 20637 13512
rect 18432 13416 18552 13444
rect 18432 13388 18460 13416
rect 19242 13404 19248 13456
rect 19300 13444 19306 13456
rect 19334 13444 19340 13456
rect 19300 13416 19340 13444
rect 19300 13404 19306 13416
rect 19334 13404 19340 13416
rect 19392 13404 19398 13456
rect 16942 13336 16948 13388
rect 17000 13376 17006 13388
rect 17000 13348 17816 13376
rect 17000 13336 17006 13348
rect 13817 13311 13875 13317
rect 13817 13308 13829 13311
rect 13556 13280 13829 13308
rect 13173 13271 13231 13277
rect 13817 13277 13829 13280
rect 13863 13277 13875 13311
rect 13817 13271 13875 13277
rect 15013 13311 15071 13317
rect 15013 13277 15025 13311
rect 15059 13308 15071 13311
rect 15102 13308 15108 13320
rect 15059 13280 15108 13308
rect 15059 13277 15071 13280
rect 15013 13271 15071 13277
rect 15102 13268 15108 13280
rect 15160 13268 15166 13320
rect 16022 13268 16028 13320
rect 16080 13308 16086 13320
rect 17788 13317 17816 13348
rect 18414 13336 18420 13388
rect 18472 13336 18478 13388
rect 19996 13376 20024 13484
rect 20625 13481 20637 13484
rect 20671 13512 20683 13515
rect 20898 13512 20904 13524
rect 20671 13484 20904 13512
rect 20671 13481 20683 13484
rect 20625 13475 20683 13481
rect 20898 13472 20904 13484
rect 20956 13472 20962 13524
rect 27433 13515 27491 13521
rect 21008 13484 27200 13512
rect 20438 13444 20444 13456
rect 18616 13348 20024 13376
rect 17773 13311 17831 13317
rect 16080 13280 16804 13308
rect 16080 13268 16086 13280
rect 11146 13240 11152 13252
rect 10704 13212 11152 13240
rect 11146 13200 11152 13212
rect 11204 13200 11210 13252
rect 11241 13243 11299 13249
rect 11241 13209 11253 13243
rect 11287 13209 11299 13243
rect 11698 13240 11704 13252
rect 11241 13203 11299 13209
rect 11624 13212 11704 13240
rect 2832 13144 6500 13172
rect 2832 13132 2838 13144
rect 6546 13132 6552 13184
rect 6604 13132 6610 13184
rect 7009 13175 7067 13181
rect 7009 13141 7021 13175
rect 7055 13172 7067 13175
rect 8018 13172 8024 13184
rect 7055 13144 8024 13172
rect 7055 13141 7067 13144
rect 7009 13135 7067 13141
rect 8018 13132 8024 13144
rect 8076 13132 8082 13184
rect 8570 13132 8576 13184
rect 8628 13132 8634 13184
rect 9398 13132 9404 13184
rect 9456 13172 9462 13184
rect 9493 13175 9551 13181
rect 9493 13172 9505 13175
rect 9456 13144 9505 13172
rect 9456 13132 9462 13144
rect 9493 13141 9505 13144
rect 9539 13141 9551 13175
rect 9493 13135 9551 13141
rect 9582 13132 9588 13184
rect 9640 13132 9646 13184
rect 10873 13175 10931 13181
rect 10873 13141 10885 13175
rect 10919 13172 10931 13175
rect 11256 13172 11284 13203
rect 10919 13144 11284 13172
rect 11624 13172 11652 13212
rect 11698 13200 11704 13212
rect 11756 13200 11762 13252
rect 12406 13212 13492 13240
rect 12406 13172 12434 13212
rect 11624 13144 12434 13172
rect 10919 13141 10931 13144
rect 10873 13135 10931 13141
rect 12710 13132 12716 13184
rect 12768 13132 12774 13184
rect 13081 13175 13139 13181
rect 13081 13141 13093 13175
rect 13127 13172 13139 13175
rect 13354 13172 13360 13184
rect 13127 13144 13360 13172
rect 13127 13141 13139 13144
rect 13081 13135 13139 13141
rect 13354 13132 13360 13144
rect 13412 13132 13418 13184
rect 13464 13172 13492 13212
rect 15194 13200 15200 13252
rect 15252 13200 15258 13252
rect 16666 13200 16672 13252
rect 16724 13200 16730 13252
rect 13538 13172 13544 13184
rect 13464 13144 13544 13172
rect 13538 13132 13544 13144
rect 13596 13132 13602 13184
rect 13630 13132 13636 13184
rect 13688 13132 13694 13184
rect 15470 13132 15476 13184
rect 15528 13172 15534 13184
rect 16485 13175 16543 13181
rect 16485 13172 16497 13175
rect 15528 13144 16497 13172
rect 15528 13132 15534 13144
rect 16485 13141 16497 13144
rect 16531 13141 16543 13175
rect 16776 13172 16804 13280
rect 17773 13277 17785 13311
rect 17819 13308 17831 13311
rect 17819 13280 18368 13308
rect 18616 13302 18644 13348
rect 19996 13320 20024 13348
rect 20088 13416 20444 13444
rect 20088 13320 20116 13416
rect 20438 13404 20444 13416
rect 20496 13404 20502 13456
rect 20180 13348 20576 13376
rect 17819 13277 17831 13280
rect 17773 13271 17831 13277
rect 16850 13200 16856 13252
rect 16908 13200 16914 13252
rect 18230 13200 18236 13252
rect 18288 13200 18294 13252
rect 18340 13240 18368 13280
rect 18524 13274 18644 13302
rect 18524 13240 18552 13274
rect 19518 13268 19524 13320
rect 19576 13268 19582 13320
rect 19978 13268 19984 13320
rect 20036 13268 20042 13320
rect 20070 13268 20076 13320
rect 20128 13268 20134 13320
rect 20180 13317 20208 13348
rect 20548 13320 20576 13348
rect 20622 13336 20628 13388
rect 20680 13376 20686 13388
rect 21008 13385 21036 13484
rect 22649 13447 22707 13453
rect 22649 13413 22661 13447
rect 22695 13444 22707 13447
rect 22738 13444 22744 13456
rect 22695 13416 22744 13444
rect 22695 13413 22707 13416
rect 22649 13407 22707 13413
rect 22738 13404 22744 13416
rect 22796 13404 22802 13456
rect 22925 13447 22983 13453
rect 22925 13413 22937 13447
rect 22971 13444 22983 13447
rect 23106 13444 23112 13456
rect 22971 13416 23112 13444
rect 22971 13413 22983 13416
rect 22925 13407 22983 13413
rect 23106 13404 23112 13416
rect 23164 13404 23170 13456
rect 27062 13444 27068 13456
rect 24504 13416 27068 13444
rect 20993 13379 21051 13385
rect 20993 13376 21005 13379
rect 20680 13348 21005 13376
rect 20680 13336 20686 13348
rect 20993 13345 21005 13348
rect 21039 13345 21051 13379
rect 20993 13339 21051 13345
rect 20165 13311 20223 13317
rect 20165 13277 20177 13311
rect 20211 13277 20223 13311
rect 20165 13271 20223 13277
rect 20349 13311 20407 13317
rect 20349 13277 20361 13311
rect 20395 13277 20407 13311
rect 20349 13271 20407 13277
rect 18874 13249 18880 13252
rect 18861 13243 18880 13249
rect 18340 13212 18552 13240
rect 18616 13212 18828 13240
rect 18414 13172 18420 13184
rect 18472 13181 18478 13184
rect 18616 13181 18644 13212
rect 18472 13175 18491 13181
rect 16776 13144 18420 13172
rect 16485 13135 16543 13141
rect 18414 13132 18420 13144
rect 18479 13141 18491 13175
rect 18472 13135 18491 13141
rect 18601 13175 18659 13181
rect 18601 13141 18613 13175
rect 18647 13141 18659 13175
rect 18601 13135 18659 13141
rect 18472 13132 18478 13135
rect 18690 13132 18696 13184
rect 18748 13132 18754 13184
rect 18800 13172 18828 13212
rect 18861 13209 18873 13243
rect 18861 13203 18880 13209
rect 18874 13200 18880 13203
rect 18932 13200 18938 13252
rect 18966 13200 18972 13252
rect 19024 13240 19030 13252
rect 19061 13243 19119 13249
rect 19061 13240 19073 13243
rect 19024 13212 19073 13240
rect 19024 13200 19030 13212
rect 19061 13209 19073 13212
rect 19107 13209 19119 13243
rect 19536 13240 19564 13268
rect 20364 13240 20392 13271
rect 20530 13268 20536 13320
rect 20588 13268 20594 13320
rect 21082 13268 21088 13320
rect 21140 13268 21146 13320
rect 21358 13268 21364 13320
rect 21416 13268 21422 13320
rect 21726 13268 21732 13320
rect 21784 13268 21790 13320
rect 21910 13268 21916 13320
rect 21968 13308 21974 13320
rect 22373 13311 22431 13317
rect 22373 13308 22385 13311
rect 21968 13280 22385 13308
rect 21968 13268 21974 13280
rect 22373 13277 22385 13280
rect 22419 13277 22431 13311
rect 22373 13271 22431 13277
rect 22557 13311 22615 13317
rect 22557 13277 22569 13311
rect 22603 13308 22615 13311
rect 22925 13311 22983 13317
rect 22925 13308 22937 13311
rect 22603 13280 22937 13308
rect 22603 13277 22615 13280
rect 22557 13271 22615 13277
rect 22925 13277 22937 13280
rect 22971 13277 22983 13311
rect 22925 13271 22983 13277
rect 20441 13243 20499 13249
rect 20441 13240 20453 13243
rect 19536 13212 20453 13240
rect 19061 13203 19119 13209
rect 20441 13209 20453 13212
rect 20487 13209 20499 13243
rect 20548 13240 20576 13268
rect 20641 13243 20699 13249
rect 20641 13240 20653 13243
rect 20548 13212 20653 13240
rect 20441 13203 20499 13209
rect 20641 13209 20653 13212
rect 20687 13209 20699 13243
rect 22572 13240 22600 13271
rect 20641 13203 20699 13209
rect 21192 13212 22600 13240
rect 22940 13240 22968 13271
rect 23198 13268 23204 13320
rect 23256 13308 23262 13320
rect 23477 13311 23535 13317
rect 23477 13308 23489 13311
rect 23256 13280 23489 13308
rect 23256 13268 23262 13280
rect 23477 13277 23489 13280
rect 23523 13277 23535 13311
rect 23477 13271 23535 13277
rect 24118 13268 24124 13320
rect 24176 13308 24182 13320
rect 24397 13311 24455 13317
rect 24397 13308 24409 13311
rect 24176 13280 24409 13308
rect 24176 13268 24182 13280
rect 24397 13277 24409 13280
rect 24443 13277 24455 13311
rect 24397 13271 24455 13277
rect 24504 13252 24532 13416
rect 24765 13379 24823 13385
rect 24765 13345 24777 13379
rect 24811 13376 24823 13379
rect 25774 13376 25780 13388
rect 24811 13348 25780 13376
rect 24811 13345 24823 13348
rect 24765 13339 24823 13345
rect 25774 13336 25780 13348
rect 25832 13336 25838 13388
rect 26050 13376 26056 13388
rect 25976 13348 26056 13376
rect 24581 13311 24639 13317
rect 24581 13277 24593 13311
rect 24627 13277 24639 13311
rect 24581 13271 24639 13277
rect 23293 13243 23351 13249
rect 23293 13240 23305 13243
rect 22940 13212 23305 13240
rect 21192 13184 21220 13212
rect 23293 13209 23305 13212
rect 23339 13209 23351 13243
rect 23293 13203 23351 13209
rect 23661 13243 23719 13249
rect 23661 13209 23673 13243
rect 23707 13240 23719 13243
rect 24486 13240 24492 13252
rect 23707 13212 24492 13240
rect 23707 13209 23719 13212
rect 23661 13203 23719 13209
rect 24486 13200 24492 13212
rect 24544 13200 24550 13252
rect 19242 13172 19248 13184
rect 18800 13144 19248 13172
rect 19242 13132 19248 13144
rect 19300 13132 19306 13184
rect 20809 13175 20867 13181
rect 20809 13141 20821 13175
rect 20855 13172 20867 13175
rect 21082 13172 21088 13184
rect 20855 13144 21088 13172
rect 20855 13141 20867 13144
rect 20809 13135 20867 13141
rect 21082 13132 21088 13144
rect 21140 13132 21146 13184
rect 21174 13132 21180 13184
rect 21232 13132 21238 13184
rect 21542 13132 21548 13184
rect 21600 13172 21606 13184
rect 22738 13172 22744 13184
rect 21600 13144 22744 13172
rect 21600 13132 21606 13144
rect 22738 13132 22744 13144
rect 22796 13132 22802 13184
rect 22922 13132 22928 13184
rect 22980 13172 22986 13184
rect 23106 13172 23112 13184
rect 22980 13144 23112 13172
rect 22980 13132 22986 13144
rect 23106 13132 23112 13144
rect 23164 13132 23170 13184
rect 24596 13172 24624 13271
rect 25590 13268 25596 13320
rect 25648 13308 25654 13320
rect 25685 13311 25743 13317
rect 25685 13308 25697 13311
rect 25648 13280 25697 13308
rect 25648 13268 25654 13280
rect 25685 13277 25697 13280
rect 25731 13277 25743 13311
rect 25685 13271 25743 13277
rect 25866 13268 25872 13320
rect 25924 13268 25930 13320
rect 25976 13317 26004 13348
rect 26050 13336 26056 13348
rect 26108 13336 26114 13388
rect 26234 13336 26240 13388
rect 26292 13336 26298 13388
rect 26344 13385 26372 13416
rect 27062 13404 27068 13416
rect 27120 13404 27126 13456
rect 27172 13444 27200 13484
rect 27433 13481 27445 13515
rect 27479 13512 27491 13515
rect 27798 13512 27804 13524
rect 27479 13484 27804 13512
rect 27479 13481 27491 13484
rect 27433 13475 27491 13481
rect 27798 13472 27804 13484
rect 27856 13472 27862 13524
rect 27890 13472 27896 13524
rect 27948 13512 27954 13524
rect 28077 13515 28135 13521
rect 28077 13512 28089 13515
rect 27948 13484 28089 13512
rect 27948 13472 27954 13484
rect 28077 13481 28089 13484
rect 28123 13481 28135 13515
rect 28077 13475 28135 13481
rect 28166 13472 28172 13524
rect 28224 13512 28230 13524
rect 28353 13515 28411 13521
rect 28353 13512 28365 13515
rect 28224 13484 28365 13512
rect 28224 13472 28230 13484
rect 28353 13481 28365 13484
rect 28399 13512 28411 13515
rect 28442 13512 28448 13524
rect 28399 13484 28448 13512
rect 28399 13481 28411 13484
rect 28353 13475 28411 13481
rect 28442 13472 28448 13484
rect 28500 13472 28506 13524
rect 28994 13472 29000 13524
rect 29052 13512 29058 13524
rect 29089 13515 29147 13521
rect 29089 13512 29101 13515
rect 29052 13484 29101 13512
rect 29052 13472 29058 13484
rect 29089 13481 29101 13484
rect 29135 13481 29147 13515
rect 29089 13475 29147 13481
rect 29178 13472 29184 13524
rect 29236 13512 29242 13524
rect 29236 13484 30328 13512
rect 29236 13472 29242 13484
rect 30300 13456 30328 13484
rect 32398 13472 32404 13524
rect 32456 13512 32462 13524
rect 33137 13515 33195 13521
rect 33137 13512 33149 13515
rect 32456 13484 33149 13512
rect 32456 13472 32462 13484
rect 33137 13481 33149 13484
rect 33183 13481 33195 13515
rect 33137 13475 33195 13481
rect 33226 13472 33232 13524
rect 33284 13472 33290 13524
rect 33410 13472 33416 13524
rect 33468 13512 33474 13524
rect 33689 13515 33747 13521
rect 33689 13512 33701 13515
rect 33468 13484 33701 13512
rect 33468 13472 33474 13484
rect 33689 13481 33701 13484
rect 33735 13481 33747 13515
rect 33689 13475 33747 13481
rect 28258 13444 28264 13456
rect 27172 13416 28264 13444
rect 28258 13404 28264 13416
rect 28316 13404 28322 13456
rect 30282 13404 30288 13456
rect 30340 13404 30346 13456
rect 33428 13444 33456 13472
rect 32968 13416 33456 13444
rect 26329 13379 26387 13385
rect 26329 13345 26341 13379
rect 26375 13345 26387 13379
rect 26329 13339 26387 13345
rect 26697 13379 26755 13385
rect 26697 13345 26709 13379
rect 26743 13376 26755 13379
rect 26743 13348 27016 13376
rect 26743 13345 26755 13348
rect 26697 13339 26755 13345
rect 25961 13311 26019 13317
rect 25961 13277 25973 13311
rect 26007 13277 26019 13311
rect 25961 13271 26019 13277
rect 26142 13268 26148 13320
rect 26200 13268 26206 13320
rect 26510 13268 26516 13320
rect 26568 13268 26574 13320
rect 26786 13268 26792 13320
rect 26844 13268 26850 13320
rect 26988 13317 27016 13348
rect 27338 13336 27344 13388
rect 27396 13376 27402 13388
rect 32968 13385 32996 13416
rect 28997 13379 29055 13385
rect 28997 13376 29009 13379
rect 27396 13348 29009 13376
rect 27396 13336 27402 13348
rect 28997 13345 29009 13348
rect 29043 13345 29055 13379
rect 32953 13379 33011 13385
rect 28997 13339 29055 13345
rect 29196 13348 29776 13376
rect 26973 13311 27031 13317
rect 26973 13277 26985 13311
rect 27019 13277 27031 13311
rect 26973 13271 27031 13277
rect 27065 13311 27123 13317
rect 27065 13277 27077 13311
rect 27111 13277 27123 13311
rect 27177 13311 27235 13317
rect 27177 13308 27189 13311
rect 27065 13271 27123 13277
rect 27172 13277 27189 13308
rect 27223 13308 27235 13311
rect 27356 13308 27384 13336
rect 27223 13280 27384 13308
rect 27223 13277 27235 13280
rect 27172 13271 27235 13277
rect 26878 13200 26884 13252
rect 26936 13240 26942 13252
rect 27080 13240 27108 13271
rect 26936 13212 27108 13240
rect 26936 13200 26942 13212
rect 24854 13172 24860 13184
rect 24596 13144 24860 13172
rect 24854 13132 24860 13144
rect 24912 13132 24918 13184
rect 25777 13175 25835 13181
rect 25777 13141 25789 13175
rect 25823 13172 25835 13175
rect 26234 13172 26240 13184
rect 25823 13144 26240 13172
rect 25823 13141 25835 13144
rect 25777 13135 25835 13141
rect 26234 13132 26240 13144
rect 26292 13132 26298 13184
rect 26694 13132 26700 13184
rect 26752 13172 26758 13184
rect 27172 13172 27200 13271
rect 27430 13268 27436 13320
rect 27488 13308 27494 13320
rect 28350 13308 28356 13320
rect 27488 13280 28356 13308
rect 27488 13268 27494 13280
rect 28350 13268 28356 13280
rect 28408 13268 28414 13320
rect 28445 13311 28503 13317
rect 28445 13277 28457 13311
rect 28491 13277 28503 13311
rect 28445 13271 28503 13277
rect 28460 13240 28488 13271
rect 28534 13268 28540 13320
rect 28592 13268 28598 13320
rect 28721 13311 28779 13317
rect 28721 13277 28733 13311
rect 28767 13308 28779 13311
rect 29196 13308 29224 13348
rect 28767 13280 29224 13308
rect 28767 13277 28779 13280
rect 28721 13271 28779 13277
rect 29270 13268 29276 13320
rect 29328 13268 29334 13320
rect 29362 13268 29368 13320
rect 29420 13308 29426 13320
rect 29748 13317 29776 13348
rect 32953 13345 32965 13379
rect 32999 13345 33011 13379
rect 34057 13379 34115 13385
rect 34057 13376 34069 13379
rect 32953 13339 33011 13345
rect 33152 13348 34069 13376
rect 33152 13320 33180 13348
rect 34057 13345 34069 13348
rect 34103 13345 34115 13379
rect 34057 13339 34115 13345
rect 29549 13311 29607 13317
rect 29549 13308 29561 13311
rect 29420 13280 29561 13308
rect 29420 13268 29426 13280
rect 29549 13277 29561 13280
rect 29595 13277 29607 13311
rect 29549 13271 29607 13277
rect 29733 13311 29791 13317
rect 29733 13277 29745 13311
rect 29779 13308 29791 13311
rect 31202 13308 31208 13320
rect 29779 13280 31208 13308
rect 29779 13277 29791 13280
rect 29733 13271 29791 13277
rect 31202 13268 31208 13280
rect 31260 13268 31266 13320
rect 32858 13268 32864 13320
rect 32916 13268 32922 13320
rect 33134 13268 33140 13320
rect 33192 13268 33198 13320
rect 33413 13311 33471 13317
rect 33413 13277 33425 13311
rect 33459 13277 33471 13311
rect 33413 13271 33471 13277
rect 28460 13212 29684 13240
rect 29656 13184 29684 13212
rect 32398 13200 32404 13252
rect 32456 13240 32462 13252
rect 32493 13243 32551 13249
rect 32493 13240 32505 13243
rect 32456 13212 32505 13240
rect 32456 13200 32462 13212
rect 32493 13209 32505 13212
rect 32539 13209 32551 13243
rect 32493 13203 32551 13209
rect 32582 13200 32588 13252
rect 32640 13200 32646 13252
rect 33042 13200 33048 13252
rect 33100 13240 33106 13252
rect 33428 13240 33456 13271
rect 33502 13268 33508 13320
rect 33560 13268 33566 13320
rect 33870 13268 33876 13320
rect 33928 13268 33934 13320
rect 33100 13212 33456 13240
rect 33100 13200 33106 13212
rect 26752 13144 27200 13172
rect 26752 13132 26758 13144
rect 29638 13132 29644 13184
rect 29696 13132 29702 13184
rect 1104 13082 38272 13104
rect 1104 13030 4874 13082
rect 4926 13030 4938 13082
rect 4990 13030 5002 13082
rect 5054 13030 5066 13082
rect 5118 13030 5130 13082
rect 5182 13030 35594 13082
rect 35646 13030 35658 13082
rect 35710 13030 35722 13082
rect 35774 13030 35786 13082
rect 35838 13030 35850 13082
rect 35902 13030 38272 13082
rect 1104 13008 38272 13030
rect 3145 12971 3203 12977
rect 3145 12937 3157 12971
rect 3191 12968 3203 12971
rect 3970 12968 3976 12980
rect 3191 12940 3976 12968
rect 3191 12937 3203 12940
rect 3145 12931 3203 12937
rect 3970 12928 3976 12940
rect 4028 12928 4034 12980
rect 4614 12928 4620 12980
rect 4672 12968 4678 12980
rect 4985 12971 5043 12977
rect 4985 12968 4997 12971
rect 4672 12940 4997 12968
rect 4672 12928 4678 12940
rect 4985 12937 4997 12940
rect 5031 12937 5043 12971
rect 4985 12931 5043 12937
rect 6546 12928 6552 12980
rect 6604 12928 6610 12980
rect 7024 12940 7788 12968
rect 4065 12903 4123 12909
rect 4065 12869 4077 12903
rect 4111 12900 4123 12903
rect 4525 12903 4583 12909
rect 4525 12900 4537 12903
rect 4111 12872 4537 12900
rect 4111 12869 4123 12872
rect 4065 12863 4123 12869
rect 4525 12869 4537 12872
rect 4571 12869 4583 12903
rect 6564 12900 6592 12928
rect 4525 12863 4583 12869
rect 6012 12872 6592 12900
rect 1394 12792 1400 12844
rect 1452 12792 1458 12844
rect 2774 12792 2780 12844
rect 2832 12792 2838 12844
rect 3970 12792 3976 12844
rect 4028 12792 4034 12844
rect 4430 12792 4436 12844
rect 4488 12792 4494 12844
rect 4617 12835 4675 12841
rect 4617 12801 4629 12835
rect 4663 12832 4675 12835
rect 4706 12832 4712 12844
rect 4663 12804 4712 12832
rect 4663 12801 4675 12804
rect 4617 12795 4675 12801
rect 1670 12724 1676 12776
rect 1728 12724 1734 12776
rect 3878 12724 3884 12776
rect 3936 12764 3942 12776
rect 4157 12767 4215 12773
rect 4157 12764 4169 12767
rect 3936 12736 4169 12764
rect 3936 12724 3942 12736
rect 4157 12733 4169 12736
rect 4203 12733 4215 12767
rect 4157 12727 4215 12733
rect 3786 12656 3792 12708
rect 3844 12696 3850 12708
rect 4632 12696 4660 12795
rect 4706 12792 4712 12804
rect 4764 12792 4770 12844
rect 5169 12835 5227 12841
rect 5169 12801 5181 12835
rect 5215 12832 5227 12835
rect 5810 12832 5816 12844
rect 5215 12804 5816 12832
rect 5215 12801 5227 12804
rect 5169 12795 5227 12801
rect 5810 12792 5816 12804
rect 5868 12792 5874 12844
rect 6012 12841 6040 12872
rect 6914 12860 6920 12912
rect 6972 12900 6978 12912
rect 7024 12900 7052 12940
rect 6972 12872 7130 12900
rect 6972 12860 6978 12872
rect 5997 12835 6055 12841
rect 5997 12801 6009 12835
rect 6043 12801 6055 12835
rect 5997 12795 6055 12801
rect 6362 12792 6368 12844
rect 6420 12792 6426 12844
rect 6641 12767 6699 12773
rect 6641 12764 6653 12767
rect 6196 12736 6653 12764
rect 6196 12705 6224 12736
rect 6641 12733 6653 12736
rect 6687 12733 6699 12767
rect 7760 12764 7788 12940
rect 8018 12928 8024 12980
rect 8076 12968 8082 12980
rect 8113 12971 8171 12977
rect 8113 12968 8125 12971
rect 8076 12940 8125 12968
rect 8076 12928 8082 12940
rect 8113 12937 8125 12940
rect 8159 12937 8171 12971
rect 9858 12968 9864 12980
rect 8113 12931 8171 12937
rect 8312 12940 9864 12968
rect 8312 12841 8340 12940
rect 9858 12928 9864 12940
rect 9916 12928 9922 12980
rect 10410 12928 10416 12980
rect 10468 12928 10474 12980
rect 10505 12971 10563 12977
rect 10505 12937 10517 12971
rect 10551 12968 10563 12971
rect 13630 12968 13636 12980
rect 10551 12940 11836 12968
rect 10551 12937 10563 12940
rect 10505 12931 10563 12937
rect 8570 12860 8576 12912
rect 8628 12860 8634 12912
rect 8297 12835 8355 12841
rect 8297 12801 8309 12835
rect 8343 12801 8355 12835
rect 8297 12795 8355 12801
rect 9674 12792 9680 12844
rect 9732 12792 9738 12844
rect 10226 12792 10232 12844
rect 10284 12832 10290 12844
rect 10321 12835 10379 12841
rect 10321 12832 10333 12835
rect 10284 12804 10333 12832
rect 10284 12792 10290 12804
rect 10321 12801 10333 12804
rect 10367 12801 10379 12835
rect 10428 12832 10456 12928
rect 10597 12835 10655 12841
rect 10597 12832 10609 12835
rect 10428 12804 10609 12832
rect 10321 12795 10379 12801
rect 10597 12801 10609 12804
rect 10643 12801 10655 12835
rect 10597 12795 10655 12801
rect 9692 12764 9720 12792
rect 7760 12736 9720 12764
rect 6641 12727 6699 12733
rect 3844 12668 4660 12696
rect 6181 12699 6239 12705
rect 3844 12656 3850 12668
rect 6181 12665 6193 12699
rect 6227 12665 6239 12699
rect 6181 12659 6239 12665
rect 9582 12656 9588 12708
rect 9640 12696 9646 12708
rect 10045 12699 10103 12705
rect 10045 12696 10057 12699
rect 9640 12668 10057 12696
rect 9640 12656 9646 12668
rect 10045 12665 10057 12668
rect 10091 12696 10103 12699
rect 10704 12696 10732 12940
rect 11808 12832 11836 12940
rect 13464 12940 13636 12968
rect 11882 12860 11888 12912
rect 11940 12900 11946 12912
rect 13464 12909 13492 12940
rect 13630 12928 13636 12940
rect 13688 12928 13694 12980
rect 14921 12971 14979 12977
rect 13832 12940 14780 12968
rect 13449 12903 13507 12909
rect 11940 12872 13216 12900
rect 11940 12860 11946 12872
rect 11808 12804 12388 12832
rect 12250 12724 12256 12776
rect 12308 12724 12314 12776
rect 12360 12764 12388 12804
rect 12710 12792 12716 12844
rect 12768 12832 12774 12844
rect 13188 12841 13216 12872
rect 13449 12869 13461 12903
rect 13495 12869 13507 12903
rect 13449 12863 13507 12869
rect 13538 12860 13544 12912
rect 13596 12900 13602 12912
rect 13832 12900 13860 12940
rect 13596 12872 13938 12900
rect 13596 12860 13602 12872
rect 13081 12835 13139 12841
rect 13081 12832 13093 12835
rect 12768 12804 13093 12832
rect 12768 12792 12774 12804
rect 13081 12801 13093 12804
rect 13127 12801 13139 12835
rect 13081 12795 13139 12801
rect 13173 12835 13231 12841
rect 13173 12801 13185 12835
rect 13219 12801 13231 12835
rect 14752 12832 14780 12940
rect 14921 12937 14933 12971
rect 14967 12968 14979 12971
rect 15194 12968 15200 12980
rect 14967 12940 15200 12968
rect 14967 12937 14979 12940
rect 14921 12931 14979 12937
rect 15194 12928 15200 12940
rect 15252 12928 15258 12980
rect 15565 12971 15623 12977
rect 15565 12968 15577 12971
rect 15304 12940 15577 12968
rect 14826 12860 14832 12912
rect 14884 12900 14890 12912
rect 15304 12900 15332 12940
rect 15565 12937 15577 12940
rect 15611 12968 15623 12971
rect 19426 12968 19432 12980
rect 15611 12940 19432 12968
rect 15611 12937 15623 12940
rect 15565 12931 15623 12937
rect 17604 12909 17632 12940
rect 19426 12928 19432 12940
rect 19484 12928 19490 12980
rect 19731 12971 19789 12977
rect 19731 12937 19743 12971
rect 19777 12968 19789 12971
rect 20070 12968 20076 12980
rect 19777 12940 20076 12968
rect 19777 12937 19789 12940
rect 19731 12931 19789 12937
rect 20070 12928 20076 12940
rect 20128 12928 20134 12980
rect 20349 12971 20407 12977
rect 20349 12937 20361 12971
rect 20395 12968 20407 12971
rect 21174 12968 21180 12980
rect 20395 12940 21180 12968
rect 20395 12937 20407 12940
rect 20349 12931 20407 12937
rect 21174 12928 21180 12940
rect 21232 12928 21238 12980
rect 21637 12971 21695 12977
rect 21637 12937 21649 12971
rect 21683 12968 21695 12971
rect 21726 12968 21732 12980
rect 21683 12940 21732 12968
rect 21683 12937 21695 12940
rect 21637 12931 21695 12937
rect 21726 12928 21732 12940
rect 21784 12928 21790 12980
rect 22005 12971 22063 12977
rect 22005 12937 22017 12971
rect 22051 12937 22063 12971
rect 22005 12931 22063 12937
rect 17589 12903 17647 12909
rect 14884 12872 15332 12900
rect 15396 12872 16988 12900
rect 14884 12860 14890 12872
rect 15286 12832 15292 12844
rect 14752 12804 15292 12832
rect 13173 12795 13231 12801
rect 15286 12792 15292 12804
rect 15344 12792 15350 12844
rect 15396 12764 15424 12872
rect 15473 12835 15531 12841
rect 15473 12801 15485 12835
rect 15519 12832 15531 12835
rect 15838 12832 15844 12844
rect 15519 12804 15844 12832
rect 15519 12801 15531 12804
rect 15473 12795 15531 12801
rect 15838 12792 15844 12804
rect 15896 12792 15902 12844
rect 16850 12792 16856 12844
rect 16908 12792 16914 12844
rect 16960 12832 16988 12872
rect 17589 12869 17601 12903
rect 17635 12869 17647 12903
rect 17589 12863 17647 12869
rect 19518 12860 19524 12912
rect 19576 12860 19582 12912
rect 18414 12832 18420 12844
rect 16960 12804 18420 12832
rect 18414 12792 18420 12804
rect 18472 12792 18478 12844
rect 15657 12767 15715 12773
rect 15657 12764 15669 12767
rect 12360 12736 15424 12764
rect 15488 12736 15669 12764
rect 15488 12696 15516 12736
rect 15657 12733 15669 12736
rect 15703 12733 15715 12767
rect 19536 12764 19564 12860
rect 20088 12832 20116 12928
rect 22020 12900 22048 12931
rect 22738 12928 22744 12980
rect 22796 12968 22802 12980
rect 22796 12940 24808 12968
rect 22796 12928 22802 12940
rect 23106 12900 23112 12912
rect 22020 12872 23112 12900
rect 23106 12860 23112 12872
rect 23164 12900 23170 12912
rect 24394 12900 24400 12912
rect 23164 12872 24400 12900
rect 23164 12860 23170 12872
rect 24394 12860 24400 12872
rect 24452 12860 24458 12912
rect 20533 12835 20591 12841
rect 20533 12832 20545 12835
rect 20088 12804 20545 12832
rect 20533 12801 20545 12804
rect 20579 12801 20591 12835
rect 20533 12795 20591 12801
rect 21082 12792 21088 12844
rect 21140 12841 21146 12844
rect 21140 12835 21165 12841
rect 21153 12832 21165 12835
rect 21153 12804 21404 12832
rect 21153 12801 21165 12804
rect 21140 12795 21165 12801
rect 21140 12792 21146 12795
rect 20165 12767 20223 12773
rect 20165 12764 20177 12767
rect 19536 12736 20177 12764
rect 15657 12727 15715 12733
rect 20165 12733 20177 12736
rect 20211 12733 20223 12767
rect 21376 12764 21404 12804
rect 21450 12792 21456 12844
rect 21508 12792 21514 12844
rect 21821 12835 21879 12841
rect 21821 12801 21833 12835
rect 21867 12832 21879 12835
rect 22094 12832 22100 12844
rect 21867 12804 22100 12832
rect 21867 12801 21879 12804
rect 21821 12795 21879 12801
rect 21836 12764 21864 12795
rect 22094 12792 22100 12804
rect 22152 12792 22158 12844
rect 22462 12832 22468 12844
rect 22296 12804 22468 12832
rect 22296 12773 22324 12804
rect 22462 12792 22468 12804
rect 22520 12832 22526 12844
rect 22520 12804 23796 12832
rect 22520 12792 22526 12804
rect 21376 12736 21864 12764
rect 22281 12767 22339 12773
rect 20165 12727 20223 12733
rect 22281 12733 22293 12767
rect 22327 12733 22339 12767
rect 22281 12727 22339 12733
rect 22373 12767 22431 12773
rect 22373 12733 22385 12767
rect 22419 12764 22431 12767
rect 23198 12764 23204 12776
rect 22419 12736 23204 12764
rect 22419 12733 22431 12736
rect 22373 12727 22431 12733
rect 10091 12668 10732 12696
rect 14660 12668 15516 12696
rect 19889 12699 19947 12705
rect 10091 12665 10103 12668
rect 10045 12659 10103 12665
rect 14660 12640 14688 12668
rect 19889 12665 19901 12699
rect 19935 12696 19947 12699
rect 20254 12696 20260 12708
rect 19935 12668 20260 12696
rect 19935 12665 19947 12668
rect 19889 12659 19947 12665
rect 20254 12656 20260 12668
rect 20312 12656 20318 12708
rect 3050 12588 3056 12640
rect 3108 12628 3114 12640
rect 3605 12631 3663 12637
rect 3605 12628 3617 12631
rect 3108 12600 3617 12628
rect 3108 12588 3114 12600
rect 3605 12597 3617 12600
rect 3651 12597 3663 12631
rect 3605 12591 3663 12597
rect 10134 12588 10140 12640
rect 10192 12588 10198 12640
rect 14642 12588 14648 12640
rect 14700 12588 14706 12640
rect 15102 12588 15108 12640
rect 15160 12588 15166 12640
rect 19610 12588 19616 12640
rect 19668 12628 19674 12640
rect 19705 12631 19763 12637
rect 19705 12628 19717 12631
rect 19668 12600 19717 12628
rect 19668 12588 19674 12600
rect 19705 12597 19717 12600
rect 19751 12597 19763 12631
rect 19705 12591 19763 12597
rect 19978 12588 19984 12640
rect 20036 12588 20042 12640
rect 21358 12588 21364 12640
rect 21416 12628 21422 12640
rect 21453 12631 21511 12637
rect 21453 12628 21465 12631
rect 21416 12600 21465 12628
rect 21416 12588 21422 12600
rect 21453 12597 21465 12600
rect 21499 12628 21511 12631
rect 22388 12628 22416 12727
rect 23198 12724 23204 12736
rect 23256 12724 23262 12776
rect 23768 12640 23796 12804
rect 24302 12792 24308 12844
rect 24360 12832 24366 12844
rect 24673 12835 24731 12841
rect 24673 12832 24685 12835
rect 24360 12804 24685 12832
rect 24360 12792 24366 12804
rect 24673 12801 24685 12804
rect 24719 12801 24731 12835
rect 24780 12832 24808 12940
rect 25866 12928 25872 12980
rect 25924 12968 25930 12980
rect 26237 12971 26295 12977
rect 26237 12968 26249 12971
rect 25924 12940 26249 12968
rect 25924 12928 25930 12940
rect 26237 12937 26249 12940
rect 26283 12937 26295 12971
rect 26694 12968 26700 12980
rect 26237 12931 26295 12937
rect 26528 12940 26700 12968
rect 26142 12860 26148 12912
rect 26200 12900 26206 12912
rect 26200 12872 26464 12900
rect 26200 12860 26206 12872
rect 24949 12835 25007 12841
rect 24949 12832 24961 12835
rect 24780 12804 24961 12832
rect 24673 12795 24731 12801
rect 24949 12801 24961 12804
rect 24995 12801 25007 12835
rect 24949 12795 25007 12801
rect 25041 12835 25099 12841
rect 25041 12801 25053 12835
rect 25087 12832 25099 12835
rect 25590 12832 25596 12844
rect 25087 12804 25596 12832
rect 25087 12801 25099 12804
rect 25041 12795 25099 12801
rect 24394 12724 24400 12776
rect 24452 12724 24458 12776
rect 24486 12724 24492 12776
rect 24544 12724 24550 12776
rect 24581 12767 24639 12773
rect 24581 12733 24593 12767
rect 24627 12764 24639 12767
rect 24854 12764 24860 12776
rect 24627 12736 24860 12764
rect 24627 12733 24639 12736
rect 24581 12727 24639 12733
rect 21499 12600 22416 12628
rect 21499 12597 21511 12600
rect 21453 12591 21511 12597
rect 23750 12588 23756 12640
rect 23808 12628 23814 12640
rect 24688 12628 24716 12736
rect 24854 12724 24860 12736
rect 24912 12724 24918 12776
rect 24762 12656 24768 12708
rect 24820 12656 24826 12708
rect 24964 12696 24992 12795
rect 25590 12792 25596 12804
rect 25648 12792 25654 12844
rect 26326 12792 26332 12844
rect 26384 12792 26390 12844
rect 26436 12841 26464 12872
rect 26528 12841 26556 12940
rect 26694 12928 26700 12940
rect 26752 12928 26758 12980
rect 26970 12928 26976 12980
rect 27028 12928 27034 12980
rect 29638 12928 29644 12980
rect 29696 12928 29702 12980
rect 31202 12928 31208 12980
rect 31260 12928 31266 12980
rect 31846 12928 31852 12980
rect 31904 12928 31910 12980
rect 32858 12928 32864 12980
rect 32916 12928 32922 12980
rect 33134 12928 33140 12980
rect 33192 12928 33198 12980
rect 26421 12835 26479 12841
rect 26421 12801 26433 12835
rect 26467 12801 26479 12835
rect 26421 12795 26479 12801
rect 26513 12835 26571 12841
rect 26513 12801 26525 12835
rect 26559 12801 26571 12835
rect 26513 12795 26571 12801
rect 26697 12835 26755 12841
rect 26697 12801 26709 12835
rect 26743 12801 26755 12835
rect 26697 12795 26755 12801
rect 26789 12835 26847 12841
rect 26789 12801 26801 12835
rect 26835 12832 26847 12835
rect 26988 12832 27016 12928
rect 26835 12804 27016 12832
rect 29089 12835 29147 12841
rect 26835 12801 26847 12804
rect 26789 12795 26847 12801
rect 29089 12801 29101 12835
rect 29135 12832 29147 12835
rect 29656 12832 29684 12928
rect 31220 12900 31248 12928
rect 31481 12903 31539 12909
rect 31481 12900 31493 12903
rect 31220 12872 31493 12900
rect 31481 12869 31493 12872
rect 31527 12869 31539 12903
rect 31481 12863 31539 12869
rect 31697 12903 31755 12909
rect 31697 12869 31709 12903
rect 31743 12900 31755 12903
rect 32493 12903 32551 12909
rect 32493 12900 32505 12903
rect 31743 12872 32505 12900
rect 31743 12869 31755 12872
rect 31697 12863 31755 12869
rect 32493 12869 32505 12872
rect 32539 12869 32551 12903
rect 32493 12863 32551 12869
rect 29135 12804 29684 12832
rect 29135 12801 29147 12804
rect 29089 12795 29147 12801
rect 25222 12724 25228 12776
rect 25280 12724 25286 12776
rect 26344 12764 26372 12792
rect 26712 12764 26740 12795
rect 30374 12792 30380 12844
rect 30432 12832 30438 12844
rect 30653 12835 30711 12841
rect 30653 12832 30665 12835
rect 30432 12804 30665 12832
rect 30432 12792 30438 12804
rect 30653 12801 30665 12804
rect 30699 12801 30711 12835
rect 30653 12795 30711 12801
rect 31205 12835 31263 12841
rect 31205 12801 31217 12835
rect 31251 12832 31263 12835
rect 31294 12832 31300 12844
rect 31251 12804 31300 12832
rect 31251 12801 31263 12804
rect 31205 12795 31263 12801
rect 26344 12736 26740 12764
rect 28442 12724 28448 12776
rect 28500 12764 28506 12776
rect 29365 12767 29423 12773
rect 29365 12764 29377 12767
rect 28500 12736 29377 12764
rect 28500 12724 28506 12736
rect 29365 12733 29377 12736
rect 29411 12764 29423 12767
rect 29411 12736 30144 12764
rect 29411 12733 29423 12736
rect 29365 12727 29423 12733
rect 24964 12668 26192 12696
rect 23808 12600 24716 12628
rect 24780 12628 24808 12656
rect 24857 12631 24915 12637
rect 24857 12628 24869 12631
rect 24780 12600 24869 12628
rect 23808 12588 23814 12600
rect 24857 12597 24869 12600
rect 24903 12597 24915 12631
rect 24857 12591 24915 12597
rect 25130 12588 25136 12640
rect 25188 12588 25194 12640
rect 26164 12628 26192 12668
rect 26234 12656 26240 12708
rect 26292 12696 26298 12708
rect 28994 12696 29000 12708
rect 26292 12668 29000 12696
rect 26292 12656 26298 12668
rect 28994 12656 29000 12668
rect 29052 12656 29058 12708
rect 29086 12656 29092 12708
rect 29144 12696 29150 12708
rect 29181 12699 29239 12705
rect 29181 12696 29193 12699
rect 29144 12668 29193 12696
rect 29144 12656 29150 12668
rect 29181 12665 29193 12668
rect 29227 12696 29239 12699
rect 29914 12696 29920 12708
rect 29227 12668 29920 12696
rect 29227 12665 29239 12668
rect 29181 12659 29239 12665
rect 29914 12656 29920 12668
rect 29972 12656 29978 12708
rect 26878 12628 26884 12640
rect 26164 12600 26884 12628
rect 26878 12588 26884 12600
rect 26936 12628 26942 12640
rect 27154 12628 27160 12640
rect 26936 12600 27160 12628
rect 26936 12588 26942 12600
rect 27154 12588 27160 12600
rect 27212 12588 27218 12640
rect 29273 12631 29331 12637
rect 29273 12597 29285 12631
rect 29319 12628 29331 12631
rect 30006 12628 30012 12640
rect 29319 12600 30012 12628
rect 29319 12597 29331 12600
rect 29273 12591 29331 12597
rect 30006 12588 30012 12600
rect 30064 12588 30070 12640
rect 30116 12628 30144 12736
rect 30282 12724 30288 12776
rect 30340 12764 30346 12776
rect 30561 12767 30619 12773
rect 30561 12764 30573 12767
rect 30340 12736 30573 12764
rect 30340 12724 30346 12736
rect 30561 12733 30573 12736
rect 30607 12733 30619 12767
rect 30561 12727 30619 12733
rect 31220 12764 31248 12795
rect 31294 12792 31300 12804
rect 31352 12792 31358 12844
rect 31386 12792 31392 12844
rect 31444 12832 31450 12844
rect 32125 12835 32183 12841
rect 32125 12832 32137 12835
rect 31444 12804 32137 12832
rect 31444 12792 31450 12804
rect 32125 12801 32137 12804
rect 32171 12801 32183 12835
rect 32125 12795 32183 12801
rect 32309 12835 32367 12841
rect 32309 12801 32321 12835
rect 32355 12832 32367 12835
rect 32398 12832 32404 12844
rect 32355 12804 32404 12832
rect 32355 12801 32367 12804
rect 32309 12795 32367 12801
rect 32324 12764 32352 12795
rect 32398 12792 32404 12804
rect 32456 12792 32462 12844
rect 33152 12841 33180 12928
rect 33137 12835 33195 12841
rect 33137 12801 33149 12835
rect 33183 12801 33195 12835
rect 33137 12795 33195 12801
rect 33870 12792 33876 12844
rect 33928 12792 33934 12844
rect 31220 12736 32352 12764
rect 31021 12699 31079 12705
rect 31021 12665 31033 12699
rect 31067 12696 31079 12699
rect 31220 12696 31248 12736
rect 32490 12724 32496 12776
rect 32548 12764 32554 12776
rect 32861 12767 32919 12773
rect 32861 12764 32873 12767
rect 32548 12736 32873 12764
rect 32548 12724 32554 12736
rect 32861 12733 32873 12736
rect 32907 12733 32919 12767
rect 32861 12727 32919 12733
rect 33045 12767 33103 12773
rect 33045 12733 33057 12767
rect 33091 12764 33103 12767
rect 33318 12764 33324 12776
rect 33091 12736 33324 12764
rect 33091 12733 33103 12736
rect 33045 12727 33103 12733
rect 33318 12724 33324 12736
rect 33376 12764 33382 12776
rect 33888 12764 33916 12792
rect 33376 12736 33916 12764
rect 33376 12724 33382 12736
rect 31067 12668 31248 12696
rect 31067 12665 31079 12668
rect 31021 12659 31079 12665
rect 31665 12631 31723 12637
rect 31665 12628 31677 12631
rect 30116 12600 31677 12628
rect 31665 12597 31677 12600
rect 31711 12597 31723 12631
rect 31665 12591 31723 12597
rect 1104 12538 38272 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 38272 12538
rect 1104 12464 38272 12486
rect 1670 12384 1676 12436
rect 1728 12424 1734 12436
rect 1949 12427 2007 12433
rect 1949 12424 1961 12427
rect 1728 12396 1961 12424
rect 1728 12384 1734 12396
rect 1949 12393 1961 12396
rect 1995 12393 2007 12427
rect 1949 12387 2007 12393
rect 3786 12384 3792 12436
rect 3844 12384 3850 12436
rect 3973 12427 4031 12433
rect 3973 12393 3985 12427
rect 4019 12424 4031 12427
rect 4062 12424 4068 12436
rect 4019 12396 4068 12424
rect 4019 12393 4031 12396
rect 3973 12387 4031 12393
rect 3988 12356 4016 12387
rect 4062 12384 4068 12396
rect 4120 12384 4126 12436
rect 4249 12427 4307 12433
rect 4249 12393 4261 12427
rect 4295 12424 4307 12427
rect 4614 12424 4620 12436
rect 4295 12396 4620 12424
rect 4295 12393 4307 12396
rect 4249 12387 4307 12393
rect 4614 12384 4620 12396
rect 4672 12384 4678 12436
rect 5810 12384 5816 12436
rect 5868 12424 5874 12436
rect 6457 12427 6515 12433
rect 6457 12424 6469 12427
rect 5868 12396 6469 12424
rect 5868 12384 5874 12396
rect 6457 12393 6469 12396
rect 6503 12393 6515 12427
rect 6457 12387 6515 12393
rect 8573 12427 8631 12433
rect 8573 12393 8585 12427
rect 8619 12424 8631 12427
rect 8846 12424 8852 12436
rect 8619 12396 8852 12424
rect 8619 12393 8631 12396
rect 8573 12387 8631 12393
rect 8846 12384 8852 12396
rect 8904 12424 8910 12436
rect 10226 12424 10232 12436
rect 8904 12396 10232 12424
rect 8904 12384 8910 12396
rect 10226 12384 10232 12396
rect 10284 12384 10290 12436
rect 11146 12384 11152 12436
rect 11204 12424 11210 12436
rect 11517 12427 11575 12433
rect 11517 12424 11529 12427
rect 11204 12396 11529 12424
rect 11204 12384 11210 12396
rect 11517 12393 11529 12396
rect 11563 12393 11575 12427
rect 11517 12387 11575 12393
rect 11624 12396 16436 12424
rect 11624 12356 11652 12396
rect 16408 12356 16436 12396
rect 16850 12384 16856 12436
rect 16908 12384 16914 12436
rect 21729 12427 21787 12433
rect 21729 12393 21741 12427
rect 21775 12424 21787 12427
rect 21910 12424 21916 12436
rect 21775 12396 21916 12424
rect 21775 12393 21787 12396
rect 21729 12387 21787 12393
rect 21910 12384 21916 12396
rect 21968 12384 21974 12436
rect 24210 12424 24216 12436
rect 23216 12396 23612 12424
rect 17589 12359 17647 12365
rect 17589 12356 17601 12359
rect 2976 12328 4016 12356
rect 2976 12229 3004 12328
rect 3050 12248 3056 12300
rect 3108 12248 3114 12300
rect 3234 12248 3240 12300
rect 3292 12248 3298 12300
rect 2133 12223 2191 12229
rect 2133 12189 2145 12223
rect 2179 12220 2191 12223
rect 2961 12223 3019 12229
rect 2179 12192 2636 12220
rect 2179 12189 2191 12192
rect 2133 12183 2191 12189
rect 2608 12093 2636 12192
rect 2961 12189 2973 12223
rect 3007 12189 3019 12223
rect 3988 12220 4016 12328
rect 4080 12328 11652 12356
rect 11716 12328 14136 12356
rect 16408 12328 17601 12356
rect 4080 12300 4108 12328
rect 4062 12248 4068 12300
rect 4120 12248 4126 12300
rect 6270 12248 6276 12300
rect 6328 12288 6334 12300
rect 6917 12291 6975 12297
rect 6917 12288 6929 12291
rect 6328 12260 6929 12288
rect 6328 12248 6334 12260
rect 6917 12257 6929 12260
rect 6963 12257 6975 12291
rect 6917 12251 6975 12257
rect 7098 12248 7104 12300
rect 7156 12248 7162 12300
rect 9769 12291 9827 12297
rect 9769 12288 9781 12291
rect 8128 12260 9781 12288
rect 4249 12223 4307 12229
rect 4249 12220 4261 12223
rect 3988 12192 4261 12220
rect 2961 12183 3019 12189
rect 4249 12189 4261 12192
rect 4295 12189 4307 12223
rect 4249 12183 4307 12189
rect 4525 12223 4583 12229
rect 4525 12189 4537 12223
rect 4571 12189 4583 12223
rect 4525 12183 4583 12189
rect 6825 12223 6883 12229
rect 6825 12189 6837 12223
rect 6871 12220 6883 12223
rect 8018 12220 8024 12232
rect 6871 12192 8024 12220
rect 6871 12189 6883 12192
rect 6825 12183 6883 12189
rect 3142 12112 3148 12164
rect 3200 12152 3206 12164
rect 4157 12155 4215 12161
rect 4157 12152 4169 12155
rect 3200 12124 4169 12152
rect 3200 12112 3206 12124
rect 4157 12121 4169 12124
rect 4203 12152 4215 12155
rect 4433 12155 4491 12161
rect 4433 12152 4445 12155
rect 4203 12124 4445 12152
rect 4203 12121 4215 12124
rect 4157 12115 4215 12121
rect 4433 12121 4445 12124
rect 4479 12121 4491 12155
rect 4433 12115 4491 12121
rect 2593 12087 2651 12093
rect 2593 12053 2605 12087
rect 2639 12053 2651 12087
rect 2593 12047 2651 12053
rect 3418 12044 3424 12096
rect 3476 12084 3482 12096
rect 3947 12087 4005 12093
rect 3947 12084 3959 12087
rect 3476 12056 3959 12084
rect 3476 12044 3482 12056
rect 3947 12053 3959 12056
rect 3993 12084 4005 12087
rect 4540 12084 4568 12183
rect 8018 12180 8024 12192
rect 8076 12220 8082 12232
rect 8128 12220 8156 12260
rect 9769 12257 9781 12260
rect 9815 12288 9827 12291
rect 11716 12288 11744 12328
rect 9815 12260 11744 12288
rect 12161 12291 12219 12297
rect 9815 12257 9827 12260
rect 9769 12251 9827 12257
rect 12161 12257 12173 12291
rect 12207 12288 12219 12291
rect 12526 12288 12532 12300
rect 12207 12260 12532 12288
rect 12207 12257 12219 12260
rect 12161 12251 12219 12257
rect 12526 12248 12532 12260
rect 12584 12248 12590 12300
rect 14108 12288 14136 12328
rect 17589 12325 17601 12328
rect 17635 12325 17647 12359
rect 17589 12319 17647 12325
rect 18064 12328 20852 12356
rect 15746 12288 15752 12300
rect 14108 12260 15752 12288
rect 15746 12248 15752 12260
rect 15804 12248 15810 12300
rect 18064 12297 18092 12328
rect 20824 12300 20852 12328
rect 22830 12316 22836 12368
rect 22888 12356 22894 12368
rect 23216 12356 23244 12396
rect 22888 12328 23244 12356
rect 23308 12328 23536 12356
rect 22888 12316 22894 12328
rect 18049 12291 18107 12297
rect 18049 12257 18061 12291
rect 18095 12257 18107 12291
rect 18049 12251 18107 12257
rect 18233 12291 18291 12297
rect 18233 12257 18245 12291
rect 18279 12257 18291 12291
rect 18233 12251 18291 12257
rect 8076 12192 8156 12220
rect 8205 12223 8263 12229
rect 8076 12180 8082 12192
rect 8205 12189 8217 12223
rect 8251 12220 8263 12223
rect 8294 12220 8300 12232
rect 8251 12192 8300 12220
rect 8251 12189 8263 12192
rect 8205 12183 8263 12189
rect 8294 12180 8300 12192
rect 8352 12180 8358 12232
rect 8389 12223 8447 12229
rect 8389 12189 8401 12223
rect 8435 12220 8447 12223
rect 8754 12220 8760 12232
rect 8435 12192 8760 12220
rect 8435 12189 8447 12192
rect 8389 12183 8447 12189
rect 8754 12180 8760 12192
rect 8812 12180 8818 12232
rect 9398 12180 9404 12232
rect 9456 12180 9462 12232
rect 9953 12223 10011 12229
rect 9953 12189 9965 12223
rect 9999 12220 10011 12223
rect 10042 12220 10048 12232
rect 9999 12192 10048 12220
rect 9999 12189 10011 12192
rect 9953 12183 10011 12189
rect 10042 12180 10048 12192
rect 10100 12180 10106 12232
rect 10137 12223 10195 12229
rect 10137 12189 10149 12223
rect 10183 12220 10195 12223
rect 10226 12220 10232 12232
rect 10183 12192 10232 12220
rect 10183 12189 10195 12192
rect 10137 12183 10195 12189
rect 10226 12180 10232 12192
rect 10284 12180 10290 12232
rect 11977 12223 12035 12229
rect 11977 12189 11989 12223
rect 12023 12220 12035 12223
rect 12250 12220 12256 12232
rect 12023 12192 12256 12220
rect 12023 12189 12035 12192
rect 11977 12183 12035 12189
rect 12250 12180 12256 12192
rect 12308 12180 12314 12232
rect 14737 12223 14795 12229
rect 14737 12189 14749 12223
rect 14783 12220 14795 12223
rect 14826 12220 14832 12232
rect 14783 12192 14832 12220
rect 14783 12189 14795 12192
rect 14737 12183 14795 12189
rect 14826 12180 14832 12192
rect 14884 12180 14890 12232
rect 15102 12180 15108 12232
rect 15160 12180 15166 12232
rect 16482 12180 16488 12232
rect 16540 12180 16546 12232
rect 8665 12155 8723 12161
rect 8665 12121 8677 12155
rect 8711 12152 8723 12155
rect 9416 12152 9444 12180
rect 11885 12155 11943 12161
rect 11885 12152 11897 12155
rect 8711 12124 11897 12152
rect 8711 12121 8723 12124
rect 8665 12115 8723 12121
rect 11885 12121 11897 12124
rect 11931 12121 11943 12155
rect 15381 12155 15439 12161
rect 15381 12152 15393 12155
rect 11885 12115 11943 12121
rect 14936 12124 15393 12152
rect 3993 12056 4568 12084
rect 3993 12053 4005 12056
rect 3947 12047 4005 12053
rect 7834 12044 7840 12096
rect 7892 12084 7898 12096
rect 14936 12093 14964 12124
rect 15381 12121 15393 12124
rect 15427 12121 15439 12155
rect 15381 12115 15439 12121
rect 8021 12087 8079 12093
rect 8021 12084 8033 12087
rect 7892 12056 8033 12084
rect 7892 12044 7898 12056
rect 8021 12053 8033 12056
rect 8067 12053 8079 12087
rect 8021 12047 8079 12053
rect 14921 12087 14979 12093
rect 14921 12053 14933 12087
rect 14967 12053 14979 12087
rect 14921 12047 14979 12053
rect 15286 12044 15292 12096
rect 15344 12084 15350 12096
rect 16500 12084 16528 12180
rect 17678 12112 17684 12164
rect 17736 12152 17742 12164
rect 18248 12152 18276 12251
rect 18414 12248 18420 12300
rect 18472 12248 18478 12300
rect 18874 12288 18880 12300
rect 18708 12260 18880 12288
rect 18322 12180 18328 12232
rect 18380 12220 18386 12232
rect 18601 12223 18659 12229
rect 18601 12220 18613 12223
rect 18380 12192 18613 12220
rect 18380 12180 18386 12192
rect 18601 12189 18613 12192
rect 18647 12189 18659 12223
rect 18601 12183 18659 12189
rect 18708 12152 18736 12260
rect 18874 12248 18880 12260
rect 18932 12248 18938 12300
rect 20806 12248 20812 12300
rect 20864 12248 20870 12300
rect 20898 12248 20904 12300
rect 20956 12288 20962 12300
rect 21542 12288 21548 12300
rect 20956 12260 21548 12288
rect 20956 12248 20962 12260
rect 21542 12248 21548 12260
rect 21600 12248 21606 12300
rect 18782 12180 18788 12232
rect 18840 12220 18846 12232
rect 18969 12223 19027 12229
rect 18969 12220 18981 12223
rect 18840 12192 18981 12220
rect 18840 12180 18846 12192
rect 18969 12189 18981 12192
rect 19015 12189 19027 12223
rect 18969 12183 19027 12189
rect 19334 12180 19340 12232
rect 19392 12180 19398 12232
rect 21450 12180 21456 12232
rect 21508 12220 21514 12232
rect 22848 12220 22876 12316
rect 23014 12248 23020 12300
rect 23072 12248 23078 12300
rect 23124 12297 23152 12328
rect 23109 12291 23167 12297
rect 23109 12257 23121 12291
rect 23155 12257 23167 12291
rect 23109 12251 23167 12257
rect 23198 12248 23204 12300
rect 23256 12248 23262 12300
rect 21508 12192 22876 12220
rect 22925 12223 22983 12229
rect 21508 12180 21514 12192
rect 17736 12124 18736 12152
rect 18877 12155 18935 12161
rect 17736 12112 17742 12124
rect 18877 12121 18889 12155
rect 18923 12152 18935 12155
rect 20070 12152 20076 12164
rect 18923 12124 20076 12152
rect 18923 12121 18935 12124
rect 18877 12115 18935 12121
rect 20070 12112 20076 12124
rect 20128 12112 20134 12164
rect 21560 12161 21588 12192
rect 22925 12189 22937 12223
rect 22971 12189 22983 12223
rect 23032 12220 23060 12248
rect 23308 12220 23336 12328
rect 23385 12291 23443 12297
rect 23385 12257 23397 12291
rect 23431 12257 23443 12291
rect 23385 12251 23443 12257
rect 23032 12192 23336 12220
rect 22925 12183 22983 12189
rect 21545 12155 21603 12161
rect 21545 12121 21557 12155
rect 21591 12121 21603 12155
rect 21545 12115 21603 12121
rect 21761 12155 21819 12161
rect 21761 12121 21773 12155
rect 21807 12152 21819 12155
rect 22094 12152 22100 12164
rect 21807 12124 22100 12152
rect 21807 12121 21819 12124
rect 21761 12115 21819 12121
rect 22094 12112 22100 12124
rect 22152 12112 22158 12164
rect 15344 12056 16528 12084
rect 15344 12044 15350 12056
rect 17586 12044 17592 12096
rect 17644 12084 17650 12096
rect 17957 12087 18015 12093
rect 17957 12084 17969 12087
rect 17644 12056 17969 12084
rect 17644 12044 17650 12056
rect 17957 12053 17969 12056
rect 18003 12053 18015 12087
rect 17957 12047 18015 12053
rect 19518 12044 19524 12096
rect 19576 12044 19582 12096
rect 21913 12087 21971 12093
rect 21913 12053 21925 12087
rect 21959 12084 21971 12087
rect 22186 12084 22192 12096
rect 21959 12056 22192 12084
rect 21959 12053 21971 12056
rect 21913 12047 21971 12053
rect 22186 12044 22192 12056
rect 22244 12044 22250 12096
rect 22940 12084 22968 12183
rect 23400 12152 23428 12251
rect 23508 12229 23536 12328
rect 23584 12229 23612 12396
rect 23952 12396 24216 12424
rect 23753 12291 23811 12297
rect 23753 12257 23765 12291
rect 23799 12288 23811 12291
rect 23952 12288 23980 12396
rect 24210 12384 24216 12396
rect 24268 12384 24274 12436
rect 24394 12384 24400 12436
rect 24452 12424 24458 12436
rect 25130 12424 25136 12436
rect 24452 12396 25136 12424
rect 24452 12384 24458 12396
rect 25130 12384 25136 12396
rect 25188 12384 25194 12436
rect 25222 12384 25228 12436
rect 25280 12384 25286 12436
rect 26786 12384 26792 12436
rect 26844 12424 26850 12436
rect 26881 12427 26939 12433
rect 26881 12424 26893 12427
rect 26844 12396 26893 12424
rect 26844 12384 26850 12396
rect 26881 12393 26893 12396
rect 26927 12393 26939 12427
rect 26881 12387 26939 12393
rect 29549 12427 29607 12433
rect 29549 12393 29561 12427
rect 29595 12424 29607 12427
rect 29730 12424 29736 12436
rect 29595 12396 29736 12424
rect 29595 12393 29607 12396
rect 29549 12387 29607 12393
rect 29730 12384 29736 12396
rect 29788 12384 29794 12436
rect 30193 12427 30251 12433
rect 30193 12393 30205 12427
rect 30239 12424 30251 12427
rect 31754 12424 31760 12436
rect 30239 12396 31760 12424
rect 30239 12393 30251 12396
rect 30193 12387 30251 12393
rect 31754 12384 31760 12396
rect 31812 12424 31818 12436
rect 32766 12424 32772 12436
rect 31812 12396 32772 12424
rect 31812 12384 31818 12396
rect 32766 12384 32772 12396
rect 32824 12384 32830 12436
rect 26510 12316 26516 12368
rect 26568 12356 26574 12368
rect 27798 12356 27804 12368
rect 26568 12328 27804 12356
rect 26568 12316 26574 12328
rect 27798 12316 27804 12328
rect 27856 12356 27862 12368
rect 32674 12356 32680 12368
rect 27856 12328 32680 12356
rect 27856 12316 27862 12328
rect 32674 12316 32680 12328
rect 32732 12316 32738 12368
rect 23799 12260 23980 12288
rect 23799 12257 23811 12260
rect 23753 12251 23811 12257
rect 24762 12248 24768 12300
rect 24820 12288 24826 12300
rect 25777 12291 25835 12297
rect 25777 12288 25789 12291
rect 24820 12260 25789 12288
rect 24820 12248 24826 12260
rect 25777 12257 25789 12260
rect 25823 12257 25835 12291
rect 25777 12251 25835 12257
rect 26142 12248 26148 12300
rect 26200 12288 26206 12300
rect 26237 12291 26295 12297
rect 26237 12288 26249 12291
rect 26200 12260 26249 12288
rect 26200 12248 26206 12260
rect 26237 12257 26249 12260
rect 26283 12257 26295 12291
rect 26237 12251 26295 12257
rect 28902 12248 28908 12300
rect 28960 12288 28966 12300
rect 28960 12260 30420 12288
rect 28960 12248 28966 12260
rect 23477 12223 23536 12229
rect 23477 12189 23489 12223
rect 23523 12192 23536 12223
rect 23569 12223 23627 12229
rect 23523 12189 23535 12192
rect 23477 12183 23535 12189
rect 23569 12189 23581 12223
rect 23615 12220 23627 12223
rect 25038 12220 25044 12232
rect 23615 12192 25044 12220
rect 23615 12189 23627 12192
rect 23569 12183 23627 12189
rect 25038 12180 25044 12192
rect 25096 12180 25102 12232
rect 25593 12223 25651 12229
rect 25593 12189 25605 12223
rect 25639 12220 25651 12223
rect 26418 12220 26424 12232
rect 25639 12192 26424 12220
rect 25639 12189 25651 12192
rect 25593 12183 25651 12189
rect 26418 12180 26424 12192
rect 26476 12180 26482 12232
rect 26786 12180 26792 12232
rect 26844 12220 26850 12232
rect 29825 12223 29883 12229
rect 29825 12220 29837 12223
rect 26844 12192 29837 12220
rect 26844 12180 26850 12192
rect 29825 12189 29837 12192
rect 29871 12189 29883 12223
rect 29825 12183 29883 12189
rect 30006 12180 30012 12232
rect 30064 12180 30070 12232
rect 30282 12180 30288 12232
rect 30340 12180 30346 12232
rect 30392 12229 30420 12260
rect 32306 12248 32312 12300
rect 32364 12288 32370 12300
rect 32364 12260 33548 12288
rect 32364 12248 32370 12260
rect 30377 12223 30435 12229
rect 30377 12189 30389 12223
rect 30423 12189 30435 12223
rect 30377 12183 30435 12189
rect 30561 12223 30619 12229
rect 30561 12189 30573 12223
rect 30607 12189 30619 12223
rect 30561 12183 30619 12189
rect 29917 12155 29975 12161
rect 29917 12152 29929 12155
rect 23400 12124 29929 12152
rect 29917 12121 29929 12124
rect 29963 12121 29975 12155
rect 29917 12115 29975 12121
rect 23753 12087 23811 12093
rect 23753 12084 23765 12087
rect 22940 12056 23765 12084
rect 23753 12053 23765 12056
rect 23799 12053 23811 12087
rect 23753 12047 23811 12053
rect 25685 12087 25743 12093
rect 25685 12053 25697 12087
rect 25731 12084 25743 12087
rect 26050 12084 26056 12096
rect 25731 12056 26056 12084
rect 25731 12053 25743 12056
rect 25685 12047 25743 12053
rect 26050 12044 26056 12056
rect 26108 12084 26114 12096
rect 26513 12087 26571 12093
rect 26513 12084 26525 12087
rect 26108 12056 26525 12084
rect 26108 12044 26114 12056
rect 26513 12053 26525 12056
rect 26559 12053 26571 12087
rect 26513 12047 26571 12053
rect 26602 12044 26608 12096
rect 26660 12084 26666 12096
rect 28166 12084 28172 12096
rect 26660 12056 28172 12084
rect 26660 12044 26666 12056
rect 28166 12044 28172 12056
rect 28224 12044 28230 12096
rect 28902 12044 28908 12096
rect 28960 12084 28966 12096
rect 30300 12084 30328 12180
rect 30576 12152 30604 12183
rect 32030 12180 32036 12232
rect 32088 12220 32094 12232
rect 32950 12220 32956 12232
rect 32088 12192 32956 12220
rect 32088 12180 32094 12192
rect 32950 12180 32956 12192
rect 33008 12220 33014 12232
rect 33520 12229 33548 12260
rect 33137 12223 33195 12229
rect 33137 12220 33149 12223
rect 33008 12192 33149 12220
rect 33008 12180 33014 12192
rect 33137 12189 33149 12192
rect 33183 12189 33195 12223
rect 33137 12183 33195 12189
rect 33505 12223 33563 12229
rect 33505 12189 33517 12223
rect 33551 12220 33563 12223
rect 33594 12220 33600 12232
rect 33551 12192 33600 12220
rect 33551 12189 33563 12192
rect 33505 12183 33563 12189
rect 33594 12180 33600 12192
rect 33652 12180 33658 12232
rect 30392 12124 30604 12152
rect 30392 12096 30420 12124
rect 28960 12056 30328 12084
rect 28960 12044 28966 12056
rect 30374 12044 30380 12096
rect 30432 12044 30438 12096
rect 30466 12044 30472 12096
rect 30524 12044 30530 12096
rect 32582 12044 32588 12096
rect 32640 12084 32646 12096
rect 33137 12087 33195 12093
rect 33137 12084 33149 12087
rect 32640 12056 33149 12084
rect 32640 12044 32646 12056
rect 33137 12053 33149 12056
rect 33183 12053 33195 12087
rect 33137 12047 33195 12053
rect 1104 11994 38272 12016
rect 1104 11942 4874 11994
rect 4926 11942 4938 11994
rect 4990 11942 5002 11994
rect 5054 11942 5066 11994
rect 5118 11942 5130 11994
rect 5182 11942 35594 11994
rect 35646 11942 35658 11994
rect 35710 11942 35722 11994
rect 35774 11942 35786 11994
rect 35838 11942 35850 11994
rect 35902 11942 38272 11994
rect 1104 11920 38272 11942
rect 1581 11883 1639 11889
rect 1581 11849 1593 11883
rect 1627 11880 1639 11883
rect 8202 11880 8208 11892
rect 1627 11852 8208 11880
rect 1627 11849 1639 11852
rect 1581 11843 1639 11849
rect 8202 11840 8208 11852
rect 8260 11840 8266 11892
rect 8754 11840 8760 11892
rect 8812 11880 8818 11892
rect 9306 11880 9312 11892
rect 8812 11852 9312 11880
rect 8812 11840 8818 11852
rect 9306 11840 9312 11852
rect 9364 11840 9370 11892
rect 12161 11883 12219 11889
rect 12161 11849 12173 11883
rect 12207 11880 12219 11883
rect 13538 11880 13544 11892
rect 12207 11852 12434 11880
rect 12207 11849 12219 11852
rect 12161 11843 12219 11849
rect 11054 11812 11060 11824
rect 10704 11784 11060 11812
rect 934 11704 940 11756
rect 992 11744 998 11756
rect 1489 11747 1547 11753
rect 1489 11744 1501 11747
rect 992 11716 1501 11744
rect 992 11704 998 11716
rect 1489 11713 1501 11716
rect 1535 11713 1547 11747
rect 1489 11707 1547 11713
rect 9306 11704 9312 11756
rect 9364 11744 9370 11756
rect 10704 11753 10732 11784
rect 11054 11772 11060 11784
rect 11112 11772 11118 11824
rect 12406 11812 12434 11852
rect 12912 11852 13544 11880
rect 12529 11815 12587 11821
rect 12529 11812 12541 11815
rect 12406 11784 12541 11812
rect 12529 11781 12541 11784
rect 12575 11781 12587 11815
rect 12912 11812 12940 11852
rect 13538 11840 13544 11852
rect 13596 11880 13602 11892
rect 15286 11880 15292 11892
rect 13596 11852 15292 11880
rect 13596 11840 13602 11852
rect 15286 11840 15292 11852
rect 15344 11840 15350 11892
rect 20346 11880 20352 11892
rect 15396 11852 20352 11880
rect 12986 11812 12992 11824
rect 12912 11784 12992 11812
rect 12529 11775 12587 11781
rect 12986 11772 12992 11784
rect 13044 11772 13050 11824
rect 14458 11772 14464 11824
rect 14516 11812 14522 11824
rect 15396 11812 15424 11852
rect 20346 11840 20352 11852
rect 20404 11840 20410 11892
rect 24210 11840 24216 11892
rect 24268 11840 24274 11892
rect 24390 11883 24448 11889
rect 24390 11849 24402 11883
rect 24436 11880 24448 11883
rect 26786 11880 26792 11892
rect 24436 11852 26792 11880
rect 24436 11849 24448 11852
rect 24390 11843 24448 11849
rect 26786 11840 26792 11852
rect 26844 11840 26850 11892
rect 27614 11840 27620 11892
rect 27672 11840 27678 11892
rect 29086 11840 29092 11892
rect 29144 11880 29150 11892
rect 29273 11883 29331 11889
rect 29273 11880 29285 11883
rect 29144 11852 29285 11880
rect 29144 11840 29150 11852
rect 29273 11849 29285 11852
rect 29319 11849 29331 11883
rect 29273 11843 29331 11849
rect 29733 11883 29791 11889
rect 29733 11849 29745 11883
rect 29779 11849 29791 11883
rect 29733 11843 29791 11849
rect 14516 11784 15424 11812
rect 14516 11772 14522 11784
rect 15838 11772 15844 11824
rect 15896 11812 15902 11824
rect 19150 11812 19156 11824
rect 15896 11784 16160 11812
rect 15896 11772 15902 11784
rect 10689 11747 10747 11753
rect 10689 11744 10701 11747
rect 9364 11716 10701 11744
rect 9364 11704 9370 11716
rect 10689 11713 10701 11716
rect 10735 11713 10747 11747
rect 10689 11707 10747 11713
rect 10778 11704 10784 11756
rect 10836 11704 10842 11756
rect 11882 11704 11888 11756
rect 11940 11704 11946 11756
rect 11974 11704 11980 11756
rect 12032 11704 12038 11756
rect 14826 11704 14832 11756
rect 14884 11744 14890 11756
rect 15933 11747 15991 11753
rect 15933 11744 15945 11747
rect 14884 11716 15945 11744
rect 14884 11704 14890 11716
rect 15933 11713 15945 11716
rect 15979 11713 15991 11747
rect 15933 11707 15991 11713
rect 10318 11636 10324 11688
rect 10376 11676 10382 11688
rect 10870 11676 10876 11688
rect 10376 11648 10876 11676
rect 10376 11636 10382 11648
rect 10870 11636 10876 11648
rect 10928 11636 10934 11688
rect 11900 11676 11928 11704
rect 12250 11676 12256 11688
rect 11900 11648 12256 11676
rect 12250 11636 12256 11648
rect 12308 11636 12314 11688
rect 12894 11636 12900 11688
rect 12952 11676 12958 11688
rect 14277 11679 14335 11685
rect 14277 11676 14289 11679
rect 12952 11648 14289 11676
rect 12952 11636 12958 11648
rect 14277 11645 14289 11648
rect 14323 11676 14335 11679
rect 14734 11676 14740 11688
rect 14323 11648 14740 11676
rect 14323 11645 14335 11648
rect 14277 11639 14335 11645
rect 14734 11636 14740 11648
rect 14792 11636 14798 11688
rect 9490 11568 9496 11620
rect 9548 11608 9554 11620
rect 9548 11580 10456 11608
rect 9548 11568 9554 11580
rect 5442 11500 5448 11552
rect 5500 11540 5506 11552
rect 8294 11540 8300 11552
rect 5500 11512 8300 11540
rect 5500 11500 5506 11512
rect 8294 11500 8300 11512
rect 8352 11500 8358 11552
rect 10318 11500 10324 11552
rect 10376 11500 10382 11552
rect 10428 11540 10456 11580
rect 14844 11540 14872 11704
rect 16132 11685 16160 11784
rect 18800 11784 19156 11812
rect 18800 11753 18828 11784
rect 19150 11772 19156 11784
rect 19208 11772 19214 11824
rect 20254 11772 20260 11824
rect 20312 11772 20318 11824
rect 24228 11812 24256 11840
rect 23492 11784 24900 11812
rect 18601 11747 18659 11753
rect 18601 11744 18613 11747
rect 17604 11716 18613 11744
rect 16025 11679 16083 11685
rect 16025 11645 16037 11679
rect 16071 11645 16083 11679
rect 16025 11639 16083 11645
rect 16117 11679 16175 11685
rect 16117 11645 16129 11679
rect 16163 11645 16175 11679
rect 16117 11639 16175 11645
rect 16040 11608 16068 11639
rect 17604 11620 17632 11716
rect 18601 11713 18613 11716
rect 18647 11713 18659 11747
rect 18601 11707 18659 11713
rect 18785 11747 18843 11753
rect 18785 11713 18797 11747
rect 18831 11713 18843 11747
rect 20272 11744 20300 11772
rect 23492 11756 23520 11784
rect 23474 11744 23480 11756
rect 20272 11716 23480 11744
rect 18785 11707 18843 11713
rect 23474 11704 23480 11716
rect 23532 11704 23538 11756
rect 23750 11704 23756 11756
rect 23808 11704 23814 11756
rect 24210 11704 24216 11756
rect 24268 11704 24274 11756
rect 24305 11747 24363 11753
rect 24305 11713 24317 11747
rect 24351 11744 24363 11747
rect 24394 11744 24400 11756
rect 24351 11716 24400 11744
rect 24351 11713 24363 11716
rect 24305 11707 24363 11713
rect 24394 11704 24400 11716
rect 24452 11704 24458 11756
rect 24489 11747 24547 11753
rect 24489 11713 24501 11747
rect 24535 11713 24547 11747
rect 24489 11707 24547 11713
rect 23566 11676 23572 11688
rect 22066 11648 23572 11676
rect 17586 11608 17592 11620
rect 16040 11580 17592 11608
rect 17586 11568 17592 11580
rect 17644 11568 17650 11620
rect 18690 11568 18696 11620
rect 18748 11568 18754 11620
rect 10428 11512 14872 11540
rect 15562 11500 15568 11552
rect 15620 11500 15626 11552
rect 18138 11500 18144 11552
rect 18196 11540 18202 11552
rect 19242 11540 19248 11552
rect 18196 11512 19248 11540
rect 18196 11500 18202 11512
rect 19242 11500 19248 11512
rect 19300 11540 19306 11552
rect 22066 11540 22094 11648
rect 23566 11636 23572 11648
rect 23624 11636 23630 11688
rect 24504 11608 24532 11707
rect 24578 11704 24584 11756
rect 24636 11704 24642 11756
rect 24762 11704 24768 11756
rect 24820 11704 24826 11756
rect 24872 11753 24900 11784
rect 25314 11772 25320 11824
rect 25372 11812 25378 11824
rect 27632 11812 27660 11840
rect 25372 11784 27476 11812
rect 27632 11784 27736 11812
rect 25372 11772 25378 11784
rect 24857 11747 24915 11753
rect 24857 11713 24869 11747
rect 24903 11713 24915 11747
rect 24857 11707 24915 11713
rect 25038 11704 25044 11756
rect 25096 11744 25102 11756
rect 26602 11744 26608 11756
rect 25096 11716 26608 11744
rect 25096 11704 25102 11716
rect 26602 11704 26608 11716
rect 26660 11704 26666 11756
rect 26988 11688 27016 11784
rect 27157 11747 27215 11753
rect 27157 11713 27169 11747
rect 27203 11713 27215 11747
rect 27157 11707 27215 11713
rect 24949 11679 25007 11685
rect 24949 11645 24961 11679
rect 24995 11676 25007 11679
rect 26418 11676 26424 11688
rect 24995 11648 26424 11676
rect 24995 11645 25007 11648
rect 24949 11639 25007 11645
rect 26418 11636 26424 11648
rect 26476 11636 26482 11688
rect 26970 11636 26976 11688
rect 27028 11636 27034 11688
rect 27172 11676 27200 11707
rect 27338 11704 27344 11756
rect 27396 11704 27402 11756
rect 27448 11753 27476 11784
rect 27663 11781 27736 11784
rect 27433 11747 27491 11753
rect 27433 11713 27445 11747
rect 27479 11713 27491 11747
rect 27663 11747 27675 11781
rect 27709 11750 27736 11781
rect 27798 11772 27804 11824
rect 27856 11812 27862 11824
rect 27893 11815 27951 11821
rect 27893 11812 27905 11815
rect 27856 11784 27905 11812
rect 27856 11772 27862 11784
rect 27893 11781 27905 11784
rect 27939 11781 27951 11815
rect 27893 11775 27951 11781
rect 27982 11772 27988 11824
rect 28040 11812 28046 11824
rect 29748 11812 29776 11843
rect 30098 11840 30104 11892
rect 30156 11880 30162 11892
rect 30193 11883 30251 11889
rect 30193 11880 30205 11883
rect 30156 11852 30205 11880
rect 30156 11840 30162 11852
rect 30193 11849 30205 11852
rect 30239 11849 30251 11883
rect 30193 11843 30251 11849
rect 30466 11840 30472 11892
rect 30524 11840 30530 11892
rect 32401 11883 32459 11889
rect 32401 11849 32413 11883
rect 32447 11880 32459 11883
rect 33042 11880 33048 11892
rect 32447 11852 33048 11880
rect 32447 11849 32459 11852
rect 32401 11843 32459 11849
rect 33042 11840 33048 11852
rect 33100 11840 33106 11892
rect 30374 11812 30380 11824
rect 28040 11784 29684 11812
rect 29748 11784 30380 11812
rect 28040 11772 28046 11784
rect 27709 11747 27721 11750
rect 27663 11741 27721 11747
rect 27433 11707 27491 11713
rect 28810 11704 28816 11756
rect 28868 11704 28874 11756
rect 28994 11704 29000 11756
rect 29052 11744 29058 11756
rect 29457 11747 29515 11753
rect 29457 11744 29469 11747
rect 29052 11716 29469 11744
rect 29052 11704 29058 11716
rect 29457 11713 29469 11716
rect 29503 11713 29515 11747
rect 29457 11707 29515 11713
rect 28828 11676 28856 11704
rect 29549 11679 29607 11685
rect 29549 11676 29561 11679
rect 27172 11648 27568 11676
rect 28828 11648 29561 11676
rect 27540 11620 27568 11648
rect 29549 11645 29561 11648
rect 29595 11645 29607 11679
rect 29549 11639 29607 11645
rect 24581 11611 24639 11617
rect 24581 11608 24593 11611
rect 23400 11580 24593 11608
rect 23400 11552 23428 11580
rect 24581 11577 24593 11580
rect 24627 11577 24639 11611
rect 24581 11571 24639 11577
rect 27522 11568 27528 11620
rect 27580 11568 27586 11620
rect 29656 11608 29684 11784
rect 30374 11772 30380 11784
rect 30432 11772 30438 11824
rect 29730 11704 29736 11756
rect 29788 11744 29794 11756
rect 29917 11747 29975 11753
rect 29917 11744 29929 11747
rect 29788 11716 29929 11744
rect 29788 11704 29794 11716
rect 29917 11713 29929 11716
rect 29963 11713 29975 11747
rect 30484 11744 30512 11840
rect 30561 11747 30619 11753
rect 30561 11744 30573 11747
rect 30484 11716 30573 11744
rect 29917 11707 29975 11713
rect 30561 11713 30573 11716
rect 30607 11713 30619 11747
rect 30561 11707 30619 11713
rect 32582 11704 32588 11756
rect 32640 11704 32646 11756
rect 32674 11704 32680 11756
rect 32732 11704 32738 11756
rect 29822 11636 29828 11688
rect 29880 11636 29886 11688
rect 30650 11636 30656 11688
rect 30708 11636 30714 11688
rect 32214 11636 32220 11688
rect 32272 11676 32278 11688
rect 32692 11676 32720 11704
rect 32272 11648 32720 11676
rect 32272 11636 32278 11648
rect 34606 11608 34612 11620
rect 27632 11580 29132 11608
rect 29656 11580 34612 11608
rect 19300 11512 22094 11540
rect 19300 11500 19306 11512
rect 23382 11500 23388 11552
rect 23440 11500 23446 11552
rect 23569 11543 23627 11549
rect 23569 11509 23581 11543
rect 23615 11540 23627 11543
rect 26050 11540 26056 11552
rect 23615 11512 26056 11540
rect 23615 11509 23627 11512
rect 23569 11503 23627 11509
rect 26050 11500 26056 11512
rect 26108 11500 26114 11552
rect 26694 11500 26700 11552
rect 26752 11540 26758 11552
rect 26973 11543 27031 11549
rect 26973 11540 26985 11543
rect 26752 11512 26985 11540
rect 26752 11500 26758 11512
rect 26973 11509 26985 11512
rect 27019 11540 27031 11543
rect 27632 11540 27660 11580
rect 29104 11552 29132 11580
rect 34606 11568 34612 11580
rect 34664 11568 34670 11620
rect 27019 11512 27660 11540
rect 27019 11509 27031 11512
rect 26973 11503 27031 11509
rect 27706 11500 27712 11552
rect 27764 11500 27770 11552
rect 29086 11500 29092 11552
rect 29144 11500 29150 11552
rect 30374 11500 30380 11552
rect 30432 11540 30438 11552
rect 30837 11543 30895 11549
rect 30837 11540 30849 11543
rect 30432 11512 30849 11540
rect 30432 11500 30438 11512
rect 30837 11509 30849 11512
rect 30883 11509 30895 11543
rect 30837 11503 30895 11509
rect 1104 11450 38272 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 38272 11450
rect 1104 11376 38272 11398
rect 3142 11296 3148 11348
rect 3200 11296 3206 11348
rect 3418 11296 3424 11348
rect 3476 11336 3482 11348
rect 5718 11336 5724 11348
rect 3476 11308 5724 11336
rect 3476 11296 3482 11308
rect 5718 11296 5724 11308
rect 5776 11296 5782 11348
rect 7834 11296 7840 11348
rect 7892 11296 7898 11348
rect 8481 11339 8539 11345
rect 8481 11305 8493 11339
rect 8527 11336 8539 11339
rect 9030 11336 9036 11348
rect 8527 11308 9036 11336
rect 8527 11305 8539 11308
rect 8481 11299 8539 11305
rect 9030 11296 9036 11308
rect 9088 11296 9094 11348
rect 10318 11336 10324 11348
rect 9784 11308 10324 11336
rect 3878 11228 3884 11280
rect 3936 11268 3942 11280
rect 3936 11240 4384 11268
rect 3936 11228 3942 11240
rect 1397 11203 1455 11209
rect 1397 11169 1409 11203
rect 1443 11200 1455 11203
rect 4062 11200 4068 11212
rect 1443 11172 4068 11200
rect 1443 11169 1455 11172
rect 1397 11163 1455 11169
rect 4062 11160 4068 11172
rect 4120 11160 4126 11212
rect 4356 11209 4384 11240
rect 4341 11203 4399 11209
rect 4341 11169 4353 11203
rect 4387 11200 4399 11203
rect 5534 11200 5540 11212
rect 4387 11172 5540 11200
rect 4387 11169 4399 11172
rect 4341 11163 4399 11169
rect 5534 11160 5540 11172
rect 5592 11160 5598 11212
rect 7852 11200 7880 11296
rect 8021 11271 8079 11277
rect 8021 11237 8033 11271
rect 8067 11237 8079 11271
rect 8021 11231 8079 11237
rect 7668 11172 7880 11200
rect 5902 11092 5908 11144
rect 5960 11092 5966 11144
rect 6086 11092 6092 11144
rect 6144 11092 6150 11144
rect 7377 11135 7435 11141
rect 7377 11101 7389 11135
rect 7423 11101 7435 11135
rect 7377 11095 7435 11101
rect 1670 11024 1676 11076
rect 1728 11024 1734 11076
rect 2958 11064 2964 11076
rect 2898 11036 2964 11064
rect 2958 11024 2964 11036
rect 3016 11064 3022 11076
rect 3878 11064 3884 11076
rect 3016 11036 3884 11064
rect 3016 11024 3022 11036
rect 3878 11024 3884 11036
rect 3936 11024 3942 11076
rect 4157 11067 4215 11073
rect 4157 11033 4169 11067
rect 4203 11064 4215 11067
rect 5810 11064 5816 11076
rect 4203 11036 5816 11064
rect 4203 11033 4215 11036
rect 4157 11027 4215 11033
rect 5810 11024 5816 11036
rect 5868 11024 5874 11076
rect 7392 11064 7420 11095
rect 7466 11092 7472 11144
rect 7524 11092 7530 11144
rect 7668 11141 7696 11172
rect 7653 11135 7711 11141
rect 7653 11101 7665 11135
rect 7699 11101 7711 11135
rect 7653 11095 7711 11101
rect 7745 11135 7803 11141
rect 7745 11101 7757 11135
rect 7791 11132 7803 11135
rect 8036 11132 8064 11231
rect 9306 11228 9312 11280
rect 9364 11228 9370 11280
rect 9490 11228 9496 11280
rect 9548 11228 9554 11280
rect 8202 11160 8208 11212
rect 8260 11200 8266 11212
rect 8297 11203 8355 11209
rect 8297 11200 8309 11203
rect 8260 11172 8309 11200
rect 8260 11160 8266 11172
rect 8297 11169 8309 11172
rect 8343 11200 8355 11203
rect 8846 11200 8852 11212
rect 8343 11172 8852 11200
rect 8343 11169 8355 11172
rect 8297 11163 8355 11169
rect 8846 11160 8852 11172
rect 8904 11160 8910 11212
rect 9217 11203 9275 11209
rect 9217 11200 9229 11203
rect 8956 11172 9229 11200
rect 7791 11104 8064 11132
rect 7791 11101 7803 11104
rect 7745 11095 7803 11101
rect 8570 11092 8576 11144
rect 8628 11132 8634 11144
rect 8956 11132 8984 11172
rect 9217 11169 9229 11172
rect 9263 11200 9275 11203
rect 9508 11200 9536 11228
rect 9263 11172 9536 11200
rect 9263 11169 9275 11172
rect 9217 11163 9275 11169
rect 8628 11104 8984 11132
rect 8628 11092 8634 11104
rect 9030 11092 9036 11144
rect 9088 11132 9094 11144
rect 9125 11135 9183 11141
rect 9125 11132 9137 11135
rect 9088 11104 9137 11132
rect 9088 11092 9094 11104
rect 9125 11101 9137 11104
rect 9171 11101 9183 11135
rect 9125 11095 9183 11101
rect 9398 11092 9404 11144
rect 9456 11092 9462 11144
rect 9784 11141 9812 11308
rect 10318 11296 10324 11308
rect 10376 11296 10382 11348
rect 11974 11296 11980 11348
rect 12032 11336 12038 11348
rect 12437 11339 12495 11345
rect 12437 11336 12449 11339
rect 12032 11308 12449 11336
rect 12032 11296 12038 11308
rect 12437 11305 12449 11308
rect 12483 11305 12495 11339
rect 14458 11336 14464 11348
rect 12437 11299 12495 11305
rect 14016 11308 14464 11336
rect 9953 11271 10011 11277
rect 9953 11237 9965 11271
rect 9999 11268 10011 11271
rect 14016 11268 14044 11308
rect 14458 11296 14464 11308
rect 14516 11296 14522 11348
rect 16114 11336 16120 11348
rect 15672 11308 16120 11336
rect 9999 11240 10180 11268
rect 9999 11237 10011 11240
rect 9953 11231 10011 11237
rect 9858 11160 9864 11212
rect 9916 11200 9922 11212
rect 10045 11203 10103 11209
rect 10045 11200 10057 11203
rect 9916 11172 10057 11200
rect 9916 11160 9922 11172
rect 10045 11169 10057 11172
rect 10091 11169 10103 11203
rect 10152 11200 10180 11240
rect 12406 11240 14044 11268
rect 14093 11271 14151 11277
rect 10321 11203 10379 11209
rect 10321 11200 10333 11203
rect 10152 11172 10333 11200
rect 10045 11163 10103 11169
rect 10321 11169 10333 11172
rect 10367 11169 10379 11203
rect 10321 11163 10379 11169
rect 10778 11160 10784 11212
rect 10836 11200 10842 11212
rect 11793 11203 11851 11209
rect 11793 11200 11805 11203
rect 10836 11172 11805 11200
rect 10836 11160 10842 11172
rect 11793 11169 11805 11172
rect 11839 11200 11851 11203
rect 12406 11200 12434 11240
rect 14093 11237 14105 11271
rect 14139 11237 14151 11271
rect 14093 11231 14151 11237
rect 11839 11172 12434 11200
rect 11839 11169 11851 11172
rect 11793 11163 11851 11169
rect 12526 11160 12532 11212
rect 12584 11200 12590 11212
rect 12989 11203 13047 11209
rect 12989 11200 13001 11203
rect 12584 11172 13001 11200
rect 12584 11160 12590 11172
rect 12989 11169 13001 11172
rect 13035 11200 13047 11203
rect 13035 11172 13676 11200
rect 13035 11169 13047 11172
rect 12989 11163 13047 11169
rect 9769 11135 9827 11141
rect 9769 11101 9781 11135
rect 9815 11101 9827 11135
rect 11698 11132 11704 11144
rect 11454 11104 11704 11132
rect 9769 11095 9827 11101
rect 11698 11092 11704 11104
rect 11756 11092 11762 11144
rect 12434 11092 12440 11144
rect 12492 11132 12498 11144
rect 12805 11135 12863 11141
rect 12805 11132 12817 11135
rect 12492 11104 12817 11132
rect 12492 11092 12498 11104
rect 12805 11101 12817 11104
rect 12851 11132 12863 11135
rect 13354 11132 13360 11144
rect 12851 11104 13360 11132
rect 12851 11101 12863 11104
rect 12805 11095 12863 11101
rect 13354 11092 13360 11104
rect 13412 11092 13418 11144
rect 7392 11036 7604 11064
rect 7576 11008 7604 11036
rect 7834 11024 7840 11076
rect 7892 11064 7898 11076
rect 7929 11067 7987 11073
rect 7929 11064 7941 11067
rect 7892 11036 7941 11064
rect 7892 11024 7898 11036
rect 7929 11033 7941 11036
rect 7975 11033 7987 11067
rect 7929 11027 7987 11033
rect 8110 11024 8116 11076
rect 8168 11064 8174 11076
rect 8941 11067 8999 11073
rect 8941 11064 8953 11067
rect 8168 11036 8953 11064
rect 8168 11024 8174 11036
rect 8941 11033 8953 11036
rect 8987 11033 8999 11067
rect 8941 11027 8999 11033
rect 12894 11024 12900 11076
rect 12952 11024 12958 11076
rect 13648 11064 13676 11172
rect 13725 11135 13783 11141
rect 13725 11101 13737 11135
rect 13771 11132 13783 11135
rect 14108 11132 14136 11231
rect 14642 11200 14648 11212
rect 13771 11104 14136 11132
rect 14200 11172 14648 11200
rect 13771 11101 13783 11104
rect 13725 11095 13783 11101
rect 14200 11064 14228 11172
rect 14642 11160 14648 11172
rect 14700 11160 14706 11212
rect 14826 11160 14832 11212
rect 14884 11160 14890 11212
rect 14461 11135 14519 11141
rect 14461 11101 14473 11135
rect 14507 11132 14519 11135
rect 14844 11132 14872 11160
rect 14507 11104 14872 11132
rect 14507 11101 14519 11104
rect 14461 11095 14519 11101
rect 15562 11092 15568 11144
rect 15620 11092 15626 11144
rect 13648 11036 14228 11064
rect 14553 11067 14611 11073
rect 14553 11033 14565 11067
rect 14599 11064 14611 11067
rect 15672 11064 15700 11308
rect 16114 11296 16120 11308
rect 16172 11296 16178 11348
rect 17586 11296 17592 11348
rect 17644 11296 17650 11348
rect 22094 11296 22100 11348
rect 22152 11336 22158 11348
rect 23382 11336 23388 11348
rect 22152 11308 23388 11336
rect 22152 11296 22158 11308
rect 23382 11296 23388 11308
rect 23440 11296 23446 11348
rect 23474 11296 23480 11348
rect 23532 11296 23538 11348
rect 26510 11296 26516 11348
rect 26568 11296 26574 11348
rect 27338 11296 27344 11348
rect 27396 11296 27402 11348
rect 27614 11296 27620 11348
rect 27672 11296 27678 11348
rect 28905 11339 28963 11345
rect 28905 11305 28917 11339
rect 28951 11336 28963 11339
rect 29178 11336 29184 11348
rect 28951 11308 29184 11336
rect 28951 11305 28963 11308
rect 28905 11299 28963 11305
rect 29178 11296 29184 11308
rect 29236 11296 29242 11348
rect 29273 11339 29331 11345
rect 29273 11305 29285 11339
rect 29319 11336 29331 11339
rect 30098 11336 30104 11348
rect 29319 11308 30104 11336
rect 29319 11305 29331 11308
rect 29273 11299 29331 11305
rect 30098 11296 30104 11308
rect 30156 11296 30162 11348
rect 30374 11296 30380 11348
rect 30432 11296 30438 11348
rect 30466 11296 30472 11348
rect 30524 11296 30530 11348
rect 30650 11296 30656 11348
rect 30708 11336 30714 11348
rect 31389 11339 31447 11345
rect 31389 11336 31401 11339
rect 30708 11308 31401 11336
rect 30708 11296 30714 11308
rect 31389 11305 31401 11308
rect 31435 11305 31447 11339
rect 31389 11299 31447 11305
rect 32122 11296 32128 11348
rect 32180 11296 32186 11348
rect 34606 11296 34612 11348
rect 34664 11296 34670 11348
rect 15749 11271 15807 11277
rect 15749 11237 15761 11271
rect 15795 11268 15807 11271
rect 15795 11240 15976 11268
rect 15795 11237 15807 11240
rect 15749 11231 15807 11237
rect 15948 11200 15976 11240
rect 19242 11228 19248 11280
rect 19300 11268 19306 11280
rect 19300 11240 19472 11268
rect 19300 11228 19306 11240
rect 19444 11209 19472 11240
rect 19886 11228 19892 11280
rect 19944 11228 19950 11280
rect 21913 11271 21971 11277
rect 21913 11237 21925 11271
rect 21959 11268 21971 11271
rect 22278 11268 22284 11280
rect 21959 11240 22284 11268
rect 21959 11237 21971 11240
rect 21913 11231 21971 11237
rect 22278 11228 22284 11240
rect 22336 11228 22342 11280
rect 22462 11228 22468 11280
rect 22520 11228 22526 11280
rect 16117 11203 16175 11209
rect 16117 11200 16129 11203
rect 15948 11172 16129 11200
rect 16117 11169 16129 11172
rect 16163 11169 16175 11203
rect 16117 11163 16175 11169
rect 19429 11203 19487 11209
rect 19429 11169 19441 11203
rect 19475 11169 19487 11203
rect 19904 11200 19932 11228
rect 20530 11200 20536 11212
rect 19904 11172 20536 11200
rect 19429 11163 19487 11169
rect 15841 11135 15899 11141
rect 15841 11132 15853 11135
rect 14599 11036 15700 11064
rect 15764 11104 15853 11132
rect 14599 11033 14611 11036
rect 14553 11027 14611 11033
rect 15764 11008 15792 11104
rect 15841 11101 15853 11104
rect 15887 11101 15899 11135
rect 15841 11095 15899 11101
rect 18322 11092 18328 11144
rect 18380 11132 18386 11144
rect 18601 11135 18659 11141
rect 18601 11132 18613 11135
rect 18380 11104 18613 11132
rect 18380 11092 18386 11104
rect 18601 11101 18613 11104
rect 18647 11101 18659 11135
rect 18601 11095 18659 11101
rect 18785 11135 18843 11141
rect 18785 11101 18797 11135
rect 18831 11132 18843 11135
rect 19245 11135 19303 11141
rect 19245 11132 19257 11135
rect 18831 11104 19257 11132
rect 18831 11101 18843 11104
rect 18785 11095 18843 11101
rect 19245 11101 19257 11104
rect 19291 11101 19303 11135
rect 19245 11095 19303 11101
rect 19518 11092 19524 11144
rect 19576 11132 19582 11144
rect 19996 11141 20024 11172
rect 20530 11160 20536 11172
rect 20588 11160 20594 11212
rect 22480 11200 22508 11228
rect 21376 11172 22508 11200
rect 19889 11135 19947 11141
rect 19889 11132 19901 11135
rect 19576 11104 19901 11132
rect 19576 11092 19582 11104
rect 19889 11101 19901 11104
rect 19935 11101 19947 11135
rect 19889 11095 19947 11101
rect 19981 11135 20039 11141
rect 19981 11101 19993 11135
rect 20027 11101 20039 11135
rect 19981 11095 20039 11101
rect 18417 11067 18475 11073
rect 16500 11036 16606 11064
rect 16500 11008 16528 11036
rect 18417 11033 18429 11067
rect 18463 11064 18475 11067
rect 18506 11064 18512 11076
rect 18463 11036 18512 11064
rect 18463 11033 18475 11036
rect 18417 11027 18475 11033
rect 18506 11024 18512 11036
rect 18564 11024 18570 11076
rect 19904 11064 19932 11095
rect 20070 11092 20076 11144
rect 20128 11092 20134 11144
rect 21376 11141 21404 11172
rect 21361 11135 21419 11141
rect 21361 11101 21373 11135
rect 21407 11101 21419 11135
rect 21637 11135 21695 11141
rect 21637 11132 21649 11135
rect 21361 11095 21419 11101
rect 21468 11104 21649 11132
rect 20257 11067 20315 11073
rect 19904 11036 20208 11064
rect 20180 11008 20208 11036
rect 20257 11033 20269 11067
rect 20303 11064 20315 11067
rect 20990 11064 20996 11076
rect 20303 11036 20996 11064
rect 20303 11033 20315 11036
rect 20257 11027 20315 11033
rect 20990 11024 20996 11036
rect 21048 11064 21054 11076
rect 21468 11064 21496 11104
rect 21637 11101 21649 11104
rect 21683 11101 21695 11135
rect 21637 11095 21695 11101
rect 21729 11135 21787 11141
rect 21729 11101 21741 11135
rect 21775 11132 21787 11135
rect 22005 11135 22063 11141
rect 22005 11132 22017 11135
rect 21775 11104 22017 11132
rect 21775 11101 21787 11104
rect 21729 11095 21787 11101
rect 22005 11101 22017 11104
rect 22051 11101 22063 11135
rect 22005 11095 22063 11101
rect 22186 11092 22192 11144
rect 22244 11092 22250 11144
rect 22465 11135 22523 11141
rect 22465 11101 22477 11135
rect 22511 11132 22523 11135
rect 23382 11132 23388 11144
rect 22511 11104 23388 11132
rect 22511 11101 22523 11104
rect 22465 11095 22523 11101
rect 23382 11092 23388 11104
rect 23440 11092 23446 11144
rect 23492 11132 23520 11296
rect 23566 11228 23572 11280
rect 23624 11268 23630 11280
rect 24578 11268 24584 11280
rect 23624 11240 24584 11268
rect 23624 11228 23630 11240
rect 24578 11228 24584 11240
rect 24636 11228 24642 11280
rect 26528 11268 26556 11296
rect 26252 11240 26556 11268
rect 23753 11203 23811 11209
rect 23753 11169 23765 11203
rect 23799 11200 23811 11203
rect 25038 11200 25044 11212
rect 23799 11172 25044 11200
rect 23799 11169 23811 11172
rect 23753 11163 23811 11169
rect 25038 11160 25044 11172
rect 25096 11160 25102 11212
rect 26252 11209 26280 11240
rect 26237 11203 26295 11209
rect 26237 11169 26249 11203
rect 26283 11169 26295 11203
rect 27157 11203 27215 11209
rect 27157 11200 27169 11203
rect 26237 11163 26295 11169
rect 26528 11172 27169 11200
rect 26528 11144 26556 11172
rect 27157 11169 27169 11172
rect 27203 11169 27215 11203
rect 27157 11163 27215 11169
rect 23569 11135 23627 11141
rect 23569 11132 23581 11135
rect 23492 11104 23581 11132
rect 23569 11101 23581 11104
rect 23615 11101 23627 11135
rect 23569 11095 23627 11101
rect 24302 11092 24308 11144
rect 24360 11132 24366 11144
rect 25409 11135 25467 11141
rect 25409 11132 25421 11135
rect 24360 11104 25421 11132
rect 24360 11092 24366 11104
rect 25409 11101 25421 11104
rect 25455 11101 25467 11135
rect 25409 11095 25467 11101
rect 25593 11135 25651 11141
rect 25593 11101 25605 11135
rect 25639 11132 25651 11135
rect 26142 11132 26148 11144
rect 25639 11104 26148 11132
rect 25639 11101 25651 11104
rect 25593 11095 25651 11101
rect 26142 11092 26148 11104
rect 26200 11092 26206 11144
rect 26418 11092 26424 11144
rect 26476 11092 26482 11144
rect 26510 11092 26516 11144
rect 26568 11092 26574 11144
rect 26881 11135 26939 11141
rect 26881 11101 26893 11135
rect 26927 11101 26939 11135
rect 26881 11095 26939 11101
rect 21048 11036 21496 11064
rect 21545 11067 21603 11073
rect 21048 11024 21054 11036
rect 21545 11033 21557 11067
rect 21591 11033 21603 11067
rect 22094 11064 22100 11076
rect 21545 11027 21603 11033
rect 21744 11036 22100 11064
rect 3786 10956 3792 11008
rect 3844 10956 3850 11008
rect 4246 10956 4252 11008
rect 4304 10956 4310 11008
rect 7558 10956 7564 11008
rect 7616 10956 7622 11008
rect 13909 10999 13967 11005
rect 13909 10965 13921 10999
rect 13955 10996 13967 10999
rect 14090 10996 14096 11008
rect 13955 10968 14096 10996
rect 13955 10965 13967 10968
rect 13909 10959 13967 10965
rect 14090 10956 14096 10968
rect 14148 10956 14154 11008
rect 15102 10956 15108 11008
rect 15160 10996 15166 11008
rect 15746 10996 15752 11008
rect 15160 10968 15752 10996
rect 15160 10956 15166 10968
rect 15746 10956 15752 10968
rect 15804 10956 15810 11008
rect 16482 10956 16488 11008
rect 16540 10956 16546 11008
rect 20162 10956 20168 11008
rect 20220 10956 20226 11008
rect 21560 10996 21588 11027
rect 21744 10996 21772 11036
rect 22094 11024 22100 11036
rect 22152 11024 22158 11076
rect 22204 11064 22232 11092
rect 24210 11064 24216 11076
rect 22204 11036 24216 11064
rect 24210 11024 24216 11036
rect 24268 11024 24274 11076
rect 25501 11067 25559 11073
rect 25501 11033 25513 11067
rect 25547 11064 25559 11067
rect 26896 11064 26924 11095
rect 27062 11092 27068 11144
rect 27120 11092 27126 11144
rect 27249 11135 27307 11141
rect 27249 11101 27261 11135
rect 27295 11101 27307 11135
rect 27356 11132 27384 11296
rect 27632 11200 27660 11296
rect 27706 11228 27712 11280
rect 27764 11268 27770 11280
rect 30392 11268 30420 11296
rect 27764 11240 28488 11268
rect 27764 11228 27770 11240
rect 27632 11172 28212 11200
rect 27433 11135 27491 11141
rect 27433 11132 27445 11135
rect 27356 11104 27445 11132
rect 27249 11095 27307 11101
rect 27433 11101 27445 11104
rect 27479 11132 27491 11135
rect 27709 11135 27767 11141
rect 27709 11132 27721 11135
rect 27479 11104 27721 11132
rect 27479 11101 27491 11104
rect 27433 11095 27491 11101
rect 27709 11101 27721 11104
rect 27755 11101 27767 11135
rect 27709 11095 27767 11101
rect 25547 11036 26924 11064
rect 25547 11033 25559 11036
rect 25501 11027 25559 11033
rect 27154 11024 27160 11076
rect 27212 11064 27218 11076
rect 27264 11064 27292 11095
rect 27798 11092 27804 11144
rect 27856 11092 27862 11144
rect 27890 11092 27896 11144
rect 27948 11092 27954 11144
rect 28184 11141 28212 11172
rect 28460 11141 28488 11240
rect 30116 11240 30420 11268
rect 30116 11209 30144 11240
rect 30101 11203 30159 11209
rect 30101 11169 30113 11203
rect 30147 11169 30159 11203
rect 30101 11163 30159 11169
rect 30377 11203 30435 11209
rect 30377 11169 30389 11203
rect 30423 11200 30435 11203
rect 30484 11200 30512 11296
rect 30561 11271 30619 11277
rect 30561 11237 30573 11271
rect 30607 11268 30619 11271
rect 31754 11268 31760 11280
rect 30607 11240 31760 11268
rect 30607 11237 30619 11240
rect 30561 11231 30619 11237
rect 31754 11228 31760 11240
rect 31812 11228 31818 11280
rect 31864 11240 33088 11268
rect 31864 11200 31892 11240
rect 30423 11172 30512 11200
rect 31726 11172 31892 11200
rect 32324 11172 32904 11200
rect 30423 11169 30435 11172
rect 30377 11163 30435 11169
rect 28169 11135 28227 11141
rect 28169 11101 28181 11135
rect 28215 11132 28227 11135
rect 28261 11135 28319 11141
rect 28261 11132 28273 11135
rect 28215 11104 28273 11132
rect 28215 11101 28227 11104
rect 28169 11095 28227 11101
rect 28261 11101 28273 11104
rect 28307 11101 28319 11135
rect 28261 11095 28319 11101
rect 28445 11135 28503 11141
rect 28445 11101 28457 11135
rect 28491 11101 28503 11135
rect 28445 11095 28503 11101
rect 29086 11092 29092 11144
rect 29144 11092 29150 11144
rect 29365 11135 29423 11141
rect 29365 11101 29377 11135
rect 29411 11132 29423 11135
rect 30193 11135 30251 11141
rect 30193 11132 30205 11135
rect 29411 11104 30205 11132
rect 29411 11101 29423 11104
rect 29365 11095 29423 11101
rect 30193 11101 30205 11104
rect 30239 11101 30251 11135
rect 30193 11095 30251 11101
rect 27212 11036 27292 11064
rect 27816 11064 27844 11092
rect 28077 11067 28135 11073
rect 28077 11064 28089 11067
rect 27816 11036 28089 11064
rect 27212 11024 27218 11036
rect 28077 11033 28089 11036
rect 28123 11033 28135 11067
rect 28077 11027 28135 11033
rect 28353 11067 28411 11073
rect 28353 11033 28365 11067
rect 28399 11064 28411 11067
rect 30006 11064 30012 11076
rect 28399 11036 30012 11064
rect 28399 11033 28411 11036
rect 28353 11027 28411 11033
rect 30006 11024 30012 11036
rect 30064 11024 30070 11076
rect 30208 11064 30236 11095
rect 30282 11092 30288 11144
rect 30340 11092 30346 11144
rect 31573 11135 31631 11141
rect 31573 11101 31585 11135
rect 31619 11132 31631 11135
rect 31726 11132 31754 11172
rect 32324 11144 32352 11172
rect 31619 11104 31754 11132
rect 31619 11101 31631 11104
rect 31573 11095 31631 11101
rect 31846 11092 31852 11144
rect 31904 11092 31910 11144
rect 32033 11135 32091 11141
rect 32033 11101 32045 11135
rect 32079 11132 32091 11135
rect 32306 11132 32312 11144
rect 32079 11104 32312 11132
rect 32079 11101 32091 11104
rect 32033 11095 32091 11101
rect 32306 11092 32312 11104
rect 32364 11092 32370 11144
rect 32490 11092 32496 11144
rect 32548 11132 32554 11144
rect 32585 11135 32643 11141
rect 32585 11132 32597 11135
rect 32548 11104 32597 11132
rect 32548 11092 32554 11104
rect 32585 11101 32597 11104
rect 32631 11101 32643 11135
rect 32585 11095 32643 11101
rect 32766 11092 32772 11144
rect 32824 11092 32830 11144
rect 32876 11141 32904 11172
rect 33060 11144 33088 11240
rect 32861 11135 32919 11141
rect 32861 11101 32873 11135
rect 32907 11101 32919 11135
rect 32861 11095 32919 11101
rect 33042 11092 33048 11144
rect 33100 11092 33106 11144
rect 34624 11132 34652 11296
rect 37553 11135 37611 11141
rect 37553 11132 37565 11135
rect 34624 11104 37565 11132
rect 37553 11101 37565 11104
rect 37599 11101 37611 11135
rect 37553 11095 37611 11101
rect 30208 11036 30328 11064
rect 21560 10968 21772 10996
rect 21818 10956 21824 11008
rect 21876 10996 21882 11008
rect 22373 10999 22431 11005
rect 22373 10996 22385 10999
rect 21876 10968 22385 10996
rect 21876 10956 21882 10968
rect 22373 10965 22385 10968
rect 22419 10965 22431 10999
rect 22373 10959 22431 10965
rect 23382 10956 23388 11008
rect 23440 10956 23446 11008
rect 26050 10956 26056 11008
rect 26108 10996 26114 11008
rect 26329 10999 26387 11005
rect 26329 10996 26341 10999
rect 26108 10968 26341 10996
rect 26108 10956 26114 10968
rect 26329 10965 26341 10968
rect 26375 10965 26387 10999
rect 26329 10959 26387 10965
rect 26786 10956 26792 11008
rect 26844 10956 26850 11008
rect 27614 10956 27620 11008
rect 27672 10956 27678 11008
rect 30300 10996 30328 11036
rect 37918 11024 37924 11076
rect 37976 11024 37982 11076
rect 30650 10996 30656 11008
rect 30300 10968 30656 10996
rect 30650 10956 30656 10968
rect 30708 10956 30714 11008
rect 32858 10956 32864 11008
rect 32916 10996 32922 11008
rect 32953 10999 33011 11005
rect 32953 10996 32965 10999
rect 32916 10968 32965 10996
rect 32916 10956 32922 10968
rect 32953 10965 32965 10968
rect 32999 10965 33011 10999
rect 32953 10959 33011 10965
rect 1104 10906 38272 10928
rect 1104 10854 4874 10906
rect 4926 10854 4938 10906
rect 4990 10854 5002 10906
rect 5054 10854 5066 10906
rect 5118 10854 5130 10906
rect 5182 10854 35594 10906
rect 35646 10854 35658 10906
rect 35710 10854 35722 10906
rect 35774 10854 35786 10906
rect 35838 10854 35850 10906
rect 35902 10854 38272 10906
rect 1104 10832 38272 10854
rect 1670 10752 1676 10804
rect 1728 10792 1734 10804
rect 1765 10795 1823 10801
rect 1765 10792 1777 10795
rect 1728 10764 1777 10792
rect 1728 10752 1734 10764
rect 1765 10761 1777 10764
rect 1811 10761 1823 10795
rect 1765 10755 1823 10761
rect 2777 10795 2835 10801
rect 2777 10761 2789 10795
rect 2823 10792 2835 10795
rect 3786 10792 3792 10804
rect 2823 10764 3792 10792
rect 2823 10761 2835 10764
rect 2777 10755 2835 10761
rect 3786 10752 3792 10764
rect 3844 10752 3850 10804
rect 3878 10752 3884 10804
rect 3936 10792 3942 10804
rect 5813 10795 5871 10801
rect 3936 10764 4384 10792
rect 3936 10752 3942 10764
rect 4246 10724 4252 10736
rect 3712 10696 4252 10724
rect 1949 10659 2007 10665
rect 1949 10625 1961 10659
rect 1995 10656 2007 10659
rect 2685 10659 2743 10665
rect 1995 10628 2360 10656
rect 1995 10625 2007 10628
rect 1949 10619 2007 10625
rect 2332 10529 2360 10628
rect 2685 10625 2697 10659
rect 2731 10656 2743 10659
rect 3142 10656 3148 10668
rect 2731 10628 3148 10656
rect 2731 10625 2743 10628
rect 2685 10619 2743 10625
rect 3142 10616 3148 10628
rect 3200 10656 3206 10668
rect 3329 10659 3387 10665
rect 3329 10656 3341 10659
rect 3200 10628 3341 10656
rect 3200 10616 3206 10628
rect 3329 10625 3341 10628
rect 3375 10625 3387 10659
rect 3329 10619 3387 10625
rect 2961 10591 3019 10597
rect 2961 10557 2973 10591
rect 3007 10557 3019 10591
rect 2961 10551 3019 10557
rect 2317 10523 2375 10529
rect 2317 10489 2329 10523
rect 2363 10489 2375 10523
rect 2317 10483 2375 10489
rect 2976 10452 3004 10551
rect 3418 10548 3424 10600
rect 3476 10548 3482 10600
rect 3712 10597 3740 10696
rect 4246 10684 4252 10696
rect 4304 10684 4310 10736
rect 4356 10724 4384 10764
rect 5813 10761 5825 10795
rect 5859 10792 5871 10795
rect 6086 10792 6092 10804
rect 5859 10764 6092 10792
rect 5859 10761 5871 10764
rect 5813 10755 5871 10761
rect 6086 10752 6092 10764
rect 6144 10792 6150 10804
rect 8665 10795 8723 10801
rect 6144 10764 7420 10792
rect 6144 10752 6150 10764
rect 7392 10733 7420 10764
rect 8665 10761 8677 10795
rect 8711 10792 8723 10795
rect 8938 10792 8944 10804
rect 8711 10764 8944 10792
rect 8711 10761 8723 10764
rect 8665 10755 8723 10761
rect 8938 10752 8944 10764
rect 8996 10752 9002 10804
rect 9033 10795 9091 10801
rect 9033 10761 9045 10795
rect 9079 10792 9091 10795
rect 9398 10792 9404 10804
rect 9079 10764 9404 10792
rect 9079 10761 9091 10764
rect 9033 10755 9091 10761
rect 9398 10752 9404 10764
rect 9456 10752 9462 10804
rect 15102 10792 15108 10804
rect 10520 10764 12434 10792
rect 7377 10727 7435 10733
rect 4356 10696 4830 10724
rect 5644 10696 6960 10724
rect 5644 10656 5672 10696
rect 5552 10628 5672 10656
rect 5552 10600 5580 10628
rect 5718 10616 5724 10668
rect 5776 10656 5782 10668
rect 5997 10659 6055 10665
rect 5997 10656 6009 10659
rect 5776 10628 6009 10656
rect 5776 10616 5782 10628
rect 5997 10625 6009 10628
rect 6043 10625 6055 10659
rect 5997 10619 6055 10625
rect 6178 10616 6184 10668
rect 6236 10616 6242 10668
rect 6730 10616 6736 10668
rect 6788 10616 6794 10668
rect 3697 10591 3755 10597
rect 3697 10557 3709 10591
rect 3743 10557 3755 10591
rect 3697 10551 3755 10557
rect 4062 10548 4068 10600
rect 4120 10548 4126 10600
rect 4341 10591 4399 10597
rect 4341 10557 4353 10591
rect 4387 10588 4399 10591
rect 4706 10588 4712 10600
rect 4387 10560 4712 10588
rect 4387 10557 4399 10560
rect 4341 10551 4399 10557
rect 4706 10548 4712 10560
rect 4764 10548 4770 10600
rect 5534 10548 5540 10600
rect 5592 10548 5598 10600
rect 5810 10548 5816 10600
rect 5868 10548 5874 10600
rect 6932 10597 6960 10696
rect 7377 10693 7389 10727
rect 7423 10693 7435 10727
rect 7377 10687 7435 10693
rect 7561 10727 7619 10733
rect 7561 10693 7573 10727
rect 7607 10724 7619 10727
rect 10520 10724 10548 10764
rect 7607 10696 10548 10724
rect 12406 10724 12434 10764
rect 13924 10764 15108 10792
rect 13814 10724 13820 10736
rect 12406 10696 13820 10724
rect 7607 10693 7619 10696
rect 7561 10687 7619 10693
rect 13814 10684 13820 10696
rect 13872 10684 13878 10736
rect 7190 10616 7196 10668
rect 7248 10616 7254 10668
rect 8573 10659 8631 10665
rect 8573 10625 8585 10659
rect 8619 10625 8631 10659
rect 8573 10619 8631 10625
rect 6089 10591 6147 10597
rect 6089 10557 6101 10591
rect 6135 10588 6147 10591
rect 6825 10591 6883 10597
rect 6825 10588 6837 10591
rect 6135 10560 6837 10588
rect 6135 10557 6147 10560
rect 6089 10551 6147 10557
rect 6825 10557 6837 10560
rect 6871 10557 6883 10591
rect 6825 10551 6883 10557
rect 6917 10591 6975 10597
rect 6917 10557 6929 10591
rect 6963 10557 6975 10591
rect 8588 10588 8616 10619
rect 8846 10616 8852 10668
rect 8904 10616 8910 10668
rect 9585 10659 9643 10665
rect 9585 10625 9597 10659
rect 9631 10625 9643 10659
rect 9585 10619 9643 10625
rect 9125 10591 9183 10597
rect 9125 10588 9137 10591
rect 8588 10560 9137 10588
rect 6917 10551 6975 10557
rect 9125 10557 9137 10560
rect 9171 10557 9183 10591
rect 9600 10588 9628 10619
rect 10778 10616 10784 10668
rect 10836 10656 10842 10668
rect 10965 10659 11023 10665
rect 10965 10656 10977 10659
rect 10836 10628 10977 10656
rect 10836 10616 10842 10628
rect 10965 10625 10977 10628
rect 11011 10625 11023 10659
rect 10965 10619 11023 10625
rect 11514 10616 11520 10668
rect 11572 10656 11578 10668
rect 12250 10656 12256 10668
rect 11572 10628 12256 10656
rect 11572 10616 11578 10628
rect 12250 10616 12256 10628
rect 12308 10656 12314 10668
rect 13924 10665 13952 10764
rect 15102 10752 15108 10764
rect 15160 10752 15166 10804
rect 19150 10752 19156 10804
rect 19208 10752 19214 10804
rect 20714 10792 20720 10804
rect 19260 10764 20720 10792
rect 14090 10684 14096 10736
rect 14148 10724 14154 10736
rect 14185 10727 14243 10733
rect 14185 10724 14197 10727
rect 14148 10696 14197 10724
rect 14148 10684 14154 10696
rect 14185 10693 14197 10696
rect 14231 10693 14243 10727
rect 14185 10687 14243 10693
rect 15933 10727 15991 10733
rect 15933 10693 15945 10727
rect 15979 10724 15991 10727
rect 16114 10724 16120 10736
rect 15979 10696 16120 10724
rect 15979 10693 15991 10696
rect 15933 10687 15991 10693
rect 16114 10684 16120 10696
rect 16172 10684 16178 10736
rect 19260 10724 19288 10764
rect 20714 10752 20720 10764
rect 20772 10752 20778 10804
rect 20824 10764 22048 10792
rect 20824 10733 20852 10764
rect 22020 10736 22048 10764
rect 22370 10752 22376 10804
rect 22428 10792 22434 10804
rect 24121 10795 24179 10801
rect 24121 10792 24133 10795
rect 22428 10764 24133 10792
rect 22428 10752 22434 10764
rect 24121 10761 24133 10764
rect 24167 10761 24179 10795
rect 24121 10755 24179 10761
rect 27614 10752 27620 10804
rect 27672 10752 27678 10804
rect 28718 10752 28724 10804
rect 28776 10792 28782 10804
rect 32122 10792 32128 10804
rect 28776 10764 32128 10792
rect 28776 10752 28782 10764
rect 32122 10752 32128 10764
rect 32180 10752 32186 10804
rect 32217 10795 32275 10801
rect 32217 10761 32229 10795
rect 32263 10792 32275 10795
rect 32306 10792 32312 10804
rect 32263 10764 32312 10792
rect 32263 10761 32275 10764
rect 32217 10755 32275 10761
rect 32306 10752 32312 10764
rect 32364 10752 32370 10804
rect 32582 10792 32588 10804
rect 32508 10764 32588 10792
rect 20809 10727 20867 10733
rect 20809 10724 20821 10727
rect 16776 10696 19288 10724
rect 20272 10696 20821 10724
rect 13909 10659 13967 10665
rect 12308 10654 13860 10656
rect 13909 10654 13921 10659
rect 12308 10628 13921 10654
rect 12308 10616 12314 10628
rect 13832 10626 13921 10628
rect 13909 10625 13921 10626
rect 13955 10625 13967 10659
rect 13909 10619 13967 10625
rect 15286 10616 15292 10668
rect 15344 10616 15350 10668
rect 10226 10588 10232 10600
rect 9600 10560 10232 10588
rect 9125 10551 9183 10557
rect 10226 10548 10232 10560
rect 10284 10548 10290 10600
rect 11057 10591 11115 10597
rect 11057 10557 11069 10591
rect 11103 10557 11115 10591
rect 11057 10551 11115 10557
rect 5828 10520 5856 10548
rect 10597 10523 10655 10529
rect 10597 10520 10609 10523
rect 5828 10492 10609 10520
rect 10597 10489 10609 10492
rect 10643 10489 10655 10523
rect 11072 10520 11100 10551
rect 11238 10548 11244 10600
rect 11296 10548 11302 10600
rect 14016 10560 15240 10588
rect 14016 10520 14044 10560
rect 11072 10492 14044 10520
rect 15212 10520 15240 10560
rect 16776 10520 16804 10696
rect 16853 10659 16911 10665
rect 16853 10625 16865 10659
rect 16899 10656 16911 10659
rect 16942 10656 16948 10668
rect 16899 10628 16948 10656
rect 16899 10625 16911 10628
rect 16853 10619 16911 10625
rect 16942 10616 16948 10628
rect 17000 10616 17006 10668
rect 17037 10659 17095 10665
rect 17037 10625 17049 10659
rect 17083 10625 17095 10659
rect 17037 10619 17095 10625
rect 15212 10492 16804 10520
rect 10597 10483 10655 10489
rect 3234 10452 3240 10464
rect 2976 10424 3240 10452
rect 3234 10412 3240 10424
rect 3292 10452 3298 10464
rect 5810 10452 5816 10464
rect 3292 10424 5816 10452
rect 3292 10412 3298 10424
rect 5810 10412 5816 10424
rect 5868 10412 5874 10464
rect 6362 10412 6368 10464
rect 6420 10412 6426 10464
rect 7926 10412 7932 10464
rect 7984 10452 7990 10464
rect 8202 10452 8208 10464
rect 7984 10424 8208 10452
rect 7984 10412 7990 10424
rect 8202 10412 8208 10424
rect 8260 10412 8266 10464
rect 8294 10412 8300 10464
rect 8352 10452 8358 10464
rect 9309 10455 9367 10461
rect 9309 10452 9321 10455
rect 8352 10424 9321 10452
rect 8352 10412 8358 10424
rect 9309 10421 9321 10424
rect 9355 10421 9367 10455
rect 9309 10415 9367 10421
rect 13814 10412 13820 10464
rect 13872 10452 13878 10464
rect 17052 10452 17080 10619
rect 17126 10616 17132 10668
rect 17184 10616 17190 10668
rect 17221 10659 17279 10665
rect 17221 10625 17233 10659
rect 17267 10656 17279 10659
rect 18141 10659 18199 10665
rect 17267 10628 18092 10656
rect 17267 10625 17279 10628
rect 17221 10619 17279 10625
rect 17494 10480 17500 10532
rect 17552 10480 17558 10532
rect 18064 10520 18092 10628
rect 18141 10625 18153 10659
rect 18187 10656 18199 10659
rect 18322 10656 18328 10668
rect 18187 10628 18328 10656
rect 18187 10625 18199 10628
rect 18141 10619 18199 10625
rect 18322 10616 18328 10628
rect 18380 10616 18386 10668
rect 18506 10616 18512 10668
rect 18564 10656 18570 10668
rect 20272 10665 20300 10696
rect 20809 10693 20821 10696
rect 20855 10693 20867 10727
rect 20809 10687 20867 10693
rect 20990 10684 20996 10736
rect 21048 10733 21054 10736
rect 21048 10727 21067 10733
rect 21055 10724 21067 10727
rect 21055 10696 21496 10724
rect 21055 10693 21067 10696
rect 21048 10687 21067 10693
rect 21048 10684 21054 10687
rect 21468 10665 21496 10696
rect 22002 10684 22008 10736
rect 22060 10684 22066 10736
rect 22204 10696 22784 10724
rect 22204 10665 22232 10696
rect 22756 10668 22784 10696
rect 22830 10684 22836 10736
rect 22888 10724 22894 10736
rect 23017 10727 23075 10733
rect 23017 10724 23029 10727
rect 22888 10696 23029 10724
rect 22888 10684 22894 10696
rect 23017 10693 23029 10696
rect 23063 10693 23075 10727
rect 23017 10687 23075 10693
rect 23106 10684 23112 10736
rect 23164 10684 23170 10736
rect 23247 10727 23305 10733
rect 23247 10693 23259 10727
rect 23293 10724 23305 10727
rect 23382 10724 23388 10736
rect 23293 10696 23388 10724
rect 23293 10693 23305 10696
rect 23247 10687 23305 10693
rect 23382 10684 23388 10696
rect 23440 10684 23446 10736
rect 27632 10724 27660 10752
rect 27172 10696 27660 10724
rect 18969 10659 19027 10665
rect 18969 10656 18981 10659
rect 18564 10628 18981 10656
rect 18564 10616 18570 10628
rect 18969 10625 18981 10628
rect 19015 10625 19027 10659
rect 18969 10619 19027 10625
rect 20257 10659 20315 10665
rect 20257 10625 20269 10659
rect 20303 10625 20315 10659
rect 20257 10619 20315 10625
rect 21453 10659 21511 10665
rect 21453 10625 21465 10659
rect 21499 10625 21511 10659
rect 22088 10659 22146 10665
rect 22088 10656 22100 10659
rect 21453 10619 21511 10625
rect 21560 10628 22100 10656
rect 21174 10548 21180 10600
rect 21232 10588 21238 10600
rect 21269 10591 21327 10597
rect 21269 10588 21281 10591
rect 21232 10560 21281 10588
rect 21232 10548 21238 10560
rect 21269 10557 21281 10560
rect 21315 10588 21327 10591
rect 21560 10588 21588 10628
rect 22088 10625 22100 10628
rect 22134 10625 22146 10659
rect 22088 10619 22146 10625
rect 22189 10659 22247 10665
rect 22189 10625 22201 10659
rect 22235 10625 22247 10659
rect 22189 10619 22247 10625
rect 22373 10659 22431 10665
rect 22373 10625 22385 10659
rect 22419 10625 22431 10659
rect 22373 10619 22431 10625
rect 22465 10659 22523 10665
rect 22465 10625 22477 10659
rect 22511 10656 22600 10659
rect 22646 10656 22652 10668
rect 22511 10631 22652 10656
rect 22511 10625 22523 10631
rect 22572 10628 22652 10631
rect 22465 10619 22523 10625
rect 21315 10560 21588 10588
rect 21315 10557 21327 10560
rect 21269 10551 21327 10557
rect 21634 10548 21640 10600
rect 21692 10548 21698 10600
rect 22112 10588 22140 10619
rect 22388 10588 22416 10619
rect 22646 10616 22652 10628
rect 22704 10616 22710 10668
rect 22738 10616 22744 10668
rect 22796 10616 22802 10668
rect 22922 10616 22928 10668
rect 22980 10616 22986 10668
rect 24213 10659 24271 10665
rect 24213 10656 24225 10659
rect 23400 10628 24225 10656
rect 22112 10560 22324 10588
rect 22388 10560 22508 10588
rect 22186 10520 22192 10532
rect 18064 10492 22192 10520
rect 22186 10480 22192 10492
rect 22244 10480 22250 10532
rect 22296 10520 22324 10560
rect 22370 10520 22376 10532
rect 22296 10492 22376 10520
rect 22370 10480 22376 10492
rect 22428 10480 22434 10532
rect 13872 10424 17080 10452
rect 13872 10412 13878 10424
rect 18046 10412 18052 10464
rect 18104 10412 18110 10464
rect 20162 10412 20168 10464
rect 20220 10412 20226 10464
rect 20993 10455 21051 10461
rect 20993 10421 21005 10455
rect 21039 10452 21051 10455
rect 21082 10452 21088 10464
rect 21039 10424 21088 10452
rect 21039 10421 21051 10424
rect 20993 10415 21051 10421
rect 21082 10412 21088 10424
rect 21140 10412 21146 10464
rect 21177 10455 21235 10461
rect 21177 10421 21189 10455
rect 21223 10452 21235 10455
rect 21450 10452 21456 10464
rect 21223 10424 21456 10452
rect 21223 10421 21235 10424
rect 21177 10415 21235 10421
rect 21450 10412 21456 10424
rect 21508 10412 21514 10464
rect 21542 10412 21548 10464
rect 21600 10452 21606 10464
rect 21913 10455 21971 10461
rect 21913 10452 21925 10455
rect 21600 10424 21925 10452
rect 21600 10412 21606 10424
rect 21913 10421 21925 10424
rect 21959 10421 21971 10455
rect 21913 10415 21971 10421
rect 22002 10412 22008 10464
rect 22060 10452 22066 10464
rect 22480 10452 22508 10560
rect 22756 10520 22784 10616
rect 23106 10548 23112 10600
rect 23164 10588 23170 10600
rect 23400 10597 23428 10628
rect 24213 10625 24225 10628
rect 24259 10656 24271 10659
rect 24394 10656 24400 10668
rect 24259 10628 24400 10656
rect 24259 10625 24271 10628
rect 24213 10619 24271 10625
rect 24394 10616 24400 10628
rect 24452 10616 24458 10668
rect 26786 10616 26792 10668
rect 26844 10656 26850 10668
rect 27172 10665 27200 10696
rect 29086 10684 29092 10736
rect 29144 10724 29150 10736
rect 29144 10696 30512 10724
rect 29144 10684 29150 10696
rect 26973 10659 27031 10665
rect 26973 10656 26985 10659
rect 26844 10628 26985 10656
rect 26844 10616 26850 10628
rect 26973 10625 26985 10628
rect 27019 10625 27031 10659
rect 26973 10619 27031 10625
rect 27157 10659 27215 10665
rect 27157 10625 27169 10659
rect 27203 10625 27215 10659
rect 27157 10619 27215 10625
rect 27246 10616 27252 10668
rect 27304 10616 27310 10668
rect 27341 10659 27399 10665
rect 27341 10625 27353 10659
rect 27387 10656 27399 10659
rect 27522 10656 27528 10668
rect 27387 10628 27528 10656
rect 27387 10625 27399 10628
rect 27341 10619 27399 10625
rect 27522 10616 27528 10628
rect 27580 10616 27586 10668
rect 28166 10616 28172 10668
rect 28224 10616 28230 10668
rect 28258 10616 28264 10668
rect 28316 10656 28322 10668
rect 28353 10659 28411 10665
rect 28353 10656 28365 10659
rect 28316 10628 28365 10656
rect 28316 10616 28322 10628
rect 28353 10625 28365 10628
rect 28399 10656 28411 10659
rect 28721 10659 28779 10665
rect 28721 10656 28733 10659
rect 28399 10628 28733 10656
rect 28399 10625 28411 10628
rect 28353 10619 28411 10625
rect 28721 10625 28733 10628
rect 28767 10625 28779 10659
rect 28721 10619 28779 10625
rect 28905 10659 28963 10665
rect 28905 10625 28917 10659
rect 28951 10625 28963 10659
rect 28905 10619 28963 10625
rect 23385 10591 23443 10597
rect 23385 10588 23397 10591
rect 23164 10560 23397 10588
rect 23164 10548 23170 10560
rect 23385 10557 23397 10560
rect 23431 10557 23443 10591
rect 23385 10551 23443 10557
rect 23658 10548 23664 10600
rect 23716 10588 23722 10600
rect 23937 10591 23995 10597
rect 23937 10588 23949 10591
rect 23716 10560 23949 10588
rect 23716 10548 23722 10560
rect 23937 10557 23949 10560
rect 23983 10588 23995 10591
rect 24486 10588 24492 10600
rect 23983 10560 24492 10588
rect 23983 10557 23995 10560
rect 23937 10551 23995 10557
rect 24486 10548 24492 10560
rect 24544 10548 24550 10600
rect 28920 10588 28948 10619
rect 30190 10616 30196 10668
rect 30248 10656 30254 10668
rect 30484 10665 30512 10696
rect 31294 10684 31300 10736
rect 31352 10724 31358 10736
rect 32508 10724 32536 10764
rect 32582 10752 32588 10764
rect 32640 10752 32646 10804
rect 32674 10752 32680 10804
rect 32732 10792 32738 10804
rect 33689 10795 33747 10801
rect 33689 10792 33701 10795
rect 32732 10764 33701 10792
rect 32732 10752 32738 10764
rect 33689 10761 33701 10764
rect 33735 10761 33747 10795
rect 33689 10755 33747 10761
rect 35069 10795 35127 10801
rect 35069 10761 35081 10795
rect 35115 10792 35127 10795
rect 35342 10792 35348 10804
rect 35115 10764 35348 10792
rect 35115 10761 35127 10764
rect 35069 10755 35127 10761
rect 35342 10752 35348 10764
rect 35400 10752 35406 10804
rect 31352 10696 32536 10724
rect 31352 10684 31358 10696
rect 30285 10659 30343 10665
rect 30285 10656 30297 10659
rect 30248 10628 30297 10656
rect 30248 10616 30254 10628
rect 30285 10625 30297 10628
rect 30331 10625 30343 10659
rect 30285 10619 30343 10625
rect 30469 10659 30527 10665
rect 30469 10625 30481 10659
rect 30515 10656 30527 10659
rect 31846 10656 31852 10668
rect 30515 10628 31852 10656
rect 30515 10625 30527 10628
rect 30469 10619 30527 10625
rect 31846 10616 31852 10628
rect 31904 10616 31910 10668
rect 32125 10659 32183 10665
rect 32125 10625 32137 10659
rect 32171 10656 32183 10659
rect 32214 10656 32220 10668
rect 32171 10628 32220 10656
rect 32171 10625 32183 10628
rect 32125 10619 32183 10625
rect 32214 10616 32220 10628
rect 32272 10616 32278 10668
rect 32324 10665 32352 10696
rect 33226 10684 33232 10736
rect 33284 10724 33290 10736
rect 33594 10724 33600 10736
rect 33284 10696 33600 10724
rect 33284 10684 33290 10696
rect 33594 10684 33600 10696
rect 33652 10724 33658 10736
rect 33652 10696 33824 10724
rect 33652 10684 33658 10696
rect 32309 10659 32367 10665
rect 32309 10625 32321 10659
rect 32355 10625 32367 10659
rect 32309 10619 32367 10625
rect 32585 10659 32643 10665
rect 32585 10625 32597 10659
rect 32631 10656 32643 10659
rect 32766 10656 32772 10668
rect 32631 10628 32772 10656
rect 32631 10625 32643 10628
rect 32585 10619 32643 10625
rect 32766 10616 32772 10628
rect 32824 10616 32830 10668
rect 33502 10616 33508 10668
rect 33560 10616 33566 10668
rect 33796 10665 33824 10696
rect 33781 10659 33839 10665
rect 33781 10625 33793 10659
rect 33827 10625 33839 10659
rect 33781 10619 33839 10625
rect 34057 10659 34115 10665
rect 34057 10625 34069 10659
rect 34103 10625 34115 10659
rect 34057 10619 34115 10625
rect 28994 10588 29000 10600
rect 24596 10560 28856 10588
rect 28920 10560 29000 10588
rect 23566 10520 23572 10532
rect 22756 10492 23572 10520
rect 23566 10480 23572 10492
rect 23624 10480 23630 10532
rect 24596 10529 24624 10560
rect 24581 10523 24639 10529
rect 24581 10489 24593 10523
rect 24627 10489 24639 10523
rect 24581 10483 24639 10489
rect 26418 10480 26424 10532
rect 26476 10520 26482 10532
rect 28445 10523 28503 10529
rect 26476 10492 28396 10520
rect 26476 10480 26482 10492
rect 22060 10424 22508 10452
rect 22060 10412 22066 10424
rect 22738 10412 22744 10464
rect 22796 10412 22802 10464
rect 23474 10412 23480 10464
rect 23532 10452 23538 10464
rect 23842 10452 23848 10464
rect 23532 10424 23848 10452
rect 23532 10412 23538 10424
rect 23842 10412 23848 10424
rect 23900 10452 23906 10464
rect 26602 10452 26608 10464
rect 23900 10424 26608 10452
rect 23900 10412 23906 10424
rect 26602 10412 26608 10424
rect 26660 10412 26666 10464
rect 27614 10412 27620 10464
rect 27672 10412 27678 10464
rect 28368 10452 28396 10492
rect 28445 10489 28457 10523
rect 28491 10520 28503 10523
rect 28534 10520 28540 10532
rect 28491 10492 28540 10520
rect 28491 10489 28503 10492
rect 28445 10483 28503 10489
rect 28534 10480 28540 10492
rect 28592 10480 28598 10532
rect 28718 10480 28724 10532
rect 28776 10480 28782 10532
rect 28828 10520 28856 10560
rect 28994 10548 29000 10560
rect 29052 10548 29058 10600
rect 30377 10591 30435 10597
rect 30377 10557 30389 10591
rect 30423 10588 30435 10591
rect 32490 10588 32496 10600
rect 30423 10560 32496 10588
rect 30423 10557 30435 10560
rect 30377 10551 30435 10557
rect 32490 10548 32496 10560
rect 32548 10548 32554 10600
rect 33965 10591 34023 10597
rect 33965 10557 33977 10591
rect 34011 10557 34023 10591
rect 33965 10551 34023 10557
rect 33980 10520 34008 10551
rect 28828 10492 34008 10520
rect 28736 10452 28764 10480
rect 28368 10424 28764 10452
rect 30282 10412 30288 10464
rect 30340 10452 30346 10464
rect 32861 10455 32919 10461
rect 32861 10452 32873 10455
rect 30340 10424 32873 10452
rect 30340 10412 30346 10424
rect 32861 10421 32873 10424
rect 32907 10452 32919 10455
rect 32950 10452 32956 10464
rect 32907 10424 32956 10452
rect 32907 10421 32919 10424
rect 32861 10415 32919 10421
rect 32950 10412 32956 10424
rect 33008 10412 33014 10464
rect 33505 10455 33563 10461
rect 33505 10421 33517 10455
rect 33551 10452 33563 10455
rect 34072 10452 34100 10619
rect 34422 10616 34428 10668
rect 34480 10656 34486 10668
rect 34701 10659 34759 10665
rect 34701 10656 34713 10659
rect 34480 10628 34713 10656
rect 34480 10616 34486 10628
rect 34701 10625 34713 10628
rect 34747 10625 34759 10659
rect 34701 10619 34759 10625
rect 34609 10591 34667 10597
rect 34609 10557 34621 10591
rect 34655 10557 34667 10591
rect 34609 10551 34667 10557
rect 34425 10523 34483 10529
rect 34425 10489 34437 10523
rect 34471 10520 34483 10523
rect 34624 10520 34652 10551
rect 34471 10492 34652 10520
rect 34471 10489 34483 10492
rect 34425 10483 34483 10489
rect 33551 10424 34100 10452
rect 33551 10421 33563 10424
rect 33505 10415 33563 10421
rect 1104 10362 38272 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 38272 10362
rect 1104 10288 38272 10310
rect 4617 10251 4675 10257
rect 4617 10217 4629 10251
rect 4663 10248 4675 10251
rect 4706 10248 4712 10260
rect 4663 10220 4712 10248
rect 4663 10217 4675 10220
rect 4617 10211 4675 10217
rect 4706 10208 4712 10220
rect 4764 10208 4770 10260
rect 6178 10208 6184 10260
rect 6236 10208 6242 10260
rect 6362 10208 6368 10260
rect 6420 10208 6426 10260
rect 7558 10208 7564 10260
rect 7616 10248 7622 10260
rect 9950 10248 9956 10260
rect 7616 10220 9956 10248
rect 7616 10208 7622 10220
rect 9950 10208 9956 10220
rect 10008 10248 10014 10260
rect 10502 10248 10508 10260
rect 10008 10220 10508 10248
rect 10008 10208 10014 10220
rect 10502 10208 10508 10220
rect 10560 10208 10566 10260
rect 13078 10208 13084 10260
rect 13136 10208 13142 10260
rect 14458 10208 14464 10260
rect 14516 10248 14522 10260
rect 17126 10248 17132 10260
rect 14516 10220 17132 10248
rect 14516 10208 14522 10220
rect 17126 10208 17132 10220
rect 17184 10208 17190 10260
rect 20441 10251 20499 10257
rect 20441 10217 20453 10251
rect 20487 10248 20499 10251
rect 20901 10251 20959 10257
rect 20487 10220 20760 10248
rect 20487 10217 20499 10220
rect 20441 10211 20499 10217
rect 6380 10180 6408 10208
rect 5644 10152 6408 10180
rect 5644 10121 5672 10152
rect 7466 10140 7472 10192
rect 7524 10180 7530 10192
rect 8386 10180 8392 10192
rect 7524 10152 8392 10180
rect 7524 10140 7530 10152
rect 8386 10140 8392 10152
rect 8444 10140 8450 10192
rect 8481 10183 8539 10189
rect 8481 10149 8493 10183
rect 8527 10180 8539 10183
rect 8527 10152 9076 10180
rect 8527 10149 8539 10152
rect 8481 10143 8539 10149
rect 5629 10115 5687 10121
rect 5629 10081 5641 10115
rect 5675 10081 5687 10115
rect 5629 10075 5687 10081
rect 5810 10072 5816 10124
rect 5868 10072 5874 10124
rect 5902 10072 5908 10124
rect 5960 10112 5966 10124
rect 5960 10084 6224 10112
rect 5960 10072 5966 10084
rect 2961 10047 3019 10053
rect 2961 10013 2973 10047
rect 3007 10044 3019 10047
rect 3142 10044 3148 10056
rect 3007 10016 3148 10044
rect 3007 10013 3019 10016
rect 2961 10007 3019 10013
rect 3142 10004 3148 10016
rect 3200 10004 3206 10056
rect 4801 10047 4859 10053
rect 4801 10013 4813 10047
rect 4847 10044 4859 10047
rect 5537 10047 5595 10053
rect 4847 10016 5212 10044
rect 4847 10013 4859 10016
rect 4801 10007 4859 10013
rect 2777 9979 2835 9985
rect 2777 9945 2789 9979
rect 2823 9976 2835 9979
rect 3050 9976 3056 9988
rect 2823 9948 3056 9976
rect 2823 9945 2835 9948
rect 2777 9939 2835 9945
rect 3050 9936 3056 9948
rect 3108 9936 3114 9988
rect 3142 9868 3148 9920
rect 3200 9868 3206 9920
rect 5184 9917 5212 10016
rect 5537 10013 5549 10047
rect 5583 10044 5595 10047
rect 5997 10047 6055 10053
rect 5997 10044 6009 10047
rect 5583 10016 6009 10044
rect 5583 10013 5595 10016
rect 5537 10007 5595 10013
rect 5997 10013 6009 10016
rect 6043 10044 6055 10047
rect 6086 10044 6092 10056
rect 6043 10016 6092 10044
rect 6043 10013 6055 10016
rect 5997 10007 6055 10013
rect 6086 10004 6092 10016
rect 6144 10004 6150 10056
rect 6196 10053 6224 10084
rect 7484 10053 7512 10140
rect 7745 10115 7803 10121
rect 7745 10081 7757 10115
rect 7791 10112 7803 10115
rect 8202 10112 8208 10124
rect 7791 10084 8208 10112
rect 7791 10081 7803 10084
rect 7745 10075 7803 10081
rect 8202 10072 8208 10084
rect 8260 10072 8266 10124
rect 8662 10072 8668 10124
rect 8720 10072 8726 10124
rect 9048 10121 9076 10152
rect 9033 10115 9091 10121
rect 9033 10081 9045 10115
rect 9079 10081 9091 10115
rect 9033 10075 9091 10081
rect 9309 10115 9367 10121
rect 9309 10081 9321 10115
rect 9355 10112 9367 10115
rect 9766 10112 9772 10124
rect 9355 10084 9772 10112
rect 9355 10081 9367 10084
rect 9309 10075 9367 10081
rect 9766 10072 9772 10084
rect 9824 10072 9830 10124
rect 13096 10112 13124 10208
rect 13188 10152 17816 10180
rect 13188 10124 13216 10152
rect 9876 10084 13124 10112
rect 6181 10047 6239 10053
rect 6181 10013 6193 10047
rect 6227 10013 6239 10047
rect 6181 10007 6239 10013
rect 7469 10047 7527 10053
rect 7469 10013 7481 10047
rect 7515 10013 7527 10047
rect 7469 10007 7527 10013
rect 7837 10047 7895 10053
rect 7837 10013 7849 10047
rect 7883 10044 7895 10047
rect 7926 10044 7932 10056
rect 7883 10016 7932 10044
rect 7883 10013 7895 10016
rect 7837 10007 7895 10013
rect 7926 10004 7932 10016
rect 7984 10004 7990 10056
rect 8018 10004 8024 10056
rect 8076 10004 8082 10056
rect 8322 10047 8380 10053
rect 8322 10013 8334 10047
rect 8368 10044 8380 10047
rect 8680 10044 8708 10072
rect 8368 10016 8708 10044
rect 8368 10013 8380 10016
rect 8322 10007 8380 10013
rect 8938 10004 8944 10056
rect 8996 10044 9002 10056
rect 9125 10047 9183 10053
rect 9125 10044 9137 10047
rect 8996 10016 9137 10044
rect 8996 10004 9002 10016
rect 9125 10013 9137 10016
rect 9171 10013 9183 10047
rect 9125 10007 9183 10013
rect 9217 10047 9275 10053
rect 9217 10013 9229 10047
rect 9263 10044 9275 10047
rect 9876 10044 9904 10084
rect 13170 10072 13176 10124
rect 13228 10072 13234 10124
rect 13262 10072 13268 10124
rect 13320 10112 13326 10124
rect 13725 10115 13783 10121
rect 13725 10112 13737 10115
rect 13320 10084 13737 10112
rect 13320 10072 13326 10084
rect 13725 10081 13737 10084
rect 13771 10081 13783 10115
rect 13725 10075 13783 10081
rect 9263 10016 9904 10044
rect 9263 10013 9275 10016
rect 9217 10007 9275 10013
rect 8036 9976 8064 10004
rect 8036 9948 8248 9976
rect 5169 9911 5227 9917
rect 5169 9877 5181 9911
rect 5215 9877 5227 9911
rect 5169 9871 5227 9877
rect 5626 9868 5632 9920
rect 5684 9908 5690 9920
rect 5810 9908 5816 9920
rect 5684 9880 5816 9908
rect 5684 9868 5690 9880
rect 5810 9868 5816 9880
rect 5868 9868 5874 9920
rect 8220 9917 8248 9948
rect 8478 9936 8484 9988
rect 8536 9976 8542 9988
rect 9232 9976 9260 10007
rect 11422 10004 11428 10056
rect 11480 10004 11486 10056
rect 11514 10004 11520 10056
rect 11572 10044 11578 10056
rect 11701 10047 11759 10053
rect 11701 10044 11713 10047
rect 11572 10016 11713 10044
rect 11572 10004 11578 10016
rect 11701 10013 11713 10016
rect 11747 10013 11759 10047
rect 11701 10007 11759 10013
rect 13446 10004 13452 10056
rect 13504 10044 13510 10056
rect 16666 10044 16672 10056
rect 13504 10016 16672 10044
rect 13504 10004 13510 10016
rect 16666 10004 16672 10016
rect 16724 10004 16730 10056
rect 17788 10053 17816 10152
rect 18138 10112 18144 10124
rect 17880 10084 18144 10112
rect 17681 10047 17739 10053
rect 17681 10013 17693 10047
rect 17727 10013 17739 10047
rect 17681 10007 17739 10013
rect 17773 10047 17831 10053
rect 17773 10013 17785 10047
rect 17819 10013 17831 10047
rect 17773 10007 17831 10013
rect 11977 9979 12035 9985
rect 11977 9976 11989 9979
rect 8536 9948 9260 9976
rect 11624 9948 11989 9976
rect 8536 9936 8542 9948
rect 7745 9911 7803 9917
rect 7745 9877 7757 9911
rect 7791 9908 7803 9911
rect 8113 9911 8171 9917
rect 8113 9908 8125 9911
rect 7791 9880 8125 9908
rect 7791 9877 7803 9880
rect 7745 9871 7803 9877
rect 8113 9877 8125 9880
rect 8159 9877 8171 9911
rect 8113 9871 8171 9877
rect 8205 9911 8263 9917
rect 8205 9877 8217 9911
rect 8251 9877 8263 9911
rect 8205 9871 8263 9877
rect 9490 9868 9496 9920
rect 9548 9868 9554 9920
rect 11624 9917 11652 9948
rect 11977 9945 11989 9948
rect 12023 9945 12035 9979
rect 11977 9939 12035 9945
rect 12986 9936 12992 9988
rect 13044 9936 13050 9988
rect 17696 9976 17724 10007
rect 17880 9976 17908 10084
rect 18138 10072 18144 10084
rect 18196 10072 18202 10124
rect 20732 10112 20760 10220
rect 20901 10217 20913 10251
rect 20947 10248 20959 10251
rect 22002 10248 22008 10260
rect 20947 10220 22008 10248
rect 20947 10217 20959 10220
rect 20901 10211 20959 10217
rect 22002 10208 22008 10220
rect 22060 10208 22066 10260
rect 22370 10208 22376 10260
rect 22428 10208 22434 10260
rect 22554 10208 22560 10260
rect 22612 10208 22618 10260
rect 22646 10208 22652 10260
rect 22704 10208 22710 10260
rect 22738 10208 22744 10260
rect 22796 10208 22802 10260
rect 27246 10208 27252 10260
rect 27304 10248 27310 10260
rect 27890 10248 27896 10260
rect 27304 10220 27896 10248
rect 27304 10208 27310 10220
rect 27890 10208 27896 10220
rect 27948 10208 27954 10260
rect 28442 10208 28448 10260
rect 28500 10248 28506 10260
rect 30558 10248 30564 10260
rect 28500 10220 30564 10248
rect 28500 10208 28506 10220
rect 30558 10208 30564 10220
rect 30616 10208 30622 10260
rect 32677 10251 32735 10257
rect 32677 10217 32689 10251
rect 32723 10248 32735 10251
rect 32766 10248 32772 10260
rect 32723 10220 32772 10248
rect 32723 10217 32735 10220
rect 32677 10211 32735 10217
rect 32766 10208 32772 10220
rect 32824 10208 32830 10260
rect 33502 10208 33508 10260
rect 33560 10208 33566 10260
rect 20809 10183 20867 10189
rect 20809 10149 20821 10183
rect 20855 10180 20867 10183
rect 21177 10183 21235 10189
rect 21177 10180 21189 10183
rect 20855 10152 21189 10180
rect 20855 10149 20867 10152
rect 20809 10143 20867 10149
rect 21177 10149 21189 10152
rect 21223 10149 21235 10183
rect 21177 10143 21235 10149
rect 21637 10183 21695 10189
rect 21637 10149 21649 10183
rect 21683 10149 21695 10183
rect 22186 10180 22192 10192
rect 21637 10143 21695 10149
rect 21836 10152 22192 10180
rect 21269 10115 21327 10121
rect 21269 10112 21281 10115
rect 18340 10084 18552 10112
rect 18046 10004 18052 10056
rect 18104 10004 18110 10056
rect 18230 10004 18236 10056
rect 18288 10004 18294 10056
rect 18340 10053 18368 10084
rect 18524 10056 18552 10084
rect 20456 10084 20668 10112
rect 20732 10084 21281 10112
rect 18325 10047 18383 10053
rect 18325 10013 18337 10047
rect 18371 10013 18383 10047
rect 18325 10007 18383 10013
rect 18414 10004 18420 10056
rect 18472 10004 18478 10056
rect 18506 10004 18512 10056
rect 18564 10004 18570 10056
rect 20162 10004 20168 10056
rect 20220 10044 20226 10056
rect 20456 10053 20484 10084
rect 20640 10056 20668 10084
rect 21269 10081 21281 10084
rect 21315 10081 21327 10115
rect 21269 10075 21327 10081
rect 21361 10115 21419 10121
rect 21361 10081 21373 10115
rect 21407 10112 21419 10115
rect 21652 10112 21680 10143
rect 21407 10084 21680 10112
rect 21407 10081 21419 10084
rect 21361 10075 21419 10081
rect 20257 10047 20315 10053
rect 20257 10044 20269 10047
rect 20220 10016 20269 10044
rect 20220 10004 20226 10016
rect 20257 10013 20269 10016
rect 20303 10013 20315 10047
rect 20257 10007 20315 10013
rect 20441 10047 20499 10053
rect 20441 10013 20453 10047
rect 20487 10013 20499 10047
rect 20441 10007 20499 10013
rect 20530 10004 20536 10056
rect 20588 10004 20594 10056
rect 20622 10004 20628 10056
rect 20680 10004 20686 10056
rect 21085 10047 21143 10053
rect 21085 10013 21097 10047
rect 21131 10044 21143 10047
rect 21174 10044 21180 10056
rect 21131 10016 21180 10044
rect 21131 10013 21143 10016
rect 21085 10007 21143 10013
rect 21174 10004 21180 10016
rect 21232 10004 21238 10056
rect 21450 10004 21456 10056
rect 21508 10004 21514 10056
rect 21545 10047 21603 10053
rect 21545 10013 21557 10047
rect 21591 10044 21603 10047
rect 21836 10044 21864 10152
rect 22186 10140 22192 10152
rect 22244 10180 22250 10192
rect 22572 10180 22600 10208
rect 22244 10152 22600 10180
rect 22244 10140 22250 10152
rect 22373 10115 22431 10121
rect 22373 10081 22385 10115
rect 22419 10112 22431 10115
rect 22756 10112 22784 10208
rect 25958 10140 25964 10192
rect 26016 10180 26022 10192
rect 28460 10180 28488 10208
rect 26016 10152 28488 10180
rect 28997 10183 29055 10189
rect 26016 10140 26022 10152
rect 28997 10149 29009 10183
rect 29043 10180 29055 10183
rect 29086 10180 29092 10192
rect 29043 10152 29092 10180
rect 29043 10149 29055 10152
rect 28997 10143 29055 10149
rect 29086 10140 29092 10152
rect 29144 10140 29150 10192
rect 30380 10140 30386 10192
rect 30438 10140 30444 10192
rect 30576 10180 30604 10208
rect 30484 10152 30604 10180
rect 24394 10112 24400 10124
rect 22419 10084 22784 10112
rect 23676 10084 24400 10112
rect 22419 10081 22431 10084
rect 22373 10075 22431 10081
rect 21591 10016 21864 10044
rect 21591 10013 21603 10016
rect 21545 10007 21603 10013
rect 21910 10004 21916 10056
rect 21968 10004 21974 10056
rect 22278 10004 22284 10056
rect 22336 10004 22342 10056
rect 17696 9948 17908 9976
rect 17957 9979 18015 9985
rect 17957 9945 17969 9979
rect 18003 9976 18015 9979
rect 19337 9979 19395 9985
rect 19337 9976 19349 9979
rect 18003 9948 19349 9976
rect 18003 9945 18015 9948
rect 17957 9939 18015 9945
rect 19337 9945 19349 9948
rect 19383 9945 19395 9979
rect 19337 9939 19395 9945
rect 19705 9979 19763 9985
rect 19705 9945 19717 9979
rect 19751 9976 19763 9979
rect 20809 9979 20867 9985
rect 19751 9948 20760 9976
rect 19751 9945 19763 9948
rect 19705 9939 19763 9945
rect 11609 9911 11667 9917
rect 11609 9877 11621 9911
rect 11655 9877 11667 9911
rect 11609 9871 11667 9877
rect 18690 9868 18696 9920
rect 18748 9868 18754 9920
rect 20070 9868 20076 9920
rect 20128 9908 20134 9920
rect 20625 9911 20683 9917
rect 20625 9908 20637 9911
rect 20128 9880 20637 9908
rect 20128 9868 20134 9880
rect 20625 9877 20637 9880
rect 20671 9877 20683 9911
rect 20732 9908 20760 9948
rect 20809 9945 20821 9979
rect 20855 9976 20867 9979
rect 20898 9976 20904 9988
rect 20855 9948 20904 9976
rect 20855 9945 20867 9948
rect 20809 9939 20867 9945
rect 20898 9936 20904 9948
rect 20956 9936 20962 9988
rect 21468 9976 21496 10004
rect 21637 9979 21695 9985
rect 21637 9976 21649 9979
rect 21468 9948 21649 9976
rect 21637 9945 21649 9948
rect 21683 9945 21695 9979
rect 23676 9976 23704 10084
rect 24394 10072 24400 10084
rect 24452 10112 24458 10124
rect 25038 10112 25044 10124
rect 24452 10084 25044 10112
rect 24452 10072 24458 10084
rect 25038 10072 25044 10084
rect 25096 10072 25102 10124
rect 27614 10072 27620 10124
rect 27672 10112 27678 10124
rect 27672 10084 30144 10112
rect 27672 10072 27678 10084
rect 23934 10004 23940 10056
rect 23992 10044 23998 10056
rect 26234 10044 26240 10056
rect 23992 10016 26240 10044
rect 23992 10004 23998 10016
rect 26234 10004 26240 10016
rect 26292 10004 26298 10056
rect 28258 10004 28264 10056
rect 28316 10044 28322 10056
rect 28629 10047 28687 10053
rect 28629 10044 28641 10047
rect 28316 10016 28641 10044
rect 28316 10004 28322 10016
rect 28629 10013 28641 10016
rect 28675 10013 28687 10047
rect 28629 10007 28687 10013
rect 28718 10004 28724 10056
rect 28776 10004 28782 10056
rect 28810 10004 28816 10056
rect 28868 10044 28874 10056
rect 30116 10053 30144 10084
rect 28905 10047 28963 10053
rect 28905 10044 28917 10047
rect 28868 10016 28917 10044
rect 28868 10004 28874 10016
rect 28905 10013 28917 10016
rect 28951 10013 28963 10047
rect 28905 10007 28963 10013
rect 30101 10047 30159 10053
rect 30101 10013 30113 10047
rect 30147 10013 30159 10047
rect 30101 10007 30159 10013
rect 30282 10004 30288 10056
rect 30340 10004 30346 10056
rect 30398 10053 30426 10140
rect 30484 10121 30512 10152
rect 30469 10115 30527 10121
rect 30469 10081 30481 10115
rect 30515 10081 30527 10115
rect 30469 10075 30527 10081
rect 32950 10072 32956 10124
rect 33008 10112 33014 10124
rect 33008 10084 33916 10112
rect 33008 10072 33014 10084
rect 30377 10047 30435 10053
rect 30377 10013 30389 10047
rect 30423 10013 30435 10047
rect 30377 10007 30435 10013
rect 30650 10004 30656 10056
rect 30708 10044 30714 10056
rect 32585 10047 32643 10053
rect 32585 10044 32597 10047
rect 30708 10016 32597 10044
rect 30708 10004 30714 10016
rect 32585 10013 32597 10016
rect 32631 10044 32643 10047
rect 32858 10044 32864 10056
rect 32631 10016 32864 10044
rect 32631 10013 32643 10016
rect 32585 10007 32643 10013
rect 32858 10004 32864 10016
rect 32916 10004 32922 10056
rect 33888 10053 33916 10084
rect 33781 10047 33839 10053
rect 33781 10013 33793 10047
rect 33827 10013 33839 10047
rect 33781 10007 33839 10013
rect 33873 10047 33931 10053
rect 33873 10013 33885 10047
rect 33919 10013 33931 10047
rect 33873 10007 33931 10013
rect 21637 9939 21695 9945
rect 21744 9948 23704 9976
rect 21744 9908 21772 9948
rect 23750 9936 23756 9988
rect 23808 9976 23814 9988
rect 28445 9979 28503 9985
rect 28445 9976 28457 9979
rect 23808 9948 28457 9976
rect 23808 9936 23814 9948
rect 28445 9945 28457 9948
rect 28491 9976 28503 9979
rect 28994 9976 29000 9988
rect 28491 9948 29000 9976
rect 28491 9945 28503 9948
rect 28445 9939 28503 9945
rect 28994 9936 29000 9948
rect 29052 9976 29058 9988
rect 33796 9976 33824 10007
rect 33962 10004 33968 10056
rect 34020 10004 34026 10056
rect 34054 10004 34060 10056
rect 34112 10044 34118 10056
rect 34149 10047 34207 10053
rect 34149 10044 34161 10047
rect 34112 10016 34161 10044
rect 34112 10004 34118 10016
rect 34149 10013 34161 10016
rect 34195 10013 34207 10047
rect 34149 10007 34207 10013
rect 29052 9948 33824 9976
rect 29052 9936 29058 9948
rect 20732 9880 21772 9908
rect 20625 9871 20683 9877
rect 21818 9868 21824 9920
rect 21876 9868 21882 9920
rect 22094 9868 22100 9920
rect 22152 9908 22158 9920
rect 26142 9908 26148 9920
rect 22152 9880 26148 9908
rect 22152 9868 22158 9880
rect 26142 9868 26148 9880
rect 26200 9868 26206 9920
rect 27890 9868 27896 9920
rect 27948 9908 27954 9920
rect 28261 9911 28319 9917
rect 28261 9908 28273 9911
rect 27948 9880 28273 9908
rect 27948 9868 27954 9880
rect 28261 9877 28273 9880
rect 28307 9877 28319 9911
rect 28261 9871 28319 9877
rect 30834 9868 30840 9920
rect 30892 9868 30898 9920
rect 1104 9818 38272 9840
rect 1104 9766 4874 9818
rect 4926 9766 4938 9818
rect 4990 9766 5002 9818
rect 5054 9766 5066 9818
rect 5118 9766 5130 9818
rect 5182 9766 35594 9818
rect 35646 9766 35658 9818
rect 35710 9766 35722 9818
rect 35774 9766 35786 9818
rect 35838 9766 35850 9818
rect 35902 9766 38272 9818
rect 1104 9744 38272 9766
rect 3142 9664 3148 9716
rect 3200 9664 3206 9716
rect 6472 9676 6868 9704
rect 3160 9636 3188 9664
rect 3160 9608 3464 9636
rect 3234 9528 3240 9580
rect 3292 9528 3298 9580
rect 3326 9528 3332 9580
rect 3384 9528 3390 9580
rect 3436 9577 3464 9608
rect 5994 9596 6000 9648
rect 6052 9636 6058 9648
rect 6365 9639 6423 9645
rect 6365 9636 6377 9639
rect 6052 9608 6377 9636
rect 6052 9596 6058 9608
rect 6365 9605 6377 9608
rect 6411 9605 6423 9639
rect 6365 9599 6423 9605
rect 3421 9571 3479 9577
rect 3421 9537 3433 9571
rect 3467 9537 3479 9571
rect 3421 9531 3479 9537
rect 3605 9571 3663 9577
rect 3605 9537 3617 9571
rect 3651 9568 3663 9571
rect 3694 9568 3700 9580
rect 3651 9540 3700 9568
rect 3651 9537 3663 9540
rect 3605 9531 3663 9537
rect 3694 9528 3700 9540
rect 3752 9568 3758 9580
rect 4614 9568 4620 9580
rect 3752 9540 4620 9568
rect 3752 9528 3758 9540
rect 4614 9528 4620 9540
rect 4672 9568 4678 9580
rect 6472 9568 6500 9676
rect 6840 9674 6868 9676
rect 8128 9676 8708 9704
rect 6840 9646 6960 9674
rect 6932 9636 6960 9646
rect 8128 9636 8156 9676
rect 6932 9608 8156 9636
rect 4672 9540 6500 9568
rect 4672 9528 4678 9540
rect 6638 9528 6644 9580
rect 6696 9528 6702 9580
rect 6730 9528 6736 9580
rect 6788 9528 6794 9580
rect 6822 9528 6828 9580
rect 6880 9528 6886 9580
rect 7024 9577 7052 9608
rect 8202 9596 8208 9648
rect 8260 9636 8266 9648
rect 8297 9639 8355 9645
rect 8297 9636 8309 9639
rect 8260 9608 8309 9636
rect 8260 9596 8266 9608
rect 8297 9605 8309 9608
rect 8343 9636 8355 9639
rect 8573 9639 8631 9645
rect 8573 9636 8585 9639
rect 8343 9608 8585 9636
rect 8343 9605 8355 9608
rect 8297 9599 8355 9605
rect 8573 9605 8585 9608
rect 8619 9605 8631 9639
rect 8680 9636 8708 9676
rect 9324 9648 9674 9674
rect 11422 9664 11428 9716
rect 11480 9704 11486 9716
rect 11793 9707 11851 9713
rect 11793 9704 11805 9707
rect 11480 9676 11805 9704
rect 11480 9664 11486 9676
rect 11793 9673 11805 9676
rect 11839 9673 11851 9707
rect 11793 9667 11851 9673
rect 13170 9664 13176 9716
rect 13228 9704 13234 9716
rect 13541 9707 13599 9713
rect 13541 9704 13553 9707
rect 13228 9676 13553 9704
rect 13228 9664 13234 9676
rect 13541 9673 13553 9676
rect 13587 9673 13599 9707
rect 13541 9667 13599 9673
rect 15286 9664 15292 9716
rect 15344 9704 15350 9716
rect 15344 9676 15516 9704
rect 15344 9664 15350 9676
rect 8680 9608 9168 9636
rect 8573 9599 8631 9605
rect 7009 9571 7067 9577
rect 7009 9537 7021 9571
rect 7055 9537 7067 9571
rect 7009 9531 7067 9537
rect 7745 9571 7803 9577
rect 7745 9537 7757 9571
rect 7791 9568 7803 9571
rect 7834 9568 7840 9580
rect 7791 9540 7840 9568
rect 7791 9537 7803 9540
rect 7745 9531 7803 9537
rect 7834 9528 7840 9540
rect 7892 9528 7898 9580
rect 8021 9571 8079 9577
rect 8021 9537 8033 9571
rect 8067 9568 8079 9571
rect 8110 9568 8116 9580
rect 8067 9540 8116 9568
rect 8067 9537 8079 9540
rect 8021 9531 8079 9537
rect 8110 9528 8116 9540
rect 8168 9528 8174 9580
rect 8478 9528 8484 9580
rect 8536 9528 8542 9580
rect 8665 9571 8723 9577
rect 8665 9537 8677 9571
rect 8711 9568 8723 9571
rect 8938 9568 8944 9580
rect 8711 9540 8944 9568
rect 8711 9537 8723 9540
rect 8665 9531 8723 9537
rect 8938 9528 8944 9540
rect 8996 9528 9002 9580
rect 9140 9500 9168 9608
rect 9306 9596 9312 9648
rect 9364 9646 9674 9648
rect 9364 9596 9370 9646
rect 9646 9636 9674 9646
rect 15488 9645 15516 9676
rect 16022 9664 16028 9716
rect 16080 9664 16086 9716
rect 18690 9664 18696 9716
rect 18748 9704 18754 9716
rect 18748 9676 22324 9704
rect 18748 9664 18754 9676
rect 15473 9639 15531 9645
rect 9646 9608 15424 9636
rect 9950 9568 9956 9580
rect 9600 9566 9956 9568
rect 9324 9540 9956 9566
rect 9324 9538 9628 9540
rect 9324 9500 9352 9538
rect 9950 9528 9956 9540
rect 10008 9528 10014 9580
rect 10229 9571 10287 9577
rect 10229 9537 10241 9571
rect 10275 9568 10287 9571
rect 10275 9540 10364 9568
rect 10275 9537 10287 9540
rect 10229 9531 10287 9537
rect 9140 9472 9352 9500
rect 7466 9392 7472 9444
rect 7524 9392 7530 9444
rect 8021 9435 8079 9441
rect 8021 9401 8033 9435
rect 8067 9432 8079 9435
rect 8202 9432 8208 9444
rect 8067 9404 8208 9432
rect 8067 9401 8079 9404
rect 8021 9395 8079 9401
rect 8202 9392 8208 9404
rect 8260 9392 8266 9444
rect 10336 9441 10364 9540
rect 10502 9528 10508 9580
rect 10560 9568 10566 9580
rect 10689 9571 10747 9577
rect 10689 9568 10701 9571
rect 10560 9540 10701 9568
rect 10560 9528 10566 9540
rect 10689 9537 10701 9540
rect 10735 9537 10747 9571
rect 10689 9531 10747 9537
rect 10781 9571 10839 9577
rect 10781 9537 10793 9571
rect 10827 9568 10839 9571
rect 11606 9568 11612 9580
rect 10827 9540 11612 9568
rect 10827 9537 10839 9540
rect 10781 9531 10839 9537
rect 10321 9435 10379 9441
rect 9646 9404 10180 9432
rect 2958 9324 2964 9376
rect 3016 9324 3022 9376
rect 6730 9324 6736 9376
rect 6788 9364 6794 9376
rect 9646 9364 9674 9404
rect 6788 9336 9674 9364
rect 6788 9324 6794 9336
rect 10042 9324 10048 9376
rect 10100 9324 10106 9376
rect 10152 9364 10180 9404
rect 10321 9401 10333 9435
rect 10367 9401 10379 9435
rect 10704 9432 10732 9531
rect 11606 9528 11612 9540
rect 11664 9528 11670 9580
rect 12161 9571 12219 9577
rect 12161 9537 12173 9571
rect 12207 9537 12219 9571
rect 12161 9531 12219 9537
rect 12253 9571 12311 9577
rect 12253 9537 12265 9571
rect 12299 9568 12311 9571
rect 13262 9568 13268 9580
rect 12299 9540 13268 9568
rect 12299 9537 12311 9540
rect 12253 9531 12311 9537
rect 10870 9460 10876 9512
rect 10928 9460 10934 9512
rect 12176 9432 12204 9531
rect 13262 9528 13268 9540
rect 13320 9528 13326 9580
rect 13449 9571 13507 9577
rect 13449 9537 13461 9571
rect 13495 9537 13507 9571
rect 13449 9531 13507 9537
rect 12437 9503 12495 9509
rect 12437 9469 12449 9503
rect 12483 9500 12495 9503
rect 12526 9500 12532 9512
rect 12483 9472 12532 9500
rect 12483 9469 12495 9472
rect 12437 9463 12495 9469
rect 12526 9460 12532 9472
rect 12584 9460 12590 9512
rect 10704 9404 12204 9432
rect 10321 9395 10379 9401
rect 13464 9376 13492 9531
rect 13633 9503 13691 9509
rect 13633 9469 13645 9503
rect 13679 9469 13691 9503
rect 13633 9463 13691 9469
rect 15289 9503 15347 9509
rect 15289 9469 15301 9503
rect 15335 9469 15347 9503
rect 15396 9500 15424 9608
rect 15473 9605 15485 9639
rect 15519 9636 15531 9639
rect 19978 9636 19984 9648
rect 15519 9608 17264 9636
rect 15519 9605 15531 9608
rect 15473 9599 15531 9605
rect 15562 9528 15568 9580
rect 15620 9528 15626 9580
rect 15930 9528 15936 9580
rect 15988 9568 15994 9580
rect 16209 9571 16267 9577
rect 16209 9568 16221 9571
rect 15988 9540 16221 9568
rect 15988 9528 15994 9540
rect 16209 9537 16221 9540
rect 16255 9537 16267 9571
rect 16209 9531 16267 9537
rect 16666 9528 16672 9580
rect 16724 9568 16730 9580
rect 16761 9571 16819 9577
rect 16761 9568 16773 9571
rect 16724 9540 16773 9568
rect 16724 9528 16730 9540
rect 16761 9537 16773 9540
rect 16807 9568 16819 9571
rect 16942 9568 16948 9580
rect 16807 9540 16948 9568
rect 16807 9537 16819 9540
rect 16761 9531 16819 9537
rect 16942 9528 16948 9540
rect 17000 9528 17006 9580
rect 15396 9472 16344 9500
rect 15289 9463 15347 9469
rect 10502 9364 10508 9376
rect 10152 9336 10508 9364
rect 10502 9324 10508 9336
rect 10560 9324 10566 9376
rect 13078 9324 13084 9376
rect 13136 9324 13142 9376
rect 13446 9324 13452 9376
rect 13504 9324 13510 9376
rect 13648 9364 13676 9463
rect 13722 9392 13728 9444
rect 13780 9432 13786 9444
rect 15304 9432 15332 9463
rect 15838 9432 15844 9444
rect 13780 9404 15844 9432
rect 13780 9392 13786 9404
rect 15838 9392 15844 9404
rect 15896 9392 15902 9444
rect 15930 9392 15936 9444
rect 15988 9392 15994 9444
rect 16316 9432 16344 9472
rect 17126 9460 17132 9512
rect 17184 9460 17190 9512
rect 17236 9500 17264 9608
rect 18064 9608 18828 9636
rect 18064 9580 18092 9608
rect 18046 9528 18052 9580
rect 18104 9528 18110 9580
rect 18417 9571 18475 9577
rect 18417 9537 18429 9571
rect 18463 9568 18475 9571
rect 18506 9568 18512 9580
rect 18463 9540 18512 9568
rect 18463 9537 18475 9540
rect 18417 9531 18475 9537
rect 18506 9528 18512 9540
rect 18564 9528 18570 9580
rect 18800 9577 18828 9608
rect 19812 9608 19984 9636
rect 19812 9577 19840 9608
rect 19978 9596 19984 9608
rect 20036 9636 20042 9648
rect 20036 9608 20576 9636
rect 20036 9596 20042 9608
rect 20548 9580 20576 9608
rect 21082 9596 21088 9648
rect 21140 9636 21146 9648
rect 21634 9636 21640 9648
rect 21140 9608 21640 9636
rect 21140 9596 21146 9608
rect 21634 9596 21640 9608
rect 21692 9596 21698 9648
rect 22296 9636 22324 9676
rect 22370 9664 22376 9716
rect 22428 9704 22434 9716
rect 22465 9707 22523 9713
rect 22465 9704 22477 9707
rect 22428 9676 22477 9704
rect 22428 9664 22434 9676
rect 22465 9673 22477 9676
rect 22511 9673 22523 9707
rect 23934 9704 23940 9716
rect 22465 9667 22523 9673
rect 22572 9676 23940 9704
rect 22572 9636 22600 9676
rect 23934 9664 23940 9676
rect 23992 9664 23998 9716
rect 24026 9664 24032 9716
rect 24084 9704 24090 9716
rect 28810 9704 28816 9716
rect 24084 9676 24716 9704
rect 24084 9664 24090 9676
rect 24688 9645 24716 9676
rect 26252 9676 28816 9704
rect 24581 9639 24639 9645
rect 24581 9636 24593 9639
rect 22296 9608 22600 9636
rect 22940 9608 24593 9636
rect 22940 9580 22968 9608
rect 24581 9605 24593 9608
rect 24627 9605 24639 9639
rect 24581 9599 24639 9605
rect 24673 9639 24731 9645
rect 24673 9605 24685 9639
rect 24719 9636 24731 9639
rect 26252 9636 26280 9676
rect 28810 9664 28816 9676
rect 28868 9664 28874 9716
rect 30374 9704 30380 9716
rect 24719 9608 26280 9636
rect 26329 9639 26387 9645
rect 24719 9605 24731 9608
rect 24673 9599 24731 9605
rect 26329 9605 26341 9639
rect 26375 9636 26387 9639
rect 26375 9608 27752 9636
rect 26375 9605 26387 9608
rect 26329 9599 26387 9605
rect 27724 9580 27752 9608
rect 18785 9571 18843 9577
rect 18785 9537 18797 9571
rect 18831 9537 18843 9571
rect 18785 9531 18843 9537
rect 19797 9571 19855 9577
rect 19797 9537 19809 9571
rect 19843 9537 19855 9571
rect 19797 9531 19855 9537
rect 20073 9571 20131 9577
rect 20073 9537 20085 9571
rect 20119 9568 20131 9571
rect 20162 9568 20168 9580
rect 20119 9540 20168 9568
rect 20119 9537 20131 9540
rect 20073 9531 20131 9537
rect 20162 9528 20168 9540
rect 20220 9528 20226 9580
rect 20254 9528 20260 9580
rect 20312 9528 20318 9580
rect 20530 9528 20536 9580
rect 20588 9528 20594 9580
rect 22649 9571 22707 9577
rect 22649 9537 22661 9571
rect 22695 9537 22707 9571
rect 22649 9531 22707 9537
rect 18230 9500 18236 9512
rect 17236 9472 18236 9500
rect 18230 9460 18236 9472
rect 18288 9460 18294 9512
rect 18874 9460 18880 9512
rect 18932 9460 18938 9512
rect 19426 9460 19432 9512
rect 19484 9460 19490 9512
rect 19889 9503 19947 9509
rect 19889 9469 19901 9503
rect 19935 9469 19947 9503
rect 19889 9463 19947 9469
rect 19981 9503 20039 9509
rect 19981 9469 19993 9503
rect 20027 9500 20039 9503
rect 20272 9500 20300 9528
rect 22664 9500 22692 9531
rect 22738 9528 22744 9580
rect 22796 9528 22802 9580
rect 22922 9528 22928 9580
rect 22980 9528 22986 9580
rect 23017 9571 23075 9577
rect 23017 9537 23029 9571
rect 23063 9568 23075 9571
rect 23063 9540 23336 9568
rect 23063 9537 23075 9540
rect 23017 9531 23075 9537
rect 23308 9512 23336 9540
rect 23382 9528 23388 9580
rect 23440 9568 23446 9580
rect 24121 9571 24179 9577
rect 24121 9568 24133 9571
rect 23440 9540 24133 9568
rect 23440 9528 23446 9540
rect 24121 9537 24133 9540
rect 24167 9537 24179 9571
rect 24121 9531 24179 9537
rect 24210 9528 24216 9580
rect 24268 9568 24274 9580
rect 24305 9571 24363 9577
rect 24305 9568 24317 9571
rect 24268 9540 24317 9568
rect 24268 9528 24274 9540
rect 24305 9537 24317 9540
rect 24351 9537 24363 9571
rect 24305 9531 24363 9537
rect 23109 9503 23167 9509
rect 20027 9472 23060 9500
rect 20027 9469 20039 9472
rect 19981 9463 20039 9469
rect 19904 9432 19932 9463
rect 23032 9444 23060 9472
rect 23109 9469 23121 9503
rect 23155 9469 23167 9503
rect 23109 9463 23167 9469
rect 20070 9432 20076 9444
rect 16316 9404 18552 9432
rect 19904 9404 20076 9432
rect 18524 9376 18552 9404
rect 20070 9392 20076 9404
rect 20128 9392 20134 9444
rect 23014 9392 23020 9444
rect 23072 9392 23078 9444
rect 23124 9432 23152 9463
rect 23290 9460 23296 9512
rect 23348 9460 23354 9512
rect 24320 9500 24348 9531
rect 24394 9528 24400 9580
rect 24452 9528 24458 9580
rect 24765 9571 24823 9577
rect 24765 9537 24777 9571
rect 24811 9537 24823 9571
rect 24765 9531 24823 9537
rect 24780 9500 24808 9531
rect 26142 9528 26148 9580
rect 26200 9568 26206 9580
rect 26421 9571 26479 9577
rect 26421 9568 26433 9571
rect 26200 9540 26433 9568
rect 26200 9528 26206 9540
rect 26421 9537 26433 9540
rect 26467 9537 26479 9571
rect 26421 9531 26479 9537
rect 26605 9571 26663 9577
rect 26605 9537 26617 9571
rect 26651 9537 26663 9571
rect 26605 9531 26663 9537
rect 25961 9503 26019 9509
rect 25961 9500 25973 9503
rect 24320 9472 24808 9500
rect 24872 9472 25973 9500
rect 24210 9432 24216 9444
rect 23124 9404 24216 9432
rect 24210 9392 24216 9404
rect 24268 9432 24274 9444
rect 24762 9432 24768 9444
rect 24268 9404 24768 9432
rect 24268 9392 24274 9404
rect 24762 9392 24768 9404
rect 24820 9392 24826 9444
rect 13906 9364 13912 9376
rect 13648 9336 13912 9364
rect 13906 9324 13912 9336
rect 13964 9324 13970 9376
rect 18506 9324 18512 9376
rect 18564 9324 18570 9376
rect 19610 9324 19616 9376
rect 19668 9324 19674 9376
rect 24302 9324 24308 9376
rect 24360 9324 24366 9376
rect 24578 9324 24584 9376
rect 24636 9364 24642 9376
rect 24872 9364 24900 9472
rect 25961 9469 25973 9472
rect 26007 9500 26019 9503
rect 26620 9500 26648 9531
rect 26970 9528 26976 9580
rect 27028 9528 27034 9580
rect 27154 9528 27160 9580
rect 27212 9568 27218 9580
rect 27338 9568 27344 9580
rect 27212 9540 27344 9568
rect 27212 9528 27218 9540
rect 27338 9528 27344 9540
rect 27396 9528 27402 9580
rect 27430 9528 27436 9580
rect 27488 9528 27494 9580
rect 27522 9528 27528 9580
rect 27580 9568 27586 9580
rect 27580 9540 27660 9568
rect 27580 9528 27586 9540
rect 26007 9472 26648 9500
rect 26988 9500 27016 9528
rect 27632 9500 27660 9540
rect 27706 9528 27712 9580
rect 27764 9528 27770 9580
rect 28828 9568 28856 9664
rect 29454 9634 29460 9686
rect 29512 9634 29518 9686
rect 29656 9676 30380 9704
rect 29656 9636 29684 9676
rect 30374 9664 30380 9676
rect 30432 9664 30438 9716
rect 33134 9664 33140 9716
rect 33192 9704 33198 9716
rect 33229 9707 33287 9713
rect 33229 9704 33241 9707
rect 33192 9676 33241 9704
rect 33192 9664 33198 9676
rect 33229 9673 33241 9676
rect 33275 9704 33287 9707
rect 33962 9704 33968 9716
rect 33275 9676 33968 9704
rect 33275 9673 33287 9676
rect 33229 9667 33287 9673
rect 33962 9664 33968 9676
rect 34020 9664 34026 9716
rect 30006 9636 30012 9648
rect 29472 9580 29500 9634
rect 29656 9608 29776 9636
rect 28997 9571 29055 9577
rect 28997 9568 29009 9571
rect 28828 9540 29009 9568
rect 28997 9537 29009 9540
rect 29043 9537 29055 9571
rect 28997 9531 29055 9537
rect 29454 9528 29460 9580
rect 29512 9528 29518 9580
rect 29546 9528 29552 9580
rect 29604 9528 29610 9580
rect 29641 9574 29699 9577
rect 29748 9574 29776 9608
rect 29840 9608 30012 9636
rect 29840 9577 29868 9608
rect 30006 9596 30012 9608
rect 30064 9596 30070 9648
rect 31496 9608 32444 9636
rect 29641 9571 29776 9574
rect 29641 9537 29653 9571
rect 29687 9546 29776 9571
rect 29825 9571 29883 9577
rect 29687 9537 29699 9546
rect 29641 9531 29699 9537
rect 29825 9537 29837 9571
rect 29871 9537 29883 9571
rect 29825 9531 29883 9537
rect 29925 9571 29983 9577
rect 29925 9537 29937 9571
rect 29971 9568 29983 9571
rect 29971 9540 30052 9568
rect 29971 9537 29983 9540
rect 29925 9531 29983 9537
rect 28718 9500 28724 9512
rect 26988 9472 27568 9500
rect 27632 9472 28724 9500
rect 26007 9469 26019 9472
rect 25961 9463 26019 9469
rect 24949 9435 25007 9441
rect 24949 9401 24961 9435
rect 24995 9432 25007 9435
rect 27430 9432 27436 9444
rect 24995 9404 27436 9432
rect 24995 9401 25007 9404
rect 24949 9395 25007 9401
rect 27430 9392 27436 9404
rect 27488 9392 27494 9444
rect 27540 9432 27568 9472
rect 28718 9460 28724 9472
rect 28776 9500 28782 9512
rect 28813 9503 28871 9509
rect 28813 9500 28825 9503
rect 28776 9472 28825 9500
rect 28776 9460 28782 9472
rect 28813 9469 28825 9472
rect 28859 9469 28871 9503
rect 29564 9500 29592 9528
rect 29733 9503 29791 9509
rect 29733 9500 29745 9503
rect 29564 9472 29745 9500
rect 28813 9463 28871 9469
rect 29733 9469 29745 9472
rect 29779 9469 29791 9503
rect 29733 9463 29791 9469
rect 30024 9432 30052 9540
rect 30101 9561 30159 9567
rect 30101 9527 30113 9561
rect 30147 9558 30159 9561
rect 30147 9530 30236 9558
rect 30147 9527 30159 9530
rect 30101 9521 30159 9527
rect 27540 9404 30052 9432
rect 30098 9392 30104 9444
rect 30156 9432 30162 9444
rect 30208 9432 30236 9530
rect 30742 9528 30748 9580
rect 30800 9528 30806 9580
rect 30834 9528 30840 9580
rect 30892 9568 30898 9580
rect 31021 9571 31079 9577
rect 31021 9568 31033 9571
rect 30892 9540 31033 9568
rect 30892 9528 30898 9540
rect 31021 9537 31033 9540
rect 31067 9537 31079 9571
rect 31021 9531 31079 9537
rect 31297 9571 31355 9577
rect 31297 9537 31309 9571
rect 31343 9568 31355 9571
rect 31386 9568 31392 9580
rect 31343 9540 31392 9568
rect 31343 9537 31355 9540
rect 31297 9531 31355 9537
rect 31386 9528 31392 9540
rect 31444 9528 31450 9580
rect 30156 9404 30236 9432
rect 30156 9392 30162 9404
rect 30926 9392 30932 9444
rect 30984 9432 30990 9444
rect 31205 9435 31263 9441
rect 31205 9432 31217 9435
rect 30984 9404 31217 9432
rect 30984 9392 30990 9404
rect 31205 9401 31217 9404
rect 31251 9401 31263 9435
rect 31205 9395 31263 9401
rect 24636 9336 24900 9364
rect 24636 9324 24642 9336
rect 26510 9324 26516 9376
rect 26568 9364 26574 9376
rect 27522 9364 27528 9376
rect 26568 9336 27528 9364
rect 26568 9324 26574 9336
rect 27522 9324 27528 9336
rect 27580 9324 27586 9376
rect 27617 9367 27675 9373
rect 27617 9333 27629 9367
rect 27663 9364 27675 9367
rect 28074 9364 28080 9376
rect 27663 9336 28080 9364
rect 27663 9333 27675 9336
rect 27617 9327 27675 9333
rect 28074 9324 28080 9336
rect 28132 9324 28138 9376
rect 29181 9367 29239 9373
rect 29181 9333 29193 9367
rect 29227 9364 29239 9367
rect 29730 9364 29736 9376
rect 29227 9336 29736 9364
rect 29227 9333 29239 9336
rect 29181 9327 29239 9333
rect 29730 9324 29736 9336
rect 29788 9324 29794 9376
rect 30009 9367 30067 9373
rect 30009 9333 30021 9367
rect 30055 9364 30067 9367
rect 31496 9364 31524 9608
rect 31573 9571 31631 9577
rect 31573 9537 31585 9571
rect 31619 9537 31631 9571
rect 31573 9531 31631 9537
rect 31588 9376 31616 9531
rect 32416 9509 32444 9608
rect 33042 9596 33048 9648
rect 33100 9596 33106 9648
rect 32493 9571 32551 9577
rect 32493 9537 32505 9571
rect 32539 9568 32551 9571
rect 32766 9568 32772 9580
rect 32539 9540 32772 9568
rect 32539 9537 32551 9540
rect 32493 9531 32551 9537
rect 32766 9528 32772 9540
rect 32824 9528 32830 9580
rect 32861 9571 32919 9577
rect 32861 9537 32873 9571
rect 32907 9537 32919 9571
rect 32861 9531 32919 9537
rect 32401 9503 32459 9509
rect 32401 9469 32413 9503
rect 32447 9469 32459 9503
rect 32401 9463 32459 9469
rect 32030 9392 32036 9444
rect 32088 9432 32094 9444
rect 32125 9435 32183 9441
rect 32125 9432 32137 9435
rect 32088 9404 32137 9432
rect 32088 9392 32094 9404
rect 32125 9401 32137 9404
rect 32171 9432 32183 9435
rect 32876 9432 32904 9531
rect 32171 9404 32904 9432
rect 32171 9401 32183 9404
rect 32125 9395 32183 9401
rect 30055 9336 31524 9364
rect 30055 9333 30067 9336
rect 30009 9327 30067 9333
rect 31570 9324 31576 9376
rect 31628 9324 31634 9376
rect 31662 9324 31668 9376
rect 31720 9364 31726 9376
rect 33226 9364 33232 9376
rect 31720 9336 33232 9364
rect 31720 9324 31726 9336
rect 33226 9324 33232 9336
rect 33284 9324 33290 9376
rect 1104 9274 38272 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 38272 9274
rect 1104 9200 38272 9222
rect 2958 9160 2964 9172
rect 2746 9132 2964 9160
rect 1765 8959 1823 8965
rect 1765 8925 1777 8959
rect 1811 8956 1823 8959
rect 2746 8956 2774 9132
rect 2958 9120 2964 9132
rect 3016 9120 3022 9172
rect 6730 9120 6736 9172
rect 6788 9120 6794 9172
rect 6914 9120 6920 9172
rect 6972 9160 6978 9172
rect 11517 9163 11575 9169
rect 6972 9132 11468 9160
rect 6972 9120 6978 9132
rect 3326 9052 3332 9104
rect 3384 9092 3390 9104
rect 6748 9092 6776 9120
rect 3384 9064 6776 9092
rect 11440 9092 11468 9132
rect 11517 9129 11529 9163
rect 11563 9160 11575 9163
rect 11606 9160 11612 9172
rect 11563 9132 11612 9160
rect 11563 9129 11575 9132
rect 11517 9123 11575 9129
rect 11606 9120 11612 9132
rect 11664 9120 11670 9172
rect 13078 9160 13084 9172
rect 12406 9132 13084 9160
rect 12406 9092 12434 9132
rect 13078 9120 13084 9132
rect 13136 9120 13142 9172
rect 13814 9120 13820 9172
rect 13872 9120 13878 9172
rect 13906 9120 13912 9172
rect 13964 9160 13970 9172
rect 17497 9163 17555 9169
rect 13964 9132 15148 9160
rect 13964 9120 13970 9132
rect 11440 9064 12434 9092
rect 3384 9052 3390 9064
rect 1811 8928 2774 8956
rect 1811 8925 1823 8928
rect 1765 8919 1823 8925
rect 3050 8916 3056 8968
rect 3108 8916 3114 8968
rect 4154 8916 4160 8968
rect 4212 8916 4218 8968
rect 4264 8965 4292 9064
rect 4617 9027 4675 9033
rect 4617 9024 4629 9027
rect 4356 8996 4629 9024
rect 4356 8965 4384 8996
rect 4617 8993 4629 8996
rect 4663 8993 4675 9027
rect 4617 8987 4675 8993
rect 5626 8984 5632 9036
rect 5684 9024 5690 9036
rect 8665 9027 8723 9033
rect 8665 9024 8677 9027
rect 5684 8996 8677 9024
rect 5684 8984 5690 8996
rect 8665 8993 8677 8996
rect 8711 9024 8723 9027
rect 8711 8996 8892 9024
rect 8711 8993 8723 8996
rect 8665 8987 8723 8993
rect 4249 8959 4307 8965
rect 4249 8925 4261 8959
rect 4295 8925 4307 8959
rect 4249 8919 4307 8925
rect 4341 8959 4399 8965
rect 4341 8925 4353 8959
rect 4387 8925 4399 8959
rect 4341 8919 4399 8925
rect 4522 8916 4528 8968
rect 4580 8916 4586 8968
rect 4985 8959 5043 8965
rect 4985 8956 4997 8959
rect 4632 8928 4997 8956
rect 934 8848 940 8900
rect 992 8888 998 8900
rect 1397 8891 1455 8897
rect 1397 8888 1409 8891
rect 992 8860 1409 8888
rect 992 8848 998 8860
rect 1397 8857 1409 8860
rect 1443 8857 1455 8891
rect 3068 8888 3096 8916
rect 4632 8888 4660 8928
rect 4985 8925 4997 8928
rect 5031 8956 5043 8959
rect 5813 8959 5871 8965
rect 5813 8956 5825 8959
rect 5031 8928 5825 8956
rect 5031 8925 5043 8928
rect 4985 8919 5043 8925
rect 5813 8925 5825 8928
rect 5859 8956 5871 8959
rect 7190 8956 7196 8968
rect 5859 8928 7196 8956
rect 5859 8925 5871 8928
rect 5813 8919 5871 8925
rect 7190 8916 7196 8928
rect 7248 8916 7254 8968
rect 3068 8860 4660 8888
rect 1397 8851 1455 8857
rect 4706 8848 4712 8900
rect 4764 8888 4770 8900
rect 4801 8891 4859 8897
rect 4801 8888 4813 8891
rect 4764 8860 4813 8888
rect 4764 8848 4770 8860
rect 4801 8857 4813 8860
rect 4847 8857 4859 8891
rect 4801 8851 4859 8857
rect 5994 8848 6000 8900
rect 6052 8848 6058 8900
rect 6181 8891 6239 8897
rect 6181 8857 6193 8891
rect 6227 8888 6239 8891
rect 6822 8888 6828 8900
rect 6227 8860 6828 8888
rect 6227 8857 6239 8860
rect 6181 8851 6239 8857
rect 6822 8848 6828 8860
rect 6880 8848 6886 8900
rect 8389 8891 8447 8897
rect 8389 8857 8401 8891
rect 8435 8888 8447 8891
rect 8435 8860 8708 8888
rect 8435 8857 8447 8860
rect 8389 8851 8447 8857
rect 8680 8832 8708 8860
rect 3878 8780 3884 8832
rect 3936 8780 3942 8832
rect 8018 8780 8024 8832
rect 8076 8780 8082 8832
rect 8478 8780 8484 8832
rect 8536 8780 8542 8832
rect 8662 8780 8668 8832
rect 8720 8780 8726 8832
rect 8864 8820 8892 8996
rect 9766 8984 9772 9036
rect 9824 8984 9830 9036
rect 10042 8984 10048 9036
rect 10100 8984 10106 9036
rect 10502 8984 10508 9036
rect 10560 9024 10566 9036
rect 10560 8996 13492 9024
rect 10560 8984 10566 8996
rect 11698 8956 11704 8968
rect 11178 8928 11704 8956
rect 11698 8916 11704 8928
rect 11756 8916 11762 8968
rect 12710 8916 12716 8968
rect 12768 8916 12774 8968
rect 12912 8965 12940 8996
rect 12897 8959 12955 8965
rect 12897 8925 12909 8959
rect 12943 8925 12955 8959
rect 12897 8919 12955 8925
rect 13354 8916 13360 8968
rect 13412 8916 13418 8968
rect 13464 8956 13492 8996
rect 13538 8984 13544 9036
rect 13596 9024 13602 9036
rect 13633 9027 13691 9033
rect 13633 9024 13645 9027
rect 13596 8996 13645 9024
rect 13596 8984 13602 8996
rect 13633 8993 13645 8996
rect 13679 9024 13691 9027
rect 13722 9024 13728 9036
rect 13679 8996 13728 9024
rect 13679 8993 13691 8996
rect 13633 8987 13691 8993
rect 13722 8984 13728 8996
rect 13780 8984 13786 9036
rect 13832 9024 13860 9120
rect 14458 9052 14464 9104
rect 14516 9052 14522 9104
rect 15120 9092 15148 9132
rect 17497 9129 17509 9163
rect 17543 9160 17555 9163
rect 18230 9160 18236 9172
rect 17543 9132 18236 9160
rect 17543 9129 17555 9132
rect 17497 9123 17555 9129
rect 18230 9120 18236 9132
rect 18288 9120 18294 9172
rect 20806 9160 20812 9172
rect 18432 9132 20812 9160
rect 15120 9064 15608 9092
rect 14476 9024 14504 9052
rect 13832 8996 14136 9024
rect 13906 8956 13912 8968
rect 13464 8928 13912 8956
rect 13906 8916 13912 8928
rect 13964 8916 13970 8968
rect 14108 8965 14136 8996
rect 14384 8996 14504 9024
rect 14384 8965 14412 8996
rect 15378 8984 15384 9036
rect 15436 8984 15442 9036
rect 15580 9033 15608 9064
rect 15565 9027 15623 9033
rect 15565 8993 15577 9027
rect 15611 9024 15623 9027
rect 17586 9024 17592 9036
rect 15611 8996 17592 9024
rect 15611 8993 15623 8996
rect 15565 8987 15623 8993
rect 17586 8984 17592 8996
rect 17644 8984 17650 9036
rect 18325 9027 18383 9033
rect 18325 8993 18337 9027
rect 18371 9024 18383 9027
rect 18432 9024 18460 9132
rect 20806 9120 20812 9132
rect 20864 9120 20870 9172
rect 20901 9163 20959 9169
rect 20901 9129 20913 9163
rect 20947 9160 20959 9163
rect 21082 9160 21088 9172
rect 20947 9132 21088 9160
rect 20947 9129 20959 9132
rect 20901 9123 20959 9129
rect 21082 9120 21088 9132
rect 21140 9120 21146 9172
rect 22094 9120 22100 9172
rect 22152 9160 22158 9172
rect 23937 9163 23995 9169
rect 23937 9160 23949 9163
rect 22152 9132 23949 9160
rect 22152 9120 22158 9132
rect 23937 9129 23949 9132
rect 23983 9160 23995 9163
rect 23983 9132 26188 9160
rect 23983 9129 23995 9132
rect 23937 9123 23995 9129
rect 18506 9052 18512 9104
rect 18564 9092 18570 9104
rect 22278 9092 22284 9104
rect 18564 9064 22284 9092
rect 18564 9052 18570 9064
rect 22278 9052 22284 9064
rect 22336 9092 22342 9104
rect 22738 9092 22744 9104
rect 22336 9064 22744 9092
rect 22336 9052 22342 9064
rect 22738 9052 22744 9064
rect 22796 9052 22802 9104
rect 22833 9095 22891 9101
rect 22833 9061 22845 9095
rect 22879 9061 22891 9095
rect 22833 9055 22891 9061
rect 20717 9027 20775 9033
rect 20717 9024 20729 9027
rect 18371 8996 18460 9024
rect 19996 8996 20729 9024
rect 18371 8993 18383 8996
rect 18325 8987 18383 8993
rect 14093 8959 14151 8965
rect 14093 8925 14105 8959
rect 14139 8925 14151 8959
rect 14093 8919 14151 8925
rect 14277 8959 14335 8965
rect 14277 8925 14289 8959
rect 14323 8925 14335 8959
rect 14277 8919 14335 8925
rect 14369 8959 14427 8965
rect 14369 8925 14381 8959
rect 14415 8925 14427 8959
rect 14369 8919 14427 8925
rect 14461 8959 14519 8965
rect 14461 8925 14473 8959
rect 14507 8956 14519 8959
rect 15010 8956 15016 8968
rect 14507 8928 15016 8956
rect 14507 8925 14519 8928
rect 14461 8919 14519 8925
rect 12805 8891 12863 8897
rect 12805 8857 12817 8891
rect 12851 8888 12863 8891
rect 14292 8888 14320 8919
rect 12851 8860 14320 8888
rect 12851 8857 12863 8860
rect 12805 8851 12863 8857
rect 11054 8820 11060 8832
rect 8864 8792 11060 8820
rect 11054 8780 11060 8792
rect 11112 8780 11118 8832
rect 12986 8780 12992 8832
rect 13044 8780 13050 8832
rect 13446 8780 13452 8832
rect 13504 8780 13510 8832
rect 13906 8780 13912 8832
rect 13964 8820 13970 8832
rect 14384 8820 14412 8919
rect 15010 8916 15016 8928
rect 15068 8916 15074 8968
rect 15286 8916 15292 8968
rect 15344 8916 15350 8968
rect 13964 8792 14412 8820
rect 13964 8780 13970 8792
rect 14734 8780 14740 8832
rect 14792 8780 14798 8832
rect 14918 8780 14924 8832
rect 14976 8780 14982 8832
rect 15396 8820 15424 8984
rect 19996 8968 20024 8996
rect 20717 8993 20729 8996
rect 20763 8993 20775 9027
rect 20717 8987 20775 8993
rect 22186 8984 22192 9036
rect 22244 8984 22250 9036
rect 22649 9027 22707 9033
rect 22649 9024 22661 9027
rect 22388 8996 22661 9024
rect 22388 8968 22416 8996
rect 22649 8993 22661 8996
rect 22695 8993 22707 9027
rect 22649 8987 22707 8993
rect 15746 8916 15752 8968
rect 15804 8916 15810 8968
rect 17957 8959 18015 8965
rect 17957 8956 17969 8959
rect 17328 8928 17969 8956
rect 16022 8848 16028 8900
rect 16080 8848 16086 8900
rect 16758 8848 16764 8900
rect 16816 8848 16822 8900
rect 17328 8820 17356 8928
rect 17957 8925 17969 8928
rect 18003 8925 18015 8959
rect 17957 8919 18015 8925
rect 18138 8916 18144 8968
rect 18196 8956 18202 8968
rect 18509 8959 18567 8965
rect 18509 8956 18521 8959
rect 18196 8928 18521 8956
rect 18196 8916 18202 8928
rect 18509 8925 18521 8928
rect 18555 8925 18567 8959
rect 18509 8919 18567 8925
rect 19518 8916 19524 8968
rect 19576 8956 19582 8968
rect 19705 8959 19763 8965
rect 19705 8956 19717 8959
rect 19576 8928 19717 8956
rect 19576 8916 19582 8928
rect 19705 8925 19717 8928
rect 19751 8956 19763 8959
rect 19751 8928 19840 8956
rect 19751 8925 19763 8928
rect 19705 8919 19763 8925
rect 15396 8792 17356 8820
rect 19521 8823 19579 8829
rect 19521 8789 19533 8823
rect 19567 8820 19579 8823
rect 19702 8820 19708 8832
rect 19567 8792 19708 8820
rect 19567 8789 19579 8792
rect 19521 8783 19579 8789
rect 19702 8780 19708 8792
rect 19760 8780 19766 8832
rect 19812 8820 19840 8928
rect 19978 8916 19984 8968
rect 20036 8916 20042 8968
rect 20070 8916 20076 8968
rect 20128 8956 20134 8968
rect 20625 8959 20683 8965
rect 20625 8956 20637 8959
rect 20128 8928 20637 8956
rect 20128 8916 20134 8928
rect 20625 8925 20637 8928
rect 20671 8925 20683 8959
rect 20625 8919 20683 8925
rect 22370 8916 22376 8968
rect 22428 8916 22434 8968
rect 22554 8916 22560 8968
rect 22612 8916 22618 8968
rect 19886 8848 19892 8900
rect 19944 8888 19950 8900
rect 20088 8888 20116 8916
rect 19944 8860 20116 8888
rect 19944 8848 19950 8860
rect 20254 8848 20260 8900
rect 20312 8848 20318 8900
rect 22278 8848 22284 8900
rect 22336 8848 22342 8900
rect 22664 8888 22692 8987
rect 22848 8956 22876 9055
rect 22922 9052 22928 9104
rect 22980 9052 22986 9104
rect 23106 9052 23112 9104
rect 23164 9092 23170 9104
rect 23566 9092 23572 9104
rect 23164 9064 23572 9092
rect 23164 9052 23170 9064
rect 23566 9052 23572 9064
rect 23624 9092 23630 9104
rect 23624 9064 24440 9092
rect 23624 9052 23630 9064
rect 22940 9024 22968 9052
rect 22940 8996 23704 9024
rect 22925 8959 22983 8965
rect 22925 8956 22937 8959
rect 22848 8928 22937 8956
rect 22925 8925 22937 8928
rect 22971 8925 22983 8959
rect 22925 8919 22983 8925
rect 23014 8916 23020 8968
rect 23072 8956 23078 8968
rect 23216 8965 23244 8996
rect 23201 8959 23259 8965
rect 23072 8928 23117 8956
rect 23072 8916 23078 8928
rect 23201 8925 23213 8959
rect 23247 8925 23259 8959
rect 23201 8919 23259 8925
rect 23382 8916 23388 8968
rect 23440 8965 23446 8968
rect 23440 8956 23448 8965
rect 23440 8928 23485 8956
rect 23440 8919 23448 8928
rect 23440 8916 23446 8919
rect 23290 8888 23296 8900
rect 22664 8860 23296 8888
rect 23290 8848 23296 8860
rect 23348 8848 23354 8900
rect 20272 8820 20300 8848
rect 19812 8792 20300 8820
rect 23566 8780 23572 8832
rect 23624 8780 23630 8832
rect 23676 8820 23704 8996
rect 24210 8984 24216 9036
rect 24268 8984 24274 9036
rect 23845 8959 23903 8965
rect 23845 8925 23857 8959
rect 23891 8956 23903 8959
rect 24228 8956 24256 8984
rect 24412 8965 24440 9064
rect 24670 9052 24676 9104
rect 24728 9092 24734 9104
rect 26160 9092 26188 9132
rect 26326 9120 26332 9172
rect 26384 9160 26390 9172
rect 29365 9163 29423 9169
rect 26384 9132 27614 9160
rect 26384 9120 26390 9132
rect 26970 9092 26976 9104
rect 24728 9064 25636 9092
rect 24728 9052 24734 9064
rect 25314 8984 25320 9036
rect 25372 8984 25378 9036
rect 23891 8928 24256 8956
rect 24397 8959 24455 8965
rect 23891 8925 23903 8928
rect 23845 8919 23903 8925
rect 24397 8925 24409 8959
rect 24443 8925 24455 8959
rect 24397 8919 24455 8925
rect 24490 8959 24548 8965
rect 24490 8925 24502 8959
rect 24536 8925 24548 8959
rect 24490 8919 24548 8925
rect 24504 8888 24532 8919
rect 24854 8916 24860 8968
rect 24912 8965 24918 8968
rect 24912 8959 24939 8965
rect 24927 8925 24939 8959
rect 24912 8919 24939 8925
rect 24912 8916 24918 8919
rect 25038 8916 25044 8968
rect 25096 8956 25102 8968
rect 25608 8965 25636 9064
rect 26160 9064 26976 9092
rect 25777 9027 25835 9033
rect 25777 8993 25789 9027
rect 25823 9024 25835 9027
rect 25823 8996 26096 9024
rect 25823 8993 25835 8996
rect 25777 8987 25835 8993
rect 25225 8959 25283 8965
rect 25225 8956 25237 8959
rect 25096 8928 25237 8956
rect 25096 8916 25102 8928
rect 25225 8925 25237 8928
rect 25271 8925 25283 8959
rect 25501 8959 25559 8965
rect 25501 8956 25513 8959
rect 25225 8919 25283 8925
rect 25424 8928 25513 8956
rect 24578 8888 24584 8900
rect 24504 8860 24584 8888
rect 24578 8848 24584 8860
rect 24636 8848 24642 8900
rect 24673 8891 24731 8897
rect 24673 8857 24685 8891
rect 24719 8857 24731 8891
rect 24673 8851 24731 8857
rect 24765 8891 24823 8897
rect 24765 8857 24777 8891
rect 24811 8888 24823 8891
rect 25056 8888 25084 8916
rect 25424 8900 25452 8928
rect 25501 8925 25513 8928
rect 25547 8925 25559 8959
rect 25501 8919 25559 8925
rect 25593 8959 25651 8965
rect 25593 8925 25605 8959
rect 25639 8925 25651 8959
rect 25593 8919 25651 8925
rect 25869 8959 25927 8965
rect 25869 8925 25881 8959
rect 25915 8956 25927 8959
rect 25958 8956 25964 8968
rect 25915 8928 25964 8956
rect 25915 8925 25927 8928
rect 25869 8919 25927 8925
rect 25958 8916 25964 8928
rect 26016 8916 26022 8968
rect 26068 8965 26096 8996
rect 26160 8965 26188 9064
rect 26970 9052 26976 9064
rect 27028 9052 27034 9104
rect 27062 9052 27068 9104
rect 27120 9092 27126 9104
rect 27586 9092 27614 9132
rect 29365 9129 29377 9163
rect 29411 9160 29423 9163
rect 29638 9160 29644 9172
rect 29411 9132 29644 9160
rect 29411 9129 29423 9132
rect 29365 9123 29423 9129
rect 29178 9092 29184 9104
rect 27120 9064 27200 9092
rect 27586 9064 29184 9092
rect 27120 9052 27126 9064
rect 26878 9024 26884 9036
rect 26804 8996 26884 9024
rect 26053 8959 26111 8965
rect 26053 8925 26065 8959
rect 26099 8925 26111 8959
rect 26053 8919 26111 8925
rect 26145 8959 26203 8965
rect 26145 8925 26157 8959
rect 26191 8925 26203 8959
rect 26145 8919 26203 8925
rect 26237 8959 26295 8965
rect 26237 8925 26249 8959
rect 26283 8956 26295 8959
rect 26510 8956 26516 8968
rect 26283 8928 26516 8956
rect 26283 8925 26295 8928
rect 26237 8919 26295 8925
rect 26510 8916 26516 8928
rect 26568 8916 26574 8968
rect 26804 8965 26832 8996
rect 26878 8984 26884 8996
rect 26936 8984 26942 9036
rect 27172 9024 27200 9064
rect 27985 9027 28043 9033
rect 27985 9024 27997 9027
rect 27172 8996 27997 9024
rect 27985 8993 27997 8996
rect 28031 8993 28043 9027
rect 27985 8987 28043 8993
rect 28074 8984 28080 9036
rect 28132 9024 28138 9036
rect 28132 8996 28212 9024
rect 28132 8984 28138 8996
rect 26789 8959 26847 8965
rect 26789 8925 26801 8959
rect 26835 8925 26847 8959
rect 26789 8919 26847 8925
rect 26973 8959 27031 8965
rect 26973 8925 26985 8959
rect 27019 8925 27031 8959
rect 26973 8919 27031 8925
rect 27065 8959 27123 8965
rect 27065 8925 27077 8959
rect 27111 8925 27123 8959
rect 27065 8919 27123 8925
rect 27157 8959 27215 8965
rect 27157 8925 27169 8959
rect 27203 8925 27215 8959
rect 27157 8919 27215 8925
rect 24811 8860 25360 8888
rect 24811 8857 24823 8860
rect 24765 8851 24823 8857
rect 24688 8820 24716 8851
rect 23676 8792 24716 8820
rect 25041 8823 25099 8829
rect 25041 8789 25053 8823
rect 25087 8820 25099 8823
rect 25130 8820 25136 8832
rect 25087 8792 25136 8820
rect 25087 8789 25099 8792
rect 25041 8783 25099 8789
rect 25130 8780 25136 8792
rect 25188 8780 25194 8832
rect 25332 8820 25360 8860
rect 25406 8848 25412 8900
rect 25464 8848 25470 8900
rect 26528 8888 26556 8916
rect 26528 8860 26832 8888
rect 26326 8820 26332 8832
rect 25332 8792 26332 8820
rect 26326 8780 26332 8792
rect 26384 8780 26390 8832
rect 26510 8780 26516 8832
rect 26568 8780 26574 8832
rect 26804 8820 26832 8860
rect 26878 8848 26884 8900
rect 26936 8888 26942 8900
rect 26988 8888 27016 8919
rect 26936 8860 27016 8888
rect 26936 8848 26942 8860
rect 27080 8820 27108 8919
rect 27172 8832 27200 8919
rect 27246 8916 27252 8968
rect 27304 8956 27310 8968
rect 27341 8959 27399 8965
rect 27341 8956 27353 8959
rect 27304 8928 27353 8956
rect 27304 8916 27310 8928
rect 27341 8925 27353 8928
rect 27387 8925 27399 8959
rect 27341 8919 27399 8925
rect 27614 8916 27620 8968
rect 27672 8916 27678 8968
rect 28184 8965 28212 8996
rect 28169 8959 28227 8965
rect 28169 8925 28181 8959
rect 28215 8925 28227 8959
rect 28169 8919 28227 8925
rect 28353 8959 28411 8965
rect 28353 8925 28365 8959
rect 28399 8925 28411 8959
rect 28353 8919 28411 8925
rect 27706 8848 27712 8900
rect 27764 8888 27770 8900
rect 27801 8891 27859 8897
rect 27801 8888 27813 8891
rect 27764 8860 27813 8888
rect 27764 8848 27770 8860
rect 27801 8857 27813 8860
rect 27847 8857 27859 8891
rect 28368 8888 28396 8919
rect 28442 8916 28448 8968
rect 28500 8916 28506 8968
rect 28920 8965 28948 9064
rect 29178 9052 29184 9064
rect 29236 9052 29242 9104
rect 29270 9024 29276 9036
rect 29104 8996 29276 9024
rect 29104 8965 29132 8996
rect 29270 8984 29276 8996
rect 29328 8984 29334 9036
rect 29564 8965 29592 9132
rect 29638 9120 29644 9132
rect 29696 9120 29702 9172
rect 29730 9120 29736 9172
rect 29788 9160 29794 9172
rect 29788 9132 30512 9160
rect 29788 9120 29794 9132
rect 29917 9095 29975 9101
rect 29917 9061 29929 9095
rect 29963 9061 29975 9095
rect 29917 9055 29975 9061
rect 28537 8959 28595 8965
rect 28537 8925 28549 8959
rect 28583 8925 28595 8959
rect 28537 8919 28595 8925
rect 28905 8959 28963 8965
rect 28905 8925 28917 8959
rect 28951 8925 28963 8959
rect 28905 8919 28963 8925
rect 29089 8959 29147 8965
rect 29089 8925 29101 8959
rect 29135 8925 29147 8959
rect 29089 8919 29147 8925
rect 29181 8959 29239 8965
rect 29181 8925 29193 8959
rect 29227 8925 29239 8959
rect 29181 8919 29239 8925
rect 29365 8959 29423 8965
rect 29365 8925 29377 8959
rect 29411 8925 29423 8959
rect 29365 8919 29423 8925
rect 29549 8959 29607 8965
rect 29549 8925 29561 8959
rect 29595 8925 29607 8959
rect 29549 8919 29607 8925
rect 29641 8959 29699 8965
rect 29641 8925 29653 8959
rect 29687 8925 29699 8959
rect 29932 8956 29960 9055
rect 30009 8959 30067 8965
rect 30009 8956 30021 8959
rect 29932 8928 30021 8956
rect 29641 8919 29699 8925
rect 30009 8925 30021 8928
rect 30055 8925 30067 8959
rect 30009 8919 30067 8925
rect 27801 8851 27859 8857
rect 27908 8860 28396 8888
rect 28552 8888 28580 8919
rect 29196 8888 29224 8919
rect 28552 8860 28948 8888
rect 26804 8792 27108 8820
rect 27154 8780 27160 8832
rect 27212 8780 27218 8832
rect 27525 8823 27583 8829
rect 27525 8789 27537 8823
rect 27571 8820 27583 8823
rect 27908 8820 27936 8860
rect 28920 8832 28948 8860
rect 29012 8860 29224 8888
rect 29012 8832 29040 8860
rect 29270 8848 29276 8900
rect 29328 8888 29334 8900
rect 29380 8888 29408 8919
rect 29328 8860 29408 8888
rect 29328 8848 29334 8860
rect 27571 8792 27936 8820
rect 27571 8789 27583 8792
rect 27525 8783 27583 8789
rect 28810 8780 28816 8832
rect 28868 8780 28874 8832
rect 28902 8780 28908 8832
rect 28960 8780 28966 8832
rect 28994 8780 29000 8832
rect 29052 8780 29058 8832
rect 29086 8780 29092 8832
rect 29144 8820 29150 8832
rect 29656 8820 29684 8919
rect 30190 8916 30196 8968
rect 30248 8916 30254 8968
rect 30374 8848 30380 8900
rect 30432 8848 30438 8900
rect 30484 8888 30512 9132
rect 30742 9120 30748 9172
rect 30800 9120 30806 9172
rect 31570 9120 31576 9172
rect 31628 9160 31634 9172
rect 31757 9163 31815 9169
rect 31757 9160 31769 9163
rect 31628 9132 31769 9160
rect 31628 9120 31634 9132
rect 31757 9129 31769 9132
rect 31803 9129 31815 9163
rect 31757 9123 31815 9129
rect 32861 9163 32919 9169
rect 32861 9129 32873 9163
rect 32907 9160 32919 9163
rect 33134 9160 33140 9172
rect 32907 9132 33140 9160
rect 32907 9129 32919 9132
rect 32861 9123 32919 9129
rect 33134 9120 33140 9132
rect 33192 9120 33198 9172
rect 33229 9163 33287 9169
rect 33229 9129 33241 9163
rect 33275 9160 33287 9163
rect 33318 9160 33324 9172
rect 33275 9132 33324 9160
rect 33275 9129 33287 9132
rect 33229 9123 33287 9129
rect 33318 9120 33324 9132
rect 33376 9120 33382 9172
rect 30760 9092 30788 9120
rect 32401 9095 32459 9101
rect 32401 9092 32413 9095
rect 30760 9064 32413 9092
rect 32401 9061 32413 9064
rect 32447 9061 32459 9095
rect 32401 9055 32459 9061
rect 31481 9027 31539 9033
rect 31481 8993 31493 9027
rect 31527 9024 31539 9027
rect 32030 9024 32036 9036
rect 31527 8996 32036 9024
rect 31527 8993 31539 8996
rect 31481 8987 31539 8993
rect 32030 8984 32036 8996
rect 32088 8984 32094 9036
rect 31573 8959 31631 8965
rect 31573 8925 31585 8959
rect 31619 8956 31631 8959
rect 31754 8956 31760 8968
rect 31619 8928 31760 8956
rect 31619 8925 31631 8928
rect 31573 8919 31631 8925
rect 31754 8916 31760 8928
rect 31812 8916 31818 8968
rect 31846 8916 31852 8968
rect 31904 8916 31910 8968
rect 32125 8959 32183 8965
rect 32125 8925 32137 8959
rect 32171 8956 32183 8959
rect 32585 8959 32643 8965
rect 32171 8928 32536 8956
rect 32171 8925 32183 8928
rect 32125 8919 32183 8925
rect 32140 8888 32168 8919
rect 30484 8860 32168 8888
rect 29144 8792 29684 8820
rect 29144 8780 29150 8792
rect 30834 8780 30840 8832
rect 30892 8820 30898 8832
rect 31113 8823 31171 8829
rect 31113 8820 31125 8823
rect 30892 8792 31125 8820
rect 30892 8780 30898 8792
rect 31113 8789 31125 8792
rect 31159 8789 31171 8823
rect 31113 8783 31171 8789
rect 31938 8780 31944 8832
rect 31996 8780 32002 8832
rect 32508 8820 32536 8928
rect 32585 8925 32597 8959
rect 32631 8925 32643 8959
rect 32585 8919 32643 8925
rect 32677 8959 32735 8965
rect 32677 8925 32689 8959
rect 32723 8956 32735 8959
rect 32766 8956 32772 8968
rect 32723 8928 32772 8956
rect 32723 8925 32735 8928
rect 32677 8919 32735 8925
rect 32600 8888 32628 8919
rect 32766 8916 32772 8928
rect 32824 8916 32830 8968
rect 32953 8959 33011 8965
rect 32953 8925 32965 8959
rect 32999 8925 33011 8959
rect 32953 8919 33011 8925
rect 32858 8888 32864 8900
rect 32600 8860 32864 8888
rect 32858 8848 32864 8860
rect 32916 8848 32922 8900
rect 32968 8888 32996 8919
rect 33042 8916 33048 8968
rect 33100 8916 33106 8968
rect 33134 8916 33140 8968
rect 33192 8916 33198 8968
rect 33229 8959 33287 8965
rect 33229 8925 33241 8959
rect 33275 8925 33287 8959
rect 33229 8919 33287 8925
rect 33152 8888 33180 8916
rect 32968 8860 33180 8888
rect 33244 8832 33272 8919
rect 33502 8916 33508 8968
rect 33560 8916 33566 8968
rect 37921 8959 37979 8965
rect 37921 8925 37933 8959
rect 37967 8956 37979 8959
rect 38286 8956 38292 8968
rect 37967 8928 38292 8956
rect 37967 8925 37979 8928
rect 37921 8919 37979 8925
rect 38286 8916 38292 8928
rect 38344 8916 38350 8968
rect 35986 8848 35992 8900
rect 36044 8888 36050 8900
rect 36814 8888 36820 8900
rect 36044 8860 36820 8888
rect 36044 8848 36050 8860
rect 36814 8848 36820 8860
rect 36872 8888 36878 8900
rect 37645 8891 37703 8897
rect 37645 8888 37657 8891
rect 36872 8860 37657 8888
rect 36872 8848 36878 8860
rect 37645 8857 37657 8860
rect 37691 8857 37703 8891
rect 37645 8851 37703 8857
rect 33226 8820 33232 8832
rect 32508 8792 33232 8820
rect 33226 8780 33232 8792
rect 33284 8780 33290 8832
rect 1104 8730 38272 8752
rect 1104 8678 4874 8730
rect 4926 8678 4938 8730
rect 4990 8678 5002 8730
rect 5054 8678 5066 8730
rect 5118 8678 5130 8730
rect 5182 8678 35594 8730
rect 35646 8678 35658 8730
rect 35710 8678 35722 8730
rect 35774 8678 35786 8730
rect 35838 8678 35850 8730
rect 35902 8678 38272 8730
rect 1104 8656 38272 8678
rect 4249 8619 4307 8625
rect 4249 8585 4261 8619
rect 4295 8616 4307 8619
rect 5077 8619 5135 8625
rect 5077 8616 5089 8619
rect 4295 8588 5089 8616
rect 4295 8585 4307 8588
rect 4249 8579 4307 8585
rect 5077 8585 5089 8588
rect 5123 8585 5135 8619
rect 5077 8579 5135 8585
rect 5920 8588 6592 8616
rect 5920 8557 5948 8588
rect 5905 8551 5963 8557
rect 5905 8548 5917 8551
rect 4724 8520 5917 8548
rect 4724 8492 4752 8520
rect 5905 8517 5917 8520
rect 5951 8517 5963 8551
rect 5905 8511 5963 8517
rect 5994 8508 6000 8560
rect 6052 8548 6058 8560
rect 6564 8557 6592 8588
rect 7098 8576 7104 8628
rect 7156 8616 7162 8628
rect 9214 8616 9220 8628
rect 7156 8588 9220 8616
rect 7156 8576 7162 8588
rect 9214 8576 9220 8588
rect 9272 8576 9278 8628
rect 9309 8619 9367 8625
rect 9309 8585 9321 8619
rect 9355 8616 9367 8619
rect 9398 8616 9404 8628
rect 9355 8588 9404 8616
rect 9355 8585 9367 8588
rect 9309 8579 9367 8585
rect 9398 8576 9404 8588
rect 9456 8616 9462 8628
rect 9858 8616 9864 8628
rect 9456 8588 9864 8616
rect 9456 8576 9462 8588
rect 9858 8576 9864 8588
rect 9916 8576 9922 8628
rect 10045 8619 10103 8625
rect 10045 8585 10057 8619
rect 10091 8616 10103 8619
rect 10134 8616 10140 8628
rect 10091 8588 10140 8616
rect 10091 8585 10103 8588
rect 10045 8579 10103 8585
rect 10134 8576 10140 8588
rect 10192 8576 10198 8628
rect 10597 8619 10655 8625
rect 10597 8585 10609 8619
rect 10643 8616 10655 8619
rect 12710 8616 12716 8628
rect 10643 8588 12716 8616
rect 10643 8585 10655 8588
rect 10597 8579 10655 8585
rect 6533 8551 6592 8557
rect 6052 8520 6500 8548
rect 6052 8508 6058 8520
rect 3421 8483 3479 8489
rect 3421 8449 3433 8483
rect 3467 8480 3479 8483
rect 4157 8483 4215 8489
rect 3467 8452 3832 8480
rect 3467 8449 3479 8452
rect 3421 8443 3479 8449
rect 3804 8353 3832 8452
rect 4157 8449 4169 8483
rect 4203 8480 4215 8483
rect 4706 8480 4712 8492
rect 4203 8452 4712 8480
rect 4203 8449 4215 8452
rect 4157 8443 4215 8449
rect 4706 8440 4712 8452
rect 4764 8440 4770 8492
rect 6104 8489 6132 8520
rect 5445 8483 5503 8489
rect 5445 8449 5457 8483
rect 5491 8480 5503 8483
rect 6089 8483 6147 8489
rect 5491 8452 6040 8480
rect 5491 8449 5503 8452
rect 5445 8443 5503 8449
rect 4433 8415 4491 8421
rect 4433 8381 4445 8415
rect 4479 8412 4491 8415
rect 4479 8384 4752 8412
rect 4479 8381 4491 8384
rect 4433 8375 4491 8381
rect 3789 8347 3847 8353
rect 3789 8313 3801 8347
rect 3835 8313 3847 8347
rect 3789 8307 3847 8313
rect 4062 8304 4068 8356
rect 4120 8344 4126 8356
rect 4724 8344 4752 8384
rect 5534 8372 5540 8424
rect 5592 8372 5598 8424
rect 5626 8372 5632 8424
rect 5684 8372 5690 8424
rect 5718 8372 5724 8424
rect 5776 8372 5782 8424
rect 6012 8412 6040 8452
rect 6089 8449 6101 8483
rect 6135 8449 6147 8483
rect 6089 8443 6147 8449
rect 6181 8483 6239 8489
rect 6181 8449 6193 8483
rect 6227 8480 6239 8483
rect 6270 8480 6276 8492
rect 6227 8452 6276 8480
rect 6227 8449 6239 8452
rect 6181 8443 6239 8449
rect 6270 8440 6276 8452
rect 6328 8440 6334 8492
rect 6472 8480 6500 8520
rect 6533 8517 6545 8551
rect 6579 8520 6592 8551
rect 6733 8551 6791 8557
rect 6579 8517 6591 8520
rect 6533 8511 6591 8517
rect 6733 8517 6745 8551
rect 6779 8517 6791 8551
rect 6733 8511 6791 8517
rect 7837 8551 7895 8557
rect 7837 8517 7849 8551
rect 7883 8548 7895 8551
rect 9582 8548 9588 8560
rect 7883 8520 9588 8548
rect 7883 8517 7895 8520
rect 7837 8511 7895 8517
rect 6748 8480 6776 8511
rect 9582 8508 9588 8520
rect 9640 8508 9646 8560
rect 10612 8548 10640 8579
rect 12710 8576 12716 8588
rect 12768 8576 12774 8628
rect 12986 8576 12992 8628
rect 13044 8576 13050 8628
rect 13357 8619 13415 8625
rect 13357 8585 13369 8619
rect 13403 8585 13415 8619
rect 13357 8579 13415 8585
rect 12437 8551 12495 8557
rect 12437 8548 12449 8551
rect 10152 8520 10640 8548
rect 11992 8520 12449 8548
rect 6472 8452 6776 8480
rect 8662 8440 8668 8492
rect 8720 8480 8726 8492
rect 10152 8489 10180 8520
rect 10137 8483 10195 8489
rect 8720 8452 9904 8480
rect 8720 8440 8726 8452
rect 9876 8412 9904 8452
rect 10137 8449 10149 8483
rect 10183 8449 10195 8483
rect 10505 8483 10563 8489
rect 10505 8480 10517 8483
rect 10137 8443 10195 8449
rect 10244 8452 10517 8480
rect 10244 8412 10272 8452
rect 10505 8449 10517 8452
rect 10551 8449 10563 8483
rect 10505 8443 10563 8449
rect 11146 8440 11152 8492
rect 11204 8480 11210 8492
rect 11517 8483 11575 8489
rect 11517 8480 11529 8483
rect 11204 8452 11529 8480
rect 11204 8440 11210 8452
rect 11517 8449 11529 8452
rect 11563 8449 11575 8483
rect 11517 8443 11575 8449
rect 11790 8440 11796 8492
rect 11848 8480 11854 8492
rect 11992 8489 12020 8520
rect 12437 8517 12449 8520
rect 12483 8517 12495 8551
rect 12437 8511 12495 8517
rect 12618 8508 12624 8560
rect 12676 8508 12682 8560
rect 13004 8548 13032 8576
rect 13372 8548 13400 8579
rect 13446 8576 13452 8628
rect 13504 8616 13510 8628
rect 15197 8619 15255 8625
rect 15197 8616 15209 8619
rect 13504 8588 15209 8616
rect 13504 8576 13510 8588
rect 15197 8585 15209 8588
rect 15243 8616 15255 8619
rect 18414 8616 18420 8628
rect 15243 8588 18420 8616
rect 15243 8585 15255 8588
rect 15197 8579 15255 8585
rect 18414 8576 18420 8588
rect 18472 8576 18478 8628
rect 18877 8619 18935 8625
rect 18877 8585 18889 8619
rect 18923 8616 18935 8619
rect 22370 8616 22376 8628
rect 18923 8588 22376 8616
rect 18923 8585 18935 8588
rect 18877 8579 18935 8585
rect 22370 8576 22376 8588
rect 22428 8576 22434 8628
rect 23566 8576 23572 8628
rect 23624 8576 23630 8628
rect 24302 8576 24308 8628
rect 24360 8616 24366 8628
rect 24949 8619 25007 8625
rect 24949 8616 24961 8619
rect 24360 8588 24961 8616
rect 24360 8576 24366 8588
rect 24949 8585 24961 8588
rect 24995 8616 25007 8619
rect 24995 8588 26464 8616
rect 24995 8585 25007 8588
rect 24949 8579 25007 8585
rect 13725 8551 13783 8557
rect 13725 8548 13737 8551
rect 13004 8520 13216 8548
rect 13372 8520 13737 8548
rect 11977 8483 12035 8489
rect 11977 8480 11989 8483
rect 11848 8452 11989 8480
rect 11848 8440 11854 8452
rect 11977 8449 11989 8452
rect 12023 8449 12035 8483
rect 11977 8443 12035 8449
rect 12342 8440 12348 8492
rect 12400 8440 12406 8492
rect 12526 8440 12532 8492
rect 12584 8440 12590 8492
rect 12986 8440 12992 8492
rect 13044 8440 13050 8492
rect 13188 8489 13216 8520
rect 13725 8517 13737 8520
rect 13771 8517 13783 8551
rect 13725 8511 13783 8517
rect 15010 8508 15016 8560
rect 15068 8548 15074 8560
rect 15068 8520 18736 8548
rect 15068 8508 15074 8520
rect 13173 8483 13231 8489
rect 13173 8449 13185 8483
rect 13219 8449 13231 8483
rect 16758 8480 16764 8492
rect 14858 8452 16764 8480
rect 13173 8443 13231 8449
rect 16758 8440 16764 8452
rect 16816 8440 16822 8492
rect 17126 8440 17132 8492
rect 17184 8440 17190 8492
rect 17402 8440 17408 8492
rect 17460 8440 17466 8492
rect 6012 8384 9812 8412
rect 9876 8384 10272 8412
rect 10321 8415 10379 8421
rect 5644 8344 5672 8372
rect 4120 8316 4660 8344
rect 4724 8316 5672 8344
rect 4120 8304 4126 8316
rect 4632 8288 4660 8316
rect 5902 8304 5908 8356
rect 5960 8304 5966 8356
rect 6365 8347 6423 8353
rect 6365 8313 6377 8347
rect 6411 8344 6423 8347
rect 6454 8344 6460 8356
rect 6411 8316 6460 8344
rect 6411 8313 6423 8316
rect 6365 8307 6423 8313
rect 6454 8304 6460 8316
rect 6512 8304 6518 8356
rect 8478 8304 8484 8356
rect 8536 8344 8542 8356
rect 9677 8347 9735 8353
rect 9677 8344 9689 8347
rect 8536 8316 9689 8344
rect 8536 8304 8542 8316
rect 9677 8313 9689 8316
rect 9723 8313 9735 8347
rect 9784 8344 9812 8384
rect 10321 8381 10333 8415
rect 10367 8412 10379 8415
rect 10410 8412 10416 8424
rect 10367 8384 10416 8412
rect 10367 8381 10379 8384
rect 10321 8375 10379 8381
rect 10410 8372 10416 8384
rect 10468 8372 10474 8424
rect 10594 8372 10600 8424
rect 10652 8412 10658 8424
rect 11885 8415 11943 8421
rect 11885 8412 11897 8415
rect 10652 8384 11897 8412
rect 10652 8372 10658 8384
rect 11885 8381 11897 8384
rect 11931 8381 11943 8415
rect 11885 8375 11943 8381
rect 12250 8372 12256 8424
rect 12308 8412 12314 8424
rect 13449 8415 13507 8421
rect 13449 8412 13461 8415
rect 12308 8384 13461 8412
rect 12308 8372 12314 8384
rect 13449 8381 13461 8384
rect 13495 8381 13507 8415
rect 14918 8412 14924 8424
rect 13449 8375 13507 8381
rect 13556 8384 14924 8412
rect 13556 8344 13584 8384
rect 14918 8372 14924 8384
rect 14976 8372 14982 8424
rect 17144 8412 17172 8440
rect 17589 8415 17647 8421
rect 17589 8412 17601 8415
rect 17144 8384 17601 8412
rect 17589 8381 17601 8384
rect 17635 8381 17647 8415
rect 18708 8412 18736 8520
rect 18800 8520 19196 8548
rect 18800 8489 18828 8520
rect 19168 8492 19196 8520
rect 19518 8508 19524 8560
rect 19576 8508 19582 8560
rect 19705 8551 19763 8557
rect 19705 8517 19717 8551
rect 19751 8548 19763 8551
rect 19886 8548 19892 8560
rect 19751 8520 19892 8548
rect 19751 8517 19763 8520
rect 19705 8511 19763 8517
rect 19886 8508 19892 8520
rect 19944 8508 19950 8560
rect 19978 8508 19984 8560
rect 20036 8508 20042 8560
rect 21450 8508 21456 8560
rect 21508 8548 21514 8560
rect 22097 8551 22155 8557
rect 22097 8548 22109 8551
rect 21508 8520 22109 8548
rect 21508 8508 21514 8520
rect 22097 8517 22109 8520
rect 22143 8517 22155 8551
rect 23584 8548 23612 8576
rect 22097 8511 22155 8517
rect 23216 8520 23612 8548
rect 24857 8551 24915 8557
rect 18785 8483 18843 8489
rect 18785 8449 18797 8483
rect 18831 8449 18843 8483
rect 18785 8443 18843 8449
rect 18966 8440 18972 8492
rect 19024 8440 19030 8492
rect 19150 8440 19156 8492
rect 19208 8440 19214 8492
rect 19797 8483 19855 8489
rect 19797 8449 19809 8483
rect 19843 8480 19855 8483
rect 19996 8480 20024 8508
rect 19843 8452 20024 8480
rect 19843 8449 19855 8452
rect 19797 8443 19855 8449
rect 20806 8440 20812 8492
rect 20864 8480 20870 8492
rect 21818 8480 21824 8492
rect 20864 8452 21824 8480
rect 20864 8440 20870 8452
rect 21818 8440 21824 8452
rect 21876 8440 21882 8492
rect 21913 8483 21971 8489
rect 21913 8449 21925 8483
rect 21959 8480 21971 8483
rect 22002 8480 22008 8492
rect 21959 8452 22008 8480
rect 21959 8449 21971 8452
rect 21913 8443 21971 8449
rect 22002 8440 22008 8452
rect 22060 8440 22066 8492
rect 23216 8489 23244 8520
rect 24857 8517 24869 8551
rect 24903 8548 24915 8551
rect 25314 8548 25320 8560
rect 24903 8520 25320 8548
rect 24903 8517 24915 8520
rect 24857 8511 24915 8517
rect 25314 8508 25320 8520
rect 25372 8508 25378 8560
rect 26436 8548 26464 8588
rect 28902 8576 28908 8628
rect 28960 8616 28966 8628
rect 29273 8619 29331 8625
rect 28960 8588 29132 8616
rect 28960 8576 28966 8588
rect 26878 8548 26884 8560
rect 26436 8520 26884 8548
rect 26878 8508 26884 8520
rect 26936 8548 26942 8560
rect 28994 8548 29000 8560
rect 26936 8520 27200 8548
rect 26936 8508 26942 8520
rect 23201 8483 23259 8489
rect 23201 8449 23213 8483
rect 23247 8449 23259 8483
rect 23201 8443 23259 8449
rect 23477 8483 23535 8489
rect 23477 8449 23489 8483
rect 23523 8480 23535 8483
rect 23566 8480 23572 8492
rect 23523 8452 23572 8480
rect 23523 8449 23535 8452
rect 23477 8443 23535 8449
rect 23566 8440 23572 8452
rect 23624 8440 23630 8492
rect 23661 8483 23719 8489
rect 23661 8449 23673 8483
rect 23707 8480 23719 8483
rect 24210 8480 24216 8492
rect 23707 8452 24216 8480
rect 23707 8449 23719 8452
rect 23661 8443 23719 8449
rect 24210 8440 24216 8452
rect 24268 8440 24274 8492
rect 25406 8480 25412 8492
rect 24780 8452 25412 8480
rect 21542 8412 21548 8424
rect 18708 8384 21548 8412
rect 17589 8375 17647 8381
rect 21542 8372 21548 8384
rect 21600 8372 21606 8424
rect 24780 8421 24808 8452
rect 25406 8440 25412 8452
rect 25464 8440 25470 8492
rect 26510 8440 26516 8492
rect 26568 8480 26574 8492
rect 27172 8489 27200 8520
rect 27264 8520 29000 8548
rect 27264 8489 27292 8520
rect 28994 8508 29000 8520
rect 29052 8508 29058 8560
rect 29104 8548 29132 8588
rect 29273 8585 29285 8619
rect 29319 8616 29331 8619
rect 30190 8616 30196 8628
rect 29319 8588 30196 8616
rect 29319 8585 29331 8588
rect 29273 8579 29331 8585
rect 30190 8576 30196 8588
rect 30248 8576 30254 8628
rect 31297 8619 31355 8625
rect 31297 8585 31309 8619
rect 31343 8616 31355 8619
rect 31386 8616 31392 8628
rect 31343 8588 31392 8616
rect 31343 8585 31355 8588
rect 31297 8579 31355 8585
rect 31386 8576 31392 8588
rect 31444 8576 31450 8628
rect 32030 8576 32036 8628
rect 32088 8576 32094 8628
rect 32766 8576 32772 8628
rect 32824 8616 32830 8628
rect 33502 8616 33508 8628
rect 32824 8588 33508 8616
rect 32824 8576 32830 8588
rect 33502 8576 33508 8588
rect 33560 8576 33566 8628
rect 30006 8548 30012 8560
rect 29104 8520 30012 8548
rect 26973 8483 27031 8489
rect 26973 8480 26985 8483
rect 26568 8452 26985 8480
rect 26568 8440 26574 8452
rect 26973 8449 26985 8452
rect 27019 8449 27031 8483
rect 26973 8443 27031 8449
rect 27157 8483 27215 8489
rect 27157 8449 27169 8483
rect 27203 8449 27215 8483
rect 27157 8443 27215 8449
rect 27249 8483 27307 8489
rect 27249 8449 27261 8483
rect 27295 8449 27307 8483
rect 27249 8443 27307 8449
rect 27338 8440 27344 8492
rect 27396 8440 27402 8492
rect 27430 8440 27436 8492
rect 27488 8480 27494 8492
rect 27525 8483 27583 8489
rect 27525 8480 27537 8483
rect 27488 8452 27537 8480
rect 27488 8440 27494 8452
rect 27525 8449 27537 8452
rect 27571 8449 27583 8483
rect 27525 8443 27583 8449
rect 27614 8440 27620 8492
rect 27672 8480 27678 8492
rect 29104 8489 29132 8520
rect 30006 8508 30012 8520
rect 30064 8548 30070 8560
rect 31938 8548 31944 8560
rect 30064 8520 31944 8548
rect 30064 8508 30070 8520
rect 31938 8508 31944 8520
rect 31996 8508 32002 8560
rect 28905 8483 28963 8489
rect 28905 8480 28917 8483
rect 27672 8452 28917 8480
rect 27672 8440 27678 8452
rect 28905 8449 28917 8452
rect 28951 8449 28963 8483
rect 28905 8443 28963 8449
rect 29089 8483 29147 8489
rect 29089 8449 29101 8483
rect 29135 8449 29147 8483
rect 29089 8443 29147 8449
rect 31573 8483 31631 8489
rect 31573 8449 31585 8483
rect 31619 8480 31631 8483
rect 31662 8480 31668 8492
rect 31619 8452 31668 8480
rect 31619 8449 31631 8452
rect 31573 8443 31631 8449
rect 24765 8415 24823 8421
rect 24765 8381 24777 8415
rect 24811 8381 24823 8415
rect 28920 8412 28948 8443
rect 31662 8440 31668 8452
rect 31720 8440 31726 8492
rect 31849 8483 31907 8489
rect 31849 8449 31861 8483
rect 31895 8480 31907 8483
rect 32048 8480 32076 8576
rect 35986 8548 35992 8560
rect 31895 8452 32076 8480
rect 32968 8520 35992 8548
rect 31895 8449 31907 8452
rect 31849 8443 31907 8449
rect 29270 8412 29276 8424
rect 24765 8375 24823 8381
rect 27448 8384 27936 8412
rect 28920 8384 29276 8412
rect 9784 8316 13584 8344
rect 9677 8307 9735 8313
rect 16942 8304 16948 8356
rect 17000 8344 17006 8356
rect 17000 8316 17172 8344
rect 17000 8304 17006 8316
rect 2958 8236 2964 8288
rect 3016 8276 3022 8288
rect 3237 8279 3295 8285
rect 3237 8276 3249 8279
rect 3016 8248 3249 8276
rect 3016 8236 3022 8248
rect 3237 8245 3249 8248
rect 3283 8245 3295 8279
rect 3237 8239 3295 8245
rect 4614 8236 4620 8288
rect 4672 8236 4678 8288
rect 6270 8236 6276 8288
rect 6328 8276 6334 8288
rect 6549 8279 6607 8285
rect 6549 8276 6561 8279
rect 6328 8248 6561 8276
rect 6328 8236 6334 8248
rect 6549 8245 6561 8248
rect 6595 8276 6607 8279
rect 6822 8276 6828 8288
rect 6595 8248 6828 8276
rect 6595 8245 6607 8248
rect 6549 8239 6607 8245
rect 6822 8236 6828 8248
rect 6880 8276 6886 8288
rect 8662 8276 8668 8288
rect 6880 8248 8668 8276
rect 6880 8236 6886 8248
rect 8662 8236 8668 8248
rect 8720 8236 8726 8288
rect 17144 8276 17172 8316
rect 17218 8304 17224 8356
rect 17276 8304 17282 8356
rect 27448 8344 27476 8384
rect 17328 8316 27476 8344
rect 27709 8347 27767 8353
rect 17328 8276 17356 8316
rect 27709 8313 27721 8347
rect 27755 8344 27767 8347
rect 27798 8344 27804 8356
rect 27755 8316 27804 8344
rect 27755 8313 27767 8316
rect 27709 8307 27767 8313
rect 27798 8304 27804 8316
rect 27856 8304 27862 8356
rect 27908 8344 27936 8384
rect 29270 8372 29276 8384
rect 29328 8372 29334 8424
rect 31018 8372 31024 8424
rect 31076 8412 31082 8424
rect 31389 8415 31447 8421
rect 31389 8412 31401 8415
rect 31076 8384 31401 8412
rect 31076 8372 31082 8384
rect 31389 8381 31401 8384
rect 31435 8381 31447 8415
rect 32968 8412 32996 8520
rect 35986 8508 35992 8520
rect 36044 8508 36050 8560
rect 33042 8440 33048 8492
rect 33100 8480 33106 8492
rect 33137 8483 33195 8489
rect 33137 8480 33149 8483
rect 33100 8452 33149 8480
rect 33100 8440 33106 8452
rect 33137 8449 33149 8452
rect 33183 8449 33195 8483
rect 33137 8443 33195 8449
rect 31389 8375 31447 8381
rect 31726 8384 32996 8412
rect 31726 8344 31754 8384
rect 33226 8372 33232 8424
rect 33284 8372 33290 8424
rect 27908 8316 31754 8344
rect 32582 8304 32588 8356
rect 32640 8344 32646 8356
rect 32769 8347 32827 8353
rect 32769 8344 32781 8347
rect 32640 8316 32781 8344
rect 32640 8304 32646 8316
rect 32769 8313 32781 8316
rect 32815 8313 32827 8347
rect 32769 8307 32827 8313
rect 17144 8248 17356 8276
rect 19518 8236 19524 8288
rect 19576 8236 19582 8288
rect 20898 8236 20904 8288
rect 20956 8276 20962 8288
rect 21910 8276 21916 8288
rect 20956 8248 21916 8276
rect 20956 8236 20962 8248
rect 21910 8236 21916 8248
rect 21968 8236 21974 8288
rect 22281 8279 22339 8285
rect 22281 8245 22293 8279
rect 22327 8276 22339 8279
rect 22370 8276 22376 8288
rect 22327 8248 22376 8276
rect 22327 8245 22339 8248
rect 22281 8239 22339 8245
rect 22370 8236 22376 8248
rect 22428 8236 22434 8288
rect 23014 8236 23020 8288
rect 23072 8236 23078 8288
rect 25314 8236 25320 8288
rect 25372 8236 25378 8288
rect 28994 8236 29000 8288
rect 29052 8236 29058 8288
rect 1104 8186 38272 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 38272 8186
rect 1104 8112 38272 8134
rect 5534 8032 5540 8084
rect 5592 8072 5598 8084
rect 5629 8075 5687 8081
rect 5629 8072 5641 8075
rect 5592 8044 5641 8072
rect 5592 8032 5598 8044
rect 5629 8041 5641 8044
rect 5675 8041 5687 8075
rect 5629 8035 5687 8041
rect 5810 8032 5816 8084
rect 5868 8072 5874 8084
rect 6362 8072 6368 8084
rect 5868 8044 6368 8072
rect 5868 8032 5874 8044
rect 6362 8032 6368 8044
rect 6420 8032 6426 8084
rect 6472 8044 8248 8072
rect 5828 7936 5856 8032
rect 5644 7908 5856 7936
rect 5644 7877 5672 7908
rect 5629 7871 5687 7877
rect 5629 7837 5641 7871
rect 5675 7837 5687 7871
rect 5629 7831 5687 7837
rect 5718 7828 5724 7880
rect 5776 7828 5782 7880
rect 5813 7871 5871 7877
rect 5813 7837 5825 7871
rect 5859 7868 5871 7871
rect 5902 7868 5908 7880
rect 5859 7840 5908 7868
rect 5859 7837 5871 7840
rect 5813 7831 5871 7837
rect 5902 7828 5908 7840
rect 5960 7828 5966 7880
rect 6472 7877 6500 8044
rect 8220 8004 8248 8044
rect 8662 8032 8668 8084
rect 8720 8032 8726 8084
rect 8846 8032 8852 8084
rect 8904 8072 8910 8084
rect 9858 8072 9864 8084
rect 8904 8044 9864 8072
rect 8904 8032 8910 8044
rect 9858 8032 9864 8044
rect 9916 8032 9922 8084
rect 12526 8032 12532 8084
rect 12584 8072 12590 8084
rect 12805 8075 12863 8081
rect 12805 8072 12817 8075
rect 12584 8044 12817 8072
rect 12584 8032 12590 8044
rect 12805 8041 12817 8044
rect 12851 8041 12863 8075
rect 12805 8035 12863 8041
rect 12986 8032 12992 8084
rect 13044 8072 13050 8084
rect 13541 8075 13599 8081
rect 13541 8072 13553 8075
rect 13044 8044 13553 8072
rect 13044 8032 13050 8044
rect 13541 8041 13553 8044
rect 13587 8041 13599 8075
rect 13541 8035 13599 8041
rect 13722 8032 13728 8084
rect 13780 8032 13786 8084
rect 20165 8075 20223 8081
rect 20165 8041 20177 8075
rect 20211 8072 20223 8075
rect 23566 8072 23572 8084
rect 20211 8044 23572 8072
rect 20211 8041 20223 8044
rect 20165 8035 20223 8041
rect 23566 8032 23572 8044
rect 23624 8032 23630 8084
rect 26234 8032 26240 8084
rect 26292 8072 26298 8084
rect 29362 8072 29368 8084
rect 26292 8044 29368 8072
rect 26292 8032 26298 8044
rect 29362 8032 29368 8044
rect 29420 8032 29426 8084
rect 29454 8032 29460 8084
rect 29512 8032 29518 8084
rect 31478 8072 31484 8084
rect 30576 8044 31484 8072
rect 17497 8007 17555 8013
rect 17497 8004 17509 8007
rect 8220 7976 17509 8004
rect 17497 7973 17509 7976
rect 17543 7973 17555 8007
rect 17497 7967 17555 7973
rect 21637 8007 21695 8013
rect 21637 7973 21649 8007
rect 21683 8004 21695 8007
rect 22646 8004 22652 8016
rect 21683 7976 22652 8004
rect 21683 7973 21695 7976
rect 21637 7967 21695 7973
rect 22646 7964 22652 7976
rect 22704 7964 22710 8016
rect 22738 7964 22744 8016
rect 22796 8004 22802 8016
rect 23293 8007 23351 8013
rect 23293 8004 23305 8007
rect 22796 7976 23305 8004
rect 22796 7964 22802 7976
rect 23293 7973 23305 7976
rect 23339 7973 23351 8007
rect 23293 7967 23351 7973
rect 6641 7939 6699 7945
rect 6641 7905 6653 7939
rect 6687 7905 6699 7939
rect 6641 7899 6699 7905
rect 6457 7871 6515 7877
rect 6457 7837 6469 7871
rect 6503 7837 6515 7871
rect 6457 7831 6515 7837
rect 5736 7800 5764 7828
rect 6656 7800 6684 7899
rect 6914 7896 6920 7948
rect 6972 7936 6978 7948
rect 9398 7936 9404 7948
rect 6972 7908 9404 7936
rect 6972 7896 6978 7908
rect 9398 7896 9404 7908
rect 9456 7896 9462 7948
rect 10594 7936 10600 7948
rect 9692 7908 10600 7936
rect 8294 7828 8300 7880
rect 8352 7868 8358 7880
rect 8846 7868 8852 7880
rect 8352 7840 8852 7868
rect 8352 7828 8358 7840
rect 8846 7828 8852 7840
rect 8904 7828 8910 7880
rect 9214 7828 9220 7880
rect 9272 7868 9278 7880
rect 9692 7877 9720 7908
rect 10594 7896 10600 7908
rect 10652 7896 10658 7948
rect 12161 7939 12219 7945
rect 12161 7905 12173 7939
rect 12207 7936 12219 7939
rect 12250 7936 12256 7948
rect 12207 7908 12256 7936
rect 12207 7905 12219 7908
rect 12161 7899 12219 7905
rect 12250 7896 12256 7908
rect 12308 7896 12314 7948
rect 12621 7939 12679 7945
rect 12621 7936 12633 7939
rect 12406 7908 12633 7936
rect 9677 7871 9735 7877
rect 9677 7868 9689 7871
rect 9272 7840 9689 7868
rect 9272 7828 9278 7840
rect 9677 7837 9689 7840
rect 9723 7837 9735 7871
rect 9677 7831 9735 7837
rect 9861 7871 9919 7877
rect 9861 7837 9873 7871
rect 9907 7868 9919 7871
rect 10870 7868 10876 7880
rect 9907 7840 10876 7868
rect 9907 7837 9919 7840
rect 9861 7831 9919 7837
rect 10870 7828 10876 7840
rect 10928 7868 10934 7880
rect 12406 7868 12434 7908
rect 12621 7905 12633 7908
rect 12667 7936 12679 7939
rect 13538 7936 13544 7948
rect 12667 7908 13544 7936
rect 12667 7905 12679 7908
rect 12621 7899 12679 7905
rect 13538 7896 13544 7908
rect 13596 7896 13602 7948
rect 13998 7896 14004 7948
rect 14056 7896 14062 7948
rect 15930 7896 15936 7948
rect 15988 7896 15994 7948
rect 17144 7908 17816 7936
rect 10928 7840 12434 7868
rect 10928 7828 10934 7840
rect 12894 7828 12900 7880
rect 12952 7868 12958 7880
rect 13357 7871 13415 7877
rect 13357 7868 13369 7871
rect 12952 7840 13369 7868
rect 12952 7828 12958 7840
rect 13357 7837 13369 7840
rect 13403 7868 13415 7871
rect 13725 7871 13783 7877
rect 13725 7868 13737 7871
rect 13403 7840 13737 7868
rect 13403 7837 13415 7840
rect 13357 7831 13415 7837
rect 13725 7837 13737 7840
rect 13771 7837 13783 7871
rect 13725 7831 13783 7837
rect 13909 7871 13967 7877
rect 13909 7837 13921 7871
rect 13955 7837 13967 7871
rect 14016 7868 14044 7896
rect 15749 7871 15807 7877
rect 15749 7868 15761 7871
rect 14016 7840 15761 7868
rect 13909 7831 13967 7837
rect 15749 7837 15761 7840
rect 15795 7837 15807 7871
rect 15749 7831 15807 7837
rect 15841 7871 15899 7877
rect 15841 7837 15853 7871
rect 15887 7868 15899 7871
rect 17144 7868 17172 7908
rect 17788 7880 17816 7908
rect 19518 7896 19524 7948
rect 19576 7896 19582 7948
rect 20622 7936 20628 7948
rect 19904 7908 20628 7936
rect 15887 7840 17172 7868
rect 17221 7871 17279 7877
rect 15887 7837 15899 7840
rect 15841 7831 15899 7837
rect 17221 7837 17233 7871
rect 17267 7868 17279 7871
rect 17586 7868 17592 7880
rect 17267 7840 17592 7868
rect 17267 7837 17279 7840
rect 17221 7831 17279 7837
rect 5736 7772 6684 7800
rect 7190 7760 7196 7812
rect 7248 7760 7254 7812
rect 10413 7803 10471 7809
rect 10413 7800 10425 7803
rect 9692 7772 10425 7800
rect 9692 7744 9720 7772
rect 10413 7769 10425 7772
rect 10459 7769 10471 7803
rect 10413 7763 10471 7769
rect 12342 7760 12348 7812
rect 12400 7760 12406 7812
rect 12526 7760 12532 7812
rect 12584 7800 12590 7812
rect 13538 7800 13544 7812
rect 12584 7772 13544 7800
rect 12584 7760 12590 7772
rect 13538 7760 13544 7772
rect 13596 7800 13602 7812
rect 13924 7800 13952 7831
rect 17586 7828 17592 7840
rect 17644 7828 17650 7880
rect 17770 7828 17776 7880
rect 17828 7828 17834 7880
rect 19536 7868 19564 7896
rect 19702 7868 19708 7880
rect 19536 7840 19708 7868
rect 19702 7828 19708 7840
rect 19760 7828 19766 7880
rect 19904 7877 19932 7908
rect 20622 7896 20628 7908
rect 20680 7936 20686 7948
rect 22278 7936 22284 7948
rect 20680 7908 22284 7936
rect 20680 7896 20686 7908
rect 19889 7871 19947 7877
rect 19889 7837 19901 7871
rect 19935 7837 19947 7871
rect 19889 7831 19947 7837
rect 20073 7871 20131 7877
rect 20073 7837 20085 7871
rect 20119 7837 20131 7871
rect 20073 7831 20131 7837
rect 20257 7871 20315 7877
rect 20257 7837 20269 7871
rect 20303 7868 20315 7871
rect 20303 7840 20576 7868
rect 20303 7837 20315 7840
rect 20257 7831 20315 7837
rect 16850 7800 16856 7812
rect 13596 7772 16856 7800
rect 13596 7760 13602 7772
rect 16850 7760 16856 7772
rect 16908 7760 16914 7812
rect 17497 7803 17555 7809
rect 17497 7769 17509 7803
rect 17543 7800 17555 7803
rect 17681 7803 17739 7809
rect 17681 7800 17693 7803
rect 17543 7772 17693 7800
rect 17543 7769 17555 7772
rect 17497 7763 17555 7769
rect 17681 7769 17693 7772
rect 17727 7769 17739 7803
rect 17681 7763 17739 7769
rect 19797 7803 19855 7809
rect 19797 7769 19809 7803
rect 19843 7800 19855 7803
rect 20088 7800 20116 7831
rect 19843 7772 20116 7800
rect 19843 7769 19855 7772
rect 19797 7763 19855 7769
rect 20548 7744 20576 7840
rect 21450 7828 21456 7880
rect 21508 7868 21514 7880
rect 21744 7877 21772 7908
rect 22278 7896 22284 7908
rect 22336 7896 22342 7948
rect 22370 7896 22376 7948
rect 22428 7896 22434 7948
rect 23014 7936 23020 7948
rect 22572 7908 23020 7936
rect 21545 7871 21603 7877
rect 21545 7868 21557 7871
rect 21508 7840 21557 7868
rect 21508 7828 21514 7840
rect 21545 7837 21557 7840
rect 21591 7837 21603 7871
rect 21545 7831 21603 7837
rect 21729 7871 21787 7877
rect 21729 7837 21741 7871
rect 21775 7837 21787 7871
rect 21729 7831 21787 7837
rect 21818 7828 21824 7880
rect 21876 7828 21882 7880
rect 21913 7871 21971 7877
rect 21913 7837 21925 7871
rect 21959 7837 21971 7871
rect 21913 7831 21971 7837
rect 22097 7871 22155 7877
rect 22097 7837 22109 7871
rect 22143 7837 22155 7871
rect 22097 7831 22155 7837
rect 22189 7871 22247 7877
rect 22189 7837 22201 7871
rect 22235 7868 22247 7871
rect 22572 7868 22600 7908
rect 23014 7896 23020 7908
rect 23072 7896 23078 7948
rect 28534 7896 28540 7948
rect 28592 7936 28598 7948
rect 28718 7936 28724 7948
rect 28592 7908 28724 7936
rect 28592 7896 28598 7908
rect 28718 7896 28724 7908
rect 28776 7896 28782 7948
rect 29472 7936 29500 8032
rect 30285 7939 30343 7945
rect 29472 7908 30236 7936
rect 22235 7840 22600 7868
rect 22235 7837 22247 7840
rect 22189 7831 22247 7837
rect 6086 7692 6092 7744
rect 6144 7692 6150 7744
rect 6546 7692 6552 7744
rect 6604 7692 6610 7744
rect 9674 7692 9680 7744
rect 9732 7692 9738 7744
rect 9766 7692 9772 7744
rect 9824 7692 9830 7744
rect 15378 7692 15384 7744
rect 15436 7692 15442 7744
rect 17310 7692 17316 7744
rect 17368 7692 17374 7744
rect 20530 7692 20536 7744
rect 20588 7692 20594 7744
rect 21928 7732 21956 7831
rect 22112 7800 22140 7831
rect 22646 7828 22652 7880
rect 22704 7828 22710 7880
rect 30006 7828 30012 7880
rect 30064 7828 30070 7880
rect 30208 7877 30236 7908
rect 30285 7905 30297 7939
rect 30331 7936 30343 7939
rect 30466 7936 30472 7948
rect 30331 7908 30472 7936
rect 30331 7905 30343 7908
rect 30285 7899 30343 7905
rect 30466 7896 30472 7908
rect 30524 7896 30530 7948
rect 30576 7880 30604 8044
rect 31478 8032 31484 8044
rect 31536 8032 31542 8084
rect 31754 8032 31760 8084
rect 31812 8072 31818 8084
rect 31849 8075 31907 8081
rect 31849 8072 31861 8075
rect 31812 8044 31861 8072
rect 31812 8032 31818 8044
rect 31849 8041 31861 8044
rect 31895 8041 31907 8075
rect 31849 8035 31907 8041
rect 30745 8007 30803 8013
rect 30745 7973 30757 8007
rect 30791 8004 30803 8007
rect 33042 8004 33048 8016
rect 30791 7976 33048 8004
rect 30791 7973 30803 7976
rect 30745 7967 30803 7973
rect 33042 7964 33048 7976
rect 33100 7964 33106 8016
rect 30193 7871 30251 7877
rect 30193 7837 30205 7871
rect 30239 7837 30251 7871
rect 30193 7831 30251 7837
rect 30374 7828 30380 7880
rect 30432 7828 30438 7880
rect 30558 7828 30564 7880
rect 30616 7828 30622 7880
rect 30834 7828 30840 7880
rect 30892 7868 30898 7880
rect 30929 7871 30987 7877
rect 30929 7868 30941 7871
rect 30892 7840 30941 7868
rect 30892 7828 30898 7840
rect 30929 7837 30941 7840
rect 30975 7837 30987 7871
rect 30929 7831 30987 7837
rect 31018 7828 31024 7880
rect 31076 7868 31082 7880
rect 31389 7871 31447 7877
rect 31389 7868 31401 7871
rect 31076 7840 31401 7868
rect 31076 7828 31082 7840
rect 31389 7837 31401 7840
rect 31435 7868 31447 7871
rect 31481 7871 31539 7877
rect 31481 7868 31493 7871
rect 31435 7840 31493 7868
rect 31435 7837 31447 7840
rect 31389 7831 31447 7837
rect 31481 7837 31493 7840
rect 31527 7837 31539 7871
rect 31481 7831 31539 7837
rect 22370 7800 22376 7812
rect 22112 7772 22376 7800
rect 22370 7760 22376 7772
rect 22428 7760 22434 7812
rect 22738 7760 22744 7812
rect 22796 7760 22802 7812
rect 23106 7760 23112 7812
rect 23164 7760 23170 7812
rect 30392 7800 30420 7828
rect 30742 7800 30748 7812
rect 30392 7772 30748 7800
rect 30742 7760 30748 7772
rect 30800 7800 30806 7812
rect 31297 7803 31355 7809
rect 31297 7800 31309 7803
rect 30800 7772 31309 7800
rect 30800 7760 30806 7772
rect 31297 7769 31309 7772
rect 31343 7769 31355 7803
rect 31297 7763 31355 7769
rect 22094 7732 22100 7744
rect 21928 7704 22100 7732
rect 22094 7692 22100 7704
rect 22152 7692 22158 7744
rect 22278 7692 22284 7744
rect 22336 7692 22342 7744
rect 22462 7692 22468 7744
rect 22520 7732 22526 7744
rect 23198 7732 23204 7744
rect 22520 7704 23204 7732
rect 22520 7692 22526 7704
rect 23198 7692 23204 7704
rect 23256 7692 23262 7744
rect 24026 7692 24032 7744
rect 24084 7732 24090 7744
rect 24302 7732 24308 7744
rect 24084 7704 24308 7732
rect 24084 7692 24090 7704
rect 24302 7692 24308 7704
rect 24360 7732 24366 7744
rect 31110 7732 31116 7744
rect 24360 7704 31116 7732
rect 24360 7692 24366 7704
rect 31110 7692 31116 7704
rect 31168 7692 31174 7744
rect 31202 7692 31208 7744
rect 31260 7692 31266 7744
rect 31312 7732 31340 7763
rect 31662 7760 31668 7812
rect 31720 7760 31726 7812
rect 31680 7732 31708 7760
rect 31312 7704 31708 7732
rect 1104 7642 38272 7664
rect 1104 7590 4874 7642
rect 4926 7590 4938 7642
rect 4990 7590 5002 7642
rect 5054 7590 5066 7642
rect 5118 7590 5130 7642
rect 5182 7590 35594 7642
rect 35646 7590 35658 7642
rect 35710 7590 35722 7642
rect 35774 7590 35786 7642
rect 35838 7590 35850 7642
rect 35902 7590 38272 7642
rect 1104 7568 38272 7590
rect 4614 7528 4620 7540
rect 2608 7500 4620 7528
rect 1486 7352 1492 7404
rect 1544 7352 1550 7404
rect 2608 7401 2636 7500
rect 4614 7488 4620 7500
rect 4672 7488 4678 7540
rect 5629 7531 5687 7537
rect 5629 7497 5641 7531
rect 5675 7528 5687 7531
rect 6086 7528 6092 7540
rect 5675 7500 6092 7528
rect 5675 7497 5687 7500
rect 5629 7491 5687 7497
rect 6086 7488 6092 7500
rect 6144 7488 6150 7540
rect 6546 7488 6552 7540
rect 6604 7488 6610 7540
rect 7190 7488 7196 7540
rect 7248 7528 7254 7540
rect 7653 7531 7711 7537
rect 7653 7528 7665 7531
rect 7248 7500 7665 7528
rect 7248 7488 7254 7500
rect 7653 7497 7665 7500
rect 7699 7497 7711 7531
rect 7653 7491 7711 7497
rect 8018 7488 8024 7540
rect 8076 7488 8082 7540
rect 9766 7528 9772 7540
rect 9692 7500 9772 7528
rect 2869 7463 2927 7469
rect 2869 7429 2881 7463
rect 2915 7460 2927 7463
rect 2958 7460 2964 7472
rect 2915 7432 2964 7460
rect 2915 7429 2927 7432
rect 2869 7423 2927 7429
rect 2958 7420 2964 7432
rect 3016 7420 3022 7472
rect 2593 7395 2651 7401
rect 2593 7361 2605 7395
rect 2639 7361 2651 7395
rect 2593 7355 2651 7361
rect 3970 7352 3976 7404
rect 4028 7352 4034 7404
rect 5442 7392 5448 7404
rect 4264 7364 5448 7392
rect 1673 7327 1731 7333
rect 1673 7293 1685 7327
rect 1719 7324 1731 7327
rect 4264 7324 4292 7364
rect 5442 7352 5448 7364
rect 5500 7352 5506 7404
rect 5537 7395 5595 7401
rect 5537 7361 5549 7395
rect 5583 7392 5595 7395
rect 5994 7392 6000 7404
rect 5583 7364 6000 7392
rect 5583 7361 5595 7364
rect 5537 7355 5595 7361
rect 5994 7352 6000 7364
rect 6052 7352 6058 7404
rect 1719 7296 4292 7324
rect 4341 7327 4399 7333
rect 1719 7293 1731 7296
rect 1673 7287 1731 7293
rect 4341 7293 4353 7327
rect 4387 7324 4399 7327
rect 4706 7324 4712 7336
rect 4387 7296 4712 7324
rect 4387 7293 4399 7296
rect 4341 7287 4399 7293
rect 4706 7284 4712 7296
rect 4764 7284 4770 7336
rect 5626 7284 5632 7336
rect 5684 7324 5690 7336
rect 5721 7327 5779 7333
rect 5721 7324 5733 7327
rect 5684 7296 5733 7324
rect 5684 7284 5690 7296
rect 5721 7293 5733 7296
rect 5767 7293 5779 7327
rect 5721 7287 5779 7293
rect 6012 7256 6040 7352
rect 6365 7327 6423 7333
rect 6365 7293 6377 7327
rect 6411 7324 6423 7327
rect 6564 7324 6592 7488
rect 6733 7395 6791 7401
rect 6733 7361 6745 7395
rect 6779 7361 6791 7395
rect 6733 7355 6791 7361
rect 7837 7395 7895 7401
rect 7837 7361 7849 7395
rect 7883 7392 7895 7395
rect 8036 7392 8064 7488
rect 9692 7469 9720 7500
rect 9766 7488 9772 7500
rect 9824 7488 9830 7540
rect 9858 7488 9864 7540
rect 9916 7488 9922 7540
rect 13630 7488 13636 7540
rect 13688 7488 13694 7540
rect 15378 7488 15384 7540
rect 15436 7488 15442 7540
rect 19150 7488 19156 7540
rect 19208 7488 19214 7540
rect 21082 7488 21088 7540
rect 21140 7488 21146 7540
rect 22278 7488 22284 7540
rect 22336 7488 22342 7540
rect 22370 7488 22376 7540
rect 22428 7488 22434 7540
rect 22756 7500 23060 7528
rect 9677 7463 9735 7469
rect 9677 7429 9689 7463
rect 9723 7429 9735 7463
rect 9876 7460 9904 7488
rect 9876 7432 10166 7460
rect 9677 7423 9735 7429
rect 11790 7420 11796 7472
rect 11848 7420 11854 7472
rect 12066 7420 12072 7472
rect 12124 7460 12130 7472
rect 13648 7460 13676 7488
rect 15286 7460 15292 7472
rect 12124 7432 12282 7460
rect 13648 7432 15292 7460
rect 12124 7420 12130 7432
rect 7883 7364 8064 7392
rect 7883 7361 7895 7364
rect 7837 7355 7895 7361
rect 6411 7296 6592 7324
rect 6411 7293 6423 7296
rect 6365 7287 6423 7293
rect 6748 7256 6776 7355
rect 9398 7352 9404 7404
rect 9456 7352 9462 7404
rect 12802 7352 12808 7404
rect 12860 7352 12866 7404
rect 14182 7352 14188 7404
rect 14240 7392 14246 7404
rect 14277 7395 14335 7401
rect 14277 7392 14289 7395
rect 14240 7364 14289 7392
rect 14240 7352 14246 7364
rect 14277 7361 14289 7364
rect 14323 7361 14335 7395
rect 14277 7355 14335 7361
rect 6822 7284 6828 7336
rect 6880 7284 6886 7336
rect 11517 7327 11575 7333
rect 11517 7293 11529 7327
rect 11563 7324 11575 7327
rect 11882 7324 11888 7336
rect 11563 7296 11888 7324
rect 11563 7293 11575 7296
rect 11517 7287 11575 7293
rect 11882 7284 11888 7296
rect 11940 7324 11946 7336
rect 12250 7324 12256 7336
rect 11940 7296 12256 7324
rect 11940 7284 11946 7296
rect 12250 7284 12256 7296
rect 12308 7284 12314 7336
rect 12820 7324 12848 7352
rect 13817 7327 13875 7333
rect 13817 7324 13829 7327
rect 12820 7296 13829 7324
rect 13817 7293 13829 7296
rect 13863 7293 13875 7327
rect 14292 7324 14320 7355
rect 14458 7352 14464 7404
rect 14516 7392 14522 7404
rect 14844 7401 14872 7432
rect 15286 7420 15292 7432
rect 15344 7420 15350 7472
rect 14553 7395 14611 7401
rect 14553 7392 14565 7395
rect 14516 7364 14565 7392
rect 14516 7352 14522 7364
rect 14553 7361 14565 7364
rect 14599 7361 14611 7395
rect 14553 7355 14611 7361
rect 14829 7395 14887 7401
rect 14829 7361 14841 7395
rect 14875 7361 14887 7395
rect 15396 7392 15424 7488
rect 18506 7460 18512 7472
rect 17972 7432 18512 7460
rect 15473 7395 15531 7401
rect 15473 7392 15485 7395
rect 15396 7364 15485 7392
rect 14829 7355 14887 7361
rect 15473 7361 15485 7364
rect 15519 7361 15531 7395
rect 15473 7355 15531 7361
rect 17770 7352 17776 7404
rect 17828 7352 17834 7404
rect 17972 7401 18000 7432
rect 18506 7420 18512 7432
rect 18564 7460 18570 7472
rect 19168 7460 19196 7488
rect 18564 7432 19196 7460
rect 19337 7463 19395 7469
rect 18564 7420 18570 7432
rect 19337 7429 19349 7463
rect 19383 7460 19395 7463
rect 20165 7463 20223 7469
rect 20165 7460 20177 7463
rect 19383 7432 20177 7460
rect 19383 7429 19395 7432
rect 19337 7423 19395 7429
rect 20165 7429 20177 7432
rect 20211 7429 20223 7463
rect 21100 7460 21128 7488
rect 20165 7423 20223 7429
rect 20916 7432 21128 7460
rect 17957 7395 18015 7401
rect 17957 7361 17969 7395
rect 18003 7361 18015 7395
rect 19153 7395 19211 7401
rect 19153 7392 19165 7395
rect 17957 7355 18015 7361
rect 18064 7364 19165 7392
rect 14645 7327 14703 7333
rect 14645 7324 14657 7327
rect 14292 7296 14657 7324
rect 13817 7287 13875 7293
rect 14645 7293 14657 7296
rect 14691 7293 14703 7327
rect 14645 7287 14703 7293
rect 15013 7327 15071 7333
rect 15013 7293 15025 7327
rect 15059 7324 15071 7327
rect 15286 7324 15292 7336
rect 15059 7296 15292 7324
rect 15059 7293 15071 7296
rect 15013 7287 15071 7293
rect 15286 7284 15292 7296
rect 15344 7284 15350 7336
rect 6012 7228 6776 7256
rect 14461 7259 14519 7265
rect 14461 7225 14473 7259
rect 14507 7256 14519 7259
rect 14918 7256 14924 7268
rect 14507 7228 14924 7256
rect 14507 7225 14519 7228
rect 14461 7219 14519 7225
rect 14918 7216 14924 7228
rect 14976 7256 14982 7268
rect 15470 7256 15476 7268
rect 14976 7228 15476 7256
rect 14976 7216 14982 7228
rect 15470 7216 15476 7228
rect 15528 7216 15534 7268
rect 18064 7200 18092 7364
rect 19153 7361 19165 7364
rect 19199 7392 19211 7395
rect 19521 7395 19579 7401
rect 19521 7392 19533 7395
rect 19199 7364 19533 7392
rect 19199 7361 19211 7364
rect 19153 7355 19211 7361
rect 19521 7361 19533 7364
rect 19567 7361 19579 7395
rect 19521 7355 19579 7361
rect 19613 7395 19671 7401
rect 19613 7361 19625 7395
rect 19659 7361 19671 7395
rect 19613 7355 19671 7361
rect 18690 7284 18696 7336
rect 18748 7324 18754 7336
rect 18969 7327 19027 7333
rect 18969 7324 18981 7327
rect 18748 7296 18981 7324
rect 18748 7284 18754 7296
rect 18969 7293 18981 7296
rect 19015 7324 19027 7327
rect 19628 7324 19656 7355
rect 19702 7352 19708 7404
rect 19760 7392 19766 7404
rect 19797 7395 19855 7401
rect 19797 7392 19809 7395
rect 19760 7364 19809 7392
rect 19760 7352 19766 7364
rect 19797 7361 19809 7364
rect 19843 7361 19855 7395
rect 19797 7355 19855 7361
rect 20349 7395 20407 7401
rect 20349 7361 20361 7395
rect 20395 7392 20407 7395
rect 20622 7392 20628 7404
rect 20395 7364 20628 7392
rect 20395 7361 20407 7364
rect 20349 7355 20407 7361
rect 20622 7352 20628 7364
rect 20680 7392 20686 7404
rect 20809 7395 20867 7401
rect 20809 7392 20821 7395
rect 20680 7364 20821 7392
rect 20680 7352 20686 7364
rect 20809 7361 20821 7364
rect 20855 7361 20867 7395
rect 20809 7355 20867 7361
rect 20916 7333 20944 7432
rect 21821 7395 21879 7401
rect 21821 7392 21833 7395
rect 21100 7364 21833 7392
rect 20901 7327 20959 7333
rect 19015 7296 20668 7324
rect 19015 7293 19027 7296
rect 18969 7287 19027 7293
rect 19981 7259 20039 7265
rect 19981 7225 19993 7259
rect 20027 7256 20039 7259
rect 20027 7228 20576 7256
rect 20027 7225 20039 7228
rect 19981 7219 20039 7225
rect 20548 7200 20576 7228
rect 4798 7148 4804 7200
rect 4856 7188 4862 7200
rect 5169 7191 5227 7197
rect 5169 7188 5181 7191
rect 4856 7160 5181 7188
rect 4856 7148 4862 7160
rect 5169 7157 5181 7160
rect 5215 7157 5227 7191
rect 5169 7151 5227 7157
rect 11146 7148 11152 7200
rect 11204 7148 11210 7200
rect 12894 7148 12900 7200
rect 12952 7188 12958 7200
rect 13265 7191 13323 7197
rect 13265 7188 13277 7191
rect 12952 7160 13277 7188
rect 12952 7148 12958 7160
rect 13265 7157 13277 7160
rect 13311 7157 13323 7191
rect 13265 7151 13323 7157
rect 15562 7148 15568 7200
rect 15620 7188 15626 7200
rect 15657 7191 15715 7197
rect 15657 7188 15669 7191
rect 15620 7160 15669 7188
rect 15620 7148 15626 7160
rect 15657 7157 15669 7160
rect 15703 7157 15715 7191
rect 15657 7151 15715 7157
rect 17862 7148 17868 7200
rect 17920 7148 17926 7200
rect 18046 7148 18052 7200
rect 18104 7148 18110 7200
rect 20530 7148 20536 7200
rect 20588 7148 20594 7200
rect 20640 7188 20668 7296
rect 20901 7293 20913 7327
rect 20947 7293 20959 7327
rect 20901 7287 20959 7293
rect 21100 7188 21128 7364
rect 21821 7361 21833 7364
rect 21867 7361 21879 7395
rect 21821 7355 21879 7361
rect 22094 7352 22100 7404
rect 22152 7352 22158 7404
rect 22186 7352 22192 7404
rect 22244 7352 22250 7404
rect 22296 7392 22324 7488
rect 22756 7401 22784 7500
rect 22922 7420 22928 7472
rect 22980 7420 22986 7472
rect 23032 7460 23060 7500
rect 23106 7488 23112 7540
rect 23164 7528 23170 7540
rect 23201 7531 23259 7537
rect 23201 7528 23213 7531
rect 23164 7500 23213 7528
rect 23164 7488 23170 7500
rect 23201 7497 23213 7500
rect 23247 7497 23259 7531
rect 26418 7528 26424 7540
rect 23201 7491 23259 7497
rect 23860 7500 26424 7528
rect 23860 7460 23888 7500
rect 26418 7488 26424 7500
rect 26476 7488 26482 7540
rect 26602 7488 26608 7540
rect 26660 7528 26666 7540
rect 27430 7528 27436 7540
rect 26660 7500 27436 7528
rect 26660 7488 26666 7500
rect 27430 7488 27436 7500
rect 27488 7488 27494 7540
rect 27614 7488 27620 7540
rect 27672 7488 27678 7540
rect 27706 7488 27712 7540
rect 27764 7528 27770 7540
rect 27764 7500 29592 7528
rect 27764 7488 27770 7500
rect 23032 7432 23888 7460
rect 23937 7463 23995 7469
rect 23937 7429 23949 7463
rect 23983 7460 23995 7463
rect 23983 7432 24164 7460
rect 23983 7429 23995 7432
rect 23937 7423 23995 7429
rect 22557 7395 22615 7401
rect 22557 7392 22569 7395
rect 22296 7364 22569 7392
rect 22557 7361 22569 7364
rect 22603 7361 22615 7395
rect 22557 7355 22615 7361
rect 22705 7395 22784 7401
rect 22705 7361 22717 7395
rect 22751 7364 22784 7395
rect 22833 7395 22891 7401
rect 22751 7361 22763 7364
rect 22705 7355 22763 7361
rect 22833 7361 22845 7395
rect 22879 7361 22891 7395
rect 22833 7355 22891 7361
rect 23063 7395 23121 7401
rect 23063 7361 23075 7395
rect 23109 7392 23121 7395
rect 23109 7364 23244 7392
rect 23109 7361 23121 7364
rect 23063 7355 23121 7361
rect 21266 7284 21272 7336
rect 21324 7324 21330 7336
rect 22848 7324 22876 7355
rect 21324 7296 22876 7324
rect 23216 7324 23244 7364
rect 23566 7352 23572 7404
rect 23624 7392 23630 7404
rect 23845 7395 23903 7401
rect 23845 7392 23857 7395
rect 23624 7364 23857 7392
rect 23624 7352 23630 7364
rect 23845 7361 23857 7364
rect 23891 7361 23903 7395
rect 23845 7355 23903 7361
rect 24026 7352 24032 7404
rect 24084 7352 24090 7404
rect 24136 7401 24164 7432
rect 24320 7432 25084 7460
rect 24320 7401 24348 7432
rect 24121 7395 24179 7401
rect 24121 7361 24133 7395
rect 24167 7361 24179 7395
rect 24121 7355 24179 7361
rect 24305 7395 24363 7401
rect 24305 7361 24317 7395
rect 24351 7361 24363 7395
rect 24305 7355 24363 7361
rect 24486 7352 24492 7404
rect 24544 7352 24550 7404
rect 24578 7352 24584 7404
rect 24636 7392 24642 7404
rect 24673 7395 24731 7401
rect 24673 7392 24685 7395
rect 24636 7364 24685 7392
rect 24636 7352 24642 7364
rect 24673 7361 24685 7364
rect 24719 7361 24731 7395
rect 24673 7355 24731 7361
rect 24397 7327 24455 7333
rect 24397 7324 24409 7327
rect 23216 7296 24409 7324
rect 21324 7284 21330 7296
rect 21177 7259 21235 7265
rect 21177 7225 21189 7259
rect 21223 7256 21235 7259
rect 22002 7256 22008 7268
rect 21223 7228 22008 7256
rect 21223 7225 21235 7228
rect 21177 7219 21235 7225
rect 22002 7216 22008 7228
rect 22060 7256 22066 7268
rect 23216 7256 23244 7296
rect 24397 7293 24409 7296
rect 24443 7293 24455 7327
rect 24397 7287 24455 7293
rect 22060 7228 23244 7256
rect 22060 7216 22066 7228
rect 23290 7216 23296 7268
rect 23348 7256 23354 7268
rect 24688 7256 24716 7355
rect 23348 7228 24716 7256
rect 25056 7256 25084 7432
rect 25314 7420 25320 7472
rect 25372 7460 25378 7472
rect 25593 7463 25651 7469
rect 25593 7460 25605 7463
rect 25372 7432 25605 7460
rect 25372 7420 25378 7432
rect 25593 7429 25605 7432
rect 25639 7429 25651 7463
rect 25593 7423 25651 7429
rect 26234 7420 26240 7472
rect 26292 7420 26298 7472
rect 26326 7420 26332 7472
rect 26384 7460 26390 7472
rect 27632 7460 27660 7488
rect 29564 7460 29592 7500
rect 30006 7488 30012 7540
rect 30064 7528 30070 7540
rect 30101 7531 30159 7537
rect 30101 7528 30113 7531
rect 30064 7500 30113 7528
rect 30064 7488 30070 7500
rect 30101 7497 30113 7500
rect 30147 7497 30159 7531
rect 30101 7491 30159 7497
rect 31202 7488 31208 7540
rect 31260 7528 31266 7540
rect 31260 7500 31754 7528
rect 31260 7488 31266 7500
rect 31570 7460 31576 7472
rect 26384 7432 26648 7460
rect 27632 7432 27844 7460
rect 26384 7420 26390 7432
rect 25133 7395 25191 7401
rect 25133 7361 25145 7395
rect 25179 7392 25191 7395
rect 25222 7392 25228 7404
rect 25179 7364 25228 7392
rect 25179 7361 25191 7364
rect 25133 7355 25191 7361
rect 25222 7352 25228 7364
rect 25280 7352 25286 7404
rect 26252 7392 26280 7420
rect 26620 7401 26648 7432
rect 27816 7401 27844 7432
rect 29012 7432 29500 7460
rect 29564 7432 30144 7460
rect 26421 7395 26479 7401
rect 26421 7392 26433 7395
rect 26252 7364 26433 7392
rect 26421 7361 26433 7364
rect 26467 7361 26479 7395
rect 26421 7355 26479 7361
rect 26605 7395 26663 7401
rect 26605 7361 26617 7395
rect 26651 7361 26663 7395
rect 26605 7355 26663 7361
rect 27617 7395 27675 7401
rect 27617 7361 27629 7395
rect 27663 7361 27675 7395
rect 27617 7355 27675 7361
rect 27801 7395 27859 7401
rect 27801 7361 27813 7395
rect 27847 7361 27859 7395
rect 27801 7355 27859 7361
rect 27893 7395 27951 7401
rect 27893 7361 27905 7395
rect 27939 7361 27951 7395
rect 27893 7355 27951 7361
rect 27985 7395 28043 7401
rect 27985 7361 27997 7395
rect 28031 7392 28043 7395
rect 28445 7395 28503 7401
rect 28445 7392 28457 7395
rect 28031 7364 28457 7392
rect 28031 7361 28043 7364
rect 27985 7355 28043 7361
rect 28445 7361 28457 7364
rect 28491 7392 28503 7395
rect 28534 7392 28540 7404
rect 28491 7364 28540 7392
rect 28491 7361 28503 7364
rect 28445 7355 28503 7361
rect 25317 7327 25375 7333
rect 25317 7293 25329 7327
rect 25363 7324 25375 7327
rect 25406 7324 25412 7336
rect 25363 7296 25412 7324
rect 25363 7293 25375 7296
rect 25317 7287 25375 7293
rect 25406 7284 25412 7296
rect 25464 7284 25470 7336
rect 25958 7284 25964 7336
rect 26016 7324 26022 7336
rect 27632 7324 27660 7355
rect 26016 7296 27660 7324
rect 26016 7284 26022 7296
rect 25976 7256 26004 7284
rect 25056 7228 26004 7256
rect 23348 7216 23354 7228
rect 21358 7188 21364 7200
rect 20640 7160 21364 7188
rect 21358 7148 21364 7160
rect 21416 7148 21422 7200
rect 21910 7148 21916 7200
rect 21968 7188 21974 7200
rect 24762 7188 24768 7200
rect 21968 7160 24768 7188
rect 21968 7148 21974 7160
rect 24762 7148 24768 7160
rect 24820 7148 24826 7200
rect 24854 7148 24860 7200
rect 24912 7148 24918 7200
rect 24949 7191 25007 7197
rect 24949 7157 24961 7191
rect 24995 7188 25007 7191
rect 25038 7188 25044 7200
rect 24995 7160 25044 7188
rect 24995 7157 25007 7160
rect 24949 7151 25007 7157
rect 25038 7148 25044 7160
rect 25096 7148 25102 7200
rect 25130 7148 25136 7200
rect 25188 7148 25194 7200
rect 27632 7188 27660 7296
rect 27709 7327 27767 7333
rect 27709 7293 27721 7327
rect 27755 7324 27767 7327
rect 27908 7324 27936 7355
rect 28534 7352 28540 7364
rect 28592 7352 28598 7404
rect 29012 7401 29040 7432
rect 29472 7404 29500 7432
rect 28997 7395 29055 7401
rect 28997 7361 29009 7395
rect 29043 7361 29055 7395
rect 28997 7355 29055 7361
rect 29089 7395 29147 7401
rect 29089 7361 29101 7395
rect 29135 7361 29147 7395
rect 29089 7355 29147 7361
rect 27755 7296 27936 7324
rect 27755 7293 27767 7296
rect 27709 7287 27767 7293
rect 28626 7284 28632 7336
rect 28684 7284 28690 7336
rect 28074 7216 28080 7268
rect 28132 7256 28138 7268
rect 29104 7256 29132 7355
rect 29178 7352 29184 7404
rect 29236 7392 29242 7404
rect 29365 7395 29423 7401
rect 29365 7392 29377 7395
rect 29236 7364 29377 7392
rect 29236 7352 29242 7364
rect 29365 7361 29377 7364
rect 29411 7361 29423 7395
rect 29365 7355 29423 7361
rect 29454 7352 29460 7404
rect 29512 7352 29518 7404
rect 30116 7401 30144 7432
rect 30392 7432 31576 7460
rect 29641 7395 29699 7401
rect 29641 7361 29653 7395
rect 29687 7361 29699 7395
rect 29641 7355 29699 7361
rect 30101 7395 30159 7401
rect 30101 7361 30113 7395
rect 30147 7361 30159 7395
rect 30101 7355 30159 7361
rect 30285 7395 30343 7401
rect 30285 7361 30297 7395
rect 30331 7392 30343 7395
rect 30392 7392 30420 7432
rect 31570 7420 31576 7432
rect 31628 7420 31634 7472
rect 31726 7460 31754 7500
rect 31726 7432 31892 7460
rect 30331 7364 30420 7392
rect 30331 7361 30343 7364
rect 30285 7355 30343 7361
rect 28132 7228 29132 7256
rect 29656 7256 29684 7355
rect 30392 7336 30420 7364
rect 30650 7352 30656 7404
rect 30708 7392 30714 7404
rect 30745 7395 30803 7401
rect 30745 7392 30757 7395
rect 30708 7364 30757 7392
rect 30708 7352 30714 7364
rect 30745 7361 30757 7364
rect 30791 7361 30803 7395
rect 30745 7355 30803 7361
rect 31386 7352 31392 7404
rect 31444 7352 31450 7404
rect 31754 7352 31760 7404
rect 31812 7352 31818 7404
rect 31864 7401 31892 7432
rect 31849 7395 31907 7401
rect 31849 7361 31861 7395
rect 31895 7361 31907 7395
rect 31849 7355 31907 7361
rect 30374 7284 30380 7336
rect 30432 7284 30438 7336
rect 31294 7284 31300 7336
rect 31352 7284 31358 7336
rect 34054 7256 34060 7268
rect 29656 7228 34060 7256
rect 28132 7216 28138 7228
rect 34054 7216 34060 7228
rect 34112 7216 34118 7268
rect 30558 7188 30564 7200
rect 27632 7160 30564 7188
rect 30558 7148 30564 7160
rect 30616 7148 30622 7200
rect 1104 7098 38272 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 38272 7098
rect 1104 7024 38272 7046
rect 3970 6944 3976 6996
rect 4028 6984 4034 6996
rect 4028 6956 5580 6984
rect 4028 6944 4034 6956
rect 4249 6851 4307 6857
rect 4249 6817 4261 6851
rect 4295 6848 4307 6851
rect 4614 6848 4620 6860
rect 4295 6820 4620 6848
rect 4295 6817 4307 6820
rect 4249 6811 4307 6817
rect 4614 6808 4620 6820
rect 4672 6808 4678 6860
rect 5552 6848 5580 6956
rect 5994 6944 6000 6996
rect 6052 6944 6058 6996
rect 12342 6944 12348 6996
rect 12400 6944 12406 6996
rect 12805 6987 12863 6993
rect 12805 6953 12817 6987
rect 12851 6984 12863 6987
rect 13538 6984 13544 6996
rect 12851 6956 13544 6984
rect 12851 6953 12863 6956
rect 12805 6947 12863 6953
rect 13538 6944 13544 6956
rect 13596 6944 13602 6996
rect 15562 6944 15568 6996
rect 15620 6984 15626 6996
rect 15730 6987 15788 6993
rect 15730 6984 15742 6987
rect 15620 6956 15742 6984
rect 15620 6944 15626 6956
rect 15730 6953 15742 6956
rect 15776 6953 15788 6987
rect 15730 6947 15788 6953
rect 17221 6987 17279 6993
rect 17221 6953 17233 6987
rect 17267 6984 17279 6987
rect 17770 6984 17776 6996
rect 17267 6956 17776 6984
rect 17267 6953 17279 6956
rect 17221 6947 17279 6953
rect 17770 6944 17776 6956
rect 17828 6944 17834 6996
rect 18046 6944 18052 6996
rect 18104 6944 18110 6996
rect 21266 6944 21272 6996
rect 21324 6944 21330 6996
rect 23198 6944 23204 6996
rect 23256 6944 23262 6996
rect 23842 6944 23848 6996
rect 23900 6944 23906 6996
rect 25406 6944 25412 6996
rect 25464 6944 25470 6996
rect 30374 6984 30380 6996
rect 27080 6956 30380 6984
rect 11146 6876 11152 6928
rect 11204 6916 11210 6928
rect 11204 6888 12434 6916
rect 11204 6876 11210 6888
rect 12406 6848 12434 6888
rect 17310 6876 17316 6928
rect 17368 6916 17374 6928
rect 17681 6919 17739 6925
rect 17681 6916 17693 6919
rect 17368 6888 17693 6916
rect 17368 6876 17374 6888
rect 17681 6885 17693 6888
rect 17727 6916 17739 6919
rect 17727 6888 18460 6916
rect 17727 6885 17739 6888
rect 17681 6879 17739 6885
rect 12621 6851 12679 6857
rect 12621 6848 12633 6851
rect 5552 6820 5764 6848
rect 12406 6820 12633 6848
rect 4522 6672 4528 6724
rect 4580 6672 4586 6724
rect 5736 6712 5764 6820
rect 12621 6817 12633 6820
rect 12667 6848 12679 6851
rect 13722 6848 13728 6860
rect 12667 6820 13728 6848
rect 12667 6817 12679 6820
rect 12621 6811 12679 6817
rect 13722 6808 13728 6820
rect 13780 6808 13786 6860
rect 15473 6851 15531 6857
rect 15473 6817 15485 6851
rect 15519 6848 15531 6851
rect 15746 6848 15752 6860
rect 15519 6820 15752 6848
rect 15519 6817 15531 6820
rect 15473 6811 15531 6817
rect 15746 6808 15752 6820
rect 15804 6808 15810 6860
rect 17862 6808 17868 6860
rect 17920 6848 17926 6860
rect 18432 6848 18460 6888
rect 17920 6820 18368 6848
rect 17920 6808 17926 6820
rect 8202 6740 8208 6792
rect 8260 6780 8266 6792
rect 8941 6783 8999 6789
rect 8941 6780 8953 6783
rect 8260 6752 8953 6780
rect 8260 6740 8266 6752
rect 8941 6749 8953 6752
rect 8987 6749 8999 6783
rect 8941 6743 8999 6749
rect 9125 6783 9183 6789
rect 9125 6749 9137 6783
rect 9171 6780 9183 6783
rect 9490 6780 9496 6792
rect 9171 6752 9496 6780
rect 9171 6749 9183 6752
rect 9125 6743 9183 6749
rect 9490 6740 9496 6752
rect 9548 6740 9554 6792
rect 10686 6740 10692 6792
rect 10744 6780 10750 6792
rect 12802 6780 12808 6792
rect 10744 6752 12808 6780
rect 10744 6740 10750 6752
rect 12802 6740 12808 6752
rect 12860 6740 12866 6792
rect 12894 6740 12900 6792
rect 12952 6740 12958 6792
rect 15194 6740 15200 6792
rect 15252 6740 15258 6792
rect 17589 6783 17647 6789
rect 17589 6749 17601 6783
rect 17635 6749 17647 6783
rect 17589 6743 17647 6749
rect 17957 6783 18015 6789
rect 17957 6749 17969 6783
rect 18003 6780 18015 6783
rect 18141 6783 18199 6789
rect 18141 6780 18153 6783
rect 18003 6752 18153 6780
rect 18003 6749 18015 6752
rect 17957 6743 18015 6749
rect 18141 6749 18153 6752
rect 18187 6780 18199 6783
rect 18230 6780 18236 6792
rect 18187 6752 18236 6780
rect 18187 6749 18199 6752
rect 18141 6743 18199 6749
rect 6454 6712 6460 6724
rect 5736 6698 6460 6712
rect 5750 6684 6460 6698
rect 6454 6672 6460 6684
rect 6512 6712 6518 6724
rect 6512 6684 8340 6712
rect 6512 6672 6518 6684
rect 8312 6656 8340 6684
rect 16758 6672 16764 6724
rect 16816 6672 16822 6724
rect 17604 6712 17632 6743
rect 18230 6740 18236 6752
rect 18288 6740 18294 6792
rect 18340 6789 18368 6820
rect 18432 6820 19012 6848
rect 18432 6789 18460 6820
rect 18984 6792 19012 6820
rect 19978 6808 19984 6860
rect 20036 6808 20042 6860
rect 20441 6851 20499 6857
rect 20441 6817 20453 6851
rect 20487 6848 20499 6851
rect 21284 6848 21312 6944
rect 23216 6916 23244 6944
rect 23860 6916 23888 6944
rect 27080 6916 27108 6956
rect 30374 6944 30380 6956
rect 30432 6944 30438 6996
rect 30834 6984 30840 6996
rect 30576 6956 30840 6984
rect 30576 6916 30604 6956
rect 30834 6944 30840 6956
rect 30892 6944 30898 6996
rect 31294 6944 31300 6996
rect 31352 6944 31358 6996
rect 31386 6944 31392 6996
rect 31444 6984 31450 6996
rect 31481 6987 31539 6993
rect 31481 6984 31493 6987
rect 31444 6956 31493 6984
rect 31444 6944 31450 6956
rect 31481 6953 31493 6956
rect 31527 6953 31539 6987
rect 31481 6947 31539 6953
rect 31938 6944 31944 6996
rect 31996 6944 32002 6996
rect 23216 6888 23612 6916
rect 23860 6888 27108 6916
rect 27172 6888 28304 6916
rect 20487 6820 21312 6848
rect 20487 6817 20499 6820
rect 20441 6811 20499 6817
rect 18325 6783 18383 6789
rect 18325 6749 18337 6783
rect 18371 6749 18383 6783
rect 18325 6743 18383 6749
rect 18417 6783 18475 6789
rect 18417 6749 18429 6783
rect 18463 6749 18475 6783
rect 18417 6743 18475 6749
rect 18506 6740 18512 6792
rect 18564 6740 18570 6792
rect 18966 6740 18972 6792
rect 19024 6740 19030 6792
rect 20073 6783 20131 6789
rect 20073 6749 20085 6783
rect 20119 6780 20131 6783
rect 20622 6780 20628 6792
rect 20119 6752 20628 6780
rect 20119 6749 20131 6752
rect 20073 6743 20131 6749
rect 20622 6740 20628 6752
rect 20680 6740 20686 6792
rect 21177 6783 21235 6789
rect 21177 6749 21189 6783
rect 21223 6749 21235 6783
rect 21177 6743 21235 6749
rect 18524 6712 18552 6740
rect 17604 6684 18552 6712
rect 18785 6715 18843 6721
rect 18785 6681 18797 6715
rect 18831 6712 18843 6715
rect 21192 6712 21220 6743
rect 21266 6740 21272 6792
rect 21324 6740 21330 6792
rect 21358 6740 21364 6792
rect 21416 6780 21422 6792
rect 21453 6783 21511 6789
rect 21453 6780 21465 6783
rect 21416 6752 21465 6780
rect 21416 6740 21422 6752
rect 21453 6749 21465 6752
rect 21499 6749 21511 6783
rect 21453 6743 21511 6749
rect 22094 6712 22100 6724
rect 18831 6684 22100 6712
rect 18831 6681 18843 6684
rect 18785 6675 18843 6681
rect 22094 6672 22100 6684
rect 22152 6672 22158 6724
rect 23584 6712 23612 6888
rect 24854 6808 24860 6860
rect 24912 6808 24918 6860
rect 26602 6848 26608 6860
rect 26160 6820 26608 6848
rect 24946 6740 24952 6792
rect 25004 6740 25010 6792
rect 25685 6783 25743 6789
rect 25685 6780 25697 6783
rect 25056 6752 25697 6780
rect 25056 6712 25084 6752
rect 25685 6749 25697 6752
rect 25731 6749 25743 6783
rect 25685 6743 25743 6749
rect 25961 6783 26019 6789
rect 25961 6749 25973 6783
rect 26007 6780 26019 6783
rect 26050 6780 26056 6792
rect 26007 6752 26056 6780
rect 26007 6749 26019 6752
rect 25961 6743 26019 6749
rect 26050 6740 26056 6752
rect 26108 6740 26114 6792
rect 26160 6789 26188 6820
rect 26602 6808 26608 6820
rect 26660 6808 26666 6860
rect 27065 6851 27123 6857
rect 27065 6848 27077 6851
rect 26896 6820 27077 6848
rect 26145 6783 26203 6789
rect 26145 6749 26157 6783
rect 26191 6749 26203 6783
rect 26145 6743 26203 6749
rect 26234 6740 26240 6792
rect 26292 6740 26298 6792
rect 26329 6783 26387 6789
rect 26329 6749 26341 6783
rect 26375 6749 26387 6783
rect 26896 6780 26924 6820
rect 27065 6817 27077 6820
rect 27111 6848 27123 6851
rect 27172 6848 27200 6888
rect 27111 6820 27200 6848
rect 27249 6851 27307 6857
rect 27111 6817 27123 6820
rect 27065 6811 27123 6817
rect 27249 6817 27261 6851
rect 27295 6848 27307 6851
rect 27798 6848 27804 6860
rect 27295 6820 27804 6848
rect 27295 6817 27307 6820
rect 27249 6811 27307 6817
rect 27798 6808 27804 6820
rect 27856 6808 27862 6860
rect 28276 6848 28304 6888
rect 30300 6888 30604 6916
rect 30653 6919 30711 6925
rect 28442 6848 28448 6860
rect 27908 6820 28212 6848
rect 28276 6820 28448 6848
rect 26329 6743 26387 6749
rect 26528 6752 26924 6780
rect 23584 6684 25084 6712
rect 25409 6715 25467 6721
rect 25409 6681 25421 6715
rect 25455 6712 25467 6715
rect 25498 6712 25504 6724
rect 25455 6684 25504 6712
rect 25455 6681 25467 6684
rect 25409 6675 25467 6681
rect 25498 6672 25504 6684
rect 25556 6712 25562 6724
rect 26344 6712 26372 6743
rect 25556 6684 26372 6712
rect 25556 6672 25562 6684
rect 8294 6604 8300 6656
rect 8352 6604 8358 6656
rect 9030 6604 9036 6656
rect 9088 6604 9094 6656
rect 14550 6604 14556 6656
rect 14608 6604 14614 6656
rect 21637 6647 21695 6653
rect 21637 6613 21649 6647
rect 21683 6644 21695 6647
rect 22370 6644 22376 6656
rect 21683 6616 22376 6644
rect 21683 6613 21695 6616
rect 21637 6607 21695 6613
rect 22370 6604 22376 6616
rect 22428 6604 22434 6656
rect 23566 6604 23572 6656
rect 23624 6644 23630 6656
rect 23842 6644 23848 6656
rect 23624 6616 23848 6644
rect 23624 6604 23630 6616
rect 23842 6604 23848 6616
rect 23900 6604 23906 6656
rect 25314 6604 25320 6656
rect 25372 6604 25378 6656
rect 25593 6647 25651 6653
rect 25593 6613 25605 6647
rect 25639 6644 25651 6647
rect 26528 6644 26556 6752
rect 26970 6740 26976 6792
rect 27028 6740 27034 6792
rect 27430 6780 27436 6792
rect 27172 6752 27436 6780
rect 27172 6712 27200 6752
rect 27430 6740 27436 6752
rect 27488 6740 27494 6792
rect 27908 6789 27936 6820
rect 28184 6792 28212 6820
rect 28442 6808 28448 6820
rect 28500 6808 28506 6860
rect 28534 6808 28540 6860
rect 28592 6808 28598 6860
rect 28626 6808 28632 6860
rect 28684 6848 28690 6860
rect 30300 6848 30328 6888
rect 30653 6885 30665 6919
rect 30699 6916 30711 6919
rect 31312 6916 31340 6944
rect 31956 6916 31984 6944
rect 30699 6888 31340 6916
rect 31772 6888 31984 6916
rect 30699 6885 30711 6888
rect 30653 6879 30711 6885
rect 28684 6820 30328 6848
rect 28684 6808 28690 6820
rect 30558 6808 30564 6860
rect 30616 6848 30622 6860
rect 30616 6820 30880 6848
rect 30616 6808 30622 6820
rect 27525 6783 27583 6789
rect 27525 6749 27537 6783
rect 27571 6749 27583 6783
rect 27525 6743 27583 6749
rect 27618 6783 27676 6789
rect 27618 6749 27630 6783
rect 27664 6749 27676 6783
rect 27618 6743 27676 6749
rect 27893 6783 27951 6789
rect 27893 6749 27905 6783
rect 27939 6749 27951 6783
rect 27893 6743 27951 6749
rect 26620 6684 27200 6712
rect 27249 6715 27307 6721
rect 26620 6653 26648 6684
rect 27249 6681 27261 6715
rect 27295 6712 27307 6715
rect 27540 6712 27568 6743
rect 27295 6684 27568 6712
rect 27295 6681 27307 6684
rect 27249 6675 27307 6681
rect 25639 6616 26556 6644
rect 26605 6647 26663 6653
rect 25639 6613 25651 6616
rect 25593 6607 25651 6613
rect 26605 6613 26617 6647
rect 26651 6613 26663 6647
rect 26605 6607 26663 6613
rect 26694 6604 26700 6656
rect 26752 6644 26758 6656
rect 27632 6644 27660 6743
rect 27982 6740 27988 6792
rect 28040 6789 28046 6792
rect 28040 6743 28048 6789
rect 28040 6740 28046 6743
rect 28166 6740 28172 6792
rect 28224 6740 28230 6792
rect 28258 6740 28264 6792
rect 28316 6740 28322 6792
rect 28353 6783 28411 6789
rect 28353 6749 28365 6783
rect 28399 6749 28411 6783
rect 28353 6743 28411 6749
rect 27801 6715 27859 6721
rect 27801 6681 27813 6715
rect 27847 6712 27859 6715
rect 28074 6712 28080 6724
rect 27847 6684 28080 6712
rect 27847 6681 27859 6684
rect 27801 6675 27859 6681
rect 28074 6672 28080 6684
rect 28132 6672 28138 6724
rect 28368 6712 28396 6743
rect 28810 6740 28816 6792
rect 28868 6780 28874 6792
rect 29917 6783 29975 6789
rect 29917 6780 29929 6783
rect 28868 6752 29929 6780
rect 28868 6740 28874 6752
rect 29917 6749 29929 6752
rect 29963 6749 29975 6783
rect 29917 6743 29975 6749
rect 30006 6740 30012 6792
rect 30064 6780 30070 6792
rect 30101 6783 30159 6789
rect 30101 6780 30113 6783
rect 30064 6752 30113 6780
rect 30064 6740 30070 6752
rect 30101 6749 30113 6752
rect 30147 6749 30159 6783
rect 30101 6743 30159 6749
rect 30377 6783 30435 6789
rect 30377 6749 30389 6783
rect 30423 6780 30435 6783
rect 30466 6780 30472 6792
rect 30423 6752 30472 6780
rect 30423 6749 30435 6752
rect 30377 6743 30435 6749
rect 30466 6740 30472 6752
rect 30524 6740 30530 6792
rect 30742 6740 30748 6792
rect 30800 6740 30806 6792
rect 30852 6789 30880 6820
rect 31772 6792 31800 6888
rect 32490 6876 32496 6928
rect 32548 6916 32554 6928
rect 32548 6888 33088 6916
rect 32548 6876 32554 6888
rect 32769 6851 32827 6857
rect 32769 6848 32781 6851
rect 31956 6820 32781 6848
rect 30837 6783 30895 6789
rect 30837 6749 30849 6783
rect 30883 6749 30895 6783
rect 30837 6743 30895 6749
rect 31754 6740 31760 6792
rect 31812 6740 31818 6792
rect 31846 6740 31852 6792
rect 31904 6740 31910 6792
rect 31956 6789 31984 6820
rect 32232 6792 32260 6820
rect 32769 6817 32781 6820
rect 32815 6817 32827 6851
rect 32769 6811 32827 6817
rect 32858 6808 32864 6860
rect 32916 6848 32922 6860
rect 32953 6851 33011 6857
rect 32953 6848 32965 6851
rect 32916 6820 32965 6848
rect 32916 6808 32922 6820
rect 32953 6817 32965 6820
rect 32999 6817 33011 6851
rect 33060 6848 33088 6888
rect 33137 6851 33195 6857
rect 33137 6848 33149 6851
rect 33060 6820 33149 6848
rect 32953 6811 33011 6817
rect 33137 6817 33149 6820
rect 33183 6817 33195 6851
rect 33137 6811 33195 6817
rect 31941 6783 31999 6789
rect 31941 6749 31953 6783
rect 31987 6749 31999 6783
rect 31941 6743 31999 6749
rect 32122 6740 32128 6792
rect 32180 6740 32186 6792
rect 32214 6740 32220 6792
rect 32272 6740 32278 6792
rect 32493 6783 32551 6789
rect 32493 6749 32505 6783
rect 32539 6749 32551 6783
rect 32493 6743 32551 6749
rect 28184 6684 28396 6712
rect 28184 6653 28212 6684
rect 28442 6672 28448 6724
rect 28500 6712 28506 6724
rect 32508 6712 32536 6743
rect 32582 6740 32588 6792
rect 32640 6740 32646 6792
rect 32677 6783 32735 6789
rect 32677 6749 32689 6783
rect 32723 6749 32735 6783
rect 32677 6743 32735 6749
rect 28500 6684 32536 6712
rect 28500 6672 28506 6684
rect 32692 6656 32720 6743
rect 33042 6740 33048 6792
rect 33100 6780 33106 6792
rect 33229 6783 33287 6789
rect 33229 6780 33241 6783
rect 33100 6752 33241 6780
rect 33100 6740 33106 6752
rect 33229 6749 33241 6752
rect 33275 6749 33287 6783
rect 33229 6743 33287 6749
rect 34422 6672 34428 6724
rect 34480 6672 34486 6724
rect 26752 6616 27660 6644
rect 28169 6647 28227 6653
rect 26752 6604 26758 6616
rect 28169 6613 28181 6647
rect 28215 6613 28227 6647
rect 28169 6607 28227 6613
rect 28350 6604 28356 6656
rect 28408 6644 28414 6656
rect 28721 6647 28779 6653
rect 28721 6644 28733 6647
rect 28408 6616 28733 6644
rect 28408 6604 28414 6616
rect 28721 6613 28733 6616
rect 28767 6613 28779 6647
rect 28721 6607 28779 6613
rect 32674 6604 32680 6656
rect 32732 6604 32738 6656
rect 33597 6647 33655 6653
rect 33597 6613 33609 6647
rect 33643 6644 33655 6647
rect 34440 6644 34468 6672
rect 33643 6616 34468 6644
rect 33643 6613 33655 6616
rect 33597 6607 33655 6613
rect 1104 6554 38272 6576
rect 1104 6502 4874 6554
rect 4926 6502 4938 6554
rect 4990 6502 5002 6554
rect 5054 6502 5066 6554
rect 5118 6502 5130 6554
rect 5182 6502 35594 6554
rect 35646 6502 35658 6554
rect 35710 6502 35722 6554
rect 35774 6502 35786 6554
rect 35838 6502 35850 6554
rect 35902 6502 38272 6554
rect 1104 6480 38272 6502
rect 4522 6400 4528 6452
rect 4580 6440 4586 6452
rect 4709 6443 4767 6449
rect 4709 6440 4721 6443
rect 4580 6412 4721 6440
rect 4580 6400 4586 6412
rect 4709 6409 4721 6412
rect 4755 6409 4767 6443
rect 4709 6403 4767 6409
rect 4798 6400 4804 6452
rect 4856 6400 4862 6452
rect 7837 6443 7895 6449
rect 7837 6409 7849 6443
rect 7883 6440 7895 6443
rect 9490 6440 9496 6452
rect 7883 6412 9496 6440
rect 7883 6409 7895 6412
rect 7837 6403 7895 6409
rect 9490 6400 9496 6412
rect 9548 6400 9554 6452
rect 14458 6440 14464 6452
rect 14016 6412 14464 6440
rect 4816 6304 4844 6400
rect 7745 6375 7803 6381
rect 7745 6341 7757 6375
rect 7791 6372 7803 6375
rect 8846 6372 8852 6384
rect 7791 6344 8852 6372
rect 7791 6341 7803 6344
rect 7745 6335 7803 6341
rect 8846 6332 8852 6344
rect 8904 6332 8910 6384
rect 9398 6332 9404 6384
rect 9456 6372 9462 6384
rect 9953 6375 10011 6381
rect 9953 6372 9965 6375
rect 9456 6344 9965 6372
rect 9456 6332 9462 6344
rect 9953 6341 9965 6344
rect 9999 6341 10011 6375
rect 9953 6335 10011 6341
rect 11054 6332 11060 6384
rect 11112 6372 11118 6384
rect 13357 6375 13415 6381
rect 13357 6372 13369 6375
rect 11112 6344 13369 6372
rect 11112 6332 11118 6344
rect 13357 6341 13369 6344
rect 13403 6341 13415 6375
rect 13357 6335 13415 6341
rect 4893 6307 4951 6313
rect 4893 6304 4905 6307
rect 4816 6276 4905 6304
rect 4893 6273 4905 6276
rect 4939 6273 4951 6307
rect 4893 6267 4951 6273
rect 8202 6264 8208 6316
rect 8260 6304 8266 6316
rect 8389 6307 8447 6313
rect 8389 6304 8401 6307
rect 8260 6276 8401 6304
rect 8260 6264 8266 6276
rect 8389 6273 8401 6276
rect 8435 6273 8447 6307
rect 8389 6267 8447 6273
rect 9493 6307 9551 6313
rect 9493 6273 9505 6307
rect 9539 6273 9551 6307
rect 9493 6267 9551 6273
rect 9677 6307 9735 6313
rect 9677 6273 9689 6307
rect 9723 6304 9735 6307
rect 10045 6307 10103 6313
rect 10045 6304 10057 6307
rect 9723 6276 10057 6304
rect 9723 6273 9735 6276
rect 9677 6267 9735 6273
rect 10045 6273 10057 6276
rect 10091 6304 10103 6307
rect 10226 6304 10232 6316
rect 10091 6276 10232 6304
rect 10091 6273 10103 6276
rect 10045 6267 10103 6273
rect 7466 6196 7472 6248
rect 7524 6236 7530 6248
rect 7929 6239 7987 6245
rect 7929 6236 7941 6239
rect 7524 6208 7941 6236
rect 7524 6196 7530 6208
rect 7929 6205 7941 6208
rect 7975 6236 7987 6239
rect 8573 6239 8631 6245
rect 8573 6236 8585 6239
rect 7975 6208 8585 6236
rect 7975 6205 7987 6208
rect 7929 6199 7987 6205
rect 8573 6205 8585 6208
rect 8619 6205 8631 6239
rect 8573 6199 8631 6205
rect 8665 6239 8723 6245
rect 8665 6205 8677 6239
rect 8711 6236 8723 6239
rect 8757 6239 8815 6245
rect 8757 6236 8769 6239
rect 8711 6208 8769 6236
rect 8711 6205 8723 6208
rect 8665 6199 8723 6205
rect 8757 6205 8769 6208
rect 8803 6205 8815 6239
rect 8757 6199 8815 6205
rect 8588 6168 8616 6199
rect 9306 6196 9312 6248
rect 9364 6196 9370 6248
rect 9508 6236 9536 6267
rect 10226 6264 10232 6276
rect 10284 6304 10290 6316
rect 12253 6307 12311 6313
rect 12253 6304 12265 6307
rect 10284 6276 12265 6304
rect 10284 6264 10290 6276
rect 12253 6273 12265 6276
rect 12299 6273 12311 6307
rect 12253 6267 12311 6273
rect 12437 6307 12495 6313
rect 12437 6273 12449 6307
rect 12483 6304 12495 6307
rect 12529 6307 12587 6313
rect 12529 6304 12541 6307
rect 12483 6276 12541 6304
rect 12483 6273 12495 6276
rect 12437 6267 12495 6273
rect 12529 6273 12541 6276
rect 12575 6273 12587 6307
rect 12529 6267 12587 6273
rect 12805 6307 12863 6313
rect 12805 6273 12817 6307
rect 12851 6304 12863 6307
rect 13538 6304 13544 6316
rect 12851 6276 13544 6304
rect 12851 6273 12863 6276
rect 12805 6267 12863 6273
rect 9766 6236 9772 6248
rect 9508 6208 9772 6236
rect 9766 6196 9772 6208
rect 9824 6236 9830 6248
rect 12069 6239 12127 6245
rect 12069 6236 12081 6239
rect 9824 6208 12081 6236
rect 9824 6196 9830 6208
rect 12069 6205 12081 6208
rect 12115 6205 12127 6239
rect 12268 6236 12296 6267
rect 13538 6264 13544 6276
rect 13596 6264 13602 6316
rect 14016 6313 14044 6412
rect 14458 6400 14464 6412
rect 14516 6440 14522 6452
rect 15289 6443 15347 6449
rect 15289 6440 15301 6443
rect 14516 6412 15301 6440
rect 14516 6400 14522 6412
rect 15289 6409 15301 6412
rect 15335 6409 15347 6443
rect 15289 6403 15347 6409
rect 15470 6400 15476 6452
rect 15528 6400 15534 6452
rect 17862 6400 17868 6452
rect 17920 6400 17926 6452
rect 18690 6400 18696 6452
rect 18748 6400 18754 6452
rect 19610 6400 19616 6452
rect 19668 6400 19674 6452
rect 19794 6400 19800 6452
rect 19852 6400 19858 6452
rect 19889 6443 19947 6449
rect 19889 6409 19901 6443
rect 19935 6440 19947 6443
rect 19978 6440 19984 6452
rect 19935 6412 19984 6440
rect 19935 6409 19947 6412
rect 19889 6403 19947 6409
rect 19978 6400 19984 6412
rect 20036 6400 20042 6452
rect 22373 6443 22431 6449
rect 22373 6409 22385 6443
rect 22419 6440 22431 6443
rect 22738 6440 22744 6452
rect 22419 6412 22744 6440
rect 22419 6409 22431 6412
rect 22373 6403 22431 6409
rect 15378 6372 15384 6384
rect 15028 6344 15384 6372
rect 15028 6313 15056 6344
rect 15378 6332 15384 6344
rect 15436 6332 15442 6384
rect 14001 6307 14059 6313
rect 14001 6273 14013 6307
rect 14047 6273 14059 6307
rect 14001 6267 14059 6273
rect 14093 6307 14151 6313
rect 14093 6273 14105 6307
rect 14139 6273 14151 6307
rect 14093 6267 14151 6273
rect 15013 6307 15071 6313
rect 15013 6273 15025 6307
rect 15059 6273 15071 6307
rect 15013 6267 15071 6273
rect 13556 6236 13584 6264
rect 14108 6236 14136 6267
rect 15194 6264 15200 6316
rect 15252 6264 15258 6316
rect 15286 6264 15292 6316
rect 15344 6264 15350 6316
rect 15488 6304 15516 6400
rect 17880 6372 17908 6400
rect 18506 6372 18512 6384
rect 17880 6344 18276 6372
rect 15565 6307 15623 6313
rect 15565 6304 15577 6307
rect 15488 6276 15577 6304
rect 15565 6273 15577 6276
rect 15611 6273 15623 6307
rect 15565 6267 15623 6273
rect 18049 6307 18107 6313
rect 18049 6273 18061 6307
rect 18095 6304 18107 6307
rect 18138 6304 18144 6316
rect 18095 6276 18144 6304
rect 18095 6273 18107 6276
rect 18049 6267 18107 6273
rect 18138 6264 18144 6276
rect 18196 6264 18202 6316
rect 18248 6313 18276 6344
rect 18432 6344 18512 6372
rect 18432 6313 18460 6344
rect 18506 6332 18512 6344
rect 18564 6372 18570 6384
rect 19061 6375 19119 6381
rect 19061 6372 19073 6375
rect 18564 6344 19073 6372
rect 18564 6332 18570 6344
rect 19061 6341 19073 6344
rect 19107 6341 19119 6375
rect 19061 6335 19119 6341
rect 18233 6307 18291 6313
rect 18233 6273 18245 6307
rect 18279 6273 18291 6307
rect 18233 6267 18291 6273
rect 18325 6307 18383 6313
rect 18325 6273 18337 6307
rect 18371 6273 18383 6307
rect 18325 6267 18383 6273
rect 18417 6307 18475 6313
rect 18417 6273 18429 6307
rect 18463 6273 18475 6307
rect 18417 6267 18475 6273
rect 18877 6307 18935 6313
rect 18877 6273 18889 6307
rect 18923 6304 18935 6307
rect 18966 6304 18972 6316
rect 18923 6276 18972 6304
rect 18923 6273 18935 6276
rect 18877 6267 18935 6273
rect 12268 6208 12572 6236
rect 13556 6208 14136 6236
rect 14829 6239 14887 6245
rect 12069 6199 12127 6205
rect 9677 6171 9735 6177
rect 9677 6168 9689 6171
rect 8588 6140 9689 6168
rect 9677 6137 9689 6140
rect 9723 6137 9735 6171
rect 12084 6168 12112 6199
rect 12342 6168 12348 6180
rect 12084 6140 12348 6168
rect 9677 6131 9735 6137
rect 12342 6128 12348 6140
rect 12400 6128 12406 6180
rect 12544 6112 12572 6208
rect 14829 6205 14841 6239
rect 14875 6236 14887 6239
rect 15212 6236 15240 6264
rect 14875 6208 15240 6236
rect 15304 6236 15332 6264
rect 15381 6239 15439 6245
rect 15381 6236 15393 6239
rect 15304 6208 15393 6236
rect 14875 6205 14887 6208
rect 14829 6199 14887 6205
rect 15381 6205 15393 6208
rect 15427 6205 15439 6239
rect 18156 6236 18184 6264
rect 18340 6236 18368 6267
rect 18156 6208 18368 6236
rect 15381 6199 15439 6205
rect 18138 6128 18144 6180
rect 18196 6128 18202 6180
rect 7374 6060 7380 6112
rect 7432 6060 7438 6112
rect 8202 6060 8208 6112
rect 8260 6060 8266 6112
rect 8846 6060 8852 6112
rect 8904 6100 8910 6112
rect 9490 6100 9496 6112
rect 8904 6072 9496 6100
rect 8904 6060 8910 6072
rect 9490 6060 9496 6072
rect 9548 6060 9554 6112
rect 12526 6060 12532 6112
rect 12584 6060 12590 6112
rect 15657 6103 15715 6109
rect 15657 6069 15669 6103
rect 15703 6100 15715 6103
rect 16482 6100 16488 6112
rect 15703 6072 16488 6100
rect 15703 6069 15715 6072
rect 15657 6063 15715 6069
rect 16482 6060 16488 6072
rect 16540 6060 16546 6112
rect 18509 6103 18567 6109
rect 18509 6069 18521 6103
rect 18555 6100 18567 6103
rect 18892 6100 18920 6267
rect 18966 6264 18972 6276
rect 19024 6264 19030 6316
rect 19628 6304 19656 6400
rect 19705 6307 19763 6313
rect 19705 6304 19717 6307
rect 19628 6276 19717 6304
rect 19705 6273 19717 6276
rect 19751 6273 19763 6307
rect 19812 6304 19840 6400
rect 19889 6307 19947 6313
rect 19889 6304 19901 6307
rect 19812 6276 19901 6304
rect 19705 6267 19763 6273
rect 19889 6273 19901 6276
rect 19935 6273 19947 6307
rect 19889 6267 19947 6273
rect 22572 6168 22600 6412
rect 22738 6400 22744 6412
rect 22796 6400 22802 6452
rect 23753 6443 23811 6449
rect 23753 6409 23765 6443
rect 23799 6409 23811 6443
rect 23753 6403 23811 6409
rect 24219 6443 24277 6449
rect 24219 6409 24231 6443
rect 24265 6440 24277 6443
rect 24946 6440 24952 6452
rect 24265 6412 24952 6440
rect 24265 6409 24277 6412
rect 24219 6403 24277 6409
rect 22922 6332 22928 6384
rect 22980 6372 22986 6384
rect 23385 6375 23443 6381
rect 23385 6372 23397 6375
rect 22980 6344 23397 6372
rect 22980 6332 22986 6344
rect 23385 6341 23397 6344
rect 23431 6341 23443 6375
rect 23385 6335 23443 6341
rect 23474 6332 23480 6384
rect 23532 6332 23538 6384
rect 23768 6372 23796 6403
rect 24946 6400 24952 6412
rect 25004 6400 25010 6452
rect 25222 6400 25228 6452
rect 25280 6440 25286 6452
rect 25501 6443 25559 6449
rect 25501 6440 25513 6443
rect 25280 6412 25513 6440
rect 25280 6400 25286 6412
rect 25501 6409 25513 6412
rect 25547 6409 25559 6443
rect 25501 6403 25559 6409
rect 27982 6400 27988 6452
rect 28040 6400 28046 6452
rect 28166 6400 28172 6452
rect 28224 6440 28230 6452
rect 31018 6440 31024 6452
rect 28224 6412 31024 6440
rect 28224 6400 28230 6412
rect 31018 6400 31024 6412
rect 31076 6400 31082 6452
rect 32490 6440 32496 6452
rect 31726 6412 32496 6440
rect 24121 6375 24179 6381
rect 24121 6372 24133 6375
rect 23768 6344 24133 6372
rect 24121 6341 24133 6344
rect 24167 6341 24179 6375
rect 24121 6335 24179 6341
rect 25314 6332 25320 6384
rect 25372 6372 25378 6384
rect 31726 6372 31754 6412
rect 32490 6400 32496 6412
rect 32548 6400 32554 6452
rect 32582 6400 32588 6452
rect 32640 6400 32646 6452
rect 25372 6344 31754 6372
rect 32600 6372 32628 6400
rect 32769 6375 32827 6381
rect 32769 6372 32781 6375
rect 32600 6344 32781 6372
rect 25372 6332 25378 6344
rect 32769 6341 32781 6344
rect 32815 6341 32827 6375
rect 32769 6335 32827 6341
rect 22646 6264 22652 6316
rect 22704 6264 22710 6316
rect 22741 6307 22799 6313
rect 22741 6273 22753 6307
rect 22787 6304 22799 6307
rect 23106 6304 23112 6316
rect 22787 6276 23112 6304
rect 22787 6273 22799 6276
rect 22741 6267 22799 6273
rect 23106 6264 23112 6276
rect 23164 6304 23170 6316
rect 23201 6307 23259 6313
rect 23201 6304 23213 6307
rect 23164 6276 23213 6304
rect 23164 6264 23170 6276
rect 23201 6273 23213 6276
rect 23247 6273 23259 6307
rect 23201 6267 23259 6273
rect 23566 6264 23572 6316
rect 23624 6264 23630 6316
rect 24302 6264 24308 6316
rect 24360 6264 24366 6316
rect 24397 6307 24455 6313
rect 24397 6273 24409 6307
rect 24443 6273 24455 6307
rect 24397 6267 24455 6273
rect 22664 6236 22692 6264
rect 22833 6239 22891 6245
rect 22833 6236 22845 6239
rect 22664 6208 22845 6236
rect 22833 6205 22845 6208
rect 22879 6205 22891 6239
rect 24412 6236 24440 6267
rect 24762 6264 24768 6316
rect 24820 6304 24826 6316
rect 25409 6307 25467 6313
rect 25409 6304 25421 6307
rect 24820 6276 25421 6304
rect 24820 6264 24826 6276
rect 25409 6273 25421 6276
rect 25455 6273 25467 6307
rect 25409 6267 25467 6273
rect 25593 6307 25651 6313
rect 25593 6273 25605 6307
rect 25639 6304 25651 6307
rect 26050 6304 26056 6316
rect 25639 6276 26056 6304
rect 25639 6273 25651 6276
rect 25593 6267 25651 6273
rect 26050 6264 26056 6276
rect 26108 6264 26114 6316
rect 27798 6304 27804 6316
rect 27448 6276 27804 6304
rect 22833 6199 22891 6205
rect 23308 6208 24440 6236
rect 23308 6180 23336 6208
rect 22572 6140 23244 6168
rect 18555 6072 18920 6100
rect 19245 6103 19303 6109
rect 18555 6069 18567 6072
rect 18509 6063 18567 6069
rect 19245 6069 19257 6103
rect 19291 6100 19303 6103
rect 19518 6100 19524 6112
rect 19291 6072 19524 6100
rect 19291 6069 19303 6072
rect 19245 6063 19303 6069
rect 19518 6060 19524 6072
rect 19576 6060 19582 6112
rect 23014 6060 23020 6112
rect 23072 6060 23078 6112
rect 23216 6100 23244 6140
rect 23290 6128 23296 6180
rect 23348 6128 23354 6180
rect 27448 6100 27476 6276
rect 27798 6264 27804 6276
rect 27856 6264 27862 6316
rect 28077 6307 28135 6313
rect 28077 6273 28089 6307
rect 28123 6273 28135 6307
rect 28077 6267 28135 6273
rect 28261 6307 28319 6313
rect 28261 6273 28273 6307
rect 28307 6273 28319 6307
rect 28261 6267 28319 6273
rect 27522 6196 27528 6248
rect 27580 6236 27586 6248
rect 27580 6208 27660 6236
rect 27580 6196 27586 6208
rect 27632 6168 27660 6208
rect 27706 6196 27712 6248
rect 27764 6236 27770 6248
rect 28092 6236 28120 6267
rect 27764 6208 28120 6236
rect 27764 6196 27770 6208
rect 28276 6168 28304 6267
rect 32214 6264 32220 6316
rect 32272 6304 32278 6316
rect 32493 6307 32551 6313
rect 32493 6304 32505 6307
rect 32272 6276 32505 6304
rect 32272 6264 32278 6276
rect 32493 6273 32505 6276
rect 32539 6273 32551 6307
rect 32493 6267 32551 6273
rect 32585 6307 32643 6313
rect 32585 6273 32597 6307
rect 32631 6304 32643 6307
rect 32674 6304 32680 6316
rect 32631 6276 32680 6304
rect 32631 6273 32643 6276
rect 32585 6267 32643 6273
rect 32600 6236 32628 6267
rect 32674 6264 32680 6276
rect 32732 6264 32738 6316
rect 27632 6140 28304 6168
rect 32048 6208 32628 6236
rect 32048 6112 32076 6208
rect 32766 6128 32772 6180
rect 32824 6128 32830 6180
rect 23216 6072 27476 6100
rect 27614 6060 27620 6112
rect 27672 6060 27678 6112
rect 32030 6060 32036 6112
rect 32088 6060 32094 6112
rect 1104 6010 38272 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 38272 6010
rect 1104 5936 38272 5958
rect 8202 5856 8208 5908
rect 8260 5856 8266 5908
rect 9306 5896 9312 5908
rect 9048 5868 9312 5896
rect 4614 5720 4620 5772
rect 4672 5760 4678 5772
rect 5077 5763 5135 5769
rect 5077 5760 5089 5763
rect 4672 5732 5089 5760
rect 4672 5720 4678 5732
rect 5077 5729 5089 5732
rect 5123 5760 5135 5763
rect 6914 5760 6920 5772
rect 5123 5732 6920 5760
rect 5123 5729 5135 5732
rect 5077 5723 5135 5729
rect 6914 5720 6920 5732
rect 6972 5720 6978 5772
rect 7193 5763 7251 5769
rect 7193 5729 7205 5763
rect 7239 5760 7251 5763
rect 8220 5760 8248 5856
rect 7239 5732 8248 5760
rect 8665 5763 8723 5769
rect 7239 5729 7251 5732
rect 7193 5723 7251 5729
rect 8665 5729 8677 5763
rect 8711 5760 8723 5763
rect 9048 5760 9076 5868
rect 9306 5856 9312 5868
rect 9364 5856 9370 5908
rect 10060 5868 10732 5896
rect 9125 5831 9183 5837
rect 9125 5797 9137 5831
rect 9171 5828 9183 5831
rect 9674 5828 9680 5840
rect 9171 5800 9680 5828
rect 9171 5797 9183 5800
rect 9125 5791 9183 5797
rect 9674 5788 9680 5800
rect 9732 5788 9738 5840
rect 8711 5732 9076 5760
rect 8711 5729 8723 5732
rect 8665 5723 8723 5729
rect 6454 5652 6460 5704
rect 6512 5652 6518 5704
rect 8294 5652 8300 5704
rect 8352 5652 8358 5704
rect 9048 5701 9076 5732
rect 9309 5763 9367 5769
rect 9309 5729 9321 5763
rect 9355 5760 9367 5763
rect 9355 5732 9812 5760
rect 9355 5729 9367 5732
rect 9309 5723 9367 5729
rect 9784 5704 9812 5732
rect 9033 5695 9091 5701
rect 9033 5661 9045 5695
rect 9079 5661 9091 5695
rect 9033 5655 9091 5661
rect 9398 5652 9404 5704
rect 9456 5652 9462 5704
rect 9490 5652 9496 5704
rect 9548 5692 9554 5704
rect 9548 5664 9593 5692
rect 9548 5652 9554 5664
rect 9766 5652 9772 5704
rect 9824 5652 9830 5704
rect 9907 5695 9965 5701
rect 9907 5661 9919 5695
rect 9953 5692 9965 5695
rect 10060 5692 10088 5868
rect 10704 5840 10732 5868
rect 10778 5856 10784 5908
rect 10836 5896 10842 5908
rect 12805 5899 12863 5905
rect 12805 5896 12817 5899
rect 10836 5868 12817 5896
rect 10836 5856 10842 5868
rect 12805 5865 12817 5868
rect 12851 5896 12863 5899
rect 14090 5896 14096 5908
rect 12851 5868 14096 5896
rect 12851 5865 12863 5868
rect 12805 5859 12863 5865
rect 14090 5856 14096 5868
rect 14148 5856 14154 5908
rect 15286 5856 15292 5908
rect 15344 5896 15350 5908
rect 15703 5899 15761 5905
rect 15703 5896 15715 5899
rect 15344 5868 15715 5896
rect 15344 5856 15350 5868
rect 15703 5865 15715 5868
rect 15749 5896 15761 5899
rect 16298 5896 16304 5908
rect 15749 5868 16304 5896
rect 15749 5865 15761 5868
rect 15703 5859 15761 5865
rect 16298 5856 16304 5868
rect 16356 5856 16362 5908
rect 18138 5856 18144 5908
rect 18196 5856 18202 5908
rect 22554 5856 22560 5908
rect 22612 5896 22618 5908
rect 22649 5899 22707 5905
rect 22649 5896 22661 5899
rect 22612 5868 22661 5896
rect 22612 5856 22618 5868
rect 22649 5865 22661 5868
rect 22695 5865 22707 5899
rect 22649 5859 22707 5865
rect 27798 5856 27804 5908
rect 27856 5896 27862 5908
rect 28626 5896 28632 5908
rect 27856 5868 28632 5896
rect 27856 5856 27862 5868
rect 28626 5856 28632 5868
rect 28684 5856 28690 5908
rect 30466 5856 30472 5908
rect 30524 5856 30530 5908
rect 32030 5856 32036 5908
rect 32088 5856 32094 5908
rect 32214 5856 32220 5908
rect 32272 5856 32278 5908
rect 10686 5788 10692 5840
rect 10744 5788 10750 5840
rect 12434 5720 12440 5772
rect 12492 5760 12498 5772
rect 12529 5763 12587 5769
rect 12529 5760 12541 5763
rect 12492 5732 12541 5760
rect 12492 5720 12498 5732
rect 12529 5729 12541 5732
rect 12575 5760 12587 5763
rect 14918 5760 14924 5772
rect 12575 5732 12940 5760
rect 12575 5729 12587 5732
rect 12529 5723 12587 5729
rect 10686 5701 10692 5704
rect 9953 5664 10088 5692
rect 10137 5695 10195 5701
rect 9953 5661 9965 5664
rect 9907 5655 9965 5661
rect 10137 5661 10149 5695
rect 10183 5661 10195 5695
rect 10137 5655 10195 5661
rect 10285 5695 10343 5701
rect 10285 5661 10297 5695
rect 10331 5661 10343 5695
rect 10285 5655 10343 5661
rect 10641 5695 10692 5701
rect 10641 5661 10653 5695
rect 10687 5661 10692 5695
rect 10641 5655 10692 5661
rect 5353 5627 5411 5633
rect 5353 5593 5365 5627
rect 5399 5624 5411 5627
rect 5626 5624 5632 5636
rect 5399 5596 5632 5624
rect 5399 5593 5411 5596
rect 5353 5587 5411 5593
rect 5626 5584 5632 5596
rect 5684 5584 5690 5636
rect 9677 5627 9735 5633
rect 9677 5593 9689 5627
rect 9723 5593 9735 5627
rect 10152 5624 10180 5655
rect 9677 5587 9735 5593
rect 9876 5596 10180 5624
rect 6825 5559 6883 5565
rect 6825 5525 6837 5559
rect 6871 5556 6883 5559
rect 8202 5556 8208 5568
rect 6871 5528 8208 5556
rect 6871 5525 6883 5528
rect 6825 5519 6883 5525
rect 8202 5516 8208 5528
rect 8260 5516 8266 5568
rect 9033 5559 9091 5565
rect 9033 5525 9045 5559
rect 9079 5556 9091 5559
rect 9692 5556 9720 5587
rect 9876 5568 9904 5596
rect 9079 5528 9720 5556
rect 9079 5525 9091 5528
rect 9033 5519 9091 5525
rect 9858 5516 9864 5568
rect 9916 5516 9922 5568
rect 10042 5516 10048 5568
rect 10100 5516 10106 5568
rect 10300 5556 10328 5655
rect 10686 5652 10692 5655
rect 10744 5652 10750 5704
rect 12912 5701 12940 5732
rect 13924 5732 14924 5760
rect 12713 5695 12771 5701
rect 12713 5661 12725 5695
rect 12759 5661 12771 5695
rect 12713 5655 12771 5661
rect 12897 5695 12955 5701
rect 12897 5661 12909 5695
rect 12943 5692 12955 5695
rect 12986 5692 12992 5704
rect 12943 5664 12992 5692
rect 12943 5661 12955 5664
rect 12897 5655 12955 5661
rect 10410 5584 10416 5636
rect 10468 5584 10474 5636
rect 10505 5627 10563 5633
rect 10505 5593 10517 5627
rect 10551 5624 10563 5627
rect 11977 5627 12035 5633
rect 11977 5624 11989 5627
rect 10551 5596 11989 5624
rect 10551 5593 10563 5596
rect 10505 5587 10563 5593
rect 11977 5593 11989 5596
rect 12023 5593 12035 5627
rect 11977 5587 12035 5593
rect 12434 5584 12440 5636
rect 12492 5624 12498 5636
rect 12728 5624 12756 5655
rect 12986 5652 12992 5664
rect 13044 5652 13050 5704
rect 13924 5701 13952 5732
rect 14918 5720 14924 5732
rect 14976 5760 14982 5772
rect 14976 5732 15424 5760
rect 14976 5720 14982 5732
rect 13633 5695 13691 5701
rect 13633 5661 13645 5695
rect 13679 5661 13691 5695
rect 13633 5655 13691 5661
rect 13909 5695 13967 5701
rect 13909 5661 13921 5695
rect 13955 5661 13967 5695
rect 13909 5655 13967 5661
rect 12492 5596 12756 5624
rect 13648 5624 13676 5655
rect 14550 5652 14556 5704
rect 14608 5652 14614 5704
rect 14737 5695 14795 5701
rect 14737 5661 14749 5695
rect 14783 5692 14795 5695
rect 15194 5692 15200 5704
rect 14783 5664 15200 5692
rect 14783 5661 14795 5664
rect 14737 5655 14795 5661
rect 15194 5652 15200 5664
rect 15252 5652 15258 5704
rect 15396 5701 15424 5732
rect 15746 5720 15752 5772
rect 15804 5760 15810 5772
rect 17497 5763 17555 5769
rect 17497 5760 17509 5763
rect 15804 5732 17509 5760
rect 15804 5720 15810 5732
rect 17497 5729 17509 5732
rect 17543 5729 17555 5763
rect 17497 5723 17555 5729
rect 15381 5695 15439 5701
rect 15381 5661 15393 5695
rect 15427 5661 15439 5695
rect 15381 5655 15439 5661
rect 17126 5652 17132 5704
rect 17184 5652 17190 5704
rect 18156 5692 18184 5856
rect 22189 5831 22247 5837
rect 19260 5800 19840 5828
rect 19260 5769 19288 5800
rect 19812 5772 19840 5800
rect 22189 5797 22201 5831
rect 22235 5828 22247 5831
rect 23198 5828 23204 5840
rect 22235 5800 23204 5828
rect 22235 5797 22247 5800
rect 22189 5791 22247 5797
rect 23198 5788 23204 5800
rect 23256 5828 23262 5840
rect 27522 5828 27528 5840
rect 23256 5800 27528 5828
rect 23256 5788 23262 5800
rect 27522 5788 27528 5800
rect 27580 5788 27586 5840
rect 29362 5788 29368 5840
rect 29420 5828 29426 5840
rect 29825 5831 29883 5837
rect 29825 5828 29837 5831
rect 29420 5800 29837 5828
rect 29420 5788 29426 5800
rect 29825 5797 29837 5800
rect 29871 5797 29883 5831
rect 29825 5791 29883 5797
rect 19245 5763 19303 5769
rect 19245 5729 19257 5763
rect 19291 5729 19303 5763
rect 19245 5723 19303 5729
rect 19334 5720 19340 5772
rect 19392 5720 19398 5772
rect 19518 5720 19524 5772
rect 19576 5760 19582 5772
rect 19705 5763 19763 5769
rect 19705 5760 19717 5763
rect 19576 5732 19717 5760
rect 19576 5720 19582 5732
rect 19705 5729 19717 5732
rect 19751 5729 19763 5763
rect 19705 5723 19763 5729
rect 19794 5720 19800 5772
rect 19852 5720 19858 5772
rect 22204 5732 22692 5760
rect 19352 5692 19380 5720
rect 19613 5695 19671 5701
rect 19613 5692 19625 5695
rect 18156 5664 19625 5692
rect 19613 5661 19625 5664
rect 19659 5661 19671 5695
rect 19613 5655 19671 5661
rect 20070 5652 20076 5704
rect 20128 5652 20134 5704
rect 20438 5652 20444 5704
rect 20496 5652 20502 5704
rect 20530 5652 20536 5704
rect 20588 5692 20594 5704
rect 22204 5701 22232 5732
rect 22664 5704 22692 5732
rect 24210 5720 24216 5772
rect 24268 5760 24274 5772
rect 24268 5732 25084 5760
rect 24268 5720 24274 5732
rect 20625 5695 20683 5701
rect 20625 5692 20637 5695
rect 20588 5664 20637 5692
rect 20588 5652 20594 5664
rect 20625 5661 20637 5664
rect 20671 5661 20683 5695
rect 20625 5655 20683 5661
rect 22189 5695 22247 5701
rect 22189 5661 22201 5695
rect 22235 5661 22247 5695
rect 22189 5655 22247 5661
rect 22373 5695 22431 5701
rect 22373 5661 22385 5695
rect 22419 5661 22431 5695
rect 22373 5655 22431 5661
rect 14182 5624 14188 5636
rect 13648 5596 14188 5624
rect 12492 5584 12498 5596
rect 14182 5584 14188 5596
rect 14240 5584 14246 5636
rect 14568 5624 14596 5652
rect 14292 5596 14596 5624
rect 15473 5627 15531 5633
rect 10686 5556 10692 5568
rect 10300 5528 10692 5556
rect 10686 5516 10692 5528
rect 10744 5516 10750 5568
rect 10781 5559 10839 5565
rect 10781 5525 10793 5559
rect 10827 5556 10839 5559
rect 11698 5556 11704 5568
rect 10827 5528 11704 5556
rect 10827 5525 10839 5528
rect 10781 5519 10839 5525
rect 11698 5516 11704 5528
rect 11756 5516 11762 5568
rect 13449 5559 13507 5565
rect 13449 5525 13461 5559
rect 13495 5556 13507 5559
rect 13630 5556 13636 5568
rect 13495 5528 13636 5556
rect 13495 5525 13507 5528
rect 13449 5519 13507 5525
rect 13630 5516 13636 5528
rect 13688 5516 13694 5568
rect 13817 5559 13875 5565
rect 13817 5525 13829 5559
rect 13863 5556 13875 5559
rect 14292 5556 14320 5596
rect 15473 5593 15485 5627
rect 15519 5624 15531 5627
rect 15930 5624 15936 5636
rect 15519 5596 15936 5624
rect 15519 5593 15531 5596
rect 15473 5587 15531 5593
rect 15930 5584 15936 5596
rect 15988 5584 15994 5636
rect 16114 5584 16120 5636
rect 16172 5584 16178 5636
rect 19337 5627 19395 5633
rect 19337 5593 19349 5627
rect 19383 5593 19395 5627
rect 22388 5624 22416 5655
rect 22646 5652 22652 5704
rect 22704 5652 22710 5704
rect 22922 5652 22928 5704
rect 22980 5652 22986 5704
rect 23106 5652 23112 5704
rect 23164 5652 23170 5704
rect 23290 5652 23296 5704
rect 23348 5652 23354 5704
rect 23566 5652 23572 5704
rect 23624 5652 23630 5704
rect 23658 5652 23664 5704
rect 23716 5652 23722 5704
rect 24581 5695 24639 5701
rect 24581 5661 24593 5695
rect 24627 5692 24639 5695
rect 24762 5692 24768 5704
rect 24627 5664 24768 5692
rect 24627 5661 24639 5664
rect 24581 5655 24639 5661
rect 24762 5652 24768 5664
rect 24820 5652 24826 5704
rect 25056 5701 25084 5732
rect 29178 5720 29184 5772
rect 29236 5760 29242 5772
rect 29549 5763 29607 5769
rect 29549 5760 29561 5763
rect 29236 5732 29561 5760
rect 29236 5720 29242 5732
rect 29549 5729 29561 5732
rect 29595 5729 29607 5763
rect 29549 5723 29607 5729
rect 24857 5695 24915 5701
rect 24857 5661 24869 5695
rect 24903 5661 24915 5695
rect 24857 5655 24915 5661
rect 25041 5695 25099 5701
rect 25041 5661 25053 5695
rect 25087 5692 25099 5695
rect 30006 5692 30012 5704
rect 25087 5664 30012 5692
rect 25087 5661 25099 5664
rect 25041 5655 25099 5661
rect 23124 5624 23152 5652
rect 19337 5587 19395 5593
rect 19904 5596 22324 5624
rect 22388 5596 23152 5624
rect 23308 5624 23336 5652
rect 24872 5624 24900 5655
rect 30006 5652 30012 5664
rect 30064 5652 30070 5704
rect 31754 5652 31760 5704
rect 31812 5652 31818 5704
rect 32122 5652 32128 5704
rect 32180 5652 32186 5704
rect 32309 5695 32367 5701
rect 32309 5661 32321 5695
rect 32355 5661 32367 5695
rect 32309 5655 32367 5661
rect 23308 5596 24900 5624
rect 30101 5627 30159 5633
rect 13863 5528 14320 5556
rect 13863 5525 13875 5528
rect 13817 5519 13875 5525
rect 14366 5516 14372 5568
rect 14424 5516 14430 5568
rect 14829 5559 14887 5565
rect 14829 5525 14841 5559
rect 14875 5556 14887 5559
rect 15378 5556 15384 5568
rect 14875 5528 15384 5556
rect 14875 5525 14887 5528
rect 14829 5519 14887 5525
rect 15378 5516 15384 5528
rect 15436 5516 15442 5568
rect 19352 5556 19380 5587
rect 19610 5556 19616 5568
rect 19352 5528 19616 5556
rect 19610 5516 19616 5528
rect 19668 5516 19674 5568
rect 19904 5565 19932 5596
rect 19889 5559 19947 5565
rect 19889 5525 19901 5559
rect 19935 5525 19947 5559
rect 19889 5519 19947 5525
rect 20441 5559 20499 5565
rect 20441 5525 20453 5559
rect 20487 5556 20499 5559
rect 20990 5556 20996 5568
rect 20487 5528 20996 5556
rect 20487 5525 20499 5528
rect 20441 5519 20499 5525
rect 20990 5516 20996 5528
rect 21048 5516 21054 5568
rect 22296 5556 22324 5596
rect 30101 5593 30113 5627
rect 30147 5624 30159 5627
rect 30190 5624 30196 5636
rect 30147 5596 30196 5624
rect 30147 5593 30159 5596
rect 30101 5587 30159 5593
rect 30190 5584 30196 5596
rect 30248 5584 30254 5636
rect 30282 5584 30288 5636
rect 30340 5584 30346 5636
rect 31665 5627 31723 5633
rect 31665 5593 31677 5627
rect 31711 5593 31723 5627
rect 31772 5624 31800 5652
rect 31849 5627 31907 5633
rect 31849 5624 31861 5627
rect 31772 5596 31861 5624
rect 31665 5587 31723 5593
rect 31849 5593 31861 5596
rect 31895 5593 31907 5627
rect 31849 5587 31907 5593
rect 22922 5556 22928 5568
rect 22296 5528 22928 5556
rect 22922 5516 22928 5528
rect 22980 5556 22986 5568
rect 23750 5556 23756 5568
rect 22980 5528 23756 5556
rect 22980 5516 22986 5528
rect 23750 5516 23756 5528
rect 23808 5516 23814 5568
rect 24394 5516 24400 5568
rect 24452 5516 24458 5568
rect 29454 5516 29460 5568
rect 29512 5556 29518 5568
rect 30009 5559 30067 5565
rect 30009 5556 30021 5559
rect 29512 5528 30021 5556
rect 29512 5516 29518 5528
rect 30009 5525 30021 5528
rect 30055 5556 30067 5559
rect 31680 5556 31708 5587
rect 31938 5584 31944 5636
rect 31996 5624 32002 5636
rect 32324 5624 32352 5655
rect 31996 5596 32352 5624
rect 31996 5584 32002 5596
rect 30055 5528 31708 5556
rect 30055 5525 30067 5528
rect 30009 5519 30067 5525
rect 1104 5466 38272 5488
rect 1104 5414 4874 5466
rect 4926 5414 4938 5466
rect 4990 5414 5002 5466
rect 5054 5414 5066 5466
rect 5118 5414 5130 5466
rect 5182 5414 35594 5466
rect 35646 5414 35658 5466
rect 35710 5414 35722 5466
rect 35774 5414 35786 5466
rect 35838 5414 35850 5466
rect 35902 5414 38272 5466
rect 1104 5392 38272 5414
rect 5626 5312 5632 5364
rect 5684 5352 5690 5364
rect 6457 5355 6515 5361
rect 6457 5352 6469 5355
rect 5684 5324 6469 5352
rect 5684 5312 5690 5324
rect 6457 5321 6469 5324
rect 6503 5321 6515 5355
rect 6457 5315 6515 5321
rect 7374 5312 7380 5364
rect 7432 5312 7438 5364
rect 8846 5312 8852 5364
rect 8904 5312 8910 5364
rect 9858 5352 9864 5364
rect 9324 5324 9864 5352
rect 6641 5219 6699 5225
rect 6641 5185 6653 5219
rect 6687 5216 6699 5219
rect 7392 5216 7420 5312
rect 6687 5188 7420 5216
rect 6687 5185 6699 5188
rect 6641 5179 6699 5185
rect 8202 5176 8208 5228
rect 8260 5176 8266 5228
rect 9030 5176 9036 5228
rect 9088 5216 9094 5228
rect 9324 5225 9352 5324
rect 9858 5312 9864 5324
rect 9916 5312 9922 5364
rect 11882 5352 11888 5364
rect 11532 5324 11888 5352
rect 9493 5287 9551 5293
rect 9493 5253 9505 5287
rect 9539 5284 9551 5287
rect 9677 5287 9735 5293
rect 9677 5284 9689 5287
rect 9539 5256 9689 5284
rect 9539 5253 9551 5256
rect 9493 5247 9551 5253
rect 9677 5253 9689 5256
rect 9723 5253 9735 5287
rect 10410 5284 10416 5296
rect 9677 5247 9735 5253
rect 9968 5256 10416 5284
rect 9309 5219 9367 5225
rect 9309 5216 9321 5219
rect 9088 5188 9321 5216
rect 9088 5176 9094 5188
rect 9309 5185 9321 5188
rect 9355 5185 9367 5219
rect 9309 5179 9367 5185
rect 9585 5219 9643 5225
rect 9585 5185 9597 5219
rect 9631 5216 9643 5219
rect 9858 5216 9864 5228
rect 9631 5188 9864 5216
rect 9631 5185 9643 5188
rect 9585 5179 9643 5185
rect 9858 5176 9864 5188
rect 9916 5216 9922 5228
rect 9968 5216 9996 5256
rect 10410 5244 10416 5256
rect 10468 5244 10474 5296
rect 9916 5188 9996 5216
rect 9916 5176 9922 5188
rect 10042 5176 10048 5228
rect 10100 5216 10106 5228
rect 11532 5225 11560 5324
rect 11882 5312 11888 5324
rect 11940 5352 11946 5364
rect 12158 5352 12164 5364
rect 11940 5324 12164 5352
rect 11940 5312 11946 5324
rect 12158 5312 12164 5324
rect 12216 5352 12222 5364
rect 12216 5324 13492 5352
rect 12216 5312 12222 5324
rect 11698 5244 11704 5296
rect 11756 5284 11762 5296
rect 11793 5287 11851 5293
rect 11793 5284 11805 5287
rect 11756 5256 11805 5284
rect 11756 5244 11762 5256
rect 11793 5253 11805 5256
rect 11839 5253 11851 5287
rect 11793 5247 11851 5253
rect 10505 5219 10563 5225
rect 10505 5216 10517 5219
rect 10100 5188 10517 5216
rect 10100 5176 10106 5188
rect 10505 5185 10517 5188
rect 10551 5185 10563 5219
rect 10505 5179 10563 5185
rect 11517 5219 11575 5225
rect 11517 5185 11529 5219
rect 11563 5185 11575 5219
rect 11517 5179 11575 5185
rect 12894 5176 12900 5228
rect 12952 5216 12958 5228
rect 13464 5225 13492 5324
rect 15194 5312 15200 5364
rect 15252 5312 15258 5364
rect 17126 5312 17132 5364
rect 17184 5352 17190 5364
rect 17313 5355 17371 5361
rect 17313 5352 17325 5355
rect 17184 5324 17325 5352
rect 17184 5312 17190 5324
rect 17313 5321 17325 5324
rect 17359 5321 17371 5355
rect 17313 5315 17371 5321
rect 19705 5355 19763 5361
rect 19705 5321 19717 5355
rect 19751 5352 19763 5355
rect 20162 5352 20168 5364
rect 19751 5324 20168 5352
rect 19751 5321 19763 5324
rect 19705 5315 19763 5321
rect 20162 5312 20168 5324
rect 20220 5352 20226 5364
rect 20438 5352 20444 5364
rect 20220 5324 20444 5352
rect 20220 5312 20226 5324
rect 20438 5312 20444 5324
rect 20496 5312 20502 5364
rect 23109 5355 23167 5361
rect 23109 5321 23121 5355
rect 23155 5352 23167 5355
rect 23566 5352 23572 5364
rect 23155 5324 23572 5352
rect 23155 5321 23167 5324
rect 23109 5315 23167 5321
rect 23566 5312 23572 5324
rect 23624 5312 23630 5364
rect 23658 5312 23664 5364
rect 23716 5312 23722 5364
rect 27525 5355 27583 5361
rect 27525 5321 27537 5355
rect 27571 5352 27583 5355
rect 27614 5352 27620 5364
rect 27571 5324 27620 5352
rect 27571 5321 27583 5324
rect 27525 5315 27583 5321
rect 27614 5312 27620 5324
rect 27672 5312 27678 5364
rect 29457 5355 29515 5361
rect 29457 5352 29469 5355
rect 28736 5324 29469 5352
rect 13630 5244 13636 5296
rect 13688 5284 13694 5296
rect 13725 5287 13783 5293
rect 13725 5284 13737 5287
rect 13688 5256 13737 5284
rect 13688 5244 13694 5256
rect 13725 5253 13737 5256
rect 13771 5253 13783 5287
rect 16114 5284 16120 5296
rect 14950 5270 16120 5284
rect 13725 5247 13783 5253
rect 14936 5256 16120 5270
rect 13449 5219 13507 5225
rect 12952 5188 13400 5216
rect 12952 5176 12958 5188
rect 9674 5108 9680 5160
rect 9732 5148 9738 5160
rect 10229 5151 10287 5157
rect 10229 5148 10241 5151
rect 9732 5120 10241 5148
rect 9732 5108 9738 5120
rect 10229 5117 10241 5120
rect 10275 5117 10287 5151
rect 10229 5111 10287 5117
rect 12986 5108 12992 5160
rect 13044 5108 13050 5160
rect 13372 5148 13400 5188
rect 13449 5185 13461 5219
rect 13495 5185 13507 5219
rect 13449 5179 13507 5185
rect 14936 5148 14964 5256
rect 16114 5244 16120 5256
rect 16172 5244 16178 5296
rect 19334 5244 19340 5296
rect 19392 5244 19398 5296
rect 19518 5244 19524 5296
rect 19576 5284 19582 5296
rect 19576 5256 20024 5284
rect 19576 5244 19582 5256
rect 19352 5216 19380 5244
rect 19996 5225 20024 5256
rect 20990 5244 20996 5296
rect 21048 5284 21054 5296
rect 21085 5287 21143 5293
rect 21085 5284 21097 5287
rect 21048 5256 21097 5284
rect 21048 5244 21054 5256
rect 21085 5253 21097 5256
rect 21131 5253 21143 5287
rect 21085 5247 21143 5253
rect 22925 5287 22983 5293
rect 22925 5253 22937 5287
rect 22971 5284 22983 5287
rect 25869 5287 25927 5293
rect 22971 5256 23152 5284
rect 22971 5253 22983 5256
rect 22925 5247 22983 5253
rect 23124 5228 23152 5256
rect 23308 5256 25728 5284
rect 19797 5219 19855 5225
rect 19797 5216 19809 5219
rect 19352 5188 19809 5216
rect 19797 5185 19809 5188
rect 19843 5185 19855 5219
rect 19797 5179 19855 5185
rect 19981 5219 20039 5225
rect 19981 5185 19993 5219
rect 20027 5185 20039 5219
rect 19981 5179 20039 5185
rect 20898 5176 20904 5228
rect 20956 5176 20962 5228
rect 22281 5219 22339 5225
rect 22281 5185 22293 5219
rect 22327 5216 22339 5219
rect 22646 5216 22652 5228
rect 22327 5188 22652 5216
rect 22327 5185 22339 5188
rect 22281 5179 22339 5185
rect 22646 5176 22652 5188
rect 22704 5176 22710 5228
rect 23014 5176 23020 5228
rect 23072 5176 23078 5228
rect 23106 5176 23112 5228
rect 23164 5176 23170 5228
rect 23198 5176 23204 5228
rect 23256 5176 23262 5228
rect 13372 5120 14964 5148
rect 15378 5108 15384 5160
rect 15436 5148 15442 5160
rect 15838 5148 15844 5160
rect 15436 5120 15844 5148
rect 15436 5108 15442 5120
rect 15838 5108 15844 5120
rect 15896 5108 15902 5160
rect 16666 5108 16672 5160
rect 16724 5108 16730 5160
rect 22370 5108 22376 5160
rect 22428 5148 22434 5160
rect 23308 5148 23336 5256
rect 23385 5219 23443 5225
rect 23385 5185 23397 5219
rect 23431 5185 23443 5219
rect 23385 5179 23443 5185
rect 22428 5120 23336 5148
rect 22428 5108 22434 5120
rect 13004 5080 13032 5108
rect 13265 5083 13323 5089
rect 13265 5080 13277 5083
rect 13004 5052 13277 5080
rect 13265 5049 13277 5052
rect 13311 5049 13323 5083
rect 13265 5043 13323 5049
rect 21269 5083 21327 5089
rect 21269 5049 21281 5083
rect 21315 5080 21327 5083
rect 23290 5080 23296 5092
rect 21315 5052 23296 5080
rect 21315 5049 21327 5052
rect 21269 5043 21327 5049
rect 23290 5040 23296 5052
rect 23348 5040 23354 5092
rect 23400 5024 23428 5179
rect 24854 5176 24860 5228
rect 24912 5216 24918 5228
rect 25498 5216 25504 5228
rect 24912 5188 25504 5216
rect 24912 5176 24918 5188
rect 25498 5176 25504 5188
rect 25556 5216 25562 5228
rect 25700 5225 25728 5256
rect 25869 5253 25881 5287
rect 25915 5284 25927 5287
rect 28442 5284 28448 5296
rect 25915 5256 27200 5284
rect 25915 5253 25927 5256
rect 25869 5247 25927 5253
rect 25593 5219 25651 5225
rect 25593 5216 25605 5219
rect 25556 5188 25605 5216
rect 25556 5176 25562 5188
rect 25593 5185 25605 5188
rect 25639 5185 25651 5219
rect 25593 5179 25651 5185
rect 25685 5219 25743 5225
rect 25685 5185 25697 5219
rect 25731 5216 25743 5219
rect 26234 5216 26240 5228
rect 25731 5188 26240 5216
rect 25731 5185 25743 5188
rect 25685 5179 25743 5185
rect 26234 5176 26240 5188
rect 26292 5176 26298 5228
rect 27172 5225 27200 5256
rect 27908 5256 28448 5284
rect 27157 5219 27215 5225
rect 27157 5185 27169 5219
rect 27203 5185 27215 5219
rect 27157 5179 27215 5185
rect 27614 5176 27620 5228
rect 27672 5176 27678 5228
rect 27706 5176 27712 5228
rect 27764 5176 27770 5228
rect 27798 5176 27804 5228
rect 27856 5216 27862 5228
rect 27908 5225 27936 5256
rect 28442 5244 28448 5256
rect 28500 5244 28506 5296
rect 28736 5225 28764 5324
rect 29457 5321 29469 5324
rect 29503 5352 29515 5355
rect 29730 5352 29736 5364
rect 29503 5324 29736 5352
rect 29503 5321 29515 5324
rect 29457 5315 29515 5321
rect 29730 5312 29736 5324
rect 29788 5312 29794 5364
rect 30193 5355 30251 5361
rect 30193 5321 30205 5355
rect 30239 5352 30251 5355
rect 30282 5352 30288 5364
rect 30239 5324 30288 5352
rect 30239 5321 30251 5324
rect 30193 5315 30251 5321
rect 30282 5312 30288 5324
rect 30340 5312 30346 5364
rect 31481 5355 31539 5361
rect 31481 5321 31493 5355
rect 31527 5352 31539 5355
rect 32122 5352 32128 5364
rect 31527 5324 32128 5352
rect 31527 5321 31539 5324
rect 31481 5315 31539 5321
rect 32122 5312 32128 5324
rect 32180 5312 32186 5364
rect 29362 5244 29368 5296
rect 29420 5244 29426 5296
rect 30374 5284 30380 5296
rect 29564 5256 30380 5284
rect 27893 5219 27951 5225
rect 27893 5216 27905 5219
rect 27856 5188 27905 5216
rect 27856 5176 27862 5188
rect 27893 5185 27905 5188
rect 27939 5185 27951 5219
rect 28537 5219 28595 5225
rect 28537 5216 28549 5219
rect 27893 5179 27951 5185
rect 28000 5188 28549 5216
rect 23661 5151 23719 5157
rect 23661 5117 23673 5151
rect 23707 5148 23719 5151
rect 24394 5148 24400 5160
rect 23707 5120 24400 5148
rect 23707 5117 23719 5120
rect 23661 5111 23719 5117
rect 24394 5108 24400 5120
rect 24452 5108 24458 5160
rect 25869 5151 25927 5157
rect 25869 5117 25881 5151
rect 25915 5148 25927 5151
rect 25915 5120 26096 5148
rect 25915 5117 25927 5120
rect 25869 5111 25927 5117
rect 26068 5092 26096 5120
rect 26970 5108 26976 5160
rect 27028 5148 27034 5160
rect 27065 5151 27123 5157
rect 27065 5148 27077 5151
rect 27028 5120 27077 5148
rect 27028 5108 27034 5120
rect 27065 5117 27077 5120
rect 27111 5148 27123 5151
rect 28000 5148 28028 5188
rect 28537 5185 28549 5188
rect 28583 5185 28595 5219
rect 28537 5179 28595 5185
rect 28721 5219 28779 5225
rect 28721 5185 28733 5219
rect 28767 5185 28779 5219
rect 28721 5179 28779 5185
rect 28905 5219 28963 5225
rect 28905 5185 28917 5219
rect 28951 5185 28963 5219
rect 28905 5179 28963 5185
rect 28997 5219 29055 5225
rect 28997 5185 29009 5219
rect 29043 5216 29055 5219
rect 29380 5216 29408 5244
rect 29043 5188 29408 5216
rect 29043 5185 29055 5188
rect 28997 5179 29055 5185
rect 27111 5120 28028 5148
rect 27111 5117 27123 5120
rect 27065 5111 27123 5117
rect 28258 5108 28264 5160
rect 28316 5108 28322 5160
rect 28920 5148 28948 5179
rect 29454 5176 29460 5228
rect 29512 5176 29518 5228
rect 29564 5225 29592 5256
rect 30374 5244 30380 5256
rect 30432 5284 30438 5296
rect 30432 5256 31156 5284
rect 30432 5244 30438 5256
rect 29549 5219 29607 5225
rect 29549 5185 29561 5219
rect 29595 5185 29607 5219
rect 29549 5179 29607 5185
rect 29733 5219 29791 5225
rect 29733 5185 29745 5219
rect 29779 5185 29791 5219
rect 29733 5179 29791 5185
rect 29472 5148 29500 5176
rect 28920 5120 29500 5148
rect 26050 5040 26056 5092
rect 26108 5040 26114 5092
rect 27893 5083 27951 5089
rect 27893 5049 27905 5083
rect 27939 5080 27951 5083
rect 28276 5080 28304 5108
rect 27939 5052 28304 5080
rect 27939 5049 27951 5052
rect 27893 5043 27951 5049
rect 29178 5040 29184 5092
rect 29236 5080 29242 5092
rect 29273 5083 29331 5089
rect 29273 5080 29285 5083
rect 29236 5052 29285 5080
rect 29236 5040 29242 5052
rect 29273 5049 29285 5052
rect 29319 5049 29331 5083
rect 29273 5043 29331 5049
rect 9122 4972 9128 5024
rect 9180 4972 9186 5024
rect 11146 4972 11152 5024
rect 11204 4972 11210 5024
rect 16390 4972 16396 5024
rect 16448 4972 16454 5024
rect 19886 4972 19892 5024
rect 19944 4972 19950 5024
rect 23382 4972 23388 5024
rect 23440 4972 23446 5024
rect 23477 5015 23535 5021
rect 23477 4981 23489 5015
rect 23523 5012 23535 5015
rect 24394 5012 24400 5024
rect 23523 4984 24400 5012
rect 23523 4981 23535 4984
rect 23477 4975 23535 4981
rect 24394 4972 24400 4984
rect 24452 4972 24458 5024
rect 29748 5012 29776 5179
rect 29822 5176 29828 5228
rect 29880 5216 29886 5228
rect 29917 5219 29975 5225
rect 29917 5216 29929 5219
rect 29880 5188 29929 5216
rect 29880 5176 29886 5188
rect 29917 5185 29929 5188
rect 29963 5185 29975 5219
rect 29917 5179 29975 5185
rect 30009 5219 30067 5225
rect 30009 5185 30021 5219
rect 30055 5216 30067 5219
rect 30098 5216 30104 5228
rect 30055 5188 30104 5216
rect 30055 5185 30067 5188
rect 30009 5179 30067 5185
rect 29932 5148 29960 5179
rect 30098 5176 30104 5188
rect 30156 5216 30162 5228
rect 31128 5225 31156 5256
rect 30469 5219 30527 5225
rect 30469 5216 30481 5219
rect 30156 5188 30481 5216
rect 30156 5176 30162 5188
rect 30469 5185 30481 5188
rect 30515 5185 30527 5219
rect 30469 5179 30527 5185
rect 30745 5219 30803 5225
rect 30745 5185 30757 5219
rect 30791 5216 30803 5219
rect 31113 5219 31171 5225
rect 30791 5188 31064 5216
rect 30791 5185 30803 5188
rect 30745 5179 30803 5185
rect 30561 5151 30619 5157
rect 30561 5148 30573 5151
rect 29932 5120 30573 5148
rect 30561 5117 30573 5120
rect 30607 5117 30619 5151
rect 30561 5111 30619 5117
rect 29822 5040 29828 5092
rect 29880 5040 29886 5092
rect 29932 5052 30420 5080
rect 29932 5012 29960 5052
rect 30006 5012 30012 5024
rect 29748 4984 30012 5012
rect 30006 4972 30012 4984
rect 30064 4972 30070 5024
rect 30282 4972 30288 5024
rect 30340 4972 30346 5024
rect 30392 5012 30420 5052
rect 30650 5040 30656 5092
rect 30708 5040 30714 5092
rect 30760 5012 30788 5179
rect 31036 5157 31064 5188
rect 31113 5185 31125 5219
rect 31159 5216 31171 5219
rect 31754 5216 31760 5228
rect 31159 5188 31760 5216
rect 31159 5185 31171 5188
rect 31113 5179 31171 5185
rect 31754 5176 31760 5188
rect 31812 5176 31818 5228
rect 31021 5151 31079 5157
rect 31021 5117 31033 5151
rect 31067 5117 31079 5151
rect 31021 5111 31079 5117
rect 30392 4984 30788 5012
rect 1104 4922 38272 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 38272 4922
rect 1104 4848 38272 4870
rect 9858 4768 9864 4820
rect 9916 4768 9922 4820
rect 10952 4811 11010 4817
rect 10952 4777 10964 4811
rect 10998 4808 11010 4811
rect 11146 4808 11152 4820
rect 10998 4780 11152 4808
rect 10998 4777 11010 4780
rect 10952 4771 11010 4777
rect 11146 4768 11152 4780
rect 11204 4768 11210 4820
rect 12434 4768 12440 4820
rect 12492 4768 12498 4820
rect 15838 4768 15844 4820
rect 15896 4808 15902 4820
rect 15933 4811 15991 4817
rect 15933 4808 15945 4811
rect 15896 4780 15945 4808
rect 15896 4768 15902 4780
rect 15933 4777 15945 4780
rect 15979 4777 15991 4811
rect 15933 4771 15991 4777
rect 16390 4768 16396 4820
rect 16448 4768 16454 4820
rect 16577 4811 16635 4817
rect 16577 4777 16589 4811
rect 16623 4808 16635 4811
rect 16666 4808 16672 4820
rect 16623 4780 16672 4808
rect 16623 4777 16635 4780
rect 16577 4771 16635 4777
rect 16666 4768 16672 4780
rect 16724 4768 16730 4820
rect 19426 4768 19432 4820
rect 19484 4768 19490 4820
rect 20162 4768 20168 4820
rect 20220 4768 20226 4820
rect 20349 4811 20407 4817
rect 20349 4777 20361 4811
rect 20395 4808 20407 4811
rect 20898 4808 20904 4820
rect 20395 4780 20904 4808
rect 20395 4777 20407 4780
rect 20349 4771 20407 4777
rect 20898 4768 20904 4780
rect 20956 4768 20962 4820
rect 23382 4768 23388 4820
rect 23440 4808 23446 4820
rect 23477 4811 23535 4817
rect 23477 4808 23489 4811
rect 23440 4780 23489 4808
rect 23440 4768 23446 4780
rect 23477 4777 23489 4780
rect 23523 4777 23535 4811
rect 23477 4771 23535 4777
rect 23566 4768 23572 4820
rect 23624 4768 23630 4820
rect 24394 4768 24400 4820
rect 24452 4768 24458 4820
rect 25498 4808 25504 4820
rect 24504 4780 25504 4808
rect 10689 4675 10747 4681
rect 10689 4641 10701 4675
rect 10735 4672 10747 4675
rect 12158 4672 12164 4684
rect 10735 4644 12164 4672
rect 10735 4641 10747 4644
rect 10689 4635 10747 4641
rect 12158 4632 12164 4644
rect 12216 4672 12222 4684
rect 14185 4675 14243 4681
rect 14185 4672 14197 4675
rect 12216 4644 14197 4672
rect 12216 4632 12222 4644
rect 14185 4641 14197 4644
rect 14231 4641 14243 4675
rect 16408 4672 16436 4768
rect 14185 4635 14243 4641
rect 16040 4644 16436 4672
rect 19444 4672 19472 4768
rect 19886 4700 19892 4752
rect 19944 4740 19950 4752
rect 23584 4740 23612 4768
rect 24504 4740 24532 4780
rect 25498 4768 25504 4780
rect 25556 4808 25562 4820
rect 25685 4811 25743 4817
rect 25685 4808 25697 4811
rect 25556 4780 25697 4808
rect 25556 4768 25562 4780
rect 25685 4777 25697 4780
rect 25731 4777 25743 4811
rect 25685 4771 25743 4777
rect 26050 4768 26056 4820
rect 26108 4768 26114 4820
rect 27525 4811 27583 4817
rect 27525 4777 27537 4811
rect 27571 4808 27583 4811
rect 27614 4808 27620 4820
rect 27571 4780 27620 4808
rect 27571 4777 27583 4780
rect 27525 4771 27583 4777
rect 27614 4768 27620 4780
rect 27672 4768 27678 4820
rect 29178 4768 29184 4820
rect 29236 4808 29242 4820
rect 29641 4811 29699 4817
rect 29641 4808 29653 4811
rect 29236 4780 29653 4808
rect 29236 4768 29242 4780
rect 29641 4777 29653 4780
rect 29687 4777 29699 4811
rect 29641 4771 29699 4777
rect 30006 4768 30012 4820
rect 30064 4768 30070 4820
rect 30282 4768 30288 4820
rect 30340 4768 30346 4820
rect 19944 4712 23428 4740
rect 23584 4712 24532 4740
rect 19944 4700 19950 4712
rect 19521 4675 19579 4681
rect 19521 4672 19533 4675
rect 19444 4644 19533 4672
rect 1765 4607 1823 4613
rect 1765 4573 1777 4607
rect 1811 4604 1823 4607
rect 3878 4604 3884 4616
rect 1811 4576 3884 4604
rect 1811 4573 1823 4576
rect 1765 4567 1823 4573
rect 3878 4564 3884 4576
rect 3936 4564 3942 4616
rect 9766 4564 9772 4616
rect 9824 4604 9830 4616
rect 10045 4607 10103 4613
rect 10045 4604 10057 4607
rect 9824 4576 10057 4604
rect 9824 4564 9830 4576
rect 10045 4573 10057 4576
rect 10091 4573 10103 4607
rect 10045 4567 10103 4573
rect 10226 4564 10232 4616
rect 10284 4564 10290 4616
rect 15930 4564 15936 4616
rect 15988 4564 15994 4616
rect 16040 4613 16068 4644
rect 19521 4641 19533 4644
rect 19567 4672 19579 4675
rect 19567 4644 21496 4672
rect 19567 4641 19579 4644
rect 19521 4635 19579 4641
rect 16025 4607 16083 4613
rect 16025 4573 16037 4607
rect 16071 4573 16083 4607
rect 16025 4567 16083 4573
rect 16298 4564 16304 4616
rect 16356 4564 16362 4616
rect 16393 4607 16451 4613
rect 16393 4573 16405 4607
rect 16439 4604 16451 4607
rect 16482 4604 16488 4616
rect 16439 4576 16488 4604
rect 16439 4573 16451 4576
rect 16393 4567 16451 4573
rect 16482 4564 16488 4576
rect 16540 4564 16546 4616
rect 19429 4607 19487 4613
rect 19429 4573 19441 4607
rect 19475 4604 19487 4607
rect 20806 4604 20812 4616
rect 19475 4576 20812 4604
rect 19475 4573 19487 4576
rect 19429 4567 19487 4573
rect 20806 4564 20812 4576
rect 20864 4604 20870 4616
rect 21269 4607 21327 4613
rect 21269 4604 21281 4607
rect 20864 4576 21281 4604
rect 20864 4564 20870 4576
rect 21269 4573 21281 4576
rect 21315 4573 21327 4607
rect 21468 4604 21496 4644
rect 22922 4632 22928 4684
rect 22980 4632 22986 4684
rect 21821 4607 21879 4613
rect 21821 4604 21833 4607
rect 21468 4576 21833 4604
rect 21269 4567 21327 4573
rect 21821 4573 21833 4576
rect 21867 4573 21879 4607
rect 22940 4604 22968 4632
rect 23192 4607 23250 4613
rect 23192 4604 23204 4607
rect 22940 4576 23204 4604
rect 21821 4567 21879 4573
rect 23192 4573 23204 4576
rect 23238 4573 23250 4607
rect 23400 4604 23428 4712
rect 24670 4700 24676 4752
rect 24728 4740 24734 4752
rect 24854 4740 24860 4752
rect 24728 4712 24860 4740
rect 24728 4700 24734 4712
rect 23750 4632 23756 4684
rect 23808 4672 23814 4684
rect 24578 4672 24584 4684
rect 23808 4644 24584 4672
rect 23808 4632 23814 4644
rect 24578 4632 24584 4644
rect 24636 4632 24642 4684
rect 24780 4613 24808 4712
rect 24854 4700 24860 4712
rect 24912 4700 24918 4752
rect 27798 4740 27804 4752
rect 25240 4712 27804 4740
rect 25240 4672 25268 4712
rect 27798 4700 27804 4712
rect 27856 4700 27862 4752
rect 29362 4700 29368 4752
rect 29420 4700 29426 4752
rect 25406 4672 25412 4684
rect 24872 4644 25268 4672
rect 25332 4644 25412 4672
rect 24872 4613 24900 4644
rect 24673 4607 24731 4613
rect 24673 4604 24685 4607
rect 23400 4582 24685 4604
rect 23192 4567 23250 4573
rect 23308 4576 24685 4582
rect 934 4496 940 4548
rect 992 4536 998 4548
rect 1397 4539 1455 4545
rect 1397 4536 1409 4539
rect 992 4508 1409 4536
rect 992 4496 998 4508
rect 1397 4505 1409 4508
rect 1443 4505 1455 4539
rect 12894 4536 12900 4548
rect 12190 4508 12900 4536
rect 1397 4499 1455 4505
rect 12894 4496 12900 4508
rect 12952 4496 12958 4548
rect 14458 4496 14464 4548
rect 14516 4496 14522 4548
rect 15948 4536 15976 4564
rect 16209 4539 16267 4545
rect 16209 4536 16221 4539
rect 15686 4508 15884 4536
rect 15948 4508 16221 4536
rect 15856 4468 15884 4508
rect 16209 4505 16221 4508
rect 16255 4505 16267 4539
rect 19981 4539 20039 4545
rect 19981 4536 19993 4539
rect 16209 4499 16267 4505
rect 19812 4508 19993 4536
rect 16758 4468 16764 4480
rect 15856 4440 16764 4468
rect 16758 4428 16764 4440
rect 16816 4428 16822 4480
rect 19812 4477 19840 4508
rect 19981 4505 19993 4508
rect 20027 4536 20039 4539
rect 20070 4536 20076 4548
rect 20027 4508 20076 4536
rect 20027 4505 20039 4508
rect 19981 4499 20039 4505
rect 20070 4496 20076 4508
rect 20128 4496 20134 4548
rect 20197 4539 20255 4545
rect 20197 4505 20209 4539
rect 20243 4536 20255 4539
rect 20530 4536 20536 4548
rect 20243 4508 20536 4536
rect 20243 4505 20255 4508
rect 20197 4499 20255 4505
rect 20530 4496 20536 4508
rect 20588 4496 20594 4548
rect 19797 4471 19855 4477
rect 19797 4437 19809 4471
rect 19843 4437 19855 4471
rect 21836 4468 21864 4567
rect 23308 4554 23428 4576
rect 24673 4573 24685 4576
rect 24719 4573 24731 4607
rect 24673 4567 24731 4573
rect 24765 4607 24823 4613
rect 24765 4573 24777 4607
rect 24811 4573 24823 4607
rect 24765 4567 24823 4573
rect 24857 4607 24915 4613
rect 24857 4573 24869 4607
rect 24903 4573 24915 4607
rect 24857 4567 24915 4573
rect 22646 4496 22652 4548
rect 22704 4496 22710 4548
rect 23198 4468 23204 4480
rect 21836 4440 23204 4468
rect 19797 4431 19855 4437
rect 23198 4428 23204 4440
rect 23256 4428 23262 4480
rect 23308 4477 23336 4554
rect 23474 4496 23480 4548
rect 23532 4536 23538 4548
rect 24578 4536 24584 4548
rect 23532 4508 24584 4536
rect 23532 4496 23538 4508
rect 24578 4496 24584 4508
rect 24636 4496 24642 4548
rect 24688 4536 24716 4567
rect 24946 4564 24952 4616
rect 25004 4604 25010 4616
rect 25332 4613 25360 4644
rect 25406 4632 25412 4644
rect 25464 4632 25470 4684
rect 26605 4675 26663 4681
rect 26605 4672 26617 4675
rect 26160 4644 26617 4672
rect 26160 4613 26188 4644
rect 26605 4641 26617 4644
rect 26651 4641 26663 4675
rect 26605 4635 26663 4641
rect 26970 4632 26976 4684
rect 27028 4672 27034 4684
rect 27065 4675 27123 4681
rect 27065 4672 27077 4675
rect 27028 4644 27077 4672
rect 27028 4632 27034 4644
rect 27065 4641 27077 4644
rect 27111 4672 27123 4675
rect 27111 4644 27384 4672
rect 27111 4641 27123 4644
rect 27065 4635 27123 4641
rect 25041 4607 25099 4613
rect 25041 4604 25053 4607
rect 25004 4576 25053 4604
rect 25004 4564 25010 4576
rect 25041 4573 25053 4576
rect 25087 4573 25099 4607
rect 25041 4567 25099 4573
rect 25317 4607 25375 4613
rect 25317 4573 25329 4607
rect 25363 4573 25375 4607
rect 25593 4607 25651 4613
rect 25593 4604 25605 4607
rect 25317 4567 25375 4573
rect 25424 4576 25605 4604
rect 25133 4539 25191 4545
rect 25133 4536 25145 4539
rect 24688 4508 25145 4536
rect 25133 4505 25145 4508
rect 25179 4505 25191 4539
rect 25133 4499 25191 4505
rect 23293 4471 23351 4477
rect 23293 4437 23305 4471
rect 23339 4437 23351 4471
rect 23293 4431 23351 4437
rect 23382 4428 23388 4480
rect 23440 4468 23446 4480
rect 25038 4468 25044 4480
rect 23440 4440 25044 4468
rect 23440 4428 23446 4440
rect 25038 4428 25044 4440
rect 25096 4468 25102 4480
rect 25424 4468 25452 4576
rect 25593 4573 25605 4576
rect 25639 4573 25651 4607
rect 25593 4567 25651 4573
rect 26145 4607 26203 4613
rect 26145 4573 26157 4607
rect 26191 4573 26203 4607
rect 26145 4567 26203 4573
rect 25501 4539 25559 4545
rect 25501 4505 25513 4539
rect 25547 4536 25559 4539
rect 26160 4536 26188 4567
rect 26326 4564 26332 4616
rect 26384 4604 26390 4616
rect 27356 4613 27384 4644
rect 27982 4632 27988 4684
rect 28040 4632 28046 4684
rect 28074 4632 28080 4684
rect 28132 4672 28138 4684
rect 28629 4675 28687 4681
rect 28629 4672 28641 4675
rect 28132 4644 28641 4672
rect 28132 4632 28138 4644
rect 28629 4641 28641 4644
rect 28675 4641 28687 4675
rect 28629 4635 28687 4641
rect 26697 4607 26755 4613
rect 26697 4604 26709 4607
rect 26384 4576 26709 4604
rect 26384 4564 26390 4576
rect 26697 4573 26709 4576
rect 26743 4573 26755 4607
rect 26697 4567 26755 4573
rect 27341 4607 27399 4613
rect 27341 4573 27353 4607
rect 27387 4604 27399 4607
rect 27893 4607 27951 4613
rect 27893 4604 27905 4607
rect 27387 4576 27905 4604
rect 27387 4573 27399 4576
rect 27341 4567 27399 4573
rect 27893 4573 27905 4576
rect 27939 4573 27951 4607
rect 29380 4604 29408 4700
rect 29549 4607 29607 4613
rect 29549 4604 29561 4607
rect 29380 4576 29561 4604
rect 27893 4567 27951 4573
rect 29549 4573 29561 4576
rect 29595 4573 29607 4607
rect 29549 4567 29607 4573
rect 30101 4607 30159 4613
rect 30101 4573 30113 4607
rect 30147 4573 30159 4607
rect 30101 4567 30159 4573
rect 25547 4508 26188 4536
rect 26237 4539 26295 4545
rect 25547 4505 25559 4508
rect 25501 4499 25559 4505
rect 26237 4505 26249 4539
rect 26283 4536 26295 4539
rect 27157 4539 27215 4545
rect 27157 4536 27169 4539
rect 26283 4508 27169 4536
rect 26283 4505 26295 4508
rect 26237 4499 26295 4505
rect 27157 4505 27169 4508
rect 27203 4505 27215 4539
rect 30116 4536 30144 4567
rect 30190 4564 30196 4616
rect 30248 4564 30254 4616
rect 30300 4613 30328 4768
rect 30285 4607 30343 4613
rect 30285 4573 30297 4607
rect 30331 4573 30343 4607
rect 30285 4567 30343 4573
rect 30374 4564 30380 4616
rect 30432 4564 30438 4616
rect 30392 4536 30420 4564
rect 30116 4508 30420 4536
rect 27157 4499 27215 4505
rect 25096 4440 25452 4468
rect 26421 4471 26479 4477
rect 25096 4428 25102 4440
rect 26421 4437 26433 4471
rect 26467 4468 26479 4471
rect 27706 4468 27712 4480
rect 26467 4440 27712 4468
rect 26467 4437 26479 4440
rect 26421 4431 26479 4437
rect 27706 4428 27712 4440
rect 27764 4468 27770 4480
rect 31938 4468 31944 4480
rect 27764 4440 31944 4468
rect 27764 4428 27770 4440
rect 31938 4428 31944 4440
rect 31996 4428 32002 4480
rect 1104 4378 38272 4400
rect 1104 4326 4874 4378
rect 4926 4326 4938 4378
rect 4990 4326 5002 4378
rect 5054 4326 5066 4378
rect 5118 4326 5130 4378
rect 5182 4326 35594 4378
rect 35646 4326 35658 4378
rect 35710 4326 35722 4378
rect 35774 4326 35786 4378
rect 35838 4326 35850 4378
rect 35902 4326 38272 4378
rect 1104 4304 38272 4326
rect 9122 4264 9128 4276
rect 8312 4236 9128 4264
rect 8312 4205 8340 4236
rect 9122 4224 9128 4236
rect 9180 4224 9186 4276
rect 9674 4224 9680 4276
rect 9732 4264 9738 4276
rect 9769 4267 9827 4273
rect 9769 4264 9781 4267
rect 9732 4236 9781 4264
rect 9732 4224 9738 4236
rect 9769 4233 9781 4236
rect 9815 4233 9827 4267
rect 9769 4227 9827 4233
rect 14458 4224 14464 4276
rect 14516 4264 14522 4276
rect 14553 4267 14611 4273
rect 14553 4264 14565 4267
rect 14516 4236 14565 4264
rect 14516 4224 14522 4236
rect 14553 4233 14565 4236
rect 14599 4233 14611 4267
rect 14553 4227 14611 4233
rect 20990 4224 20996 4276
rect 21048 4264 21054 4276
rect 25409 4267 25467 4273
rect 21048 4236 25360 4264
rect 21048 4224 21054 4236
rect 8297 4199 8355 4205
rect 8297 4165 8309 4199
rect 8343 4165 8355 4199
rect 8297 4159 8355 4165
rect 8386 4156 8392 4208
rect 8444 4196 8450 4208
rect 8444 4168 8786 4196
rect 8444 4156 8450 4168
rect 22646 4156 22652 4208
rect 22704 4196 22710 4208
rect 23474 4196 23480 4208
rect 22704 4168 23480 4196
rect 22704 4156 22710 4168
rect 23474 4156 23480 4168
rect 23532 4156 23538 4208
rect 25038 4156 25044 4208
rect 25096 4156 25102 4208
rect 25332 4196 25360 4236
rect 25409 4233 25421 4267
rect 25455 4264 25467 4267
rect 26326 4264 26332 4276
rect 25455 4236 26332 4264
rect 25455 4233 25467 4236
rect 25409 4227 25467 4233
rect 26326 4224 26332 4236
rect 26384 4224 26390 4276
rect 27893 4267 27951 4273
rect 27893 4233 27905 4267
rect 27939 4264 27951 4267
rect 27982 4264 27988 4276
rect 27939 4236 27988 4264
rect 27939 4233 27951 4236
rect 27893 4227 27951 4233
rect 27982 4224 27988 4236
rect 28040 4224 28046 4276
rect 29822 4196 29828 4208
rect 25332 4168 29828 4196
rect 6914 4088 6920 4140
rect 6972 4128 6978 4140
rect 8021 4131 8079 4137
rect 8021 4128 8033 4131
rect 6972 4100 8033 4128
rect 6972 4088 6978 4100
rect 8021 4097 8033 4100
rect 8067 4097 8079 4131
rect 8021 4091 8079 4097
rect 14366 4088 14372 4140
rect 14424 4088 14430 4140
rect 24949 4131 25007 4137
rect 24949 4097 24961 4131
rect 24995 4097 25007 4131
rect 25056 4128 25084 4156
rect 25133 4134 25191 4137
rect 25225 4134 25283 4137
rect 25133 4131 25283 4134
rect 25133 4128 25145 4131
rect 25056 4100 25145 4128
rect 24949 4091 25007 4097
rect 25133 4097 25145 4100
rect 25179 4106 25237 4131
rect 25179 4097 25191 4106
rect 25133 4091 25191 4097
rect 25225 4097 25237 4106
rect 25271 4097 25283 4131
rect 25225 4091 25283 4097
rect 25409 4131 25467 4137
rect 25409 4097 25421 4131
rect 25455 4128 25467 4131
rect 25498 4128 25504 4140
rect 25455 4100 25504 4128
rect 25455 4097 25467 4100
rect 25409 4091 25467 4097
rect 24964 3924 24992 4091
rect 25498 4088 25504 4100
rect 25556 4088 25562 4140
rect 28000 4137 28028 4168
rect 29822 4156 29828 4168
rect 29880 4196 29886 4208
rect 30650 4196 30656 4208
rect 29880 4168 30656 4196
rect 29880 4156 29886 4168
rect 30650 4156 30656 4168
rect 30708 4156 30714 4208
rect 27801 4131 27859 4137
rect 27801 4097 27813 4131
rect 27847 4097 27859 4131
rect 27801 4091 27859 4097
rect 27985 4131 28043 4137
rect 27985 4097 27997 4131
rect 28031 4097 28043 4131
rect 27985 4091 28043 4097
rect 27816 4060 27844 4091
rect 30098 4088 30104 4140
rect 30156 4088 30162 4140
rect 30116 4060 30144 4088
rect 27816 4032 30144 4060
rect 25133 3995 25191 4001
rect 25133 3961 25145 3995
rect 25179 3992 25191 3995
rect 25406 3992 25412 4004
rect 25179 3964 25412 3992
rect 25179 3961 25191 3964
rect 25133 3955 25191 3961
rect 25406 3952 25412 3964
rect 25464 3992 25470 4004
rect 27816 3992 27844 4032
rect 25464 3964 27844 3992
rect 25464 3952 25470 3964
rect 25498 3924 25504 3936
rect 24964 3896 25504 3924
rect 25498 3884 25504 3896
rect 25556 3884 25562 3936
rect 1104 3834 38272 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 38272 3834
rect 1104 3760 38272 3782
rect 1104 3290 38272 3312
rect 1104 3238 4874 3290
rect 4926 3238 4938 3290
rect 4990 3238 5002 3290
rect 5054 3238 5066 3290
rect 5118 3238 5130 3290
rect 5182 3238 35594 3290
rect 35646 3238 35658 3290
rect 35710 3238 35722 3290
rect 35774 3238 35786 3290
rect 35838 3238 35850 3290
rect 35902 3238 38272 3290
rect 1104 3216 38272 3238
rect 17218 3136 17224 3188
rect 17276 3136 17282 3188
rect 1946 3000 1952 3052
rect 2004 3000 2010 3052
rect 2406 3000 2412 3052
rect 2464 3000 2470 3052
rect 12526 3000 12532 3052
rect 12584 3000 12590 3052
rect 13170 3000 13176 3052
rect 13228 3000 13234 3052
rect 15102 3000 15108 3052
rect 15160 3000 15166 3052
rect 17236 3049 17264 3136
rect 37550 3068 37556 3120
rect 37608 3068 37614 3120
rect 17221 3043 17279 3049
rect 17221 3009 17233 3043
rect 17267 3009 17279 3043
rect 17221 3003 17279 3009
rect 19981 3043 20039 3049
rect 19981 3009 19993 3043
rect 20027 3040 20039 3043
rect 25590 3040 25596 3052
rect 20027 3012 25596 3040
rect 20027 3009 20039 3012
rect 19981 3003 20039 3009
rect 25590 3000 25596 3012
rect 25648 3000 25654 3052
rect 1762 2796 1768 2848
rect 1820 2796 1826 2848
rect 2222 2796 2228 2848
rect 2280 2796 2286 2848
rect 8386 2796 8392 2848
rect 8444 2836 8450 2848
rect 12345 2839 12403 2845
rect 12345 2836 12357 2839
rect 8444 2808 12357 2836
rect 8444 2796 8450 2808
rect 12345 2805 12357 2808
rect 12391 2805 12403 2839
rect 12345 2799 12403 2805
rect 12986 2796 12992 2848
rect 13044 2796 13050 2848
rect 14918 2796 14924 2848
rect 14976 2796 14982 2848
rect 17402 2796 17408 2848
rect 17460 2796 17466 2848
rect 19794 2796 19800 2848
rect 19852 2796 19858 2848
rect 37182 2796 37188 2848
rect 37240 2836 37246 2848
rect 37645 2839 37703 2845
rect 37645 2836 37657 2839
rect 37240 2808 37657 2836
rect 37240 2796 37246 2808
rect 37645 2805 37657 2808
rect 37691 2805 37703 2839
rect 37645 2799 37703 2805
rect 1104 2746 38272 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 38272 2746
rect 1104 2672 38272 2694
rect 8665 2635 8723 2641
rect 8665 2601 8677 2635
rect 8711 2632 8723 2635
rect 8754 2632 8760 2644
rect 8711 2604 8760 2632
rect 8711 2601 8723 2604
rect 8665 2595 8723 2601
rect 8754 2592 8760 2604
rect 8812 2592 8818 2644
rect 10134 2592 10140 2644
rect 10192 2632 10198 2644
rect 11149 2635 11207 2641
rect 11149 2632 11161 2635
rect 10192 2604 11161 2632
rect 10192 2592 10198 2604
rect 11149 2601 11161 2604
rect 11195 2601 11207 2635
rect 11149 2595 11207 2601
rect 37645 2567 37703 2573
rect 37645 2564 37657 2567
rect 26206 2536 37657 2564
rect 8938 2456 8944 2508
rect 8996 2496 9002 2508
rect 26206 2496 26234 2536
rect 37645 2533 37657 2536
rect 37691 2533 37703 2567
rect 37645 2527 37703 2533
rect 8996 2468 26234 2496
rect 8996 2456 9002 2468
rect 1762 2388 1768 2440
rect 1820 2388 1826 2440
rect 2222 2388 2228 2440
rect 2280 2428 2286 2440
rect 2409 2431 2467 2437
rect 2409 2428 2421 2431
rect 2280 2400 2421 2428
rect 2280 2388 2286 2400
rect 2409 2397 2421 2400
rect 2455 2397 2467 2431
rect 2409 2391 2467 2397
rect 4341 2431 4399 2437
rect 4341 2397 4353 2431
rect 4387 2428 4399 2431
rect 5442 2428 5448 2440
rect 4387 2400 5448 2428
rect 4387 2397 4399 2400
rect 4341 2391 4399 2397
rect 5442 2388 5448 2400
rect 5500 2388 5506 2440
rect 6917 2431 6975 2437
rect 6917 2397 6929 2431
rect 6963 2428 6975 2431
rect 8386 2428 8392 2440
rect 6963 2400 8392 2428
rect 6963 2397 6975 2400
rect 6917 2391 6975 2397
rect 8386 2388 8392 2400
rect 8444 2388 8450 2440
rect 8478 2388 8484 2440
rect 8536 2388 8542 2440
rect 12986 2388 12992 2440
rect 13044 2428 13050 2440
rect 13081 2431 13139 2437
rect 13081 2428 13093 2431
rect 13044 2400 13093 2428
rect 13044 2388 13050 2400
rect 13081 2397 13093 2400
rect 13127 2397 13139 2431
rect 13081 2391 13139 2397
rect 14918 2388 14924 2440
rect 14976 2428 14982 2440
rect 15013 2431 15071 2437
rect 15013 2428 15025 2431
rect 14976 2400 15025 2428
rect 14976 2388 14982 2400
rect 15013 2397 15025 2400
rect 15059 2397 15071 2431
rect 15013 2391 15071 2397
rect 17402 2388 17408 2440
rect 17460 2428 17466 2440
rect 17589 2431 17647 2437
rect 17589 2428 17601 2431
rect 17460 2400 17601 2428
rect 17460 2388 17466 2400
rect 17589 2397 17601 2400
rect 17635 2397 17647 2431
rect 17589 2391 17647 2397
rect 19794 2388 19800 2440
rect 19852 2388 19858 2440
rect 37458 2388 37464 2440
rect 37516 2388 37522 2440
rect 14 2320 20 2372
rect 72 2360 78 2372
rect 1397 2363 1455 2369
rect 1397 2360 1409 2363
rect 72 2332 1409 2360
rect 72 2320 78 2332
rect 1397 2329 1409 2332
rect 1443 2329 1455 2363
rect 1397 2323 1455 2329
rect 2038 2320 2044 2372
rect 2096 2320 2102 2372
rect 3970 2320 3976 2372
rect 4028 2320 4034 2372
rect 6546 2320 6552 2372
rect 6604 2320 6610 2372
rect 10962 2320 10968 2372
rect 11020 2360 11026 2372
rect 11241 2363 11299 2369
rect 11241 2360 11253 2363
rect 11020 2332 11253 2360
rect 11020 2320 11026 2332
rect 11241 2329 11253 2332
rect 11287 2329 11299 2363
rect 11241 2323 11299 2329
rect 14642 2320 14648 2372
rect 14700 2360 14706 2372
rect 14700 2332 19380 2360
rect 14700 2320 14706 2332
rect 12894 2252 12900 2304
rect 12952 2292 12958 2304
rect 13173 2295 13231 2301
rect 13173 2292 13185 2295
rect 12952 2264 13185 2292
rect 12952 2252 12958 2264
rect 13173 2261 13185 2264
rect 13219 2261 13231 2295
rect 13173 2255 13231 2261
rect 15010 2252 15016 2304
rect 15068 2292 15074 2304
rect 15289 2295 15347 2301
rect 15289 2292 15301 2295
rect 15068 2264 15301 2292
rect 15068 2252 15074 2264
rect 15289 2261 15301 2264
rect 15335 2261 15347 2295
rect 15289 2255 15347 2261
rect 17402 2252 17408 2304
rect 17460 2292 17466 2304
rect 17681 2295 17739 2301
rect 17681 2292 17693 2295
rect 17460 2264 17693 2292
rect 17460 2252 17466 2264
rect 17681 2261 17693 2264
rect 17727 2261 17739 2295
rect 19352 2292 19380 2332
rect 19426 2320 19432 2372
rect 19484 2320 19490 2372
rect 27065 2363 27123 2369
rect 27065 2360 27077 2363
rect 26206 2332 27077 2360
rect 26206 2292 26234 2332
rect 27065 2329 27077 2332
rect 27111 2329 27123 2363
rect 27065 2323 27123 2329
rect 19352 2264 26234 2292
rect 17681 2255 17739 2261
rect 26418 2252 26424 2304
rect 26476 2292 26482 2304
rect 27157 2295 27215 2301
rect 27157 2292 27169 2295
rect 26476 2264 27169 2292
rect 26476 2252 26482 2264
rect 27157 2261 27169 2264
rect 27203 2261 27215 2295
rect 27157 2255 27215 2261
rect 1104 2202 38272 2224
rect 1104 2150 4874 2202
rect 4926 2150 4938 2202
rect 4990 2150 5002 2202
rect 5054 2150 5066 2202
rect 5118 2150 5130 2202
rect 5182 2150 35594 2202
rect 35646 2150 35658 2202
rect 35710 2150 35722 2202
rect 35774 2150 35786 2202
rect 35838 2150 35850 2202
rect 35902 2150 38272 2202
rect 1104 2128 38272 2150
<< via1 >>
rect 4874 39142 4926 39194
rect 4938 39142 4990 39194
rect 5002 39142 5054 39194
rect 5066 39142 5118 39194
rect 5130 39142 5182 39194
rect 35594 39142 35646 39194
rect 35658 39142 35710 39194
rect 35722 39142 35774 39194
rect 35786 39142 35838 39194
rect 35850 39142 35902 39194
rect 20 39040 72 39092
rect 4528 39040 4580 39092
rect 9036 39040 9088 39092
rect 11060 39040 11112 39092
rect 13176 39083 13228 39092
rect 13176 39049 13185 39083
rect 13185 39049 13219 39083
rect 13219 39049 13228 39083
rect 13176 39040 13228 39049
rect 17408 39040 17460 39092
rect 21916 39040 21968 39092
rect 26424 39040 26476 39092
rect 33140 39083 33192 39092
rect 33140 39049 33149 39083
rect 33149 39049 33183 39083
rect 33183 39049 33192 39083
rect 33140 39040 33192 39049
rect 35440 39040 35492 39092
rect 12348 38972 12400 39024
rect 15476 38972 15528 39024
rect 30932 38972 30984 39024
rect 1768 38947 1820 38956
rect 1768 38913 1777 38947
rect 1777 38913 1811 38947
rect 1811 38913 1820 38947
rect 1768 38904 1820 38913
rect 5080 38947 5132 38956
rect 5080 38913 5089 38947
rect 5089 38913 5123 38947
rect 5123 38913 5132 38947
rect 5080 38904 5132 38913
rect 9220 38947 9272 38956
rect 9220 38913 9229 38947
rect 9229 38913 9263 38947
rect 9263 38913 9272 38947
rect 9220 38904 9272 38913
rect 12072 38947 12124 38956
rect 12072 38913 12081 38947
rect 12081 38913 12115 38947
rect 12115 38913 12124 38947
rect 12072 38904 12124 38913
rect 12532 38904 12584 38956
rect 17960 38947 18012 38956
rect 17960 38913 17969 38947
rect 17969 38913 18003 38947
rect 18003 38913 18012 38947
rect 17960 38904 18012 38913
rect 19432 38947 19484 38956
rect 19432 38913 19441 38947
rect 19441 38913 19475 38947
rect 19475 38913 19484 38947
rect 19432 38904 19484 38913
rect 20076 38947 20128 38956
rect 20076 38913 20085 38947
rect 20085 38913 20119 38947
rect 20119 38913 20128 38947
rect 20076 38904 20128 38913
rect 22376 38947 22428 38956
rect 22376 38913 22385 38947
rect 22385 38913 22419 38947
rect 22419 38913 22428 38947
rect 22376 38904 22428 38913
rect 27068 38947 27120 38956
rect 27068 38913 27077 38947
rect 27077 38913 27111 38947
rect 27111 38913 27120 38947
rect 27068 38904 27120 38913
rect 27712 38947 27764 38956
rect 27712 38913 27721 38947
rect 27721 38913 27755 38947
rect 27755 38913 27764 38947
rect 27712 38904 27764 38913
rect 33048 38947 33100 38956
rect 33048 38913 33057 38947
rect 33057 38913 33091 38947
rect 33091 38913 33100 38947
rect 33048 38904 33100 38913
rect 35624 38947 35676 38956
rect 35624 38913 35633 38947
rect 35633 38913 35667 38947
rect 35667 38913 35676 38947
rect 35624 38904 35676 38913
rect 37372 38904 37424 38956
rect 14004 38836 14056 38888
rect 15568 38811 15620 38820
rect 15568 38777 15577 38811
rect 15577 38777 15611 38811
rect 15611 38777 15620 38811
rect 15568 38768 15620 38777
rect 29736 38768 29788 38820
rect 37648 38811 37700 38820
rect 37648 38777 37657 38811
rect 37657 38777 37691 38811
rect 37691 38777 37700 38811
rect 37648 38768 37700 38777
rect 12808 38700 12860 38752
rect 19616 38743 19668 38752
rect 19616 38709 19625 38743
rect 19625 38709 19659 38743
rect 19659 38709 19668 38743
rect 19616 38700 19668 38709
rect 27620 38743 27672 38752
rect 27620 38709 27629 38743
rect 27629 38709 27663 38743
rect 27663 38709 27672 38743
rect 27620 38700 27672 38709
rect 4214 38598 4266 38650
rect 4278 38598 4330 38650
rect 4342 38598 4394 38650
rect 4406 38598 4458 38650
rect 4470 38598 4522 38650
rect 34934 38598 34986 38650
rect 34998 38598 35050 38650
rect 35062 38598 35114 38650
rect 35126 38598 35178 38650
rect 35190 38598 35242 38650
rect 5080 38496 5132 38548
rect 9220 38496 9272 38548
rect 17960 38496 18012 38548
rect 13636 38428 13688 38480
rect 22468 38496 22520 38548
rect 12716 38360 12768 38412
rect 5172 38335 5224 38344
rect 5172 38301 5181 38335
rect 5181 38301 5215 38335
rect 5215 38301 5224 38335
rect 5172 38292 5224 38301
rect 8576 38335 8628 38344
rect 8576 38301 8585 38335
rect 8585 38301 8619 38335
rect 8619 38301 8628 38335
rect 8576 38292 8628 38301
rect 9036 38335 9088 38344
rect 9036 38301 9045 38335
rect 9045 38301 9079 38335
rect 9079 38301 9088 38335
rect 9036 38292 9088 38301
rect 13452 38292 13504 38344
rect 9588 38267 9640 38276
rect 9588 38233 9597 38267
rect 9597 38233 9631 38267
rect 9631 38233 9640 38267
rect 9588 38224 9640 38233
rect 10232 38224 10284 38276
rect 9128 38156 9180 38208
rect 12808 38267 12860 38276
rect 12808 38233 12817 38267
rect 12817 38233 12851 38267
rect 12851 38233 12860 38267
rect 12808 38224 12860 38233
rect 11244 38156 11296 38208
rect 11336 38199 11388 38208
rect 11336 38165 11345 38199
rect 11345 38165 11379 38199
rect 11379 38165 11388 38199
rect 11336 38156 11388 38165
rect 18512 38335 18564 38344
rect 18512 38301 18521 38335
rect 18521 38301 18555 38335
rect 18555 38301 18564 38335
rect 18512 38292 18564 38301
rect 19616 38360 19668 38412
rect 21180 38292 21232 38344
rect 21272 38335 21324 38344
rect 21272 38301 21281 38335
rect 21281 38301 21315 38335
rect 21315 38301 21324 38335
rect 21272 38292 21324 38301
rect 27712 38496 27764 38548
rect 26056 38360 26108 38412
rect 20996 38199 21048 38208
rect 20996 38165 21005 38199
rect 21005 38165 21039 38199
rect 21039 38165 21048 38199
rect 20996 38156 21048 38165
rect 23480 38156 23532 38208
rect 25596 38267 25648 38276
rect 25596 38233 25605 38267
rect 25605 38233 25639 38267
rect 25639 38233 25648 38267
rect 25596 38224 25648 38233
rect 26056 38224 26108 38276
rect 26516 38156 26568 38208
rect 27620 38360 27672 38412
rect 33048 38496 33100 38548
rect 35624 38496 35676 38548
rect 37924 38496 37976 38548
rect 29644 38403 29696 38412
rect 29644 38369 29653 38403
rect 29653 38369 29687 38403
rect 29687 38369 29696 38403
rect 29644 38360 29696 38369
rect 29552 38335 29604 38344
rect 29552 38301 29561 38335
rect 29561 38301 29595 38335
rect 29595 38301 29604 38335
rect 29552 38292 29604 38301
rect 27528 38267 27580 38276
rect 27528 38233 27537 38267
rect 27537 38233 27571 38267
rect 27571 38233 27580 38267
rect 27528 38224 27580 38233
rect 29276 38267 29328 38276
rect 29276 38233 29285 38267
rect 29285 38233 29319 38267
rect 29319 38233 29328 38267
rect 29276 38224 29328 38233
rect 29460 38224 29512 38276
rect 31668 38224 31720 38276
rect 28540 38156 28592 38208
rect 30380 38156 30432 38208
rect 31116 38156 31168 38208
rect 4874 38054 4926 38106
rect 4938 38054 4990 38106
rect 5002 38054 5054 38106
rect 5066 38054 5118 38106
rect 5130 38054 5182 38106
rect 35594 38054 35646 38106
rect 35658 38054 35710 38106
rect 35722 38054 35774 38106
rect 35786 38054 35838 38106
rect 35850 38054 35902 38106
rect 9588 37952 9640 38004
rect 11336 37952 11388 38004
rect 11888 37995 11940 38004
rect 11888 37961 11897 37995
rect 11897 37961 11931 37995
rect 11931 37961 11940 37995
rect 11888 37952 11940 37961
rect 12072 37952 12124 38004
rect 12348 37995 12400 38004
rect 12348 37961 12357 37995
rect 12357 37961 12391 37995
rect 12391 37961 12400 37995
rect 12348 37952 12400 37961
rect 13636 37952 13688 38004
rect 11244 37816 11296 37868
rect 10784 37791 10836 37800
rect 10784 37757 10793 37791
rect 10793 37757 10827 37791
rect 10827 37757 10836 37791
rect 10784 37748 10836 37757
rect 13176 37816 13228 37868
rect 10600 37612 10652 37664
rect 11888 37748 11940 37800
rect 13084 37748 13136 37800
rect 13820 37859 13872 37868
rect 13820 37825 13829 37859
rect 13829 37825 13863 37859
rect 13863 37825 13872 37859
rect 13820 37816 13872 37825
rect 14096 37816 14148 37868
rect 14372 37859 14424 37868
rect 14372 37825 14376 37859
rect 14376 37825 14410 37859
rect 14410 37825 14424 37859
rect 14372 37816 14424 37825
rect 13268 37680 13320 37732
rect 15292 37816 15344 37868
rect 15936 37859 15988 37868
rect 15936 37825 15945 37859
rect 15945 37825 15979 37859
rect 15979 37825 15988 37859
rect 15936 37816 15988 37825
rect 16120 37859 16172 37868
rect 16120 37825 16129 37859
rect 16129 37825 16163 37859
rect 16163 37825 16172 37859
rect 16120 37816 16172 37825
rect 16212 37859 16264 37868
rect 16212 37825 16221 37859
rect 16221 37825 16255 37859
rect 16255 37825 16264 37859
rect 16212 37816 16264 37825
rect 16948 37884 17000 37936
rect 16396 37816 16448 37868
rect 16856 37859 16908 37868
rect 16856 37825 16865 37859
rect 16865 37825 16899 37859
rect 16899 37825 16908 37859
rect 16856 37816 16908 37825
rect 17316 37816 17368 37868
rect 17776 37816 17828 37868
rect 17868 37816 17920 37868
rect 12440 37612 12492 37664
rect 15384 37680 15436 37732
rect 16856 37680 16908 37732
rect 16488 37655 16540 37664
rect 16488 37621 16497 37655
rect 16497 37621 16531 37655
rect 16531 37621 16540 37655
rect 16488 37612 16540 37621
rect 17776 37655 17828 37664
rect 17776 37621 17785 37655
rect 17785 37621 17819 37655
rect 17819 37621 17828 37655
rect 17776 37612 17828 37621
rect 18512 37952 18564 38004
rect 19432 37995 19484 38004
rect 19432 37961 19441 37995
rect 19441 37961 19475 37995
rect 19475 37961 19484 37995
rect 19432 37952 19484 37961
rect 20996 37952 21048 38004
rect 21272 37952 21324 38004
rect 20352 37859 20404 37868
rect 20352 37825 20361 37859
rect 20361 37825 20395 37859
rect 20395 37825 20404 37859
rect 20352 37816 20404 37825
rect 20536 37884 20588 37936
rect 19340 37748 19392 37800
rect 19984 37791 20036 37800
rect 19984 37757 19993 37791
rect 19993 37757 20027 37791
rect 20027 37757 20036 37791
rect 19984 37748 20036 37757
rect 21180 37748 21232 37800
rect 20536 37680 20588 37732
rect 25596 37952 25648 38004
rect 27528 37952 27580 38004
rect 29460 37952 29512 38004
rect 29644 37952 29696 38004
rect 23020 37816 23072 37868
rect 23480 37816 23532 37868
rect 23664 37859 23716 37868
rect 23664 37825 23673 37859
rect 23673 37825 23707 37859
rect 23707 37825 23716 37859
rect 23664 37816 23716 37825
rect 23940 37816 23992 37868
rect 24124 37816 24176 37868
rect 22468 37791 22520 37800
rect 22468 37757 22477 37791
rect 22477 37757 22511 37791
rect 22511 37757 22520 37791
rect 22468 37748 22520 37757
rect 22560 37791 22612 37800
rect 22560 37757 22569 37791
rect 22569 37757 22603 37791
rect 22603 37757 22612 37791
rect 22560 37748 22612 37757
rect 25320 37859 25372 37868
rect 25320 37825 25329 37859
rect 25329 37825 25363 37859
rect 25363 37825 25372 37859
rect 25320 37816 25372 37825
rect 25780 37927 25832 37936
rect 25780 37893 25789 37927
rect 25789 37893 25823 37927
rect 25823 37893 25832 37927
rect 25780 37884 25832 37893
rect 25872 37816 25924 37868
rect 25228 37791 25280 37800
rect 25228 37757 25237 37791
rect 25237 37757 25271 37791
rect 25271 37757 25280 37791
rect 25228 37748 25280 37757
rect 26424 37859 26476 37868
rect 26424 37825 26433 37859
rect 26433 37825 26467 37859
rect 26467 37825 26476 37859
rect 26424 37816 26476 37825
rect 26608 37859 26660 37868
rect 26608 37825 26617 37859
rect 26617 37825 26651 37859
rect 26651 37825 26660 37859
rect 26608 37816 26660 37825
rect 29000 37816 29052 37868
rect 30380 37884 30432 37936
rect 31208 37859 31260 37868
rect 31208 37825 31217 37859
rect 31217 37825 31251 37859
rect 31251 37825 31260 37859
rect 31208 37816 31260 37825
rect 26148 37748 26200 37800
rect 27068 37748 27120 37800
rect 27988 37791 28040 37800
rect 27988 37757 27997 37791
rect 27997 37757 28031 37791
rect 28031 37757 28040 37791
rect 27988 37748 28040 37757
rect 29460 37748 29512 37800
rect 31668 37748 31720 37800
rect 23848 37612 23900 37664
rect 24584 37612 24636 37664
rect 25964 37612 26016 37664
rect 30932 37612 30984 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 16488 37408 16540 37460
rect 20352 37408 20404 37460
rect 24676 37408 24728 37460
rect 26424 37408 26476 37460
rect 26608 37408 26660 37460
rect 8392 37272 8444 37324
rect 17776 37272 17828 37324
rect 17960 37272 18012 37324
rect 22836 37315 22888 37324
rect 22836 37281 22845 37315
rect 22845 37281 22879 37315
rect 22879 37281 22888 37315
rect 22836 37272 22888 37281
rect 22928 37315 22980 37324
rect 22928 37281 22937 37315
rect 22937 37281 22971 37315
rect 22971 37281 22980 37315
rect 22928 37272 22980 37281
rect 23848 37272 23900 37324
rect 24860 37272 24912 37324
rect 8300 37247 8352 37256
rect 8300 37213 8309 37247
rect 8309 37213 8343 37247
rect 8343 37213 8352 37247
rect 8300 37204 8352 37213
rect 940 37136 992 37188
rect 6920 37136 6972 37188
rect 10232 37204 10284 37256
rect 17776 37179 17828 37188
rect 17776 37145 17785 37179
rect 17785 37145 17819 37179
rect 17819 37145 17828 37179
rect 17776 37136 17828 37145
rect 18604 37247 18656 37256
rect 18604 37213 18613 37247
rect 18613 37213 18647 37247
rect 18647 37213 18656 37247
rect 18604 37204 18656 37213
rect 20168 37247 20220 37256
rect 20168 37213 20177 37247
rect 20177 37213 20211 37247
rect 20211 37213 20220 37247
rect 20168 37204 20220 37213
rect 22468 37204 22520 37256
rect 23388 37204 23440 37256
rect 24032 37204 24084 37256
rect 24308 37204 24360 37256
rect 26516 37272 26568 37324
rect 10692 37111 10744 37120
rect 10692 37077 10701 37111
rect 10701 37077 10735 37111
rect 10735 37077 10744 37111
rect 10692 37068 10744 37077
rect 17224 37068 17276 37120
rect 19892 37136 19944 37188
rect 20720 37179 20772 37188
rect 20720 37145 20729 37179
rect 20729 37145 20763 37179
rect 20763 37145 20772 37179
rect 20720 37136 20772 37145
rect 21180 37136 21232 37188
rect 18972 37068 19024 37120
rect 22376 37111 22428 37120
rect 22376 37077 22385 37111
rect 22385 37077 22419 37111
rect 22419 37077 22428 37111
rect 22376 37068 22428 37077
rect 23756 37136 23808 37188
rect 28632 37272 28684 37324
rect 28908 37272 28960 37324
rect 29552 37272 29604 37324
rect 27344 37204 27396 37256
rect 29276 37204 29328 37256
rect 30932 37272 30984 37324
rect 32588 37247 32640 37256
rect 32588 37213 32597 37247
rect 32597 37213 32631 37247
rect 32631 37213 32640 37247
rect 32588 37204 32640 37213
rect 27896 37136 27948 37188
rect 30104 37136 30156 37188
rect 30472 37136 30524 37188
rect 31484 37136 31536 37188
rect 24400 37068 24452 37120
rect 27528 37068 27580 37120
rect 30012 37068 30064 37120
rect 32496 37111 32548 37120
rect 32496 37077 32505 37111
rect 32505 37077 32539 37111
rect 32539 37077 32548 37111
rect 32496 37068 32548 37077
rect 37832 37111 37884 37120
rect 37832 37077 37841 37111
rect 37841 37077 37875 37111
rect 37875 37077 37884 37111
rect 37832 37068 37884 37077
rect 4874 36966 4926 37018
rect 4938 36966 4990 37018
rect 5002 36966 5054 37018
rect 5066 36966 5118 37018
rect 5130 36966 5182 37018
rect 35594 36966 35646 37018
rect 35658 36966 35710 37018
rect 35722 36966 35774 37018
rect 35786 36966 35838 37018
rect 35850 36966 35902 37018
rect 8300 36864 8352 36916
rect 10692 36864 10744 36916
rect 20720 36864 20772 36916
rect 8392 36796 8444 36848
rect 10600 36728 10652 36780
rect 16948 36728 17000 36780
rect 18696 36728 18748 36780
rect 22376 36864 22428 36916
rect 22468 36864 22520 36916
rect 23388 36864 23440 36916
rect 9128 36660 9180 36712
rect 9864 36703 9916 36712
rect 9864 36669 9873 36703
rect 9873 36669 9907 36703
rect 9907 36669 9916 36703
rect 9864 36660 9916 36669
rect 15568 36660 15620 36712
rect 17960 36660 18012 36712
rect 17040 36592 17092 36644
rect 19708 36592 19760 36644
rect 22284 36660 22336 36712
rect 24492 36771 24544 36780
rect 24492 36737 24501 36771
rect 24501 36737 24535 36771
rect 24535 36737 24544 36771
rect 24492 36728 24544 36737
rect 24584 36728 24636 36780
rect 27804 36864 27856 36916
rect 29000 36864 29052 36916
rect 30012 36864 30064 36916
rect 31208 36864 31260 36916
rect 31484 36864 31536 36916
rect 32496 36864 32548 36916
rect 25136 36796 25188 36848
rect 25596 36728 25648 36780
rect 27712 36771 27764 36780
rect 27712 36737 27721 36771
rect 27721 36737 27755 36771
rect 27755 36737 27764 36771
rect 27712 36728 27764 36737
rect 28172 36728 28224 36780
rect 28264 36771 28316 36780
rect 28264 36737 28273 36771
rect 28273 36737 28307 36771
rect 28307 36737 28316 36771
rect 28264 36728 28316 36737
rect 29368 36728 29420 36780
rect 29644 36703 29696 36712
rect 29644 36669 29653 36703
rect 29653 36669 29687 36703
rect 29687 36669 29696 36703
rect 29644 36660 29696 36669
rect 7656 36524 7708 36576
rect 12992 36524 13044 36576
rect 13728 36524 13780 36576
rect 14096 36524 14148 36576
rect 14832 36524 14884 36576
rect 15752 36524 15804 36576
rect 23296 36524 23348 36576
rect 24216 36592 24268 36644
rect 24032 36524 24084 36576
rect 24676 36567 24728 36576
rect 24676 36533 24685 36567
rect 24685 36533 24719 36567
rect 24719 36533 24728 36567
rect 24676 36524 24728 36533
rect 24952 36567 25004 36576
rect 24952 36533 24961 36567
rect 24961 36533 24995 36567
rect 24995 36533 25004 36567
rect 24952 36524 25004 36533
rect 27436 36524 27488 36576
rect 28448 36567 28500 36576
rect 28448 36533 28457 36567
rect 28457 36533 28491 36567
rect 28491 36533 28500 36567
rect 28448 36524 28500 36533
rect 28632 36524 28684 36576
rect 30104 36660 30156 36712
rect 33692 36728 33744 36780
rect 32220 36660 32272 36712
rect 33140 36524 33192 36576
rect 34060 36567 34112 36576
rect 34060 36533 34069 36567
rect 34069 36533 34103 36567
rect 34103 36533 34112 36567
rect 34060 36524 34112 36533
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 10692 36320 10744 36372
rect 13820 36320 13872 36372
rect 9036 36184 9088 36236
rect 4712 36116 4764 36168
rect 9772 36159 9824 36168
rect 9772 36125 9781 36159
rect 9781 36125 9815 36159
rect 9815 36125 9824 36159
rect 9772 36116 9824 36125
rect 11244 36159 11296 36168
rect 11244 36125 11253 36159
rect 11253 36125 11287 36159
rect 11287 36125 11296 36159
rect 11244 36116 11296 36125
rect 11520 36159 11572 36168
rect 11520 36125 11529 36159
rect 11529 36125 11563 36159
rect 11563 36125 11572 36159
rect 11520 36116 11572 36125
rect 11796 36116 11848 36168
rect 13268 36159 13320 36168
rect 6276 36091 6328 36100
rect 6276 36057 6285 36091
rect 6285 36057 6319 36091
rect 6319 36057 6328 36091
rect 6276 36048 6328 36057
rect 6644 35980 6696 36032
rect 7656 36048 7708 36100
rect 10232 36048 10284 36100
rect 11428 36091 11480 36100
rect 11428 36057 11437 36091
rect 11437 36057 11471 36091
rect 11471 36057 11480 36091
rect 11428 36048 11480 36057
rect 11704 36048 11756 36100
rect 12440 36048 12492 36100
rect 12808 36048 12860 36100
rect 13268 36125 13276 36159
rect 13276 36125 13310 36159
rect 13310 36125 13320 36159
rect 13268 36116 13320 36125
rect 13820 36116 13872 36168
rect 14280 36159 14332 36168
rect 14280 36125 14289 36159
rect 14289 36125 14323 36159
rect 14323 36125 14332 36159
rect 14280 36116 14332 36125
rect 15936 36320 15988 36372
rect 17776 36320 17828 36372
rect 19892 36320 19944 36372
rect 14832 36184 14884 36236
rect 12992 36091 13044 36100
rect 12992 36057 13001 36091
rect 13001 36057 13035 36091
rect 13035 36057 13044 36091
rect 12992 36048 13044 36057
rect 15200 36116 15252 36168
rect 15568 36184 15620 36236
rect 15752 36159 15804 36168
rect 15752 36125 15761 36159
rect 15761 36125 15795 36159
rect 15795 36125 15804 36159
rect 15752 36116 15804 36125
rect 7748 36023 7800 36032
rect 7748 35989 7757 36023
rect 7757 35989 7791 36023
rect 7791 35989 7800 36023
rect 7748 35980 7800 35989
rect 9220 35980 9272 36032
rect 9588 36023 9640 36032
rect 9588 35989 9597 36023
rect 9597 35989 9631 36023
rect 9631 35989 9640 36023
rect 9588 35980 9640 35989
rect 11336 35980 11388 36032
rect 12624 35980 12676 36032
rect 13820 35980 13872 36032
rect 14464 35980 14516 36032
rect 15476 36048 15528 36100
rect 15292 36023 15344 36032
rect 15292 35989 15301 36023
rect 15301 35989 15335 36023
rect 15335 35989 15344 36023
rect 15292 35980 15344 35989
rect 15660 35980 15712 36032
rect 16212 36159 16264 36168
rect 16212 36125 16221 36159
rect 16221 36125 16255 36159
rect 16255 36125 16264 36159
rect 16212 36116 16264 36125
rect 16672 36116 16724 36168
rect 16856 36159 16908 36168
rect 16856 36125 16866 36159
rect 16866 36125 16900 36159
rect 16900 36125 16908 36159
rect 16856 36116 16908 36125
rect 18604 36252 18656 36304
rect 24492 36320 24544 36372
rect 28264 36320 28316 36372
rect 30104 36320 30156 36372
rect 17316 36116 17368 36168
rect 16948 36048 17000 36100
rect 17040 36091 17092 36100
rect 17040 36057 17049 36091
rect 17049 36057 17083 36091
rect 17083 36057 17092 36091
rect 17040 36048 17092 36057
rect 17592 36116 17644 36168
rect 18052 36116 18104 36168
rect 18696 36159 18748 36168
rect 18696 36125 18705 36159
rect 18705 36125 18739 36159
rect 18739 36125 18748 36159
rect 18696 36116 18748 36125
rect 19800 36227 19852 36236
rect 19800 36193 19809 36227
rect 19809 36193 19843 36227
rect 19843 36193 19852 36227
rect 19800 36184 19852 36193
rect 22100 36116 22152 36168
rect 22836 36116 22888 36168
rect 23204 36116 23256 36168
rect 24216 36252 24268 36304
rect 25688 36252 25740 36304
rect 26148 36252 26200 36304
rect 25228 36184 25280 36236
rect 29828 36252 29880 36304
rect 24676 36116 24728 36168
rect 25596 36116 25648 36168
rect 26332 36116 26384 36168
rect 26516 36116 26568 36168
rect 17684 36091 17736 36100
rect 17684 36057 17693 36091
rect 17693 36057 17727 36091
rect 17727 36057 17736 36091
rect 17684 36048 17736 36057
rect 17960 36048 18012 36100
rect 17408 36023 17460 36032
rect 17408 35989 17417 36023
rect 17417 35989 17451 36023
rect 17451 35989 17460 36023
rect 17408 35980 17460 35989
rect 18604 36023 18656 36032
rect 18604 35989 18613 36023
rect 18613 35989 18647 36023
rect 18647 35989 18656 36023
rect 18604 35980 18656 35989
rect 18788 36048 18840 36100
rect 19892 36048 19944 36100
rect 20536 36048 20588 36100
rect 21364 36048 21416 36100
rect 22652 35980 22704 36032
rect 23572 35980 23624 36032
rect 24124 36048 24176 36100
rect 24492 36048 24544 36100
rect 25044 36048 25096 36100
rect 25412 36048 25464 36100
rect 27160 36116 27212 36168
rect 27252 36159 27304 36168
rect 27252 36125 27261 36159
rect 27261 36125 27295 36159
rect 27295 36125 27304 36159
rect 27252 36116 27304 36125
rect 27344 36159 27396 36168
rect 27344 36125 27354 36159
rect 27354 36125 27388 36159
rect 27388 36125 27396 36159
rect 28724 36227 28776 36236
rect 28724 36193 28733 36227
rect 28733 36193 28767 36227
rect 28767 36193 28776 36227
rect 28724 36184 28776 36193
rect 32220 36363 32272 36372
rect 32220 36329 32229 36363
rect 32229 36329 32263 36363
rect 32263 36329 32272 36363
rect 32220 36320 32272 36329
rect 34060 36320 34112 36372
rect 32404 36184 32456 36236
rect 27344 36116 27396 36125
rect 27988 36116 28040 36168
rect 28540 36159 28592 36168
rect 28540 36125 28549 36159
rect 28549 36125 28583 36159
rect 28583 36125 28592 36159
rect 28540 36116 28592 36125
rect 28816 36116 28868 36168
rect 30012 36116 30064 36168
rect 25872 35980 25924 36032
rect 31852 36048 31904 36100
rect 30748 35980 30800 36032
rect 33140 35980 33192 36032
rect 33600 35980 33652 36032
rect 4874 35878 4926 35930
rect 4938 35878 4990 35930
rect 5002 35878 5054 35930
rect 5066 35878 5118 35930
rect 5130 35878 5182 35930
rect 35594 35878 35646 35930
rect 35658 35878 35710 35930
rect 35722 35878 35774 35930
rect 35786 35878 35838 35930
rect 35850 35878 35902 35930
rect 6276 35776 6328 35828
rect 7748 35776 7800 35828
rect 8208 35776 8260 35828
rect 9036 35776 9088 35828
rect 12716 35776 12768 35828
rect 9588 35708 9640 35760
rect 10232 35708 10284 35760
rect 14280 35776 14332 35828
rect 20996 35776 21048 35828
rect 22468 35776 22520 35828
rect 22652 35776 22704 35828
rect 18604 35708 18656 35760
rect 20444 35708 20496 35760
rect 9128 35683 9180 35692
rect 9128 35649 9137 35683
rect 9137 35649 9171 35683
rect 9171 35649 9180 35683
rect 9128 35640 9180 35649
rect 13176 35640 13228 35692
rect 13360 35640 13412 35692
rect 13728 35683 13780 35692
rect 13728 35649 13737 35683
rect 13737 35649 13771 35683
rect 13771 35649 13780 35683
rect 13728 35640 13780 35649
rect 13820 35640 13872 35692
rect 7840 35615 7892 35624
rect 7840 35581 7849 35615
rect 7849 35581 7883 35615
rect 7883 35581 7892 35615
rect 7840 35572 7892 35581
rect 8116 35572 8168 35624
rect 8300 35615 8352 35624
rect 8300 35581 8309 35615
rect 8309 35581 8343 35615
rect 8343 35581 8352 35615
rect 8300 35572 8352 35581
rect 9220 35615 9272 35624
rect 9220 35581 9229 35615
rect 9229 35581 9263 35615
rect 9263 35581 9272 35615
rect 9220 35572 9272 35581
rect 16212 35572 16264 35624
rect 11060 35504 11112 35556
rect 11244 35504 11296 35556
rect 12440 35436 12492 35488
rect 18696 35479 18748 35488
rect 18696 35445 18705 35479
rect 18705 35445 18739 35479
rect 18739 35445 18748 35479
rect 18696 35436 18748 35445
rect 18880 35683 18932 35692
rect 18880 35649 18889 35683
rect 18889 35649 18923 35683
rect 18923 35649 18932 35683
rect 18880 35640 18932 35649
rect 20076 35640 20128 35692
rect 21088 35683 21140 35692
rect 21088 35649 21097 35683
rect 21097 35649 21131 35683
rect 21131 35649 21140 35683
rect 21088 35640 21140 35649
rect 21180 35683 21232 35692
rect 21180 35649 21189 35683
rect 21189 35649 21223 35683
rect 21223 35649 21232 35683
rect 21180 35640 21232 35649
rect 22192 35683 22244 35692
rect 22192 35649 22201 35683
rect 22201 35649 22235 35683
rect 22235 35649 22244 35683
rect 22192 35640 22244 35649
rect 22284 35683 22336 35692
rect 22284 35649 22293 35683
rect 22293 35649 22327 35683
rect 22327 35649 22336 35683
rect 22284 35640 22336 35649
rect 22376 35683 22428 35692
rect 22376 35649 22390 35683
rect 22390 35649 22424 35683
rect 22424 35649 22428 35683
rect 22376 35640 22428 35649
rect 22744 35640 22796 35692
rect 23664 35708 23716 35760
rect 23112 35683 23164 35692
rect 23112 35649 23121 35683
rect 23121 35649 23155 35683
rect 23155 35649 23164 35683
rect 23112 35640 23164 35649
rect 23204 35683 23256 35692
rect 23204 35649 23213 35683
rect 23213 35649 23247 35683
rect 23247 35649 23256 35683
rect 23204 35640 23256 35649
rect 23296 35683 23348 35692
rect 23296 35649 23310 35683
rect 23310 35649 23344 35683
rect 23344 35649 23348 35683
rect 23296 35640 23348 35649
rect 23572 35640 23624 35692
rect 21548 35572 21600 35624
rect 19800 35504 19852 35556
rect 22836 35504 22888 35556
rect 23388 35504 23440 35556
rect 23940 35683 23992 35692
rect 23940 35649 23949 35683
rect 23949 35649 23983 35683
rect 23983 35649 23992 35683
rect 23940 35640 23992 35649
rect 24860 35683 24912 35692
rect 24860 35649 24869 35683
rect 24869 35649 24903 35683
rect 24903 35649 24912 35683
rect 24860 35640 24912 35649
rect 27804 35776 27856 35828
rect 25044 35751 25096 35760
rect 25044 35717 25053 35751
rect 25053 35717 25087 35751
rect 25087 35717 25096 35751
rect 25044 35708 25096 35717
rect 25228 35683 25280 35692
rect 25228 35649 25237 35683
rect 25237 35649 25271 35683
rect 25271 35649 25280 35683
rect 25228 35640 25280 35649
rect 25596 35708 25648 35760
rect 28724 35708 28776 35760
rect 21456 35436 21508 35488
rect 21824 35436 21876 35488
rect 23020 35436 23072 35488
rect 23480 35479 23532 35488
rect 23480 35445 23489 35479
rect 23489 35445 23523 35479
rect 23523 35445 23532 35479
rect 23480 35436 23532 35445
rect 24124 35436 24176 35488
rect 25504 35615 25556 35624
rect 25504 35581 25513 35615
rect 25513 35581 25547 35615
rect 25547 35581 25556 35615
rect 25504 35572 25556 35581
rect 25596 35572 25648 35624
rect 25872 35640 25924 35692
rect 26056 35683 26108 35692
rect 26056 35649 26065 35683
rect 26065 35649 26099 35683
rect 26099 35649 26108 35683
rect 26056 35640 26108 35649
rect 26240 35683 26292 35692
rect 26240 35649 26249 35683
rect 26249 35649 26283 35683
rect 26283 35649 26292 35683
rect 26240 35640 26292 35649
rect 26516 35683 26568 35692
rect 26516 35649 26525 35683
rect 26525 35649 26559 35683
rect 26559 35649 26568 35683
rect 26516 35640 26568 35649
rect 27344 35640 27396 35692
rect 30472 35708 30524 35760
rect 27436 35615 27488 35624
rect 27436 35581 27445 35615
rect 27445 35581 27479 35615
rect 27479 35581 27488 35615
rect 27436 35572 27488 35581
rect 28172 35572 28224 35624
rect 28264 35572 28316 35624
rect 29828 35640 29880 35692
rect 30012 35683 30064 35692
rect 30012 35649 30021 35683
rect 30021 35649 30055 35683
rect 30055 35649 30064 35683
rect 30012 35640 30064 35649
rect 30196 35640 30248 35692
rect 30748 35819 30800 35828
rect 30748 35785 30757 35819
rect 30757 35785 30791 35819
rect 30791 35785 30800 35819
rect 30748 35776 30800 35785
rect 32588 35708 32640 35760
rect 31392 35683 31444 35692
rect 31392 35649 31401 35683
rect 31401 35649 31435 35683
rect 31435 35649 31444 35683
rect 31392 35640 31444 35649
rect 33508 35683 33560 35692
rect 33508 35649 33517 35683
rect 33517 35649 33551 35683
rect 33551 35649 33560 35683
rect 33508 35640 33560 35649
rect 31484 35572 31536 35624
rect 26148 35436 26200 35488
rect 26608 35436 26660 35488
rect 26884 35436 26936 35488
rect 29644 35436 29696 35488
rect 30104 35436 30156 35488
rect 31024 35436 31076 35488
rect 32772 35436 32824 35488
rect 33324 35479 33376 35488
rect 33324 35445 33333 35479
rect 33333 35445 33367 35479
rect 33367 35445 33376 35479
rect 33324 35436 33376 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 9772 35232 9824 35284
rect 18880 35232 18932 35284
rect 27988 35232 28040 35284
rect 30196 35232 30248 35284
rect 30656 35232 30708 35284
rect 6920 35164 6972 35216
rect 22836 35164 22888 35216
rect 7932 35096 7984 35148
rect 8300 35028 8352 35080
rect 9680 35096 9732 35148
rect 10784 35096 10836 35148
rect 23572 35139 23624 35148
rect 23572 35105 23581 35139
rect 23581 35105 23615 35139
rect 23615 35105 23624 35139
rect 23572 35096 23624 35105
rect 24124 35164 24176 35216
rect 11152 35028 11204 35080
rect 7196 35003 7248 35012
rect 7196 34969 7205 35003
rect 7205 34969 7239 35003
rect 7239 34969 7248 35003
rect 7196 34960 7248 34969
rect 12440 34960 12492 35012
rect 17316 35071 17368 35080
rect 17316 35037 17325 35071
rect 17325 35037 17359 35071
rect 17359 35037 17368 35071
rect 17316 35028 17368 35037
rect 21824 34960 21876 35012
rect 8484 34892 8536 34944
rect 15936 34892 15988 34944
rect 19340 34892 19392 34944
rect 20720 34892 20772 34944
rect 25320 35071 25372 35080
rect 25320 35037 25329 35071
rect 25329 35037 25363 35071
rect 25363 35037 25372 35071
rect 25320 35028 25372 35037
rect 25504 35071 25556 35080
rect 25504 35037 25513 35071
rect 25513 35037 25547 35071
rect 25547 35037 25556 35071
rect 25504 35028 25556 35037
rect 26608 35096 26660 35148
rect 25872 35028 25924 35080
rect 26332 35071 26384 35080
rect 26332 35037 26341 35071
rect 26341 35037 26375 35071
rect 26375 35037 26384 35071
rect 26332 35028 26384 35037
rect 26424 35071 26476 35080
rect 26424 35037 26433 35071
rect 26433 35037 26467 35071
rect 26467 35037 26476 35071
rect 26424 35028 26476 35037
rect 28172 35207 28224 35216
rect 28172 35173 28181 35207
rect 28181 35173 28215 35207
rect 28215 35173 28224 35207
rect 28172 35164 28224 35173
rect 28356 35164 28408 35216
rect 32772 35232 32824 35284
rect 32312 35164 32364 35216
rect 23480 34892 23532 34944
rect 23572 34892 23624 34944
rect 25688 34892 25740 34944
rect 27528 34960 27580 35012
rect 28908 35071 28960 35080
rect 28908 35037 28917 35071
rect 28917 35037 28951 35071
rect 28951 35037 28960 35071
rect 28908 35028 28960 35037
rect 25964 34935 26016 34944
rect 25964 34901 25973 34935
rect 25973 34901 26007 34935
rect 26007 34901 26016 34935
rect 25964 34892 26016 34901
rect 27344 34892 27396 34944
rect 27804 34892 27856 34944
rect 28816 34935 28868 34944
rect 28816 34901 28825 34935
rect 28825 34901 28859 34935
rect 28859 34901 28868 34935
rect 28816 34892 28868 34901
rect 31024 35096 31076 35148
rect 33324 35096 33376 35148
rect 33416 35096 33468 35148
rect 33692 35096 33744 35148
rect 30380 35071 30432 35080
rect 30380 35037 30389 35071
rect 30389 35037 30423 35071
rect 30423 35037 30432 35071
rect 30380 35028 30432 35037
rect 32496 34960 32548 35012
rect 33416 34960 33468 35012
rect 31668 34892 31720 34944
rect 31760 34892 31812 34944
rect 33324 34892 33376 34944
rect 4874 34790 4926 34842
rect 4938 34790 4990 34842
rect 5002 34790 5054 34842
rect 5066 34790 5118 34842
rect 5130 34790 5182 34842
rect 35594 34790 35646 34842
rect 35658 34790 35710 34842
rect 35722 34790 35774 34842
rect 35786 34790 35838 34842
rect 35850 34790 35902 34842
rect 7196 34688 7248 34740
rect 5632 34595 5684 34604
rect 5632 34561 5641 34595
rect 5641 34561 5675 34595
rect 5675 34561 5684 34595
rect 5632 34552 5684 34561
rect 8208 34620 8260 34672
rect 8392 34595 8444 34604
rect 8392 34561 8401 34595
rect 8401 34561 8435 34595
rect 8435 34561 8444 34595
rect 8392 34552 8444 34561
rect 8208 34484 8260 34536
rect 12164 34688 12216 34740
rect 12624 34688 12676 34740
rect 17316 34688 17368 34740
rect 11428 34620 11480 34672
rect 11888 34663 11940 34672
rect 11888 34629 11897 34663
rect 11897 34629 11931 34663
rect 11931 34629 11940 34663
rect 11888 34620 11940 34629
rect 16488 34620 16540 34672
rect 16948 34620 17000 34672
rect 17960 34620 18012 34672
rect 20904 34620 20956 34672
rect 21272 34620 21324 34672
rect 21824 34620 21876 34672
rect 22284 34663 22336 34672
rect 22284 34629 22293 34663
rect 22293 34629 22327 34663
rect 22327 34629 22336 34663
rect 22284 34620 22336 34629
rect 12256 34552 12308 34604
rect 12716 34552 12768 34604
rect 16580 34552 16632 34604
rect 12440 34484 12492 34536
rect 17316 34595 17368 34604
rect 17316 34561 17325 34595
rect 17325 34561 17359 34595
rect 17359 34561 17368 34595
rect 17316 34552 17368 34561
rect 17684 34552 17736 34604
rect 17776 34484 17828 34536
rect 9496 34416 9548 34468
rect 9864 34416 9916 34468
rect 13636 34416 13688 34468
rect 22100 34595 22152 34604
rect 22100 34561 22107 34595
rect 22107 34561 22152 34595
rect 22100 34552 22152 34561
rect 22836 34552 22888 34604
rect 23756 34688 23808 34740
rect 25228 34688 25280 34740
rect 25964 34688 26016 34740
rect 28816 34688 28868 34740
rect 31392 34688 31444 34740
rect 33324 34731 33376 34740
rect 33324 34697 33333 34731
rect 33333 34697 33367 34731
rect 33367 34697 33376 34731
rect 33324 34688 33376 34697
rect 33508 34688 33560 34740
rect 23204 34620 23256 34672
rect 28540 34620 28592 34672
rect 24124 34552 24176 34604
rect 28264 34552 28316 34604
rect 27160 34484 27212 34536
rect 31760 34620 31812 34672
rect 30932 34552 30984 34604
rect 34152 34552 34204 34604
rect 36912 34552 36964 34604
rect 23480 34416 23532 34468
rect 27988 34416 28040 34468
rect 31852 34527 31904 34536
rect 31852 34493 31861 34527
rect 31861 34493 31895 34527
rect 31895 34493 31904 34527
rect 31852 34484 31904 34493
rect 32404 34484 32456 34536
rect 30196 34416 30248 34468
rect 37924 34484 37976 34536
rect 5356 34348 5408 34400
rect 11520 34391 11572 34400
rect 11520 34357 11529 34391
rect 11529 34357 11563 34391
rect 11563 34357 11572 34391
rect 11520 34348 11572 34357
rect 16856 34391 16908 34400
rect 16856 34357 16865 34391
rect 16865 34357 16899 34391
rect 16899 34357 16908 34391
rect 16856 34348 16908 34357
rect 16948 34391 17000 34400
rect 16948 34357 16957 34391
rect 16957 34357 16991 34391
rect 16991 34357 17000 34391
rect 16948 34348 17000 34357
rect 17040 34391 17092 34400
rect 17040 34357 17049 34391
rect 17049 34357 17083 34391
rect 17083 34357 17092 34391
rect 17040 34348 17092 34357
rect 18052 34348 18104 34400
rect 20628 34348 20680 34400
rect 22008 34348 22060 34400
rect 22652 34348 22704 34400
rect 23756 34348 23808 34400
rect 24768 34348 24820 34400
rect 27252 34348 27304 34400
rect 28080 34348 28132 34400
rect 30012 34348 30064 34400
rect 30564 34348 30616 34400
rect 33324 34348 33376 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 6736 34187 6788 34196
rect 6736 34153 6745 34187
rect 6745 34153 6779 34187
rect 6779 34153 6788 34187
rect 6736 34144 6788 34153
rect 12072 34144 12124 34196
rect 14648 34187 14700 34196
rect 14648 34153 14657 34187
rect 14657 34153 14691 34187
rect 14691 34153 14700 34187
rect 14648 34144 14700 34153
rect 14832 34187 14884 34196
rect 14832 34153 14841 34187
rect 14841 34153 14875 34187
rect 14875 34153 14884 34187
rect 14832 34144 14884 34153
rect 16856 34144 16908 34196
rect 16948 34144 17000 34196
rect 17040 34144 17092 34196
rect 20536 34144 20588 34196
rect 22100 34144 22152 34196
rect 22468 34144 22520 34196
rect 23112 34144 23164 34196
rect 15016 34076 15068 34128
rect 5356 34008 5408 34060
rect 6920 34008 6972 34060
rect 4712 33983 4764 33992
rect 4712 33949 4721 33983
rect 4721 33949 4755 33983
rect 4755 33949 4764 33983
rect 4712 33940 4764 33949
rect 6368 33940 6420 33992
rect 6644 33940 6696 33992
rect 8392 34008 8444 34060
rect 7564 33940 7616 33992
rect 9036 33940 9088 33992
rect 9588 33872 9640 33924
rect 11796 34008 11848 34060
rect 13636 34008 13688 34060
rect 9864 33983 9916 33992
rect 9864 33949 9873 33983
rect 9873 33949 9907 33983
rect 9907 33949 9916 33983
rect 9864 33940 9916 33949
rect 11520 33940 11572 33992
rect 14464 33940 14516 33992
rect 7196 33847 7248 33856
rect 7196 33813 7205 33847
rect 7205 33813 7239 33847
rect 7239 33813 7248 33847
rect 7196 33804 7248 33813
rect 8668 33847 8720 33856
rect 8668 33813 8677 33847
rect 8677 33813 8711 33847
rect 8711 33813 8720 33847
rect 8668 33804 8720 33813
rect 8944 33847 8996 33856
rect 8944 33813 8953 33847
rect 8953 33813 8987 33847
rect 8987 33813 8996 33847
rect 8944 33804 8996 33813
rect 9404 33804 9456 33856
rect 11980 33804 12032 33856
rect 13268 33804 13320 33856
rect 13360 33847 13412 33856
rect 13360 33813 13369 33847
rect 13369 33813 13403 33847
rect 13403 33813 13412 33847
rect 13360 33804 13412 33813
rect 13728 33804 13780 33856
rect 15752 33983 15804 33992
rect 15752 33949 15761 33983
rect 15761 33949 15795 33983
rect 15795 33949 15804 33983
rect 15752 33940 15804 33949
rect 16212 33983 16264 33992
rect 16212 33949 16221 33983
rect 16221 33949 16255 33983
rect 16255 33949 16264 33983
rect 16212 33940 16264 33949
rect 16304 33983 16356 33992
rect 16304 33949 16313 33983
rect 16313 33949 16347 33983
rect 16347 33949 16356 33983
rect 16304 33940 16356 33949
rect 16488 33940 16540 33992
rect 17684 33983 17736 33992
rect 17684 33949 17693 33983
rect 17693 33949 17727 33983
rect 17727 33949 17736 33983
rect 17684 33940 17736 33949
rect 17776 33983 17828 33992
rect 17776 33949 17786 33983
rect 17786 33949 17820 33983
rect 17820 33949 17828 33983
rect 17776 33940 17828 33949
rect 18052 33983 18104 33992
rect 18052 33949 18061 33983
rect 18061 33949 18095 33983
rect 18095 33949 18104 33983
rect 18052 33940 18104 33949
rect 18144 33983 18196 33992
rect 18144 33949 18158 33983
rect 18158 33949 18192 33983
rect 18192 33949 18196 33983
rect 18144 33940 18196 33949
rect 18420 33983 18472 33992
rect 18420 33949 18429 33983
rect 18429 33949 18463 33983
rect 18463 33949 18472 33983
rect 18420 33940 18472 33949
rect 15476 33872 15528 33924
rect 16672 33872 16724 33924
rect 17960 33915 18012 33924
rect 17960 33881 17969 33915
rect 17969 33881 18003 33915
rect 18003 33881 18012 33915
rect 17960 33872 18012 33881
rect 14924 33804 14976 33856
rect 16948 33804 17000 33856
rect 17040 33847 17092 33856
rect 17040 33813 17049 33847
rect 17049 33813 17083 33847
rect 17083 33813 17092 33847
rect 17040 33804 17092 33813
rect 17132 33847 17184 33856
rect 17132 33813 17141 33847
rect 17141 33813 17175 33847
rect 17175 33813 17184 33847
rect 17132 33804 17184 33813
rect 17500 33804 17552 33856
rect 18604 33915 18656 33924
rect 18604 33881 18613 33915
rect 18613 33881 18647 33915
rect 18647 33881 18656 33915
rect 18604 33872 18656 33881
rect 18328 33847 18380 33856
rect 18328 33813 18337 33847
rect 18337 33813 18371 33847
rect 18371 33813 18380 33847
rect 18328 33804 18380 33813
rect 18512 33804 18564 33856
rect 18788 33804 18840 33856
rect 20168 34008 20220 34060
rect 23664 34144 23716 34196
rect 24768 34144 24820 34196
rect 25412 34144 25464 34196
rect 20260 33983 20312 33992
rect 20260 33949 20269 33983
rect 20269 33949 20303 33983
rect 20303 33949 20312 33983
rect 20260 33940 20312 33949
rect 20536 33940 20588 33992
rect 20628 33940 20680 33992
rect 20904 33940 20956 33992
rect 21916 33983 21968 33992
rect 21916 33949 21925 33983
rect 21925 33949 21959 33983
rect 21959 33949 21968 33983
rect 21916 33940 21968 33949
rect 22468 33940 22520 33992
rect 22284 33872 22336 33924
rect 22652 33983 22704 33992
rect 22652 33949 22661 33983
rect 22661 33949 22695 33983
rect 22695 33949 22704 33983
rect 22652 33940 22704 33949
rect 22928 33983 22980 33992
rect 22928 33949 22937 33983
rect 22937 33949 22971 33983
rect 22971 33949 22980 33983
rect 22928 33940 22980 33949
rect 23388 33940 23440 33992
rect 23480 33915 23532 33924
rect 23480 33881 23489 33915
rect 23489 33881 23523 33915
rect 23523 33881 23532 33915
rect 23480 33872 23532 33881
rect 23664 33983 23716 33992
rect 23664 33949 23678 33983
rect 23678 33949 23712 33983
rect 23712 33949 23716 33983
rect 23664 33940 23716 33949
rect 23848 33940 23900 33992
rect 25596 33983 25648 33992
rect 25596 33949 25605 33983
rect 25605 33949 25639 33983
rect 25639 33949 25648 33983
rect 25596 33940 25648 33949
rect 20352 33804 20404 33856
rect 20812 33804 20864 33856
rect 22928 33804 22980 33856
rect 23388 33804 23440 33856
rect 23848 33847 23900 33856
rect 23848 33813 23857 33847
rect 23857 33813 23891 33847
rect 23891 33813 23900 33847
rect 23848 33804 23900 33813
rect 24584 33804 24636 33856
rect 25412 33847 25464 33856
rect 25412 33813 25421 33847
rect 25421 33813 25455 33847
rect 25455 33813 25464 33847
rect 25412 33804 25464 33813
rect 25964 33983 26016 33992
rect 25964 33949 25973 33983
rect 25973 33949 26007 33983
rect 26007 33949 26016 33983
rect 25964 33940 26016 33949
rect 26240 33983 26292 33992
rect 26240 33949 26249 33983
rect 26249 33949 26283 33983
rect 26283 33949 26292 33983
rect 26240 33940 26292 33949
rect 26792 34144 26844 34196
rect 28080 34187 28132 34196
rect 28080 34153 28089 34187
rect 28089 34153 28123 34187
rect 28123 34153 28132 34187
rect 28080 34144 28132 34153
rect 26148 33872 26200 33924
rect 26976 33940 27028 33992
rect 28816 34076 28868 34128
rect 30932 34076 30984 34128
rect 28632 34008 28684 34060
rect 30748 34008 30800 34060
rect 26516 33872 26568 33924
rect 30012 33940 30064 33992
rect 30472 33983 30524 33992
rect 30472 33949 30481 33983
rect 30481 33949 30515 33983
rect 30515 33949 30524 33983
rect 30472 33940 30524 33949
rect 30564 33983 30616 33992
rect 30564 33949 30601 33983
rect 30601 33949 30616 33983
rect 30564 33940 30616 33949
rect 29828 33872 29880 33924
rect 31484 33983 31536 33992
rect 31484 33949 31493 33983
rect 31493 33949 31527 33983
rect 31527 33949 31536 33983
rect 31484 33940 31536 33949
rect 33416 33940 33468 33992
rect 33876 33983 33928 33992
rect 33876 33949 33885 33983
rect 33885 33949 33919 33983
rect 33919 33949 33928 33983
rect 33876 33940 33928 33949
rect 27160 33847 27212 33856
rect 27160 33813 27169 33847
rect 27169 33813 27203 33847
rect 27203 33813 27212 33847
rect 27160 33804 27212 33813
rect 28816 33847 28868 33856
rect 28816 33813 28825 33847
rect 28825 33813 28859 33847
rect 28859 33813 28868 33847
rect 28816 33804 28868 33813
rect 35992 33872 36044 33924
rect 36636 33872 36688 33924
rect 31576 33847 31628 33856
rect 31576 33813 31585 33847
rect 31585 33813 31619 33847
rect 31619 33813 31628 33847
rect 31576 33804 31628 33813
rect 32220 33804 32272 33856
rect 34336 33804 34388 33856
rect 4874 33702 4926 33754
rect 4938 33702 4990 33754
rect 5002 33702 5054 33754
rect 5066 33702 5118 33754
rect 5130 33702 5182 33754
rect 35594 33702 35646 33754
rect 35658 33702 35710 33754
rect 35722 33702 35774 33754
rect 35786 33702 35838 33754
rect 35850 33702 35902 33754
rect 5632 33600 5684 33652
rect 6736 33600 6788 33652
rect 7196 33600 7248 33652
rect 8668 33600 8720 33652
rect 8300 33532 8352 33584
rect 9404 33600 9456 33652
rect 13176 33600 13228 33652
rect 14648 33600 14700 33652
rect 16488 33600 16540 33652
rect 10232 33532 10284 33584
rect 13360 33532 13412 33584
rect 11980 33464 12032 33516
rect 16580 33532 16632 33584
rect 16856 33600 16908 33652
rect 17040 33600 17092 33652
rect 17684 33600 17736 33652
rect 19340 33600 19392 33652
rect 18420 33532 18472 33584
rect 14372 33507 14424 33516
rect 14372 33473 14381 33507
rect 14381 33473 14415 33507
rect 14415 33473 14424 33507
rect 14372 33464 14424 33473
rect 14740 33464 14792 33516
rect 18604 33464 18656 33516
rect 19708 33507 19760 33516
rect 19708 33473 19742 33507
rect 19742 33473 19760 33507
rect 19708 33464 19760 33473
rect 20260 33600 20312 33652
rect 21272 33643 21324 33652
rect 21272 33609 21281 33643
rect 21281 33609 21315 33643
rect 21315 33609 21324 33643
rect 21272 33600 21324 33609
rect 21916 33600 21968 33652
rect 22100 33600 22152 33652
rect 26148 33600 26200 33652
rect 31576 33600 31628 33652
rect 21364 33532 21416 33584
rect 21548 33532 21600 33584
rect 23204 33532 23256 33584
rect 20352 33507 20404 33516
rect 20352 33473 20361 33507
rect 20361 33473 20395 33507
rect 20395 33473 20404 33507
rect 20352 33464 20404 33473
rect 5908 33439 5960 33448
rect 5908 33405 5917 33439
rect 5917 33405 5951 33439
rect 5951 33405 5960 33439
rect 5908 33396 5960 33405
rect 7288 33439 7340 33448
rect 7288 33405 7297 33439
rect 7297 33405 7331 33439
rect 7331 33405 7340 33439
rect 7288 33396 7340 33405
rect 9588 33396 9640 33448
rect 18420 33396 18472 33448
rect 19064 33439 19116 33448
rect 19064 33405 19073 33439
rect 19073 33405 19107 33439
rect 19107 33405 19116 33439
rect 19064 33396 19116 33405
rect 19340 33396 19392 33448
rect 19616 33396 19668 33448
rect 20720 33507 20772 33516
rect 20720 33473 20729 33507
rect 20729 33473 20763 33507
rect 20763 33473 20772 33507
rect 20720 33464 20772 33473
rect 21824 33507 21876 33516
rect 21824 33473 21833 33507
rect 21833 33473 21867 33507
rect 21867 33473 21876 33507
rect 21824 33464 21876 33473
rect 17040 33328 17092 33380
rect 17960 33328 18012 33380
rect 19524 33328 19576 33380
rect 19892 33328 19944 33380
rect 20628 33328 20680 33380
rect 23480 33439 23532 33448
rect 23480 33405 23489 33439
rect 23489 33405 23523 33439
rect 23523 33405 23532 33439
rect 23480 33396 23532 33405
rect 23572 33439 23624 33448
rect 23572 33405 23581 33439
rect 23581 33405 23615 33439
rect 23615 33405 23624 33439
rect 23572 33396 23624 33405
rect 23756 33507 23808 33516
rect 23756 33473 23765 33507
rect 23765 33473 23799 33507
rect 23799 33473 23808 33507
rect 23756 33464 23808 33473
rect 23848 33507 23900 33516
rect 23848 33473 23857 33507
rect 23857 33473 23891 33507
rect 23891 33473 23900 33507
rect 23848 33464 23900 33473
rect 25320 33532 25372 33584
rect 25504 33532 25556 33584
rect 26516 33464 26568 33516
rect 26608 33507 26660 33516
rect 26608 33473 26617 33507
rect 26617 33473 26651 33507
rect 26651 33473 26660 33507
rect 26608 33464 26660 33473
rect 27160 33532 27212 33584
rect 28540 33532 28592 33584
rect 29000 33532 29052 33584
rect 20904 33328 20956 33380
rect 7012 33260 7064 33312
rect 7840 33260 7892 33312
rect 11612 33260 11664 33312
rect 16212 33260 16264 33312
rect 18144 33260 18196 33312
rect 20352 33260 20404 33312
rect 20444 33260 20496 33312
rect 21456 33260 21508 33312
rect 22928 33260 22980 33312
rect 23756 33260 23808 33312
rect 24032 33303 24084 33312
rect 24032 33269 24041 33303
rect 24041 33269 24075 33303
rect 24075 33269 24084 33303
rect 24032 33260 24084 33269
rect 25320 33328 25372 33380
rect 25412 33303 25464 33312
rect 25412 33269 25421 33303
rect 25421 33269 25455 33303
rect 25455 33269 25464 33303
rect 25412 33260 25464 33269
rect 27804 33396 27856 33448
rect 33232 33600 33284 33652
rect 33600 33600 33652 33652
rect 33876 33600 33928 33652
rect 34152 33643 34204 33652
rect 34152 33609 34161 33643
rect 34161 33609 34195 33643
rect 34195 33609 34204 33643
rect 34152 33600 34204 33609
rect 32312 33464 32364 33516
rect 36912 33643 36964 33652
rect 36912 33609 36921 33643
rect 36921 33609 36955 33643
rect 36955 33609 36964 33643
rect 36912 33600 36964 33609
rect 34060 33439 34112 33448
rect 34060 33405 34069 33439
rect 34069 33405 34103 33439
rect 34103 33405 34112 33439
rect 34060 33396 34112 33405
rect 36636 33464 36688 33516
rect 36728 33507 36780 33516
rect 36728 33473 36737 33507
rect 36737 33473 36771 33507
rect 36771 33473 36780 33507
rect 36728 33464 36780 33473
rect 28540 33260 28592 33312
rect 28724 33260 28776 33312
rect 30196 33260 30248 33312
rect 35992 33328 36044 33380
rect 34796 33260 34848 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 7288 33056 7340 33108
rect 4620 32920 4672 32972
rect 6736 32963 6788 32972
rect 6736 32929 6745 32963
rect 6745 32929 6779 32963
rect 6779 32929 6788 32963
rect 6736 32920 6788 32929
rect 6828 32963 6880 32972
rect 6828 32929 6837 32963
rect 6837 32929 6871 32963
rect 6871 32929 6880 32963
rect 6828 32920 6880 32929
rect 5908 32852 5960 32904
rect 6644 32895 6696 32904
rect 6644 32861 6653 32895
rect 6653 32861 6687 32895
rect 6687 32861 6696 32895
rect 6644 32852 6696 32861
rect 8944 33056 8996 33108
rect 9864 33056 9916 33108
rect 11612 33056 11664 33108
rect 9680 32920 9732 32972
rect 11704 32988 11756 33040
rect 12164 32988 12216 33040
rect 4712 32784 4764 32836
rect 6368 32784 6420 32836
rect 8208 32895 8260 32904
rect 8208 32861 8217 32895
rect 8217 32861 8251 32895
rect 8251 32861 8260 32895
rect 8208 32852 8260 32861
rect 8484 32895 8536 32904
rect 8484 32861 8493 32895
rect 8493 32861 8527 32895
rect 8527 32861 8536 32895
rect 8484 32852 8536 32861
rect 11428 32852 11480 32904
rect 11888 32852 11940 32904
rect 8392 32784 8444 32836
rect 8576 32784 8628 32836
rect 10968 32784 11020 32836
rect 12072 32827 12124 32836
rect 12072 32793 12081 32827
rect 12081 32793 12115 32827
rect 12115 32793 12124 32827
rect 12072 32784 12124 32793
rect 6276 32759 6328 32768
rect 6276 32725 6285 32759
rect 6285 32725 6319 32759
rect 6319 32725 6328 32759
rect 6276 32716 6328 32725
rect 8852 32716 8904 32768
rect 11612 32716 11664 32768
rect 12256 32716 12308 32768
rect 12348 32759 12400 32768
rect 12348 32725 12357 32759
rect 12357 32725 12391 32759
rect 12391 32725 12400 32759
rect 12348 32716 12400 32725
rect 17408 33056 17460 33108
rect 16764 32988 16816 33040
rect 17684 32988 17736 33040
rect 18144 32988 18196 33040
rect 18328 33056 18380 33108
rect 20352 33056 20404 33108
rect 15844 32852 15896 32904
rect 16212 32895 16264 32904
rect 16212 32861 16221 32895
rect 16221 32861 16255 32895
rect 16255 32861 16264 32895
rect 16212 32852 16264 32861
rect 17960 32852 18012 32904
rect 18604 32920 18656 32972
rect 19340 32920 19392 32972
rect 18420 32895 18472 32904
rect 18420 32861 18429 32895
rect 18429 32861 18463 32895
rect 18463 32861 18472 32895
rect 18420 32852 18472 32861
rect 18880 32852 18932 32904
rect 19708 33031 19760 33040
rect 19708 32997 19717 33031
rect 19717 32997 19751 33031
rect 19751 32997 19760 33031
rect 19708 32988 19760 32997
rect 20536 32988 20588 33040
rect 19616 32963 19668 32972
rect 19616 32929 19625 32963
rect 19625 32929 19659 32963
rect 19659 32929 19668 32963
rect 19616 32920 19668 32929
rect 20904 33056 20956 33108
rect 23480 33056 23532 33108
rect 26608 33099 26660 33108
rect 26608 33065 26617 33099
rect 26617 33065 26651 33099
rect 26651 33065 26660 33099
rect 26608 33056 26660 33065
rect 30012 33056 30064 33108
rect 30472 33056 30524 33108
rect 31852 33056 31904 33108
rect 34796 33056 34848 33108
rect 20720 33031 20772 33040
rect 20720 32997 20729 33031
rect 20729 32997 20763 33031
rect 20763 32997 20772 33031
rect 20720 32988 20772 32997
rect 30656 32988 30708 33040
rect 19984 32852 20036 32904
rect 20168 32895 20220 32904
rect 20168 32861 20177 32895
rect 20177 32861 20211 32895
rect 20211 32861 20220 32895
rect 20168 32852 20220 32861
rect 24584 32920 24636 32972
rect 26056 32920 26108 32972
rect 27252 32963 27304 32972
rect 27252 32929 27261 32963
rect 27261 32929 27295 32963
rect 27295 32929 27304 32963
rect 27252 32920 27304 32929
rect 21456 32895 21508 32904
rect 21456 32861 21465 32895
rect 21465 32861 21499 32895
rect 21499 32861 21508 32895
rect 21456 32852 21508 32861
rect 21916 32852 21968 32904
rect 22192 32852 22244 32904
rect 23388 32895 23440 32904
rect 23388 32861 23397 32895
rect 23397 32861 23431 32895
rect 23431 32861 23440 32895
rect 23388 32852 23440 32861
rect 24492 32852 24544 32904
rect 27804 32920 27856 32972
rect 16856 32784 16908 32836
rect 17592 32784 17644 32836
rect 18788 32827 18840 32836
rect 18788 32793 18797 32827
rect 18797 32793 18831 32827
rect 18831 32793 18840 32827
rect 18788 32784 18840 32793
rect 19340 32784 19392 32836
rect 19524 32784 19576 32836
rect 19984 32716 20036 32768
rect 21548 32784 21600 32836
rect 22008 32716 22060 32768
rect 23572 32759 23624 32768
rect 23572 32725 23581 32759
rect 23581 32725 23615 32759
rect 23615 32725 23624 32759
rect 23572 32716 23624 32725
rect 23756 32716 23808 32768
rect 25044 32716 25096 32768
rect 25964 32716 26016 32768
rect 26332 32716 26384 32768
rect 26700 32716 26752 32768
rect 27528 32895 27580 32904
rect 27528 32861 27537 32895
rect 27537 32861 27571 32895
rect 27571 32861 27580 32895
rect 27528 32852 27580 32861
rect 28080 32784 28132 32836
rect 28540 32784 28592 32836
rect 30932 32895 30984 32904
rect 30932 32861 30941 32895
rect 30941 32861 30975 32895
rect 30975 32861 30984 32895
rect 30932 32852 30984 32861
rect 31208 32895 31260 32904
rect 31208 32861 31217 32895
rect 31217 32861 31251 32895
rect 31251 32861 31260 32895
rect 31208 32852 31260 32861
rect 32496 32852 32548 32904
rect 32956 32852 33008 32904
rect 34336 32895 34388 32904
rect 34336 32861 34345 32895
rect 34345 32861 34379 32895
rect 34379 32861 34388 32895
rect 34336 32852 34388 32861
rect 35992 32852 36044 32904
rect 27344 32716 27396 32768
rect 28724 32716 28776 32768
rect 30196 32759 30248 32768
rect 30196 32725 30205 32759
rect 30205 32725 30239 32759
rect 30239 32725 30248 32759
rect 30196 32716 30248 32725
rect 30288 32716 30340 32768
rect 31852 32716 31904 32768
rect 36268 32716 36320 32768
rect 4874 32614 4926 32666
rect 4938 32614 4990 32666
rect 5002 32614 5054 32666
rect 5066 32614 5118 32666
rect 5130 32614 5182 32666
rect 35594 32614 35646 32666
rect 35658 32614 35710 32666
rect 35722 32614 35774 32666
rect 35786 32614 35838 32666
rect 35850 32614 35902 32666
rect 4712 32512 4764 32564
rect 6276 32512 6328 32564
rect 6736 32512 6788 32564
rect 11612 32512 11664 32564
rect 11796 32512 11848 32564
rect 12348 32512 12400 32564
rect 11612 32376 11664 32428
rect 16764 32444 16816 32496
rect 17868 32512 17920 32564
rect 18696 32512 18748 32564
rect 18880 32512 18932 32564
rect 19984 32555 20036 32564
rect 19984 32521 19993 32555
rect 19993 32521 20027 32555
rect 20027 32521 20036 32555
rect 19984 32512 20036 32521
rect 15476 32376 15528 32428
rect 15752 32376 15804 32428
rect 17592 32444 17644 32496
rect 17960 32444 18012 32496
rect 22284 32512 22336 32564
rect 18420 32419 18472 32428
rect 18420 32385 18429 32419
rect 18429 32385 18463 32419
rect 18463 32385 18472 32419
rect 18420 32376 18472 32385
rect 21088 32444 21140 32496
rect 18880 32419 18932 32428
rect 18880 32385 18889 32419
rect 18889 32385 18923 32419
rect 18923 32385 18932 32419
rect 18880 32376 18932 32385
rect 5724 32240 5776 32292
rect 8300 32240 8352 32292
rect 12624 32283 12676 32292
rect 12624 32249 12633 32283
rect 12633 32249 12667 32283
rect 12667 32249 12676 32283
rect 12624 32240 12676 32249
rect 16120 32240 16172 32292
rect 17132 32240 17184 32292
rect 18236 32308 18288 32360
rect 20444 32376 20496 32428
rect 21640 32444 21692 32496
rect 23388 32512 23440 32564
rect 23572 32512 23624 32564
rect 21364 32376 21416 32428
rect 23204 32487 23256 32496
rect 23204 32453 23213 32487
rect 23213 32453 23247 32487
rect 23247 32453 23256 32487
rect 23204 32444 23256 32453
rect 27528 32512 27580 32564
rect 28080 32512 28132 32564
rect 31208 32512 31260 32564
rect 36728 32512 36780 32564
rect 22744 32376 22796 32428
rect 22928 32376 22980 32428
rect 23020 32419 23072 32428
rect 23020 32385 23029 32419
rect 23029 32385 23063 32419
rect 23063 32385 23072 32419
rect 23020 32376 23072 32385
rect 22284 32308 22336 32360
rect 6552 32172 6604 32224
rect 11612 32172 11664 32224
rect 16672 32172 16724 32224
rect 16948 32172 17000 32224
rect 19064 32240 19116 32292
rect 23204 32240 23256 32292
rect 23756 32419 23808 32428
rect 23756 32385 23765 32419
rect 23765 32385 23799 32419
rect 23799 32385 23808 32419
rect 23756 32376 23808 32385
rect 27712 32444 27764 32496
rect 24124 32419 24176 32428
rect 24124 32385 24133 32419
rect 24133 32385 24167 32419
rect 24167 32385 24176 32419
rect 24124 32376 24176 32385
rect 24400 32308 24452 32360
rect 26516 32308 26568 32360
rect 28724 32376 28776 32428
rect 27896 32240 27948 32292
rect 28448 32351 28500 32360
rect 28448 32317 28457 32351
rect 28457 32317 28491 32351
rect 28491 32317 28500 32351
rect 28448 32308 28500 32317
rect 30840 32419 30892 32428
rect 30840 32385 30849 32419
rect 30849 32385 30883 32419
rect 30883 32385 30892 32419
rect 30840 32376 30892 32385
rect 30932 32376 30984 32428
rect 32588 32444 32640 32496
rect 34612 32444 34664 32496
rect 32128 32376 32180 32428
rect 32220 32376 32272 32428
rect 33140 32419 33192 32428
rect 33140 32385 33149 32419
rect 33149 32385 33183 32419
rect 33183 32385 33192 32419
rect 33140 32376 33192 32385
rect 33232 32376 33284 32428
rect 36268 32444 36320 32496
rect 30656 32351 30708 32360
rect 30656 32317 30665 32351
rect 30665 32317 30699 32351
rect 30699 32317 30708 32351
rect 30656 32308 30708 32317
rect 20168 32172 20220 32224
rect 20904 32172 20956 32224
rect 22192 32215 22244 32224
rect 22192 32181 22201 32215
rect 22201 32181 22235 32215
rect 22235 32181 22244 32215
rect 22192 32172 22244 32181
rect 22836 32215 22888 32224
rect 22836 32181 22845 32215
rect 22845 32181 22879 32215
rect 22879 32181 22888 32215
rect 22836 32172 22888 32181
rect 24308 32215 24360 32224
rect 24308 32181 24317 32215
rect 24317 32181 24351 32215
rect 24351 32181 24360 32215
rect 24308 32172 24360 32181
rect 24952 32172 25004 32224
rect 26240 32172 26292 32224
rect 31852 32240 31904 32292
rect 32128 32283 32180 32292
rect 32128 32249 32137 32283
rect 32137 32249 32171 32283
rect 32171 32249 32180 32283
rect 32128 32240 32180 32249
rect 32312 32308 32364 32360
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 4620 31968 4672 32020
rect 7196 31968 7248 32020
rect 17408 31968 17460 32020
rect 7472 31900 7524 31952
rect 8484 31900 8536 31952
rect 18696 31943 18748 31952
rect 18696 31909 18705 31943
rect 18705 31909 18739 31943
rect 18739 31909 18748 31943
rect 18696 31900 18748 31909
rect 19064 32011 19116 32020
rect 19064 31977 19073 32011
rect 19073 31977 19107 32011
rect 19107 31977 19116 32011
rect 19064 31968 19116 31977
rect 20812 31968 20864 32020
rect 22008 31968 22060 32020
rect 20260 31900 20312 31952
rect 20628 31900 20680 31952
rect 22284 31900 22336 31952
rect 22744 31900 22796 31952
rect 23020 31900 23072 31952
rect 23940 31900 23992 31952
rect 24308 31968 24360 32020
rect 24400 31900 24452 31952
rect 26976 31968 27028 32020
rect 30288 31968 30340 32020
rect 31852 31968 31904 32020
rect 5816 31764 5868 31816
rect 6552 31807 6604 31816
rect 6552 31773 6561 31807
rect 6561 31773 6595 31807
rect 6595 31773 6604 31807
rect 6552 31764 6604 31773
rect 6644 31764 6696 31816
rect 7472 31807 7524 31816
rect 7472 31773 7481 31807
rect 7481 31773 7515 31807
rect 7515 31773 7524 31807
rect 7472 31764 7524 31773
rect 7656 31807 7708 31816
rect 7656 31773 7665 31807
rect 7665 31773 7699 31807
rect 7699 31773 7708 31807
rect 7656 31764 7708 31773
rect 11612 31832 11664 31884
rect 8116 31807 8168 31816
rect 8116 31773 8125 31807
rect 8125 31773 8159 31807
rect 8159 31773 8168 31807
rect 8116 31764 8168 31773
rect 8484 31807 8536 31816
rect 8484 31773 8493 31807
rect 8493 31773 8527 31807
rect 8527 31773 8536 31807
rect 8484 31764 8536 31773
rect 8852 31764 8904 31816
rect 9036 31764 9088 31816
rect 9772 31739 9824 31748
rect 9772 31705 9781 31739
rect 9781 31705 9815 31739
rect 9815 31705 9824 31739
rect 9772 31696 9824 31705
rect 10232 31696 10284 31748
rect 11796 31696 11848 31748
rect 13176 31696 13228 31748
rect 13636 31807 13688 31816
rect 13636 31773 13645 31807
rect 13645 31773 13679 31807
rect 13679 31773 13688 31807
rect 13636 31764 13688 31773
rect 17592 31764 17644 31816
rect 18788 31764 18840 31816
rect 18880 31807 18932 31816
rect 18880 31773 18889 31807
rect 18889 31773 18923 31807
rect 18923 31773 18932 31807
rect 18880 31764 18932 31773
rect 21732 31764 21784 31816
rect 21916 31807 21968 31816
rect 21916 31773 21925 31807
rect 21925 31773 21959 31807
rect 21959 31773 21968 31807
rect 21916 31764 21968 31773
rect 22008 31807 22060 31816
rect 22008 31773 22018 31807
rect 22018 31773 22052 31807
rect 22052 31773 22060 31807
rect 22008 31764 22060 31773
rect 22100 31764 22152 31816
rect 22284 31807 22336 31816
rect 22284 31773 22293 31807
rect 22293 31773 22327 31807
rect 22327 31773 22336 31807
rect 22284 31764 22336 31773
rect 22376 31807 22428 31816
rect 22376 31773 22390 31807
rect 22390 31773 22424 31807
rect 22424 31773 22428 31807
rect 22376 31764 22428 31773
rect 14556 31696 14608 31748
rect 16488 31696 16540 31748
rect 18144 31696 18196 31748
rect 19156 31696 19208 31748
rect 21824 31696 21876 31748
rect 22652 31807 22704 31816
rect 22652 31773 22661 31807
rect 22661 31773 22695 31807
rect 22695 31773 22704 31807
rect 22652 31764 22704 31773
rect 23204 31764 23256 31816
rect 23388 31807 23440 31816
rect 23388 31773 23397 31807
rect 23397 31773 23431 31807
rect 23431 31773 23440 31807
rect 23388 31764 23440 31773
rect 23572 31832 23624 31884
rect 24216 31764 24268 31816
rect 25412 31900 25464 31952
rect 28724 31900 28776 31952
rect 24492 31764 24544 31816
rect 7840 31628 7892 31680
rect 8300 31671 8352 31680
rect 8300 31637 8309 31671
rect 8309 31637 8343 31671
rect 8343 31637 8352 31671
rect 8300 31628 8352 31637
rect 11520 31628 11572 31680
rect 12992 31628 13044 31680
rect 13912 31628 13964 31680
rect 14372 31628 14424 31680
rect 16948 31628 17000 31680
rect 19616 31628 19668 31680
rect 19892 31628 19944 31680
rect 20444 31628 20496 31680
rect 21364 31628 21416 31680
rect 22008 31628 22060 31680
rect 22560 31671 22612 31680
rect 22560 31637 22569 31671
rect 22569 31637 22603 31671
rect 22603 31637 22612 31671
rect 22560 31628 22612 31637
rect 22652 31628 22704 31680
rect 23664 31739 23716 31748
rect 23664 31705 23673 31739
rect 23673 31705 23707 31739
rect 23707 31705 23716 31739
rect 23664 31696 23716 31705
rect 23756 31739 23808 31748
rect 23756 31705 23765 31739
rect 23765 31705 23799 31739
rect 23799 31705 23808 31739
rect 23756 31696 23808 31705
rect 24768 31807 24820 31816
rect 24768 31773 24777 31807
rect 24777 31773 24811 31807
rect 24811 31773 24820 31807
rect 24768 31764 24820 31773
rect 24952 31764 25004 31816
rect 25136 31807 25188 31816
rect 25136 31773 25145 31807
rect 25145 31773 25179 31807
rect 25179 31773 25188 31807
rect 25136 31764 25188 31773
rect 23204 31628 23256 31680
rect 25320 31764 25372 31816
rect 26148 31807 26200 31816
rect 26148 31773 26157 31807
rect 26157 31773 26191 31807
rect 26191 31773 26200 31807
rect 26148 31764 26200 31773
rect 26240 31807 26292 31816
rect 26240 31773 26249 31807
rect 26249 31773 26283 31807
rect 26283 31773 26292 31807
rect 26240 31764 26292 31773
rect 26516 31807 26568 31816
rect 26516 31773 26525 31807
rect 26525 31773 26559 31807
rect 26559 31773 26568 31807
rect 26516 31764 26568 31773
rect 26976 31807 27028 31816
rect 26976 31773 26985 31807
rect 26985 31773 27019 31807
rect 27019 31773 27028 31807
rect 26976 31764 27028 31773
rect 28908 31832 28960 31884
rect 28264 31807 28316 31816
rect 28264 31773 28273 31807
rect 28273 31773 28307 31807
rect 28307 31773 28316 31807
rect 28264 31764 28316 31773
rect 29460 31764 29512 31816
rect 25596 31671 25648 31680
rect 25596 31637 25605 31671
rect 25605 31637 25639 31671
rect 25639 31637 25648 31671
rect 25596 31628 25648 31637
rect 26148 31628 26200 31680
rect 26240 31628 26292 31680
rect 26792 31696 26844 31748
rect 27712 31628 27764 31680
rect 27988 31628 28040 31680
rect 29092 31628 29144 31680
rect 29828 31807 29880 31816
rect 29828 31773 29837 31807
rect 29837 31773 29871 31807
rect 29871 31773 29880 31807
rect 29828 31764 29880 31773
rect 30288 31832 30340 31884
rect 30748 31764 30800 31816
rect 31484 31807 31536 31816
rect 31484 31773 31493 31807
rect 31493 31773 31527 31807
rect 31527 31773 31536 31807
rect 31484 31764 31536 31773
rect 30012 31628 30064 31680
rect 31944 31807 31996 31816
rect 31944 31773 31953 31807
rect 31953 31773 31987 31807
rect 31987 31773 31996 31807
rect 31944 31764 31996 31773
rect 34612 31764 34664 31816
rect 35440 31807 35492 31816
rect 35440 31773 35449 31807
rect 35449 31773 35483 31807
rect 35483 31773 35492 31807
rect 35440 31764 35492 31773
rect 34520 31696 34572 31748
rect 30380 31671 30432 31680
rect 30380 31637 30389 31671
rect 30389 31637 30423 31671
rect 30423 31637 30432 31671
rect 30380 31628 30432 31637
rect 34796 31671 34848 31680
rect 34796 31637 34805 31671
rect 34805 31637 34839 31671
rect 34839 31637 34848 31671
rect 34796 31628 34848 31637
rect 35256 31671 35308 31680
rect 35256 31637 35265 31671
rect 35265 31637 35299 31671
rect 35299 31637 35308 31671
rect 35256 31628 35308 31637
rect 4874 31526 4926 31578
rect 4938 31526 4990 31578
rect 5002 31526 5054 31578
rect 5066 31526 5118 31578
rect 5130 31526 5182 31578
rect 35594 31526 35646 31578
rect 35658 31526 35710 31578
rect 35722 31526 35774 31578
rect 35786 31526 35838 31578
rect 35850 31526 35902 31578
rect 8300 31424 8352 31476
rect 9772 31424 9824 31476
rect 8576 31356 8628 31408
rect 10876 31424 10928 31476
rect 11612 31424 11664 31476
rect 11980 31424 12032 31476
rect 12992 31424 13044 31476
rect 13360 31424 13412 31476
rect 13452 31467 13504 31476
rect 13452 31433 13461 31467
rect 13461 31433 13495 31467
rect 13495 31433 13504 31467
rect 13452 31424 13504 31433
rect 11796 31399 11848 31408
rect 7840 31263 7892 31272
rect 7840 31229 7849 31263
rect 7849 31229 7883 31263
rect 7883 31229 7892 31263
rect 7840 31220 7892 31229
rect 9404 31220 9456 31272
rect 11796 31365 11805 31399
rect 11805 31365 11839 31399
rect 11839 31365 11848 31399
rect 11796 31356 11848 31365
rect 11520 31331 11572 31340
rect 11520 31297 11529 31331
rect 11529 31297 11563 31331
rect 11563 31297 11572 31331
rect 11520 31288 11572 31297
rect 11612 31288 11664 31340
rect 11888 31331 11940 31340
rect 11888 31297 11897 31331
rect 11897 31297 11931 31331
rect 11931 31297 11940 31331
rect 11888 31288 11940 31297
rect 12348 31288 12400 31340
rect 16212 31424 16264 31476
rect 10784 31263 10836 31272
rect 10784 31229 10793 31263
rect 10793 31229 10827 31263
rect 10827 31229 10836 31263
rect 10784 31220 10836 31229
rect 15476 31331 15528 31340
rect 15476 31297 15485 31331
rect 15485 31297 15519 31331
rect 15519 31297 15528 31331
rect 15476 31288 15528 31297
rect 15752 31288 15804 31340
rect 16028 31288 16080 31340
rect 16120 31331 16172 31340
rect 16120 31297 16129 31331
rect 16129 31297 16163 31331
rect 16163 31297 16172 31331
rect 16120 31288 16172 31297
rect 16212 31331 16264 31340
rect 16212 31297 16221 31331
rect 16221 31297 16255 31331
rect 16255 31297 16264 31331
rect 16212 31288 16264 31297
rect 16488 31288 16540 31340
rect 13360 31220 13412 31272
rect 9680 31152 9732 31204
rect 16948 31399 17000 31408
rect 16948 31365 16957 31399
rect 16957 31365 16991 31399
rect 16991 31365 17000 31399
rect 16948 31356 17000 31365
rect 17684 31424 17736 31476
rect 18696 31467 18748 31476
rect 18696 31433 18705 31467
rect 18705 31433 18739 31467
rect 18739 31433 18748 31467
rect 18696 31424 18748 31433
rect 18788 31424 18840 31476
rect 19432 31424 19484 31476
rect 19800 31424 19852 31476
rect 20352 31424 20404 31476
rect 20812 31424 20864 31476
rect 19984 31356 20036 31408
rect 17408 31331 17460 31340
rect 17408 31297 17417 31331
rect 17417 31297 17451 31331
rect 17451 31297 17460 31331
rect 17408 31288 17460 31297
rect 17592 31331 17644 31340
rect 17592 31297 17601 31331
rect 17601 31297 17635 31331
rect 17635 31297 17644 31331
rect 17592 31288 17644 31297
rect 17868 31288 17920 31340
rect 18420 31288 18472 31340
rect 18144 31152 18196 31204
rect 18788 31331 18840 31340
rect 18788 31297 18797 31331
rect 18797 31297 18831 31331
rect 18831 31297 18840 31331
rect 18788 31288 18840 31297
rect 19248 31288 19300 31340
rect 19616 31288 19668 31340
rect 20628 31331 20680 31340
rect 20628 31297 20637 31331
rect 20637 31297 20671 31331
rect 20671 31297 20680 31331
rect 20628 31288 20680 31297
rect 20720 31288 20772 31340
rect 21456 31424 21508 31476
rect 22192 31467 22244 31476
rect 22192 31433 22201 31467
rect 22201 31433 22235 31467
rect 22235 31433 22244 31467
rect 22192 31424 22244 31433
rect 23296 31424 23348 31476
rect 21180 31331 21232 31340
rect 21180 31297 21189 31331
rect 21189 31297 21223 31331
rect 21223 31297 21232 31331
rect 21180 31288 21232 31297
rect 20352 31220 20404 31272
rect 21548 31288 21600 31340
rect 22284 31356 22336 31408
rect 25504 31356 25556 31408
rect 27620 31356 27672 31408
rect 21364 31263 21416 31272
rect 21364 31229 21373 31263
rect 21373 31229 21407 31263
rect 21407 31229 21416 31263
rect 21364 31220 21416 31229
rect 21732 31220 21784 31272
rect 22652 31288 22704 31340
rect 22836 31331 22888 31340
rect 22836 31297 22845 31331
rect 22845 31297 22879 31331
rect 22879 31297 22888 31331
rect 22836 31288 22888 31297
rect 23204 31288 23256 31340
rect 23296 31331 23348 31340
rect 23296 31297 23305 31331
rect 23305 31297 23339 31331
rect 23339 31297 23348 31331
rect 23296 31288 23348 31297
rect 25412 31331 25464 31340
rect 25412 31297 25421 31331
rect 25421 31297 25455 31331
rect 25455 31297 25464 31331
rect 25412 31288 25464 31297
rect 25596 31331 25648 31340
rect 25596 31297 25605 31331
rect 25605 31297 25639 31331
rect 25639 31297 25648 31331
rect 25596 31288 25648 31297
rect 20904 31152 20956 31204
rect 22560 31220 22612 31272
rect 23388 31220 23440 31272
rect 24584 31220 24636 31272
rect 26332 31331 26384 31340
rect 26332 31297 26341 31331
rect 26341 31297 26375 31331
rect 26375 31297 26384 31331
rect 26332 31288 26384 31297
rect 27160 31331 27212 31340
rect 27160 31297 27169 31331
rect 27169 31297 27203 31331
rect 27203 31297 27212 31331
rect 27160 31288 27212 31297
rect 13544 31084 13596 31136
rect 14648 31084 14700 31136
rect 16488 31127 16540 31136
rect 16488 31093 16497 31127
rect 16497 31093 16531 31127
rect 16531 31093 16540 31127
rect 16488 31084 16540 31093
rect 16764 31084 16816 31136
rect 18052 31084 18104 31136
rect 18328 31127 18380 31136
rect 18328 31093 18337 31127
rect 18337 31093 18371 31127
rect 18371 31093 18380 31127
rect 18328 31084 18380 31093
rect 18788 31084 18840 31136
rect 22652 31127 22704 31136
rect 22652 31093 22661 31127
rect 22661 31093 22695 31127
rect 22695 31093 22704 31127
rect 22652 31084 22704 31093
rect 25412 31084 25464 31136
rect 25964 31084 26016 31136
rect 26516 31220 26568 31272
rect 26700 31195 26752 31204
rect 26700 31161 26709 31195
rect 26709 31161 26743 31195
rect 26743 31161 26752 31195
rect 26700 31152 26752 31161
rect 27528 31288 27580 31340
rect 27988 31399 28040 31408
rect 27988 31365 27997 31399
rect 27997 31365 28031 31399
rect 28031 31365 28040 31399
rect 27988 31356 28040 31365
rect 29000 31424 29052 31476
rect 34796 31424 34848 31476
rect 29644 31331 29696 31340
rect 29644 31297 29653 31331
rect 29653 31297 29687 31331
rect 29687 31297 29696 31331
rect 29644 31288 29696 31297
rect 27712 31263 27764 31272
rect 27712 31229 27721 31263
rect 27721 31229 27755 31263
rect 27755 31229 27764 31263
rect 27712 31220 27764 31229
rect 26332 31084 26384 31136
rect 26608 31084 26660 31136
rect 26792 31084 26844 31136
rect 27712 31084 27764 31136
rect 29460 31127 29512 31136
rect 29460 31093 29469 31127
rect 29469 31093 29503 31127
rect 29503 31093 29512 31127
rect 29460 31084 29512 31093
rect 31668 31288 31720 31340
rect 32864 31288 32916 31340
rect 34520 31331 34572 31340
rect 34520 31297 34529 31331
rect 34529 31297 34563 31331
rect 34563 31297 34572 31331
rect 34520 31288 34572 31297
rect 32496 31220 32548 31272
rect 34152 31263 34204 31272
rect 34152 31229 34161 31263
rect 34161 31229 34195 31263
rect 34195 31229 34204 31263
rect 34152 31220 34204 31229
rect 35256 31220 35308 31272
rect 30380 31084 30432 31136
rect 31760 31084 31812 31136
rect 32036 31084 32088 31136
rect 35992 31084 36044 31136
rect 36544 31084 36596 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 7840 30923 7892 30932
rect 7840 30889 7849 30923
rect 7849 30889 7883 30923
rect 7883 30889 7892 30923
rect 7840 30880 7892 30889
rect 8484 30880 8536 30932
rect 13360 30880 13412 30932
rect 13636 30880 13688 30932
rect 14556 30880 14608 30932
rect 17592 30880 17644 30932
rect 18512 30880 18564 30932
rect 19156 30880 19208 30932
rect 7380 30744 7432 30796
rect 8576 30744 8628 30796
rect 9404 30787 9456 30796
rect 9404 30753 9413 30787
rect 9413 30753 9447 30787
rect 9447 30753 9456 30787
rect 9404 30744 9456 30753
rect 9496 30787 9548 30796
rect 9496 30753 9505 30787
rect 9505 30753 9539 30787
rect 9539 30753 9548 30787
rect 9496 30744 9548 30753
rect 4804 30676 4856 30728
rect 5632 30719 5684 30728
rect 5632 30685 5641 30719
rect 5641 30685 5675 30719
rect 5675 30685 5684 30719
rect 5632 30676 5684 30685
rect 6184 30651 6236 30660
rect 6184 30617 6193 30651
rect 6193 30617 6227 30651
rect 6227 30617 6236 30651
rect 6184 30608 6236 30617
rect 4252 30540 4304 30592
rect 4620 30540 4672 30592
rect 6368 30540 6420 30592
rect 11704 30608 11756 30660
rect 12992 30608 13044 30660
rect 13176 30608 13228 30660
rect 7748 30540 7800 30592
rect 10876 30540 10928 30592
rect 13728 30651 13780 30660
rect 13728 30617 13737 30651
rect 13737 30617 13771 30651
rect 13771 30617 13780 30651
rect 14464 30676 14516 30728
rect 14648 30719 14700 30728
rect 14648 30685 14657 30719
rect 14657 30685 14691 30719
rect 14691 30685 14700 30719
rect 14648 30676 14700 30685
rect 14740 30676 14792 30728
rect 16580 30719 16632 30728
rect 16580 30685 16589 30719
rect 16589 30685 16623 30719
rect 16623 30685 16632 30719
rect 16580 30676 16632 30685
rect 16764 30812 16816 30864
rect 17316 30812 17368 30864
rect 18880 30812 18932 30864
rect 20720 30855 20772 30864
rect 20720 30821 20729 30855
rect 20729 30821 20763 30855
rect 20763 30821 20772 30855
rect 20720 30812 20772 30821
rect 21916 30880 21968 30932
rect 22008 30880 22060 30932
rect 16948 30744 17000 30796
rect 17132 30676 17184 30728
rect 17960 30676 18012 30728
rect 19248 30676 19300 30728
rect 20076 30676 20128 30728
rect 20352 30719 20404 30728
rect 20352 30685 20361 30719
rect 20361 30685 20395 30719
rect 20395 30685 20404 30719
rect 20352 30676 20404 30685
rect 20536 30676 20588 30728
rect 21364 30719 21416 30728
rect 21364 30685 21373 30719
rect 21373 30685 21407 30719
rect 21407 30685 21416 30719
rect 21364 30676 21416 30685
rect 22560 30744 22612 30796
rect 23296 30744 23348 30796
rect 23388 30676 23440 30728
rect 24492 30923 24544 30932
rect 24492 30889 24501 30923
rect 24501 30889 24535 30923
rect 24535 30889 24544 30923
rect 24492 30880 24544 30889
rect 25136 30880 25188 30932
rect 26056 30812 26108 30864
rect 27160 30880 27212 30932
rect 28264 30880 28316 30932
rect 29644 30880 29696 30932
rect 30656 30880 30708 30932
rect 26792 30812 26844 30864
rect 24584 30787 24636 30796
rect 24584 30753 24593 30787
rect 24593 30753 24627 30787
rect 24627 30753 24636 30787
rect 24584 30744 24636 30753
rect 27804 30744 27856 30796
rect 28632 30787 28684 30796
rect 28632 30753 28641 30787
rect 28641 30753 28675 30787
rect 28675 30753 28684 30787
rect 28632 30744 28684 30753
rect 24400 30676 24452 30728
rect 13728 30608 13780 30617
rect 13360 30540 13412 30592
rect 13636 30583 13688 30592
rect 13636 30549 13645 30583
rect 13645 30549 13679 30583
rect 13679 30549 13688 30583
rect 13636 30540 13688 30549
rect 14096 30583 14148 30592
rect 14096 30549 14105 30583
rect 14105 30549 14139 30583
rect 14139 30549 14148 30583
rect 14096 30540 14148 30549
rect 14372 30540 14424 30592
rect 14464 30540 14516 30592
rect 14832 30540 14884 30592
rect 16304 30540 16356 30592
rect 16672 30540 16724 30592
rect 18144 30608 18196 30660
rect 18604 30608 18656 30660
rect 19064 30651 19116 30660
rect 19064 30617 19073 30651
rect 19073 30617 19107 30651
rect 19107 30617 19116 30651
rect 19064 30608 19116 30617
rect 19892 30608 19944 30660
rect 17224 30583 17276 30592
rect 17224 30549 17233 30583
rect 17233 30549 17267 30583
rect 17267 30549 17276 30583
rect 17224 30540 17276 30549
rect 17960 30540 18012 30592
rect 20168 30540 20220 30592
rect 20628 30608 20680 30660
rect 21180 30608 21232 30660
rect 20720 30540 20772 30592
rect 20996 30583 21048 30592
rect 20996 30549 21005 30583
rect 21005 30549 21039 30583
rect 21039 30549 21048 30583
rect 20996 30540 21048 30549
rect 21088 30583 21140 30592
rect 21088 30549 21097 30583
rect 21097 30549 21131 30583
rect 21131 30549 21140 30583
rect 23572 30608 23624 30660
rect 21088 30540 21140 30549
rect 21640 30540 21692 30592
rect 24032 30540 24084 30592
rect 25044 30608 25096 30660
rect 26148 30719 26200 30728
rect 26148 30685 26157 30719
rect 26157 30685 26191 30719
rect 26191 30685 26200 30719
rect 26148 30676 26200 30685
rect 26424 30719 26476 30728
rect 26424 30685 26433 30719
rect 26433 30685 26467 30719
rect 26467 30685 26476 30719
rect 26424 30676 26476 30685
rect 27252 30676 27304 30728
rect 27436 30676 27488 30728
rect 32496 30812 32548 30864
rect 33140 30787 33192 30796
rect 33140 30753 33149 30787
rect 33149 30753 33183 30787
rect 33183 30753 33192 30787
rect 33140 30744 33192 30753
rect 33508 30744 33560 30796
rect 29460 30608 29512 30660
rect 30380 30608 30432 30660
rect 30932 30651 30984 30660
rect 30932 30617 30941 30651
rect 30941 30617 30975 30651
rect 30975 30617 30984 30651
rect 30932 30608 30984 30617
rect 31116 30676 31168 30728
rect 31668 30676 31720 30728
rect 34152 30880 34204 30932
rect 35440 30923 35492 30932
rect 35440 30889 35449 30923
rect 35449 30889 35483 30923
rect 35483 30889 35492 30923
rect 35440 30880 35492 30889
rect 33968 30744 34020 30796
rect 31576 30608 31628 30660
rect 36544 30608 36596 30660
rect 28448 30583 28500 30592
rect 28448 30549 28457 30583
rect 28457 30549 28491 30583
rect 28491 30549 28500 30583
rect 28448 30540 28500 30549
rect 31024 30540 31076 30592
rect 31300 30540 31352 30592
rect 33324 30583 33376 30592
rect 33324 30549 33333 30583
rect 33333 30549 33367 30583
rect 33367 30549 33376 30583
rect 33324 30540 33376 30549
rect 4874 30438 4926 30490
rect 4938 30438 4990 30490
rect 5002 30438 5054 30490
rect 5066 30438 5118 30490
rect 5130 30438 5182 30490
rect 35594 30438 35646 30490
rect 35658 30438 35710 30490
rect 35722 30438 35774 30490
rect 35786 30438 35838 30490
rect 35850 30438 35902 30490
rect 5264 30268 5316 30320
rect 6184 30336 6236 30388
rect 4252 30175 4304 30184
rect 4252 30141 4261 30175
rect 4261 30141 4295 30175
rect 4295 30141 4304 30175
rect 4252 30132 4304 30141
rect 7840 30336 7892 30388
rect 9588 30336 9640 30388
rect 13452 30336 13504 30388
rect 13636 30336 13688 30388
rect 14556 30336 14608 30388
rect 14924 30336 14976 30388
rect 18880 30336 18932 30388
rect 7472 30200 7524 30252
rect 7748 30243 7800 30252
rect 7748 30209 7757 30243
rect 7757 30209 7791 30243
rect 7791 30209 7800 30243
rect 7748 30200 7800 30209
rect 7932 30200 7984 30252
rect 8392 30268 8444 30320
rect 9956 30268 10008 30320
rect 8576 30243 8628 30252
rect 8576 30209 8585 30243
rect 8585 30209 8619 30243
rect 8619 30209 8628 30243
rect 8576 30200 8628 30209
rect 9496 30200 9548 30252
rect 10048 30200 10100 30252
rect 11428 30200 11480 30252
rect 11704 30243 11756 30252
rect 11704 30209 11714 30243
rect 11714 30209 11748 30243
rect 11748 30209 11756 30243
rect 11704 30200 11756 30209
rect 11888 30243 11940 30252
rect 11888 30209 11897 30243
rect 11897 30209 11931 30243
rect 11931 30209 11940 30243
rect 11888 30200 11940 30209
rect 12256 30200 12308 30252
rect 16488 30200 16540 30252
rect 18052 30200 18104 30252
rect 18144 30200 18196 30252
rect 18512 30243 18564 30252
rect 18512 30209 18521 30243
rect 18521 30209 18555 30243
rect 18555 30209 18564 30243
rect 18512 30200 18564 30209
rect 18604 30243 18656 30252
rect 18604 30209 18613 30243
rect 18613 30209 18647 30243
rect 18647 30209 18656 30243
rect 18604 30200 18656 30209
rect 18788 30243 18840 30252
rect 18788 30209 18797 30243
rect 18797 30209 18831 30243
rect 18831 30209 18840 30243
rect 18788 30200 18840 30209
rect 19156 30268 19208 30320
rect 19892 30311 19944 30320
rect 19892 30277 19901 30311
rect 19901 30277 19935 30311
rect 19935 30277 19944 30311
rect 19892 30268 19944 30277
rect 20076 30311 20128 30320
rect 20076 30277 20085 30311
rect 20085 30277 20119 30311
rect 20119 30277 20128 30311
rect 20076 30268 20128 30277
rect 23848 30336 23900 30388
rect 24492 30336 24544 30388
rect 20628 30311 20680 30320
rect 20628 30277 20637 30311
rect 20637 30277 20671 30311
rect 20671 30277 20680 30311
rect 20628 30268 20680 30277
rect 20812 30268 20864 30320
rect 24216 30268 24268 30320
rect 20260 30200 20312 30252
rect 30656 30268 30708 30320
rect 31116 30268 31168 30320
rect 14832 30132 14884 30184
rect 16672 30132 16724 30184
rect 17224 30132 17276 30184
rect 5264 29996 5316 30048
rect 5724 29996 5776 30048
rect 6828 29996 6880 30048
rect 9496 30064 9548 30116
rect 14280 30064 14332 30116
rect 14740 30064 14792 30116
rect 18696 30132 18748 30184
rect 25596 30132 25648 30184
rect 7932 29996 7984 30048
rect 9404 29996 9456 30048
rect 12256 30039 12308 30048
rect 12256 30005 12265 30039
rect 12265 30005 12299 30039
rect 12299 30005 12308 30039
rect 12256 29996 12308 30005
rect 12348 29996 12400 30048
rect 13728 29996 13780 30048
rect 15016 29996 15068 30048
rect 15844 29996 15896 30048
rect 16120 29996 16172 30048
rect 16948 29996 17000 30048
rect 18604 30064 18656 30116
rect 20260 30107 20312 30116
rect 20260 30073 20269 30107
rect 20269 30073 20303 30107
rect 20303 30073 20312 30107
rect 20260 30064 20312 30073
rect 18052 30039 18104 30048
rect 18052 30005 18061 30039
rect 18061 30005 18095 30039
rect 18095 30005 18104 30039
rect 18052 29996 18104 30005
rect 18328 29996 18380 30048
rect 19432 29996 19484 30048
rect 25320 30064 25372 30116
rect 25872 30064 25924 30116
rect 20444 29996 20496 30048
rect 20812 30039 20864 30048
rect 20812 30005 20821 30039
rect 20821 30005 20855 30039
rect 20855 30005 20864 30039
rect 20812 29996 20864 30005
rect 20996 29996 21048 30048
rect 26148 30200 26200 30252
rect 31300 30200 31352 30252
rect 29828 30132 29880 30184
rect 30564 30132 30616 30184
rect 30288 30064 30340 30116
rect 31116 30064 31168 30116
rect 32864 30336 32916 30388
rect 32128 30243 32180 30252
rect 32128 30209 32137 30243
rect 32137 30209 32171 30243
rect 32171 30209 32180 30243
rect 32128 30200 32180 30209
rect 32312 30243 32364 30252
rect 32312 30209 32321 30243
rect 32321 30209 32355 30243
rect 32355 30209 32364 30243
rect 32312 30200 32364 30209
rect 33048 30268 33100 30320
rect 33232 30268 33284 30320
rect 35992 30268 36044 30320
rect 32496 30243 32548 30252
rect 32496 30209 32505 30243
rect 32505 30209 32539 30243
rect 32539 30209 32548 30243
rect 32496 30200 32548 30209
rect 26240 30039 26292 30048
rect 26240 30005 26249 30039
rect 26249 30005 26283 30039
rect 26283 30005 26292 30039
rect 26240 29996 26292 30005
rect 26608 29996 26660 30048
rect 32496 29996 32548 30048
rect 32956 29996 33008 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 12256 29792 12308 29844
rect 6828 29656 6880 29708
rect 16580 29792 16632 29844
rect 15384 29724 15436 29776
rect 8300 29631 8352 29640
rect 8300 29597 8309 29631
rect 8309 29597 8343 29631
rect 8343 29597 8352 29631
rect 8300 29588 8352 29597
rect 4620 29520 4672 29572
rect 6828 29520 6880 29572
rect 4068 29495 4120 29504
rect 4068 29461 4077 29495
rect 4077 29461 4111 29495
rect 4111 29461 4120 29495
rect 4068 29452 4120 29461
rect 5448 29495 5500 29504
rect 5448 29461 5457 29495
rect 5457 29461 5491 29495
rect 5491 29461 5500 29495
rect 5448 29452 5500 29461
rect 5908 29495 5960 29504
rect 5908 29461 5917 29495
rect 5917 29461 5951 29495
rect 5951 29461 5960 29495
rect 5908 29452 5960 29461
rect 8392 29452 8444 29504
rect 10968 29588 11020 29640
rect 12716 29631 12768 29640
rect 12716 29597 12725 29631
rect 12725 29597 12759 29631
rect 12759 29597 12768 29631
rect 12716 29588 12768 29597
rect 14832 29656 14884 29708
rect 9680 29520 9732 29572
rect 13544 29631 13596 29640
rect 13544 29597 13553 29631
rect 13553 29597 13587 29631
rect 13587 29597 13596 29631
rect 13544 29588 13596 29597
rect 13820 29631 13872 29640
rect 13820 29597 13829 29631
rect 13829 29597 13863 29631
rect 13863 29597 13872 29631
rect 13820 29588 13872 29597
rect 14096 29588 14148 29640
rect 15200 29588 15252 29640
rect 15568 29588 15620 29640
rect 15660 29631 15712 29640
rect 15660 29597 15669 29631
rect 15669 29597 15703 29631
rect 15703 29597 15712 29631
rect 15660 29588 15712 29597
rect 14832 29520 14884 29572
rect 14924 29520 14976 29572
rect 18696 29792 18748 29844
rect 20352 29792 20404 29844
rect 20628 29792 20680 29844
rect 18052 29724 18104 29776
rect 15844 29588 15896 29640
rect 16028 29631 16080 29640
rect 16028 29597 16045 29631
rect 16045 29597 16079 29631
rect 16079 29597 16080 29631
rect 16028 29588 16080 29597
rect 17500 29588 17552 29640
rect 18144 29588 18196 29640
rect 18328 29631 18380 29640
rect 18328 29597 18337 29631
rect 18337 29597 18371 29631
rect 18371 29597 18380 29631
rect 18328 29588 18380 29597
rect 18972 29724 19024 29776
rect 19984 29724 20036 29776
rect 20260 29724 20312 29776
rect 19708 29656 19760 29708
rect 23112 29792 23164 29844
rect 24492 29792 24544 29844
rect 28080 29792 28132 29844
rect 22928 29724 22980 29776
rect 18696 29631 18748 29640
rect 18696 29597 18705 29631
rect 18705 29597 18739 29631
rect 18739 29597 18748 29631
rect 18696 29588 18748 29597
rect 18880 29588 18932 29640
rect 20812 29588 20864 29640
rect 20996 29588 21048 29640
rect 9036 29452 9088 29504
rect 9956 29452 10008 29504
rect 10692 29495 10744 29504
rect 10692 29461 10701 29495
rect 10701 29461 10735 29495
rect 10735 29461 10744 29495
rect 10692 29452 10744 29461
rect 13176 29452 13228 29504
rect 13268 29495 13320 29504
rect 13268 29461 13277 29495
rect 13277 29461 13311 29495
rect 13311 29461 13320 29495
rect 13268 29452 13320 29461
rect 16764 29452 16816 29504
rect 17040 29495 17092 29504
rect 17040 29461 17049 29495
rect 17049 29461 17083 29495
rect 17083 29461 17092 29495
rect 17040 29452 17092 29461
rect 18512 29563 18564 29572
rect 18512 29529 18521 29563
rect 18521 29529 18555 29563
rect 18555 29529 18564 29563
rect 18512 29520 18564 29529
rect 22100 29588 22152 29640
rect 23204 29588 23256 29640
rect 24400 29724 24452 29776
rect 24768 29724 24820 29776
rect 23480 29656 23532 29708
rect 23756 29631 23808 29640
rect 23756 29597 23765 29631
rect 23765 29597 23799 29631
rect 23799 29597 23808 29631
rect 23756 29588 23808 29597
rect 24032 29631 24084 29640
rect 24032 29597 24041 29631
rect 24041 29597 24075 29631
rect 24075 29597 24084 29631
rect 24032 29588 24084 29597
rect 24584 29588 24636 29640
rect 24768 29631 24820 29640
rect 24768 29597 24777 29631
rect 24777 29597 24811 29631
rect 24811 29597 24820 29631
rect 24768 29588 24820 29597
rect 24860 29588 24912 29640
rect 25780 29631 25832 29640
rect 25780 29597 25803 29631
rect 25803 29597 25832 29631
rect 25780 29588 25832 29597
rect 26516 29724 26568 29776
rect 26608 29724 26660 29776
rect 26332 29656 26384 29708
rect 21548 29520 21600 29572
rect 23112 29563 23164 29572
rect 23112 29529 23121 29563
rect 23121 29529 23155 29563
rect 23155 29529 23164 29563
rect 23112 29520 23164 29529
rect 26056 29588 26108 29640
rect 26424 29631 26476 29640
rect 26424 29597 26433 29631
rect 26433 29597 26467 29631
rect 26467 29597 26476 29631
rect 26424 29588 26476 29597
rect 26884 29724 26936 29776
rect 28908 29724 28960 29776
rect 29092 29724 29144 29776
rect 27620 29699 27672 29708
rect 27620 29665 27629 29699
rect 27629 29665 27663 29699
rect 27663 29665 27672 29699
rect 27620 29656 27672 29665
rect 29000 29656 29052 29708
rect 18420 29452 18472 29504
rect 18880 29495 18932 29504
rect 18880 29461 18889 29495
rect 18889 29461 18923 29495
rect 18923 29461 18932 29495
rect 18880 29452 18932 29461
rect 19064 29452 19116 29504
rect 20720 29452 20772 29504
rect 21088 29452 21140 29504
rect 21180 29495 21232 29504
rect 21180 29461 21189 29495
rect 21189 29461 21223 29495
rect 21223 29461 21232 29495
rect 21180 29452 21232 29461
rect 22744 29495 22796 29504
rect 22744 29461 22753 29495
rect 22753 29461 22787 29495
rect 22787 29461 22796 29495
rect 22744 29452 22796 29461
rect 22836 29452 22888 29504
rect 23296 29452 23348 29504
rect 23572 29495 23624 29504
rect 23572 29461 23581 29495
rect 23581 29461 23615 29495
rect 23615 29461 23624 29495
rect 23572 29452 23624 29461
rect 25412 29452 25464 29504
rect 26332 29520 26384 29572
rect 27344 29495 27396 29504
rect 27344 29461 27353 29495
rect 27353 29461 27387 29495
rect 27387 29461 27396 29495
rect 27344 29452 27396 29461
rect 27620 29452 27672 29504
rect 27804 29452 27856 29504
rect 28080 29452 28132 29504
rect 28908 29588 28960 29640
rect 29828 29631 29880 29640
rect 29828 29597 29837 29631
rect 29837 29597 29871 29631
rect 29871 29597 29880 29631
rect 29828 29588 29880 29597
rect 28448 29520 28500 29572
rect 30012 29631 30064 29640
rect 30012 29597 30021 29631
rect 30021 29597 30055 29631
rect 30055 29597 30064 29631
rect 30012 29588 30064 29597
rect 30104 29520 30156 29572
rect 28356 29495 28408 29504
rect 28356 29461 28365 29495
rect 28365 29461 28399 29495
rect 28399 29461 28408 29495
rect 28356 29452 28408 29461
rect 29276 29495 29328 29504
rect 29276 29461 29285 29495
rect 29285 29461 29319 29495
rect 29319 29461 29328 29495
rect 29276 29452 29328 29461
rect 29368 29452 29420 29504
rect 30656 29631 30708 29640
rect 30656 29597 30665 29631
rect 30665 29597 30699 29631
rect 30699 29597 30708 29631
rect 30656 29588 30708 29597
rect 30840 29588 30892 29640
rect 31300 29588 31352 29640
rect 30564 29563 30616 29572
rect 30564 29529 30573 29563
rect 30573 29529 30607 29563
rect 30607 29529 30616 29563
rect 30564 29520 30616 29529
rect 30288 29452 30340 29504
rect 30380 29452 30432 29504
rect 31300 29452 31352 29504
rect 33508 29724 33560 29776
rect 34244 29724 34296 29776
rect 34152 29631 34204 29640
rect 34152 29597 34161 29631
rect 34161 29597 34195 29631
rect 34195 29597 34204 29631
rect 34152 29588 34204 29597
rect 34796 29631 34848 29640
rect 34796 29597 34805 29631
rect 34805 29597 34839 29631
rect 34839 29597 34848 29631
rect 34796 29588 34848 29597
rect 34336 29520 34388 29572
rect 34980 29520 35032 29572
rect 33324 29452 33376 29504
rect 34520 29495 34572 29504
rect 34520 29461 34529 29495
rect 34529 29461 34563 29495
rect 34563 29461 34572 29495
rect 34520 29452 34572 29461
rect 35992 29452 36044 29504
rect 4874 29350 4926 29402
rect 4938 29350 4990 29402
rect 5002 29350 5054 29402
rect 5066 29350 5118 29402
rect 5130 29350 5182 29402
rect 35594 29350 35646 29402
rect 35658 29350 35710 29402
rect 35722 29350 35774 29402
rect 35786 29350 35838 29402
rect 35850 29350 35902 29402
rect 4068 29248 4120 29300
rect 5908 29248 5960 29300
rect 5264 29112 5316 29164
rect 7472 29248 7524 29300
rect 7564 29248 7616 29300
rect 14832 29248 14884 29300
rect 7932 29180 7984 29232
rect 10692 29180 10744 29232
rect 17960 29180 18012 29232
rect 18696 29248 18748 29300
rect 6828 29044 6880 29096
rect 4712 28908 4764 28960
rect 5356 28908 5408 28960
rect 6552 28908 6604 28960
rect 8300 29044 8352 29096
rect 12716 29112 12768 29164
rect 16120 29112 16172 29164
rect 16856 29112 16908 29164
rect 17408 29112 17460 29164
rect 18604 29112 18656 29164
rect 18972 29180 19024 29232
rect 9128 29044 9180 29096
rect 10784 29044 10836 29096
rect 8300 28908 8352 28960
rect 13728 29044 13780 29096
rect 22468 29248 22520 29300
rect 22560 29248 22612 29300
rect 22744 29248 22796 29300
rect 23204 29248 23256 29300
rect 12900 29019 12952 29028
rect 12900 28985 12909 29019
rect 12909 28985 12943 29019
rect 12943 28985 12952 29019
rect 12900 28976 12952 28985
rect 13176 28976 13228 29028
rect 19800 29112 19852 29164
rect 20812 29112 20864 29164
rect 20904 29155 20956 29164
rect 20904 29121 20913 29155
rect 20913 29121 20947 29155
rect 20947 29121 20956 29155
rect 20904 29112 20956 29121
rect 21640 29180 21692 29232
rect 22100 29223 22152 29232
rect 22100 29189 22109 29223
rect 22109 29189 22143 29223
rect 22143 29189 22152 29223
rect 22100 29180 22152 29189
rect 21180 29112 21232 29164
rect 22008 29155 22060 29164
rect 22008 29121 22015 29155
rect 22015 29121 22060 29155
rect 22008 29112 22060 29121
rect 22192 29155 22244 29164
rect 22192 29121 22201 29155
rect 22201 29121 22235 29155
rect 22235 29121 22244 29155
rect 22192 29112 22244 29121
rect 22284 29155 22336 29164
rect 22284 29121 22298 29155
rect 22298 29121 22332 29155
rect 22332 29121 22336 29155
rect 22284 29112 22336 29121
rect 23020 29155 23072 29164
rect 23020 29121 23029 29155
rect 23029 29121 23063 29155
rect 23063 29121 23072 29155
rect 23020 29112 23072 29121
rect 23664 29223 23716 29232
rect 23664 29189 23673 29223
rect 23673 29189 23707 29223
rect 23707 29189 23716 29223
rect 23664 29180 23716 29189
rect 24032 29180 24084 29232
rect 24216 29112 24268 29164
rect 21548 29044 21600 29096
rect 11520 28908 11572 28960
rect 11612 28908 11664 28960
rect 12624 28908 12676 28960
rect 14648 28908 14700 28960
rect 18328 28908 18380 28960
rect 18604 28951 18656 28960
rect 18604 28917 18613 28951
rect 18613 28917 18647 28951
rect 18647 28917 18656 28951
rect 18604 28908 18656 28917
rect 19156 28908 19208 28960
rect 19616 28908 19668 28960
rect 19984 28908 20036 28960
rect 20076 28908 20128 28960
rect 23204 28951 23256 28960
rect 23204 28917 23213 28951
rect 23213 28917 23247 28951
rect 23247 28917 23256 28951
rect 23204 28908 23256 28917
rect 25044 29044 25096 29096
rect 25596 29155 25648 29164
rect 25596 29121 25605 29155
rect 25605 29121 25639 29155
rect 25639 29121 25648 29155
rect 25596 29112 25648 29121
rect 26424 29248 26476 29300
rect 26516 29248 26568 29300
rect 27344 29248 27396 29300
rect 26240 29112 26292 29164
rect 26516 29155 26568 29164
rect 26516 29121 26525 29155
rect 26525 29121 26559 29155
rect 26559 29121 26568 29155
rect 26516 29112 26568 29121
rect 28356 29248 28408 29300
rect 29000 29291 29052 29300
rect 29000 29257 29009 29291
rect 29009 29257 29043 29291
rect 29043 29257 29052 29291
rect 29000 29248 29052 29257
rect 29276 29248 29328 29300
rect 29828 29248 29880 29300
rect 30288 29248 30340 29300
rect 28632 29112 28684 29164
rect 31116 29180 31168 29232
rect 30012 29044 30064 29096
rect 31300 29248 31352 29300
rect 31484 29180 31536 29232
rect 31576 29223 31628 29232
rect 31576 29189 31585 29223
rect 31585 29189 31619 29223
rect 31619 29189 31628 29223
rect 31576 29180 31628 29189
rect 32312 29248 32364 29300
rect 32496 29248 32548 29300
rect 34152 29248 34204 29300
rect 34796 29248 34848 29300
rect 33232 29180 33284 29232
rect 34336 29180 34388 29232
rect 33048 29155 33100 29164
rect 33048 29121 33057 29155
rect 33057 29121 33091 29155
rect 33091 29121 33100 29155
rect 33048 29112 33100 29121
rect 34520 29112 34572 29164
rect 34980 29112 35032 29164
rect 36636 29155 36688 29164
rect 36636 29121 36645 29155
rect 36645 29121 36679 29155
rect 36679 29121 36688 29155
rect 36636 29112 36688 29121
rect 36820 29155 36872 29164
rect 36820 29121 36829 29155
rect 36829 29121 36863 29155
rect 36863 29121 36872 29155
rect 36820 29112 36872 29121
rect 24216 28976 24268 29028
rect 24860 28976 24912 29028
rect 26516 28976 26568 29028
rect 27068 28976 27120 29028
rect 23940 28908 23992 28960
rect 26976 28908 27028 28960
rect 29092 28976 29144 29028
rect 29276 28908 29328 28960
rect 30104 28908 30156 28960
rect 31668 28976 31720 29028
rect 34704 28976 34756 29028
rect 37280 28976 37332 29028
rect 32404 28908 32456 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 4712 28704 4764 28756
rect 8024 28704 8076 28756
rect 14648 28704 14700 28756
rect 8300 28636 8352 28688
rect 9496 28636 9548 28688
rect 11520 28636 11572 28688
rect 12072 28636 12124 28688
rect 20260 28704 20312 28756
rect 21548 28704 21600 28756
rect 23572 28704 23624 28756
rect 24308 28704 24360 28756
rect 24768 28704 24820 28756
rect 25596 28704 25648 28756
rect 6552 28568 6604 28620
rect 19340 28636 19392 28688
rect 20076 28636 20128 28688
rect 22008 28636 22060 28688
rect 29092 28704 29144 28756
rect 5448 28500 5500 28552
rect 5632 28500 5684 28552
rect 4252 28407 4304 28416
rect 4252 28373 4261 28407
rect 4261 28373 4295 28407
rect 4295 28373 4304 28407
rect 4252 28364 4304 28373
rect 7196 28432 7248 28484
rect 8116 28432 8168 28484
rect 9956 28543 10008 28552
rect 9956 28509 9965 28543
rect 9965 28509 9999 28543
rect 9999 28509 10008 28543
rect 9956 28500 10008 28509
rect 16120 28543 16172 28552
rect 16120 28509 16129 28543
rect 16129 28509 16163 28543
rect 16163 28509 16172 28543
rect 16120 28500 16172 28509
rect 16212 28500 16264 28552
rect 16488 28543 16540 28552
rect 16488 28509 16497 28543
rect 16497 28509 16531 28543
rect 16531 28509 16540 28543
rect 16488 28500 16540 28509
rect 17868 28500 17920 28552
rect 18328 28568 18380 28620
rect 19616 28568 19668 28620
rect 18052 28500 18104 28552
rect 10416 28432 10468 28484
rect 10508 28475 10560 28484
rect 10508 28441 10517 28475
rect 10517 28441 10551 28475
rect 10551 28441 10560 28475
rect 10508 28432 10560 28441
rect 11060 28432 11112 28484
rect 16580 28432 16632 28484
rect 19800 28543 19852 28552
rect 19800 28509 19809 28543
rect 19809 28509 19843 28543
rect 19843 28509 19852 28543
rect 19800 28500 19852 28509
rect 19616 28432 19668 28484
rect 20168 28500 20220 28552
rect 20996 28500 21048 28552
rect 25320 28568 25372 28620
rect 25596 28568 25648 28620
rect 22744 28500 22796 28552
rect 24492 28500 24544 28552
rect 24676 28543 24728 28552
rect 24676 28509 24685 28543
rect 24685 28509 24719 28543
rect 24719 28509 24728 28543
rect 24676 28500 24728 28509
rect 24860 28500 24912 28552
rect 29276 28679 29328 28688
rect 29276 28645 29285 28679
rect 29285 28645 29319 28679
rect 29319 28645 29328 28679
rect 29276 28636 29328 28645
rect 30012 28611 30064 28620
rect 30012 28577 30021 28611
rect 30021 28577 30055 28611
rect 30055 28577 30064 28611
rect 30012 28568 30064 28577
rect 30288 28568 30340 28620
rect 8208 28407 8260 28416
rect 8208 28373 8217 28407
rect 8217 28373 8251 28407
rect 8251 28373 8260 28407
rect 8208 28364 8260 28373
rect 11980 28407 12032 28416
rect 11980 28373 11989 28407
rect 11989 28373 12023 28407
rect 12023 28373 12032 28407
rect 11980 28364 12032 28373
rect 17224 28364 17276 28416
rect 19432 28364 19484 28416
rect 22376 28364 22428 28416
rect 23940 28364 23992 28416
rect 24400 28407 24452 28416
rect 24400 28373 24409 28407
rect 24409 28373 24443 28407
rect 24443 28373 24452 28407
rect 24400 28364 24452 28373
rect 24768 28475 24820 28484
rect 24768 28441 24777 28475
rect 24777 28441 24811 28475
rect 24811 28441 24820 28475
rect 24768 28432 24820 28441
rect 26148 28475 26200 28484
rect 26148 28441 26157 28475
rect 26157 28441 26191 28475
rect 26191 28441 26200 28475
rect 26148 28432 26200 28441
rect 31484 28636 31536 28688
rect 30380 28543 30432 28552
rect 30380 28509 30389 28543
rect 30389 28509 30423 28543
rect 30423 28509 30432 28543
rect 30380 28500 30432 28509
rect 30564 28500 30616 28552
rect 30748 28543 30800 28552
rect 30748 28509 30757 28543
rect 30757 28509 30791 28543
rect 30791 28509 30800 28543
rect 30748 28500 30800 28509
rect 30840 28543 30892 28552
rect 30840 28509 30854 28543
rect 30854 28509 30888 28543
rect 30888 28509 30892 28543
rect 30840 28500 30892 28509
rect 30196 28364 30248 28416
rect 31392 28500 31444 28552
rect 32404 28568 32456 28620
rect 33324 28568 33376 28620
rect 33968 28568 34020 28620
rect 31760 28543 31812 28552
rect 31760 28509 31769 28543
rect 31769 28509 31803 28543
rect 31803 28509 31812 28543
rect 31760 28500 31812 28509
rect 34704 28543 34756 28552
rect 34704 28509 34713 28543
rect 34713 28509 34747 28543
rect 34747 28509 34756 28543
rect 34704 28500 34756 28509
rect 34060 28432 34112 28484
rect 34428 28432 34480 28484
rect 35992 28432 36044 28484
rect 31116 28407 31168 28416
rect 31116 28373 31125 28407
rect 31125 28373 31159 28407
rect 31159 28373 31168 28407
rect 31116 28364 31168 28373
rect 32680 28364 32732 28416
rect 34152 28407 34204 28416
rect 34152 28373 34161 28407
rect 34161 28373 34195 28407
rect 34195 28373 34204 28407
rect 34152 28364 34204 28373
rect 34520 28407 34572 28416
rect 34520 28373 34529 28407
rect 34529 28373 34563 28407
rect 34563 28373 34572 28407
rect 34520 28364 34572 28373
rect 4874 28262 4926 28314
rect 4938 28262 4990 28314
rect 5002 28262 5054 28314
rect 5066 28262 5118 28314
rect 5130 28262 5182 28314
rect 35594 28262 35646 28314
rect 35658 28262 35710 28314
rect 35722 28262 35774 28314
rect 35786 28262 35838 28314
rect 35850 28262 35902 28314
rect 4252 28160 4304 28212
rect 8024 28160 8076 28212
rect 8208 28160 8260 28212
rect 10508 28160 10560 28212
rect 6828 28135 6880 28144
rect 6828 28101 6837 28135
rect 6837 28101 6871 28135
rect 6871 28101 6880 28135
rect 6828 28092 6880 28101
rect 5448 28024 5500 28076
rect 9496 28092 9548 28144
rect 11244 28092 11296 28144
rect 4712 27956 4764 28008
rect 7012 27999 7064 28008
rect 7012 27965 7021 27999
rect 7021 27965 7055 27999
rect 7055 27965 7064 27999
rect 7012 27956 7064 27965
rect 8300 27956 8352 28008
rect 6368 27863 6420 27872
rect 6368 27829 6377 27863
rect 6377 27829 6411 27863
rect 6411 27829 6420 27863
rect 6368 27820 6420 27829
rect 7196 27820 7248 27872
rect 9680 28024 9732 28076
rect 9772 28024 9824 28076
rect 13360 28160 13412 28212
rect 13912 28203 13964 28212
rect 13912 28169 13921 28203
rect 13921 28169 13955 28203
rect 13955 28169 13964 28203
rect 13912 28160 13964 28169
rect 15752 28160 15804 28212
rect 16120 28160 16172 28212
rect 17500 28160 17552 28212
rect 17592 28160 17644 28212
rect 18788 28160 18840 28212
rect 11980 28092 12032 28144
rect 14096 28092 14148 28144
rect 12624 28067 12676 28076
rect 12624 28033 12633 28067
rect 12633 28033 12667 28067
rect 12667 28033 12676 28067
rect 12624 28024 12676 28033
rect 10140 27999 10192 28008
rect 10140 27965 10149 27999
rect 10149 27965 10183 27999
rect 10183 27965 10192 27999
rect 10140 27956 10192 27965
rect 11980 27999 12032 28008
rect 11980 27965 11989 27999
rect 11989 27965 12023 27999
rect 12023 27965 12032 27999
rect 11980 27956 12032 27965
rect 12072 27999 12124 28008
rect 12072 27965 12081 27999
rect 12081 27965 12115 27999
rect 12115 27965 12124 27999
rect 12072 27956 12124 27965
rect 13452 28024 13504 28076
rect 14556 28024 14608 28076
rect 14648 28067 14700 28076
rect 14648 28033 14657 28067
rect 14657 28033 14691 28067
rect 14691 28033 14700 28067
rect 14648 28024 14700 28033
rect 16580 28092 16632 28144
rect 17408 28092 17460 28144
rect 19248 28135 19300 28144
rect 15016 28024 15068 28076
rect 16028 28024 16080 28076
rect 16672 28067 16724 28076
rect 16672 28033 16681 28067
rect 16681 28033 16715 28067
rect 16715 28033 16724 28067
rect 16672 28024 16724 28033
rect 16764 28067 16816 28076
rect 16764 28033 16774 28067
rect 16774 28033 16808 28067
rect 16808 28033 16816 28067
rect 16764 28024 16816 28033
rect 9496 27820 9548 27872
rect 9772 27820 9824 27872
rect 11980 27820 12032 27872
rect 17868 28024 17920 28076
rect 18328 28024 18380 28076
rect 18880 28024 18932 28076
rect 19248 28101 19273 28135
rect 19273 28101 19300 28135
rect 19248 28092 19300 28101
rect 19524 28024 19576 28076
rect 19616 28067 19668 28076
rect 19616 28033 19625 28067
rect 19625 28033 19659 28067
rect 19659 28033 19668 28067
rect 19616 28024 19668 28033
rect 19800 28067 19852 28076
rect 19800 28033 19809 28067
rect 19809 28033 19843 28067
rect 19843 28033 19852 28067
rect 19800 28024 19852 28033
rect 19984 28092 20036 28144
rect 20628 28067 20680 28076
rect 20628 28033 20637 28067
rect 20637 28033 20671 28067
rect 20671 28033 20680 28067
rect 21088 28135 21140 28144
rect 21088 28101 21097 28135
rect 21097 28101 21131 28135
rect 21131 28101 21140 28135
rect 21088 28092 21140 28101
rect 22192 28160 22244 28212
rect 23020 28160 23072 28212
rect 23572 28160 23624 28212
rect 24676 28160 24728 28212
rect 30748 28160 30800 28212
rect 31760 28160 31812 28212
rect 21548 28092 21600 28144
rect 20628 28024 20680 28033
rect 15568 27888 15620 27940
rect 13636 27820 13688 27872
rect 14188 27863 14240 27872
rect 14188 27829 14197 27863
rect 14197 27829 14231 27863
rect 14231 27829 14240 27863
rect 14188 27820 14240 27829
rect 14464 27863 14516 27872
rect 14464 27829 14473 27863
rect 14473 27829 14507 27863
rect 14507 27829 14516 27863
rect 14464 27820 14516 27829
rect 15476 27820 15528 27872
rect 15844 27820 15896 27872
rect 19248 27863 19300 27872
rect 19248 27829 19257 27863
rect 19257 27829 19291 27863
rect 19291 27829 19300 27863
rect 19248 27820 19300 27829
rect 20260 27956 20312 28008
rect 20444 27999 20496 28008
rect 20444 27965 20453 27999
rect 20453 27965 20487 27999
rect 20487 27965 20496 27999
rect 20444 27956 20496 27965
rect 20352 27820 20404 27872
rect 20444 27820 20496 27872
rect 21456 28024 21508 28076
rect 22376 28024 22428 28076
rect 22468 28067 22520 28076
rect 22468 28033 22477 28067
rect 22477 28033 22511 28067
rect 22511 28033 22520 28067
rect 22468 28024 22520 28033
rect 23204 28024 23256 28076
rect 21916 27999 21968 28008
rect 21916 27965 21925 27999
rect 21925 27965 21959 27999
rect 21959 27965 21968 27999
rect 21916 27956 21968 27965
rect 22928 27956 22980 28008
rect 23388 28067 23440 28076
rect 23388 28033 23397 28067
rect 23397 28033 23431 28067
rect 23431 28033 23440 28067
rect 23388 28024 23440 28033
rect 32680 28160 32732 28212
rect 33048 28160 33100 28212
rect 34428 28203 34480 28212
rect 34428 28169 34437 28203
rect 34437 28169 34471 28203
rect 34471 28169 34480 28203
rect 34428 28160 34480 28169
rect 34704 28160 34756 28212
rect 37280 28160 37332 28212
rect 23572 27956 23624 28008
rect 24216 28024 24268 28076
rect 24400 28024 24452 28076
rect 24676 28024 24728 28076
rect 31852 28024 31904 28076
rect 31944 28067 31996 28076
rect 31944 28033 31953 28067
rect 31953 28033 31987 28067
rect 31987 28033 31996 28067
rect 31944 28024 31996 28033
rect 23756 27888 23808 27940
rect 30196 27956 30248 28008
rect 34152 28024 34204 28076
rect 34520 28024 34572 28076
rect 33140 27956 33192 28008
rect 33876 27956 33928 28008
rect 33692 27888 33744 27940
rect 34612 27888 34664 27940
rect 23388 27820 23440 27872
rect 24216 27863 24268 27872
rect 24216 27829 24225 27863
rect 24225 27829 24259 27863
rect 24259 27829 24268 27863
rect 24216 27820 24268 27829
rect 24492 27863 24544 27872
rect 24492 27829 24501 27863
rect 24501 27829 24535 27863
rect 24535 27829 24544 27863
rect 24492 27820 24544 27829
rect 37556 27863 37608 27872
rect 37556 27829 37565 27863
rect 37565 27829 37599 27863
rect 37599 27829 37608 27863
rect 37556 27820 37608 27829
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 4712 27616 4764 27668
rect 8300 27659 8352 27668
rect 8300 27625 8309 27659
rect 8309 27625 8343 27659
rect 8343 27625 8352 27659
rect 8300 27616 8352 27625
rect 9496 27616 9548 27668
rect 12624 27616 12676 27668
rect 13176 27616 13228 27668
rect 14188 27616 14240 27668
rect 14464 27616 14516 27668
rect 14648 27659 14700 27668
rect 14648 27625 14657 27659
rect 14657 27625 14691 27659
rect 14691 27625 14700 27659
rect 14648 27616 14700 27625
rect 7564 27480 7616 27532
rect 6368 27412 6420 27464
rect 9588 27548 9640 27600
rect 11980 27480 12032 27532
rect 13912 27548 13964 27600
rect 14096 27591 14148 27600
rect 14096 27557 14105 27591
rect 14105 27557 14139 27591
rect 14139 27557 14148 27591
rect 16580 27616 16632 27668
rect 16672 27616 16724 27668
rect 14096 27548 14148 27557
rect 15016 27548 15068 27600
rect 15292 27548 15344 27600
rect 11060 27412 11112 27464
rect 13728 27480 13780 27532
rect 16304 27480 16356 27532
rect 16580 27480 16632 27532
rect 21456 27616 21508 27668
rect 22008 27616 22060 27668
rect 23572 27616 23624 27668
rect 24216 27616 24268 27668
rect 25044 27616 25096 27668
rect 26608 27616 26660 27668
rect 26700 27616 26752 27668
rect 27896 27616 27948 27668
rect 28448 27616 28500 27668
rect 29736 27616 29788 27668
rect 10048 27387 10100 27396
rect 10048 27353 10057 27387
rect 10057 27353 10091 27387
rect 10091 27353 10100 27387
rect 10048 27344 10100 27353
rect 6828 27319 6880 27328
rect 6828 27285 6837 27319
rect 6837 27285 6871 27319
rect 6871 27285 6880 27319
rect 6828 27276 6880 27285
rect 9864 27276 9916 27328
rect 13452 27412 13504 27464
rect 14372 27412 14424 27464
rect 14832 27412 14884 27464
rect 12348 27344 12400 27396
rect 15844 27455 15896 27464
rect 15844 27421 15853 27455
rect 15853 27421 15887 27455
rect 15887 27421 15896 27455
rect 15844 27412 15896 27421
rect 16212 27412 16264 27464
rect 16672 27455 16724 27464
rect 16672 27421 16681 27455
rect 16681 27421 16715 27455
rect 16715 27421 16724 27455
rect 16672 27412 16724 27421
rect 16764 27455 16816 27464
rect 16764 27421 16774 27455
rect 16774 27421 16808 27455
rect 16808 27421 16816 27455
rect 16764 27412 16816 27421
rect 18328 27548 18380 27600
rect 18512 27548 18564 27600
rect 23664 27548 23716 27600
rect 25504 27548 25556 27600
rect 29000 27548 29052 27600
rect 17132 27455 17184 27464
rect 17132 27421 17146 27455
rect 17146 27421 17180 27455
rect 17180 27421 17184 27455
rect 17132 27412 17184 27421
rect 17316 27412 17368 27464
rect 17408 27455 17460 27464
rect 17408 27421 17417 27455
rect 17417 27421 17451 27455
rect 17451 27421 17460 27455
rect 17408 27412 17460 27421
rect 17500 27412 17552 27464
rect 18696 27480 18748 27532
rect 20352 27480 20404 27532
rect 21548 27480 21600 27532
rect 18144 27455 18196 27464
rect 18144 27421 18153 27455
rect 18153 27421 18187 27455
rect 18187 27421 18196 27455
rect 18144 27412 18196 27421
rect 11612 27319 11664 27328
rect 11612 27285 11621 27319
rect 11621 27285 11655 27319
rect 11655 27285 11664 27319
rect 11612 27276 11664 27285
rect 13360 27276 13412 27328
rect 14096 27276 14148 27328
rect 14556 27276 14608 27328
rect 15384 27276 15436 27328
rect 17960 27344 18012 27396
rect 17316 27319 17368 27328
rect 17316 27285 17325 27319
rect 17325 27285 17359 27319
rect 17359 27285 17368 27319
rect 17316 27276 17368 27285
rect 17776 27276 17828 27328
rect 18972 27412 19024 27464
rect 21272 27412 21324 27464
rect 23388 27480 23440 27532
rect 18512 27387 18564 27396
rect 18512 27353 18521 27387
rect 18521 27353 18555 27387
rect 18555 27353 18564 27387
rect 18512 27344 18564 27353
rect 20628 27344 20680 27396
rect 21824 27344 21876 27396
rect 18788 27319 18840 27328
rect 18788 27285 18797 27319
rect 18797 27285 18831 27319
rect 18831 27285 18840 27319
rect 18788 27276 18840 27285
rect 20168 27276 20220 27328
rect 23572 27455 23624 27464
rect 23572 27421 23581 27455
rect 23581 27421 23615 27455
rect 23615 27421 23624 27455
rect 23572 27412 23624 27421
rect 24124 27412 24176 27464
rect 25044 27412 25096 27464
rect 26424 27480 26476 27532
rect 31852 27548 31904 27600
rect 33784 27591 33836 27600
rect 33784 27557 33793 27591
rect 33793 27557 33827 27591
rect 33827 27557 33836 27591
rect 33784 27548 33836 27557
rect 34336 27548 34388 27600
rect 28172 27455 28224 27464
rect 28172 27421 28181 27455
rect 28181 27421 28215 27455
rect 28215 27421 28224 27455
rect 28172 27412 28224 27421
rect 22192 27276 22244 27328
rect 25688 27344 25740 27396
rect 26332 27344 26384 27396
rect 26792 27344 26844 27396
rect 30012 27455 30064 27464
rect 30012 27421 30021 27455
rect 30021 27421 30055 27455
rect 30055 27421 30064 27455
rect 30012 27412 30064 27421
rect 30380 27455 30432 27464
rect 30380 27421 30389 27455
rect 30389 27421 30423 27455
rect 30423 27421 30432 27455
rect 30380 27412 30432 27421
rect 30564 27412 30616 27464
rect 30840 27412 30892 27464
rect 31024 27412 31076 27464
rect 31944 27412 31996 27464
rect 33692 27455 33744 27464
rect 33692 27421 33701 27455
rect 33701 27421 33735 27455
rect 33735 27421 33744 27455
rect 33692 27412 33744 27421
rect 27804 27319 27856 27328
rect 27804 27285 27813 27319
rect 27813 27285 27847 27319
rect 27847 27285 27856 27319
rect 27804 27276 27856 27285
rect 27896 27276 27948 27328
rect 29644 27319 29696 27328
rect 29644 27285 29653 27319
rect 29653 27285 29687 27319
rect 29687 27285 29696 27319
rect 29644 27276 29696 27285
rect 29828 27319 29880 27328
rect 29828 27285 29837 27319
rect 29837 27285 29871 27319
rect 29871 27285 29880 27319
rect 29828 27276 29880 27285
rect 30104 27276 30156 27328
rect 30748 27276 30800 27328
rect 31760 27276 31812 27328
rect 33600 27319 33652 27328
rect 33600 27285 33609 27319
rect 33609 27285 33643 27319
rect 33643 27285 33652 27319
rect 33600 27276 33652 27285
rect 4874 27174 4926 27226
rect 4938 27174 4990 27226
rect 5002 27174 5054 27226
rect 5066 27174 5118 27226
rect 5130 27174 5182 27226
rect 35594 27174 35646 27226
rect 35658 27174 35710 27226
rect 35722 27174 35774 27226
rect 35786 27174 35838 27226
rect 35850 27174 35902 27226
rect 6828 27072 6880 27124
rect 7012 27072 7064 27124
rect 9864 27072 9916 27124
rect 10048 27072 10100 27124
rect 11612 27072 11664 27124
rect 12256 27072 12308 27124
rect 7196 27004 7248 27056
rect 6920 26911 6972 26920
rect 6920 26877 6929 26911
rect 6929 26877 6963 26911
rect 6963 26877 6972 26911
rect 6920 26868 6972 26877
rect 11428 26868 11480 26920
rect 11980 26868 12032 26920
rect 12348 26979 12400 26988
rect 12348 26945 12358 26979
rect 12358 26945 12392 26979
rect 12392 26945 12400 26979
rect 12348 26936 12400 26945
rect 16580 27072 16632 27124
rect 16672 27115 16724 27124
rect 16672 27081 16681 27115
rect 16681 27081 16715 27115
rect 16715 27081 16724 27115
rect 16672 27072 16724 27081
rect 16948 27115 17000 27124
rect 16948 27081 16957 27115
rect 16957 27081 16991 27115
rect 16991 27081 17000 27115
rect 16948 27072 17000 27081
rect 17224 27072 17276 27124
rect 17316 27072 17368 27124
rect 18512 27072 18564 27124
rect 18696 27072 18748 27124
rect 18972 27072 19024 27124
rect 15476 27047 15528 27056
rect 15476 27013 15485 27047
rect 15485 27013 15519 27047
rect 15519 27013 15528 27047
rect 15476 27004 15528 27013
rect 14464 26967 14495 26988
rect 14495 26967 14516 26988
rect 7656 26732 7708 26784
rect 8576 26800 8628 26852
rect 11888 26800 11940 26852
rect 12348 26800 12400 26852
rect 14464 26936 14516 26967
rect 14924 26979 14976 26988
rect 14924 26945 14933 26979
rect 14933 26945 14967 26979
rect 14967 26945 14976 26979
rect 14924 26936 14976 26945
rect 15660 26979 15712 26988
rect 15660 26945 15669 26979
rect 15669 26945 15703 26979
rect 15703 26945 15712 26979
rect 15660 26936 15712 26945
rect 8392 26775 8444 26784
rect 8392 26741 8401 26775
rect 8401 26741 8435 26775
rect 8435 26741 8444 26775
rect 8392 26732 8444 26741
rect 12900 26775 12952 26784
rect 12900 26741 12909 26775
rect 12909 26741 12943 26775
rect 12943 26741 12952 26775
rect 12900 26732 12952 26741
rect 14280 26775 14332 26784
rect 14280 26741 14289 26775
rect 14289 26741 14323 26775
rect 14323 26741 14332 26775
rect 14280 26732 14332 26741
rect 14648 26911 14700 26920
rect 14648 26877 14657 26911
rect 14657 26877 14691 26911
rect 14691 26877 14700 26911
rect 14648 26868 14700 26877
rect 14740 26911 14792 26920
rect 14740 26877 14749 26911
rect 14749 26877 14783 26911
rect 14783 26877 14792 26911
rect 14740 26868 14792 26877
rect 15108 26800 15160 26852
rect 15384 26800 15436 26852
rect 17040 26979 17092 26988
rect 17040 26945 17049 26979
rect 17049 26945 17083 26979
rect 17083 26945 17092 26979
rect 17040 26936 17092 26945
rect 21732 26936 21784 26988
rect 22376 26979 22428 26988
rect 22376 26945 22385 26979
rect 22385 26945 22419 26979
rect 22419 26945 22428 26979
rect 22376 26936 22428 26945
rect 23480 27004 23532 27056
rect 26332 27072 26384 27124
rect 27804 27072 27856 27124
rect 28632 27072 28684 27124
rect 26424 27047 26476 27056
rect 26424 27013 26433 27047
rect 26433 27013 26467 27047
rect 26467 27013 26476 27047
rect 26424 27004 26476 27013
rect 16948 26868 17000 26920
rect 18512 26868 18564 26920
rect 18972 26868 19024 26920
rect 20076 26868 20128 26920
rect 24952 26936 25004 26988
rect 24860 26868 24912 26920
rect 26700 26936 26752 26988
rect 17132 26800 17184 26852
rect 17224 26843 17276 26852
rect 17224 26809 17233 26843
rect 17233 26809 17267 26843
rect 17267 26809 17276 26843
rect 17224 26800 17276 26809
rect 21916 26800 21968 26852
rect 17684 26775 17736 26784
rect 17684 26741 17693 26775
rect 17693 26741 17727 26775
rect 17727 26741 17736 26775
rect 17684 26732 17736 26741
rect 18144 26732 18196 26784
rect 18604 26732 18656 26784
rect 19616 26732 19668 26784
rect 20720 26732 20772 26784
rect 22192 26775 22244 26784
rect 22192 26741 22201 26775
rect 22201 26741 22235 26775
rect 22235 26741 22244 26775
rect 22192 26732 22244 26741
rect 27896 26868 27948 26920
rect 29644 27072 29696 27124
rect 29828 27072 29880 27124
rect 31576 27072 31628 27124
rect 34060 27072 34112 27124
rect 32128 26936 32180 26988
rect 33140 26979 33192 26988
rect 33140 26945 33149 26979
rect 33149 26945 33183 26979
rect 33183 26945 33192 26979
rect 33140 26936 33192 26945
rect 33600 27004 33652 27056
rect 35992 26936 36044 26988
rect 29460 26800 29512 26852
rect 35440 26911 35492 26920
rect 35440 26877 35449 26911
rect 35449 26877 35483 26911
rect 35483 26877 35492 26911
rect 35440 26868 35492 26877
rect 27344 26732 27396 26784
rect 28264 26732 28316 26784
rect 30104 26732 30156 26784
rect 31392 26732 31444 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 6920 26528 6972 26580
rect 7656 26460 7708 26512
rect 4528 26367 4580 26376
rect 4528 26333 4537 26367
rect 4537 26333 4571 26367
rect 4571 26333 4580 26367
rect 4528 26324 4580 26333
rect 11152 26528 11204 26580
rect 12900 26528 12952 26580
rect 14280 26528 14332 26580
rect 14648 26528 14700 26580
rect 15108 26571 15160 26580
rect 15108 26537 15117 26571
rect 15117 26537 15151 26571
rect 15151 26537 15160 26571
rect 15108 26528 15160 26537
rect 15292 26528 15344 26580
rect 8392 26460 8444 26512
rect 9588 26460 9640 26512
rect 8576 26435 8628 26444
rect 8576 26401 8585 26435
rect 8585 26401 8619 26435
rect 8619 26401 8628 26435
rect 8576 26392 8628 26401
rect 12348 26324 12400 26376
rect 12624 26324 12676 26376
rect 14280 26392 14332 26444
rect 13636 26367 13688 26376
rect 13636 26333 13645 26367
rect 13645 26333 13679 26367
rect 13679 26333 13688 26367
rect 13636 26324 13688 26333
rect 13820 26324 13872 26376
rect 14832 26392 14884 26444
rect 5356 26256 5408 26308
rect 3884 26188 3936 26240
rect 5540 26256 5592 26308
rect 6000 26188 6052 26240
rect 7196 26256 7248 26308
rect 6920 26231 6972 26240
rect 6920 26197 6929 26231
rect 6929 26197 6963 26231
rect 6963 26197 6972 26231
rect 6920 26188 6972 26197
rect 8484 26299 8536 26308
rect 8484 26265 8493 26299
rect 8493 26265 8527 26299
rect 8527 26265 8536 26299
rect 8484 26256 8536 26265
rect 11152 26256 11204 26308
rect 14464 26256 14516 26308
rect 17224 26460 17276 26512
rect 17684 26528 17736 26580
rect 18052 26528 18104 26580
rect 17592 26460 17644 26512
rect 18328 26460 18380 26512
rect 19340 26460 19392 26512
rect 20904 26460 20956 26512
rect 22652 26460 22704 26512
rect 15108 26392 15160 26444
rect 15384 26392 15436 26444
rect 15568 26324 15620 26376
rect 8668 26188 8720 26240
rect 14648 26188 14700 26240
rect 15108 26188 15160 26240
rect 16856 26367 16908 26376
rect 16856 26333 16865 26367
rect 16865 26333 16899 26367
rect 16899 26333 16908 26367
rect 16856 26324 16908 26333
rect 20352 26392 20404 26444
rect 17224 26367 17276 26376
rect 17224 26333 17233 26367
rect 17233 26333 17267 26367
rect 17267 26333 17276 26367
rect 17224 26324 17276 26333
rect 18696 26324 18748 26376
rect 18972 26324 19024 26376
rect 19248 26324 19300 26376
rect 19340 26324 19392 26376
rect 19708 26324 19760 26376
rect 16488 26188 16540 26240
rect 16764 26188 16816 26240
rect 20168 26256 20220 26308
rect 20352 26256 20404 26308
rect 18972 26188 19024 26240
rect 21272 26392 21324 26444
rect 22008 26324 22060 26376
rect 22376 26324 22428 26376
rect 23756 26324 23808 26376
rect 24492 26324 24544 26376
rect 24584 26324 24636 26376
rect 25504 26392 25556 26444
rect 26792 26460 26844 26512
rect 27528 26460 27580 26512
rect 28172 26528 28224 26580
rect 30012 26528 30064 26580
rect 30748 26460 30800 26512
rect 33140 26528 33192 26580
rect 35440 26528 35492 26580
rect 20812 26188 20864 26240
rect 23020 26256 23072 26308
rect 24860 26256 24912 26308
rect 25688 26367 25740 26376
rect 25688 26333 25697 26367
rect 25697 26333 25731 26367
rect 25731 26333 25740 26367
rect 25688 26324 25740 26333
rect 26332 26367 26384 26376
rect 26332 26333 26341 26367
rect 26341 26333 26375 26367
rect 26375 26333 26384 26367
rect 26332 26324 26384 26333
rect 27620 26392 27672 26444
rect 27988 26392 28040 26444
rect 30288 26392 30340 26444
rect 30472 26392 30524 26444
rect 31392 26392 31444 26444
rect 31852 26392 31904 26444
rect 26608 26367 26660 26376
rect 26608 26333 26617 26367
rect 26617 26333 26651 26367
rect 26651 26333 26660 26367
rect 26608 26324 26660 26333
rect 21548 26188 21600 26240
rect 23756 26231 23808 26240
rect 23756 26197 23765 26231
rect 23765 26197 23799 26231
rect 23799 26197 23808 26231
rect 23756 26188 23808 26197
rect 26148 26256 26200 26308
rect 26240 26256 26292 26308
rect 30104 26324 30156 26376
rect 33876 26435 33928 26444
rect 33876 26401 33885 26435
rect 33885 26401 33919 26435
rect 33919 26401 33928 26435
rect 33876 26392 33928 26401
rect 34704 26367 34756 26376
rect 34704 26333 34713 26367
rect 34713 26333 34747 26367
rect 34747 26333 34756 26367
rect 34704 26324 34756 26333
rect 34980 26367 35032 26376
rect 34980 26333 34989 26367
rect 34989 26333 35023 26367
rect 35023 26333 35032 26367
rect 34980 26324 35032 26333
rect 28264 26299 28316 26308
rect 28264 26265 28273 26299
rect 28273 26265 28307 26299
rect 28307 26265 28316 26299
rect 28264 26256 28316 26265
rect 25688 26188 25740 26240
rect 26056 26231 26108 26240
rect 26056 26197 26065 26231
rect 26065 26197 26099 26231
rect 26099 26197 26108 26231
rect 26056 26188 26108 26197
rect 27344 26188 27396 26240
rect 28172 26231 28224 26240
rect 28172 26197 28181 26231
rect 28181 26197 28215 26231
rect 28215 26197 28224 26231
rect 28172 26188 28224 26197
rect 29092 26188 29144 26240
rect 31576 26256 31628 26308
rect 35992 26256 36044 26308
rect 36636 26256 36688 26308
rect 30012 26188 30064 26240
rect 30288 26188 30340 26240
rect 31668 26188 31720 26240
rect 33232 26188 33284 26240
rect 33692 26231 33744 26240
rect 33692 26197 33701 26231
rect 33701 26197 33735 26231
rect 33735 26197 33744 26231
rect 33692 26188 33744 26197
rect 4874 26086 4926 26138
rect 4938 26086 4990 26138
rect 5002 26086 5054 26138
rect 5066 26086 5118 26138
rect 5130 26086 5182 26138
rect 35594 26086 35646 26138
rect 35658 26086 35710 26138
rect 35722 26086 35774 26138
rect 35786 26086 35838 26138
rect 35850 26086 35902 26138
rect 5356 25984 5408 26036
rect 6920 25984 6972 26036
rect 14740 25984 14792 26036
rect 15568 25984 15620 26036
rect 15936 25984 15988 26036
rect 17132 25984 17184 26036
rect 19432 25984 19484 26036
rect 3884 25916 3936 25968
rect 1768 25891 1820 25900
rect 1768 25857 1777 25891
rect 1777 25857 1811 25891
rect 1811 25857 1820 25891
rect 1768 25848 1820 25857
rect 3056 25891 3108 25900
rect 3056 25857 3065 25891
rect 3065 25857 3099 25891
rect 3099 25857 3108 25891
rect 3056 25848 3108 25857
rect 3240 25848 3292 25900
rect 18328 25916 18380 25968
rect 18972 25916 19024 25968
rect 19156 25916 19208 25968
rect 10048 25848 10100 25900
rect 13820 25848 13872 25900
rect 17132 25848 17184 25900
rect 17868 25848 17920 25900
rect 18052 25848 18104 25900
rect 18696 25891 18748 25900
rect 18696 25857 18705 25891
rect 18705 25857 18739 25891
rect 18739 25857 18748 25891
rect 18696 25848 18748 25857
rect 1860 25780 1912 25832
rect 3608 25823 3660 25832
rect 3608 25789 3617 25823
rect 3617 25789 3651 25823
rect 3651 25789 3660 25823
rect 3608 25780 3660 25789
rect 8668 25823 8720 25832
rect 8668 25789 8677 25823
rect 8677 25789 8711 25823
rect 8711 25789 8720 25823
rect 8668 25780 8720 25789
rect 8944 25823 8996 25832
rect 8944 25789 8953 25823
rect 8953 25789 8987 25823
rect 8987 25789 8996 25823
rect 8944 25780 8996 25789
rect 11980 25780 12032 25832
rect 13544 25780 13596 25832
rect 14648 25780 14700 25832
rect 17408 25780 17460 25832
rect 19340 25848 19392 25900
rect 19432 25891 19484 25900
rect 19432 25857 19441 25891
rect 19441 25857 19475 25891
rect 19475 25857 19484 25891
rect 19432 25848 19484 25857
rect 20076 25984 20128 26036
rect 20812 25984 20864 26036
rect 23112 25984 23164 26036
rect 23756 25984 23808 26036
rect 25320 25984 25372 26036
rect 25872 25984 25924 26036
rect 26148 25984 26200 26036
rect 20168 25916 20220 25968
rect 20628 25959 20680 25968
rect 20628 25925 20637 25959
rect 20637 25925 20671 25959
rect 20671 25925 20680 25959
rect 20628 25916 20680 25925
rect 20904 25916 20956 25968
rect 19800 25891 19852 25900
rect 19800 25857 19809 25891
rect 19809 25857 19843 25891
rect 19843 25857 19852 25891
rect 19800 25848 19852 25857
rect 19892 25848 19944 25900
rect 20352 25848 20404 25900
rect 20076 25780 20128 25832
rect 20996 25848 21048 25900
rect 22192 25848 22244 25900
rect 22652 25891 22704 25900
rect 22652 25857 22661 25891
rect 22661 25857 22695 25891
rect 22695 25857 22704 25891
rect 22652 25848 22704 25857
rect 14832 25712 14884 25764
rect 18236 25712 18288 25764
rect 940 25644 992 25696
rect 2872 25687 2924 25696
rect 2872 25653 2881 25687
rect 2881 25653 2915 25687
rect 2915 25653 2924 25687
rect 2872 25644 2924 25653
rect 4712 25644 4764 25696
rect 9680 25644 9732 25696
rect 12992 25644 13044 25696
rect 15016 25644 15068 25696
rect 18604 25712 18656 25764
rect 19340 25712 19392 25764
rect 21180 25712 21232 25764
rect 22560 25755 22612 25764
rect 22560 25721 22569 25755
rect 22569 25721 22603 25755
rect 22603 25721 22612 25755
rect 22560 25712 22612 25721
rect 22652 25712 22704 25764
rect 23112 25891 23164 25900
rect 23112 25857 23121 25891
rect 23121 25857 23155 25891
rect 23155 25857 23164 25891
rect 23112 25848 23164 25857
rect 23388 25891 23440 25900
rect 23388 25857 23397 25891
rect 23397 25857 23431 25891
rect 23431 25857 23440 25891
rect 23388 25848 23440 25857
rect 24308 25891 24360 25900
rect 24308 25857 24317 25891
rect 24317 25857 24351 25891
rect 24351 25857 24360 25891
rect 24308 25848 24360 25857
rect 24676 25848 24728 25900
rect 24768 25891 24820 25900
rect 24768 25857 24777 25891
rect 24777 25857 24811 25891
rect 24811 25857 24820 25891
rect 24768 25848 24820 25857
rect 24032 25780 24084 25832
rect 24492 25712 24544 25764
rect 25320 25848 25372 25900
rect 25504 25891 25556 25900
rect 25504 25857 25513 25891
rect 25513 25857 25547 25891
rect 25547 25857 25556 25891
rect 25504 25848 25556 25857
rect 25688 25891 25740 25900
rect 25688 25857 25697 25891
rect 25697 25857 25731 25891
rect 25731 25857 25740 25891
rect 25688 25848 25740 25857
rect 26056 25848 26108 25900
rect 32036 25984 32088 26036
rect 32128 26027 32180 26036
rect 32128 25993 32137 26027
rect 32137 25993 32171 26027
rect 32171 25993 32180 26027
rect 32128 25984 32180 25993
rect 32680 25984 32732 26036
rect 33324 25984 33376 26036
rect 34336 25984 34388 26036
rect 34704 25984 34756 26036
rect 34980 25984 35032 26036
rect 30012 25916 30064 25968
rect 26516 25848 26568 25900
rect 27896 25848 27948 25900
rect 19156 25687 19208 25696
rect 19156 25653 19165 25687
rect 19165 25653 19199 25687
rect 19199 25653 19208 25687
rect 19156 25644 19208 25653
rect 19432 25644 19484 25696
rect 20168 25644 20220 25696
rect 20996 25687 21048 25696
rect 20996 25653 21005 25687
rect 21005 25653 21039 25687
rect 21039 25653 21048 25687
rect 20996 25644 21048 25653
rect 21088 25644 21140 25696
rect 21640 25644 21692 25696
rect 22284 25687 22336 25696
rect 22284 25653 22293 25687
rect 22293 25653 22327 25687
rect 22327 25653 22336 25687
rect 22284 25644 22336 25653
rect 23848 25687 23900 25696
rect 23848 25653 23857 25687
rect 23857 25653 23891 25687
rect 23891 25653 23900 25687
rect 23848 25644 23900 25653
rect 24308 25644 24360 25696
rect 26424 25780 26476 25832
rect 31760 25891 31812 25900
rect 31760 25857 31769 25891
rect 31769 25857 31803 25891
rect 31803 25857 31812 25891
rect 31760 25848 31812 25857
rect 31852 25780 31904 25832
rect 32680 25823 32732 25832
rect 32680 25789 32689 25823
rect 32689 25789 32723 25823
rect 32723 25789 32732 25823
rect 32680 25780 32732 25789
rect 33692 25916 33744 25968
rect 26332 25712 26384 25764
rect 25320 25687 25372 25696
rect 25320 25653 25329 25687
rect 25329 25653 25363 25687
rect 25363 25653 25372 25687
rect 25320 25644 25372 25653
rect 25504 25644 25556 25696
rect 29092 25712 29144 25764
rect 33232 25891 33284 25900
rect 33232 25857 33241 25891
rect 33241 25857 33275 25891
rect 33275 25857 33284 25891
rect 33232 25848 33284 25857
rect 34152 25823 34204 25832
rect 34152 25789 34161 25823
rect 34161 25789 34195 25823
rect 34195 25789 34204 25823
rect 34152 25780 34204 25789
rect 36636 25848 36688 25900
rect 26608 25687 26660 25696
rect 26608 25653 26617 25687
rect 26617 25653 26651 25687
rect 26651 25653 26660 25687
rect 26608 25644 26660 25653
rect 27804 25644 27856 25696
rect 28724 25644 28776 25696
rect 31300 25644 31352 25696
rect 32036 25644 32088 25696
rect 34704 25712 34756 25764
rect 34796 25644 34848 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 3608 25440 3660 25492
rect 8944 25440 8996 25492
rect 9680 25440 9732 25492
rect 12992 25440 13044 25492
rect 17224 25440 17276 25492
rect 2872 25304 2924 25356
rect 1400 25236 1452 25288
rect 1860 25279 1912 25288
rect 1860 25245 1869 25279
rect 1869 25245 1903 25279
rect 1903 25245 1912 25279
rect 1860 25236 1912 25245
rect 3240 25236 3292 25288
rect 4344 25236 4396 25288
rect 7564 25279 7616 25288
rect 7564 25245 7573 25279
rect 7573 25245 7607 25279
rect 7607 25245 7616 25279
rect 7564 25236 7616 25245
rect 8668 25236 8720 25288
rect 12072 25372 12124 25424
rect 12348 25372 12400 25424
rect 9864 25347 9916 25356
rect 9864 25313 9873 25347
rect 9873 25313 9907 25347
rect 9907 25313 9916 25347
rect 9864 25304 9916 25313
rect 18972 25372 19024 25424
rect 19892 25372 19944 25424
rect 2964 25100 3016 25152
rect 4620 25100 4672 25152
rect 7288 25100 7340 25152
rect 10140 25279 10192 25288
rect 10140 25245 10149 25279
rect 10149 25245 10183 25279
rect 10183 25245 10192 25279
rect 10140 25236 10192 25245
rect 10508 25168 10560 25220
rect 11060 25168 11112 25220
rect 11796 25168 11848 25220
rect 12624 25236 12676 25288
rect 13728 25304 13780 25356
rect 13176 25279 13228 25288
rect 13176 25245 13185 25279
rect 13185 25245 13219 25279
rect 13219 25245 13228 25279
rect 13176 25236 13228 25245
rect 13544 25236 13596 25288
rect 14832 25347 14884 25356
rect 14832 25313 14841 25347
rect 14841 25313 14875 25347
rect 14875 25313 14884 25347
rect 14832 25304 14884 25313
rect 15660 25304 15712 25356
rect 15016 25236 15068 25288
rect 15936 25279 15988 25288
rect 15936 25245 15945 25279
rect 15945 25245 15979 25279
rect 15979 25245 15988 25279
rect 15936 25236 15988 25245
rect 16028 25236 16080 25288
rect 19064 25304 19116 25356
rect 20996 25347 21048 25356
rect 20996 25313 21005 25347
rect 21005 25313 21039 25347
rect 21039 25313 21048 25347
rect 20996 25304 21048 25313
rect 9588 25100 9640 25152
rect 11980 25143 12032 25152
rect 11980 25109 11989 25143
rect 11989 25109 12023 25143
rect 12023 25109 12032 25143
rect 11980 25100 12032 25109
rect 12808 25143 12860 25152
rect 12808 25109 12817 25143
rect 12817 25109 12851 25143
rect 12851 25109 12860 25143
rect 12808 25100 12860 25109
rect 16672 25100 16724 25152
rect 16856 25100 16908 25152
rect 17316 25236 17368 25288
rect 18420 25279 18472 25288
rect 18420 25245 18429 25279
rect 18429 25245 18463 25279
rect 18463 25245 18472 25279
rect 18420 25236 18472 25245
rect 18512 25279 18564 25288
rect 18512 25245 18521 25279
rect 18521 25245 18555 25279
rect 18555 25245 18564 25279
rect 18512 25236 18564 25245
rect 19340 25236 19392 25288
rect 20260 25236 20312 25288
rect 20720 25279 20772 25288
rect 20720 25245 20729 25279
rect 20729 25245 20763 25279
rect 20763 25245 20772 25279
rect 20720 25236 20772 25245
rect 21272 25279 21324 25288
rect 21272 25245 21276 25279
rect 21276 25245 21310 25279
rect 21310 25245 21324 25279
rect 21272 25236 21324 25245
rect 21456 25279 21508 25288
rect 21456 25245 21465 25279
rect 21465 25245 21499 25279
rect 21499 25245 21508 25279
rect 21456 25236 21508 25245
rect 21548 25279 21600 25288
rect 21548 25245 21593 25279
rect 21593 25245 21600 25279
rect 21548 25236 21600 25245
rect 21824 25236 21876 25288
rect 22008 25236 22060 25288
rect 22192 25279 22244 25288
rect 22192 25245 22201 25279
rect 22201 25245 22235 25279
rect 22235 25245 22244 25279
rect 22192 25236 22244 25245
rect 19524 25168 19576 25220
rect 17500 25100 17552 25152
rect 17684 25100 17736 25152
rect 17960 25100 18012 25152
rect 19432 25100 19484 25152
rect 20628 25100 20680 25152
rect 20904 25168 20956 25220
rect 22560 25440 22612 25492
rect 24952 25440 25004 25492
rect 25136 25440 25188 25492
rect 25320 25440 25372 25492
rect 22652 25372 22704 25424
rect 22928 25304 22980 25356
rect 23664 25347 23716 25356
rect 23664 25313 23673 25347
rect 23673 25313 23707 25347
rect 23707 25313 23716 25347
rect 23664 25304 23716 25313
rect 21732 25100 21784 25152
rect 22560 25211 22612 25220
rect 22560 25177 22569 25211
rect 22569 25177 22603 25211
rect 22603 25177 22612 25211
rect 22560 25168 22612 25177
rect 24400 25236 24452 25288
rect 24768 25279 24820 25288
rect 24768 25245 24777 25279
rect 24777 25245 24811 25279
rect 24811 25245 24820 25279
rect 24768 25236 24820 25245
rect 24952 25279 25004 25288
rect 24952 25245 24961 25279
rect 24961 25245 24995 25279
rect 24995 25245 25004 25279
rect 24952 25236 25004 25245
rect 23940 25168 23992 25220
rect 26424 25236 26476 25288
rect 26976 25236 27028 25288
rect 31024 25440 31076 25492
rect 27804 25415 27856 25424
rect 27804 25381 27813 25415
rect 27813 25381 27847 25415
rect 27847 25381 27856 25415
rect 27804 25372 27856 25381
rect 30564 25372 30616 25424
rect 34704 25372 34756 25424
rect 27344 25168 27396 25220
rect 23572 25100 23624 25152
rect 27896 25236 27948 25288
rect 28724 25279 28776 25288
rect 28724 25245 28733 25279
rect 28733 25245 28767 25279
rect 28767 25245 28776 25279
rect 28724 25236 28776 25245
rect 29000 25236 29052 25288
rect 29736 25236 29788 25288
rect 27804 25168 27856 25220
rect 30288 25279 30340 25288
rect 30288 25245 30297 25279
rect 30297 25245 30331 25279
rect 30331 25245 30340 25279
rect 30288 25236 30340 25245
rect 30380 25279 30432 25288
rect 30380 25245 30389 25279
rect 30389 25245 30423 25279
rect 30423 25245 30432 25279
rect 30380 25236 30432 25245
rect 34336 25279 34388 25288
rect 34336 25245 34345 25279
rect 34345 25245 34379 25279
rect 34379 25245 34388 25279
rect 34336 25236 34388 25245
rect 28264 25100 28316 25152
rect 29092 25143 29144 25152
rect 29092 25109 29101 25143
rect 29101 25109 29135 25143
rect 29135 25109 29144 25143
rect 29092 25100 29144 25109
rect 30656 25143 30708 25152
rect 30656 25109 30665 25143
rect 30665 25109 30699 25143
rect 30699 25109 30708 25143
rect 30656 25100 30708 25109
rect 31392 25100 31444 25152
rect 35992 25168 36044 25220
rect 36728 25211 36780 25220
rect 36728 25177 36737 25211
rect 36737 25177 36771 25211
rect 36771 25177 36780 25211
rect 36728 25168 36780 25177
rect 4874 24998 4926 25050
rect 4938 24998 4990 25050
rect 5002 24998 5054 25050
rect 5066 24998 5118 25050
rect 5130 24998 5182 25050
rect 35594 24998 35646 25050
rect 35658 24998 35710 25050
rect 35722 24998 35774 25050
rect 35786 24998 35838 25050
rect 35850 24998 35902 25050
rect 4344 24939 4396 24948
rect 4344 24905 4353 24939
rect 4353 24905 4387 24939
rect 4387 24905 4396 24939
rect 4344 24896 4396 24905
rect 4712 24939 4764 24948
rect 4712 24905 4721 24939
rect 4721 24905 4755 24939
rect 4755 24905 4764 24939
rect 4712 24896 4764 24905
rect 5816 24896 5868 24948
rect 9588 24939 9640 24948
rect 9588 24905 9597 24939
rect 9597 24905 9631 24939
rect 9631 24905 9640 24939
rect 9588 24896 9640 24905
rect 10140 24896 10192 24948
rect 10508 24896 10560 24948
rect 11980 24896 12032 24948
rect 9680 24828 9732 24880
rect 10048 24828 10100 24880
rect 2964 24760 3016 24812
rect 5908 24803 5960 24812
rect 5908 24769 5917 24803
rect 5917 24769 5951 24803
rect 5951 24769 5960 24803
rect 5908 24760 5960 24769
rect 1400 24735 1452 24744
rect 1400 24701 1409 24735
rect 1409 24701 1443 24735
rect 1443 24701 1452 24735
rect 1400 24692 1452 24701
rect 1676 24735 1728 24744
rect 1676 24701 1685 24735
rect 1685 24701 1719 24735
rect 1719 24701 1728 24735
rect 1676 24692 1728 24701
rect 4804 24735 4856 24744
rect 4804 24701 4813 24735
rect 4813 24701 4847 24735
rect 4847 24701 4856 24735
rect 4804 24692 4856 24701
rect 2688 24556 2740 24608
rect 3976 24556 4028 24608
rect 7288 24735 7340 24744
rect 7288 24701 7297 24735
rect 7297 24701 7331 24735
rect 7331 24701 7340 24735
rect 7288 24692 7340 24701
rect 7932 24692 7984 24744
rect 5632 24556 5684 24608
rect 7288 24556 7340 24608
rect 10416 24803 10468 24812
rect 10416 24769 10425 24803
rect 10425 24769 10459 24803
rect 10459 24769 10468 24803
rect 10416 24760 10468 24769
rect 12440 24896 12492 24948
rect 12808 24896 12860 24948
rect 12256 24828 12308 24880
rect 13728 24896 13780 24948
rect 9220 24599 9272 24608
rect 9220 24565 9229 24599
rect 9229 24565 9263 24599
rect 9263 24565 9272 24599
rect 9220 24556 9272 24565
rect 9864 24735 9916 24744
rect 9864 24701 9873 24735
rect 9873 24701 9907 24735
rect 9907 24701 9916 24735
rect 9864 24692 9916 24701
rect 13452 24760 13504 24812
rect 14188 24760 14240 24812
rect 15016 24896 15068 24948
rect 15844 24896 15896 24948
rect 17684 24896 17736 24948
rect 18144 24896 18196 24948
rect 14924 24803 14976 24812
rect 14924 24769 14933 24803
rect 14933 24769 14967 24803
rect 14967 24769 14976 24803
rect 14924 24760 14976 24769
rect 15384 24803 15436 24812
rect 15384 24769 15393 24803
rect 15393 24769 15427 24803
rect 15427 24769 15436 24803
rect 15384 24760 15436 24769
rect 16120 24760 16172 24812
rect 16580 24760 16632 24812
rect 16856 24803 16908 24812
rect 16856 24769 16865 24803
rect 16865 24769 16899 24803
rect 16899 24769 16908 24803
rect 16856 24760 16908 24769
rect 17316 24828 17368 24880
rect 18052 24828 18104 24880
rect 18512 24871 18564 24880
rect 18512 24837 18521 24871
rect 18521 24837 18555 24871
rect 18555 24837 18564 24871
rect 18512 24828 18564 24837
rect 17592 24760 17644 24812
rect 18788 24760 18840 24812
rect 20904 24828 20956 24880
rect 19248 24760 19300 24812
rect 20076 24760 20128 24812
rect 14372 24692 14424 24744
rect 16672 24735 16724 24744
rect 16672 24701 16681 24735
rect 16681 24701 16715 24735
rect 16715 24701 16724 24735
rect 16672 24692 16724 24701
rect 17500 24692 17552 24744
rect 21456 24939 21508 24948
rect 21456 24905 21465 24939
rect 21465 24905 21499 24939
rect 21499 24905 21508 24939
rect 21456 24896 21508 24905
rect 21824 24896 21876 24948
rect 22928 24896 22980 24948
rect 23388 24939 23440 24948
rect 23388 24905 23397 24939
rect 23397 24905 23431 24939
rect 23431 24905 23440 24939
rect 23388 24896 23440 24905
rect 21180 24828 21232 24880
rect 21640 24828 21692 24880
rect 22560 24828 22612 24880
rect 24308 24828 24360 24880
rect 24492 24828 24544 24880
rect 26884 24828 26936 24880
rect 23480 24803 23532 24812
rect 23480 24769 23489 24803
rect 23489 24769 23523 24803
rect 23523 24769 23532 24803
rect 23480 24760 23532 24769
rect 23664 24760 23716 24812
rect 23848 24803 23900 24812
rect 23848 24769 23857 24803
rect 23857 24769 23891 24803
rect 23891 24769 23900 24803
rect 23848 24760 23900 24769
rect 29092 24896 29144 24948
rect 29828 24896 29880 24948
rect 31300 24896 31352 24948
rect 31392 24896 31444 24948
rect 24124 24735 24176 24744
rect 17132 24624 17184 24676
rect 17224 24624 17276 24676
rect 13176 24599 13228 24608
rect 13176 24565 13185 24599
rect 13185 24565 13219 24599
rect 13219 24565 13228 24599
rect 13176 24556 13228 24565
rect 14188 24556 14240 24608
rect 15200 24556 15252 24608
rect 17684 24624 17736 24676
rect 19892 24624 19944 24676
rect 24124 24701 24133 24735
rect 24133 24701 24167 24735
rect 24167 24701 24176 24735
rect 24124 24692 24176 24701
rect 27160 24760 27212 24812
rect 28172 24760 28224 24812
rect 28632 24803 28684 24812
rect 28632 24769 28641 24803
rect 28641 24769 28675 24803
rect 28675 24769 28684 24803
rect 28632 24760 28684 24769
rect 29460 24828 29512 24880
rect 30472 24828 30524 24880
rect 31116 24803 31168 24812
rect 31116 24769 31125 24803
rect 31125 24769 31159 24803
rect 31159 24769 31168 24803
rect 31116 24760 31168 24769
rect 34336 24896 34388 24948
rect 36728 24896 36780 24948
rect 31576 24803 31628 24812
rect 31576 24769 31585 24803
rect 31585 24769 31619 24803
rect 31619 24769 31628 24803
rect 31576 24760 31628 24769
rect 33048 24803 33100 24812
rect 33048 24769 33057 24803
rect 33057 24769 33091 24803
rect 33091 24769 33100 24803
rect 33048 24760 33100 24769
rect 33140 24760 33192 24812
rect 33784 24760 33836 24812
rect 26700 24692 26752 24744
rect 27344 24692 27396 24744
rect 23940 24624 23992 24676
rect 29276 24692 29328 24744
rect 30196 24692 30248 24744
rect 18420 24556 18472 24608
rect 18880 24556 18932 24608
rect 20812 24556 20864 24608
rect 22192 24556 22244 24608
rect 24032 24556 24084 24608
rect 25688 24556 25740 24608
rect 25964 24599 26016 24608
rect 25964 24565 25973 24599
rect 25973 24565 26007 24599
rect 26007 24565 26016 24599
rect 25964 24556 26016 24565
rect 31208 24599 31260 24608
rect 31208 24565 31217 24599
rect 31217 24565 31251 24599
rect 31251 24565 31260 24599
rect 31208 24556 31260 24565
rect 33232 24624 33284 24676
rect 33600 24624 33652 24676
rect 34152 24624 34204 24676
rect 32680 24556 32732 24608
rect 33324 24556 33376 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 1676 24352 1728 24404
rect 3056 24352 3108 24404
rect 4068 24352 4120 24404
rect 7840 24352 7892 24404
rect 7932 24395 7984 24404
rect 7932 24361 7941 24395
rect 7941 24361 7975 24395
rect 7975 24361 7984 24395
rect 7932 24352 7984 24361
rect 9220 24352 9272 24404
rect 1400 24284 1452 24336
rect 4068 24216 4120 24268
rect 6644 24284 6696 24336
rect 15384 24352 15436 24404
rect 15752 24352 15804 24404
rect 5632 24216 5684 24268
rect 4620 24148 4672 24200
rect 14924 24284 14976 24336
rect 15200 24327 15252 24336
rect 15200 24293 15209 24327
rect 15209 24293 15243 24327
rect 15243 24293 15252 24327
rect 15200 24284 15252 24293
rect 8668 24216 8720 24268
rect 12716 24216 12768 24268
rect 9128 24191 9180 24200
rect 9128 24157 9137 24191
rect 9137 24157 9171 24191
rect 9171 24157 9180 24191
rect 9128 24148 9180 24157
rect 12992 24259 13044 24268
rect 12992 24225 13001 24259
rect 13001 24225 13035 24259
rect 13035 24225 13044 24259
rect 12992 24216 13044 24225
rect 14096 24216 14148 24268
rect 14556 24216 14608 24268
rect 14372 24191 14424 24200
rect 6000 24080 6052 24132
rect 14372 24157 14381 24191
rect 14381 24157 14415 24191
rect 14415 24157 14424 24191
rect 14372 24148 14424 24157
rect 14924 24148 14976 24200
rect 15476 24216 15528 24268
rect 16396 24327 16448 24336
rect 16396 24293 16405 24327
rect 16405 24293 16439 24327
rect 16439 24293 16448 24327
rect 16396 24284 16448 24293
rect 17224 24284 17276 24336
rect 15384 24148 15436 24200
rect 2504 24012 2556 24064
rect 2688 24055 2740 24064
rect 2688 24021 2697 24055
rect 2697 24021 2731 24055
rect 2731 24021 2740 24055
rect 2688 24012 2740 24021
rect 2780 24055 2832 24064
rect 2780 24021 2789 24055
rect 2789 24021 2823 24055
rect 2823 24021 2832 24055
rect 2780 24012 2832 24021
rect 4620 24012 4672 24064
rect 9036 24055 9088 24064
rect 9036 24021 9045 24055
rect 9045 24021 9079 24055
rect 9079 24021 9088 24055
rect 9036 24012 9088 24021
rect 12624 24055 12676 24064
rect 12624 24021 12633 24055
rect 12633 24021 12667 24055
rect 12667 24021 12676 24055
rect 12624 24012 12676 24021
rect 15016 24080 15068 24132
rect 15844 24148 15896 24200
rect 16672 24148 16724 24200
rect 17224 24191 17276 24200
rect 17224 24157 17233 24191
rect 17233 24157 17267 24191
rect 17267 24157 17276 24191
rect 17224 24148 17276 24157
rect 17408 24352 17460 24404
rect 19156 24352 19208 24404
rect 20536 24352 20588 24404
rect 21456 24352 21508 24404
rect 22192 24352 22244 24404
rect 17868 24284 17920 24336
rect 17408 24216 17460 24268
rect 17684 24216 17736 24268
rect 20260 24284 20312 24336
rect 20352 24284 20404 24336
rect 21088 24284 21140 24336
rect 21364 24284 21416 24336
rect 17592 24148 17644 24200
rect 18420 24148 18472 24200
rect 18696 24191 18748 24200
rect 18696 24157 18705 24191
rect 18705 24157 18739 24191
rect 18739 24157 18748 24191
rect 18696 24148 18748 24157
rect 18880 24191 18932 24200
rect 18880 24157 18889 24191
rect 18889 24157 18923 24191
rect 18923 24157 18932 24191
rect 18880 24148 18932 24157
rect 19064 24191 19116 24200
rect 19064 24157 19073 24191
rect 19073 24157 19107 24191
rect 19107 24157 19116 24191
rect 19064 24148 19116 24157
rect 19524 24191 19576 24200
rect 19524 24157 19533 24191
rect 19533 24157 19567 24191
rect 19567 24157 19576 24191
rect 19524 24148 19576 24157
rect 20076 24216 20128 24268
rect 17960 24080 18012 24132
rect 15568 24012 15620 24064
rect 19156 24080 19208 24132
rect 22560 24216 22612 24268
rect 20720 24148 20772 24200
rect 18144 24055 18196 24064
rect 18144 24021 18153 24055
rect 18153 24021 18187 24055
rect 18187 24021 18196 24055
rect 18144 24012 18196 24021
rect 19064 24012 19116 24064
rect 19248 24055 19300 24064
rect 19248 24021 19257 24055
rect 19257 24021 19291 24055
rect 19291 24021 19300 24055
rect 19248 24012 19300 24021
rect 19892 24012 19944 24064
rect 19984 24012 20036 24064
rect 22192 24012 22244 24064
rect 23112 24216 23164 24268
rect 23664 24352 23716 24404
rect 25688 24352 25740 24404
rect 26332 24352 26384 24404
rect 27344 24395 27396 24404
rect 27344 24361 27353 24395
rect 27353 24361 27387 24395
rect 27387 24361 27396 24395
rect 27344 24352 27396 24361
rect 31208 24352 31260 24404
rect 24032 24327 24084 24336
rect 24032 24293 24041 24327
rect 24041 24293 24075 24327
rect 24075 24293 24084 24327
rect 24032 24284 24084 24293
rect 24676 24284 24728 24336
rect 23480 24148 23532 24200
rect 23756 24148 23808 24200
rect 23940 24191 23992 24200
rect 23940 24157 23949 24191
rect 23949 24157 23983 24191
rect 23983 24157 23992 24191
rect 23940 24148 23992 24157
rect 24860 24259 24912 24268
rect 24860 24225 24869 24259
rect 24869 24225 24903 24259
rect 24903 24225 24912 24259
rect 24860 24216 24912 24225
rect 26884 24284 26936 24336
rect 28724 24284 28776 24336
rect 30380 24284 30432 24336
rect 25964 24216 26016 24268
rect 26424 24216 26476 24268
rect 27160 24216 27212 24268
rect 25320 24191 25372 24200
rect 25320 24157 25329 24191
rect 25329 24157 25363 24191
rect 25363 24157 25372 24191
rect 25320 24148 25372 24157
rect 27896 24148 27948 24200
rect 28356 24148 28408 24200
rect 29552 24191 29604 24200
rect 29552 24157 29561 24191
rect 29561 24157 29595 24191
rect 29595 24157 29604 24191
rect 29552 24148 29604 24157
rect 30288 24216 30340 24268
rect 31576 24284 31628 24336
rect 29736 24191 29788 24200
rect 29736 24157 29740 24191
rect 29740 24157 29774 24191
rect 29774 24157 29788 24191
rect 29736 24148 29788 24157
rect 29828 24191 29880 24200
rect 29828 24157 29837 24191
rect 29837 24157 29871 24191
rect 29871 24157 29880 24191
rect 29828 24148 29880 24157
rect 29920 24191 29972 24200
rect 29920 24157 29929 24191
rect 29929 24157 29963 24191
rect 29963 24157 29972 24191
rect 29920 24148 29972 24157
rect 32956 24352 33008 24404
rect 33048 24327 33100 24336
rect 33048 24293 33057 24327
rect 33057 24293 33091 24327
rect 33091 24293 33100 24327
rect 33048 24284 33100 24293
rect 33508 24327 33560 24336
rect 33508 24293 33517 24327
rect 33517 24293 33551 24327
rect 33551 24293 33560 24327
rect 33508 24284 33560 24293
rect 26884 24080 26936 24132
rect 27620 24080 27672 24132
rect 32864 24191 32916 24200
rect 32864 24157 32873 24191
rect 32873 24157 32907 24191
rect 32907 24157 32916 24191
rect 32864 24148 32916 24157
rect 33140 24191 33192 24200
rect 33140 24157 33149 24191
rect 33149 24157 33183 24191
rect 33183 24157 33192 24191
rect 33140 24148 33192 24157
rect 33324 24191 33376 24200
rect 33324 24157 33333 24191
rect 33333 24157 33367 24191
rect 33367 24157 33376 24191
rect 33324 24148 33376 24157
rect 33784 24148 33836 24200
rect 29828 24012 29880 24064
rect 30196 24055 30248 24064
rect 30196 24021 30205 24055
rect 30205 24021 30239 24055
rect 30239 24021 30248 24055
rect 30196 24012 30248 24021
rect 31484 24055 31536 24064
rect 31484 24021 31493 24055
rect 31493 24021 31527 24055
rect 31527 24021 31536 24055
rect 31484 24012 31536 24021
rect 32404 24055 32456 24064
rect 32404 24021 32413 24055
rect 32413 24021 32447 24055
rect 32447 24021 32456 24055
rect 32404 24012 32456 24021
rect 32588 24055 32640 24064
rect 32588 24021 32597 24055
rect 32597 24021 32631 24055
rect 32631 24021 32640 24055
rect 32588 24012 32640 24021
rect 33140 24012 33192 24064
rect 4874 23910 4926 23962
rect 4938 23910 4990 23962
rect 5002 23910 5054 23962
rect 5066 23910 5118 23962
rect 5130 23910 5182 23962
rect 35594 23910 35646 23962
rect 35658 23910 35710 23962
rect 35722 23910 35774 23962
rect 35786 23910 35838 23962
rect 35850 23910 35902 23962
rect 1952 23808 2004 23860
rect 5908 23808 5960 23860
rect 12900 23808 12952 23860
rect 5632 23715 5684 23724
rect 5632 23681 5641 23715
rect 5641 23681 5675 23715
rect 5675 23681 5684 23715
rect 5632 23672 5684 23681
rect 6644 23672 6696 23724
rect 7012 23672 7064 23724
rect 9036 23740 9088 23792
rect 9680 23740 9732 23792
rect 13544 23740 13596 23792
rect 14280 23783 14332 23792
rect 14280 23749 14289 23783
rect 14289 23749 14323 23783
rect 14323 23749 14332 23783
rect 14280 23740 14332 23749
rect 14464 23740 14516 23792
rect 15016 23783 15068 23792
rect 15016 23749 15025 23783
rect 15025 23749 15059 23783
rect 15059 23749 15068 23783
rect 15016 23740 15068 23749
rect 4068 23604 4120 23656
rect 9312 23604 9364 23656
rect 12716 23672 12768 23724
rect 12900 23715 12952 23724
rect 12900 23681 12909 23715
rect 12909 23681 12943 23715
rect 12943 23681 12952 23715
rect 12900 23672 12952 23681
rect 13084 23715 13136 23724
rect 13084 23681 13093 23715
rect 13093 23681 13127 23715
rect 13127 23681 13136 23715
rect 13084 23672 13136 23681
rect 14188 23715 14240 23724
rect 14188 23681 14197 23715
rect 14197 23681 14231 23715
rect 14231 23681 14240 23715
rect 14188 23672 14240 23681
rect 14372 23672 14424 23724
rect 14924 23672 14976 23724
rect 15660 23808 15712 23860
rect 16028 23740 16080 23792
rect 15568 23672 15620 23724
rect 17868 23740 17920 23792
rect 18604 23808 18656 23860
rect 18696 23851 18748 23860
rect 18696 23817 18705 23851
rect 18705 23817 18739 23851
rect 18739 23817 18748 23851
rect 18696 23808 18748 23817
rect 18972 23808 19024 23860
rect 19248 23808 19300 23860
rect 19892 23851 19944 23860
rect 19892 23817 19901 23851
rect 19901 23817 19935 23851
rect 19935 23817 19944 23851
rect 19892 23808 19944 23817
rect 20168 23808 20220 23860
rect 6000 23536 6052 23588
rect 7288 23536 7340 23588
rect 5264 23468 5316 23520
rect 7472 23468 7524 23520
rect 10048 23468 10100 23520
rect 15384 23536 15436 23588
rect 16120 23604 16172 23656
rect 16672 23604 16724 23656
rect 17224 23647 17276 23656
rect 17224 23613 17233 23647
rect 17233 23613 17267 23647
rect 17267 23613 17276 23647
rect 17224 23604 17276 23613
rect 17684 23604 17736 23656
rect 19156 23715 19208 23724
rect 19156 23681 19165 23715
rect 19165 23681 19199 23715
rect 19199 23681 19208 23715
rect 19156 23672 19208 23681
rect 19432 23715 19484 23724
rect 19432 23681 19441 23715
rect 19441 23681 19475 23715
rect 19475 23681 19484 23715
rect 19432 23672 19484 23681
rect 12808 23468 12860 23520
rect 13728 23468 13780 23520
rect 15108 23511 15160 23520
rect 15108 23477 15117 23511
rect 15117 23477 15151 23511
rect 15151 23477 15160 23511
rect 15108 23468 15160 23477
rect 15936 23511 15988 23520
rect 15936 23477 15945 23511
rect 15945 23477 15979 23511
rect 15979 23477 15988 23511
rect 15936 23468 15988 23477
rect 16212 23468 16264 23520
rect 17316 23468 17368 23520
rect 17500 23468 17552 23520
rect 17868 23468 17920 23520
rect 18052 23468 18104 23520
rect 19984 23715 20036 23724
rect 19984 23681 19993 23715
rect 19993 23681 20027 23715
rect 20027 23681 20036 23715
rect 19984 23672 20036 23681
rect 20260 23715 20312 23724
rect 20260 23681 20269 23715
rect 20269 23681 20303 23715
rect 20303 23681 20312 23715
rect 20260 23672 20312 23681
rect 20720 23672 20772 23724
rect 20812 23715 20864 23724
rect 20812 23681 20821 23715
rect 20821 23681 20855 23715
rect 20855 23681 20864 23715
rect 20812 23672 20864 23681
rect 21088 23783 21140 23792
rect 21088 23749 21097 23783
rect 21097 23749 21131 23783
rect 21131 23749 21140 23783
rect 21088 23740 21140 23749
rect 22008 23672 22060 23724
rect 23112 23740 23164 23792
rect 24492 23740 24544 23792
rect 22928 23672 22980 23724
rect 23388 23672 23440 23724
rect 23756 23672 23808 23724
rect 21456 23604 21508 23656
rect 20352 23536 20404 23588
rect 22192 23579 22244 23588
rect 22192 23545 22201 23579
rect 22201 23545 22235 23579
rect 22235 23545 22244 23579
rect 23572 23604 23624 23656
rect 24124 23672 24176 23724
rect 25320 23740 25372 23792
rect 26976 23740 27028 23792
rect 28172 23808 28224 23860
rect 28632 23808 28684 23860
rect 31484 23808 31536 23860
rect 24768 23672 24820 23724
rect 25136 23715 25188 23724
rect 25136 23681 25145 23715
rect 25145 23681 25179 23715
rect 25179 23681 25188 23715
rect 25136 23672 25188 23681
rect 26056 23715 26108 23724
rect 26056 23681 26065 23715
rect 26065 23681 26099 23715
rect 26099 23681 26108 23715
rect 26056 23672 26108 23681
rect 27068 23715 27120 23724
rect 27068 23681 27077 23715
rect 27077 23681 27111 23715
rect 27111 23681 27120 23715
rect 27068 23672 27120 23681
rect 24400 23604 24452 23656
rect 22192 23536 22244 23545
rect 24308 23579 24360 23588
rect 24308 23545 24317 23579
rect 24317 23545 24351 23579
rect 24351 23545 24360 23579
rect 24308 23536 24360 23545
rect 24492 23536 24544 23588
rect 26700 23536 26752 23588
rect 19708 23468 19760 23520
rect 27436 23715 27488 23724
rect 27436 23681 27445 23715
rect 27445 23681 27479 23715
rect 27479 23681 27488 23715
rect 27436 23672 27488 23681
rect 27712 23715 27764 23724
rect 27712 23681 27721 23715
rect 27721 23681 27755 23715
rect 27755 23681 27764 23715
rect 27712 23672 27764 23681
rect 28724 23783 28776 23792
rect 28724 23749 28733 23783
rect 28733 23749 28767 23783
rect 28767 23749 28776 23783
rect 28724 23740 28776 23749
rect 32864 23808 32916 23860
rect 33140 23808 33192 23860
rect 34612 23808 34664 23860
rect 27896 23604 27948 23656
rect 35532 23715 35584 23724
rect 35532 23681 35541 23715
rect 35541 23681 35575 23715
rect 35575 23681 35584 23715
rect 35532 23672 35584 23681
rect 27528 23536 27580 23588
rect 27620 23579 27672 23588
rect 27620 23545 27629 23579
rect 27629 23545 27663 23579
rect 27663 23545 27672 23579
rect 27620 23536 27672 23545
rect 33600 23604 33652 23656
rect 34704 23604 34756 23656
rect 33048 23536 33100 23588
rect 35440 23536 35492 23588
rect 33232 23511 33284 23520
rect 33232 23477 33241 23511
rect 33241 23477 33275 23511
rect 33275 23477 33284 23511
rect 33232 23468 33284 23477
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 1768 23264 1820 23316
rect 2780 23264 2832 23316
rect 4620 23264 4672 23316
rect 4804 23264 4856 23316
rect 5632 23264 5684 23316
rect 6460 23307 6512 23316
rect 5816 23196 5868 23248
rect 6460 23273 6478 23307
rect 6478 23273 6512 23307
rect 6460 23264 6512 23273
rect 7012 23307 7064 23316
rect 7012 23273 7021 23307
rect 7021 23273 7055 23307
rect 7055 23273 7064 23307
rect 7012 23264 7064 23273
rect 7656 23264 7708 23316
rect 1952 23103 2004 23112
rect 1952 23069 1961 23103
rect 1961 23069 1995 23103
rect 1995 23069 2004 23103
rect 1952 23060 2004 23069
rect 2504 23103 2556 23112
rect 2504 23069 2513 23103
rect 2513 23069 2547 23103
rect 2547 23069 2556 23103
rect 2504 23060 2556 23069
rect 1860 22924 1912 22976
rect 2688 23103 2740 23112
rect 2688 23069 2697 23103
rect 2697 23069 2731 23103
rect 2731 23069 2740 23103
rect 2688 23060 2740 23069
rect 3056 23060 3108 23112
rect 3148 23103 3200 23112
rect 3148 23069 3157 23103
rect 3157 23069 3191 23103
rect 3191 23069 3200 23103
rect 3148 23060 3200 23069
rect 3608 23103 3660 23112
rect 3608 23069 3617 23103
rect 3617 23069 3651 23103
rect 3651 23069 3660 23103
rect 3608 23060 3660 23069
rect 4436 23103 4488 23112
rect 4436 23069 4445 23103
rect 4445 23069 4479 23103
rect 4479 23069 4488 23103
rect 4436 23060 4488 23069
rect 4896 23103 4948 23112
rect 4896 23069 4905 23103
rect 4905 23069 4939 23103
rect 4939 23069 4948 23103
rect 4896 23060 4948 23069
rect 5356 23103 5408 23112
rect 5356 23069 5365 23103
rect 5365 23069 5399 23103
rect 5399 23069 5408 23103
rect 5356 23060 5408 23069
rect 5816 23060 5868 23112
rect 6644 23128 6696 23180
rect 8024 23196 8076 23248
rect 9312 23307 9364 23316
rect 9312 23273 9321 23307
rect 9321 23273 9355 23307
rect 9355 23273 9364 23307
rect 9312 23264 9364 23273
rect 14188 23264 14240 23316
rect 20168 23264 20220 23316
rect 20720 23264 20772 23316
rect 20812 23307 20864 23316
rect 20812 23273 20821 23307
rect 20821 23273 20855 23307
rect 20855 23273 20864 23307
rect 20812 23264 20864 23273
rect 23296 23264 23348 23316
rect 26056 23264 26108 23316
rect 26332 23264 26384 23316
rect 29184 23264 29236 23316
rect 30472 23264 30524 23316
rect 35440 23264 35492 23316
rect 2872 22924 2924 22976
rect 3332 23035 3384 23044
rect 3332 23001 3341 23035
rect 3341 23001 3375 23035
rect 3375 23001 3384 23035
rect 3332 22992 3384 23001
rect 4344 22992 4396 23044
rect 4528 23035 4580 23044
rect 4528 23001 4537 23035
rect 4537 23001 4571 23035
rect 4571 23001 4580 23035
rect 4528 22992 4580 23001
rect 4620 23035 4672 23044
rect 4620 23001 4629 23035
rect 4629 23001 4663 23035
rect 4663 23001 4672 23035
rect 4620 22992 4672 23001
rect 3976 22924 4028 22976
rect 5264 23035 5316 23044
rect 5264 23001 5273 23035
rect 5273 23001 5307 23035
rect 5307 23001 5316 23035
rect 5264 22992 5316 23001
rect 9128 23128 9180 23180
rect 5724 22924 5776 22976
rect 7380 23035 7432 23044
rect 7380 23001 7389 23035
rect 7389 23001 7423 23035
rect 7423 23001 7432 23035
rect 7380 22992 7432 23001
rect 7472 23035 7524 23044
rect 7472 23001 7507 23035
rect 7507 23001 7524 23035
rect 7472 22992 7524 23001
rect 8024 22992 8076 23044
rect 9404 23060 9456 23112
rect 9680 23035 9732 23044
rect 9680 23001 9689 23035
rect 9689 23001 9723 23035
rect 9723 23001 9732 23035
rect 9680 22992 9732 23001
rect 9864 23103 9916 23112
rect 9864 23069 9873 23103
rect 9873 23069 9907 23103
rect 9907 23069 9916 23103
rect 9864 23060 9916 23069
rect 10048 23060 10100 23112
rect 12440 23128 12492 23180
rect 13912 23128 13964 23180
rect 11060 23035 11112 23044
rect 11060 23001 11069 23035
rect 11069 23001 11103 23035
rect 11103 23001 11112 23035
rect 11060 22992 11112 23001
rect 11152 22992 11204 23044
rect 11520 22992 11572 23044
rect 14280 23035 14332 23044
rect 14280 23001 14289 23035
rect 14289 23001 14323 23035
rect 14323 23001 14332 23035
rect 14280 22992 14332 23001
rect 14464 23035 14516 23044
rect 14464 23001 14473 23035
rect 14473 23001 14507 23035
rect 14507 23001 14516 23035
rect 14464 22992 14516 23001
rect 8944 22924 8996 22976
rect 19708 23196 19760 23248
rect 20076 23196 20128 23248
rect 14740 23171 14792 23180
rect 14740 23137 14749 23171
rect 14749 23137 14783 23171
rect 14783 23137 14792 23171
rect 14740 23128 14792 23137
rect 16304 23128 16356 23180
rect 15384 23103 15436 23112
rect 15384 23069 15393 23103
rect 15393 23069 15427 23103
rect 15427 23069 15436 23103
rect 15384 23060 15436 23069
rect 15292 22992 15344 23044
rect 15844 23103 15896 23112
rect 15844 23069 15853 23103
rect 15853 23069 15887 23103
rect 15887 23069 15896 23103
rect 15844 23060 15896 23069
rect 15936 23060 15988 23112
rect 17960 23128 18012 23180
rect 19984 23128 20036 23180
rect 23480 23239 23532 23248
rect 23480 23205 23489 23239
rect 23489 23205 23523 23239
rect 23523 23205 23532 23239
rect 23480 23196 23532 23205
rect 27528 23196 27580 23248
rect 22376 23128 22428 23180
rect 22468 23128 22520 23180
rect 17132 23103 17184 23112
rect 17132 23069 17141 23103
rect 17141 23069 17175 23103
rect 17175 23069 17184 23103
rect 17132 23060 17184 23069
rect 17316 23103 17368 23112
rect 17316 23069 17325 23103
rect 17325 23069 17359 23103
rect 17359 23069 17368 23103
rect 17316 23060 17368 23069
rect 17592 23060 17644 23112
rect 17684 23103 17736 23112
rect 17684 23069 17693 23103
rect 17693 23069 17727 23103
rect 17727 23069 17736 23103
rect 17684 23060 17736 23069
rect 17868 23060 17920 23112
rect 16948 22992 17000 23044
rect 17224 22992 17276 23044
rect 20352 23060 20404 23112
rect 20628 23060 20680 23112
rect 22284 23060 22336 23112
rect 19892 22992 19944 23044
rect 22652 22992 22704 23044
rect 22928 23103 22980 23112
rect 22928 23069 22937 23103
rect 22937 23069 22971 23103
rect 22971 23069 22980 23103
rect 22928 23060 22980 23069
rect 23112 23060 23164 23112
rect 23388 23103 23440 23112
rect 23388 23069 23397 23103
rect 23397 23069 23431 23103
rect 23431 23069 23440 23103
rect 23388 23060 23440 23069
rect 23572 23060 23624 23112
rect 23848 23128 23900 23180
rect 25136 23128 25188 23180
rect 16120 22924 16172 22976
rect 22008 22924 22060 22976
rect 22284 22924 22336 22976
rect 22836 22924 22888 22976
rect 24032 23060 24084 23112
rect 24400 23060 24452 23112
rect 24124 22924 24176 22976
rect 27620 23128 27672 23180
rect 35164 23196 35216 23248
rect 25688 23103 25740 23112
rect 25688 23069 25697 23103
rect 25697 23069 25731 23103
rect 25731 23069 25740 23103
rect 25688 23060 25740 23069
rect 26148 23060 26200 23112
rect 26976 23060 27028 23112
rect 29736 23103 29788 23112
rect 29736 23069 29745 23103
rect 29745 23069 29779 23103
rect 29779 23069 29788 23103
rect 29736 23060 29788 23069
rect 29920 23103 29972 23112
rect 29920 23069 29929 23103
rect 29929 23069 29963 23103
rect 29963 23069 29972 23103
rect 29920 23060 29972 23069
rect 32312 23060 32364 23112
rect 32404 23060 32456 23112
rect 32496 23103 32548 23112
rect 32496 23069 32505 23103
rect 32505 23069 32539 23103
rect 32539 23069 32548 23103
rect 32496 23060 32548 23069
rect 32772 23103 32824 23112
rect 32772 23069 32781 23103
rect 32781 23069 32815 23103
rect 32815 23069 32824 23103
rect 32772 23060 32824 23069
rect 25964 23035 26016 23044
rect 25964 23001 25973 23035
rect 25973 23001 26007 23035
rect 26007 23001 26016 23035
rect 25964 22992 26016 23001
rect 27160 22992 27212 23044
rect 30012 23035 30064 23044
rect 30012 23001 30021 23035
rect 30021 23001 30055 23035
rect 30055 23001 30064 23035
rect 30012 22992 30064 23001
rect 34612 23060 34664 23112
rect 34980 23103 35032 23112
rect 34980 23069 34989 23103
rect 34989 23069 35023 23103
rect 35023 23069 35032 23103
rect 34980 23060 35032 23069
rect 26056 22924 26108 22976
rect 26240 22967 26292 22976
rect 26240 22933 26249 22967
rect 26249 22933 26283 22967
rect 26283 22933 26292 22967
rect 26240 22924 26292 22933
rect 31852 22924 31904 22976
rect 33324 22992 33376 23044
rect 34796 22924 34848 22976
rect 34888 22924 34940 22976
rect 35256 23035 35308 23044
rect 35256 23001 35265 23035
rect 35265 23001 35299 23035
rect 35299 23001 35308 23035
rect 35256 22992 35308 23001
rect 35532 23060 35584 23112
rect 36084 23196 36136 23248
rect 35992 23128 36044 23180
rect 35440 22924 35492 22976
rect 36084 22967 36136 22976
rect 36084 22933 36093 22967
rect 36093 22933 36127 22967
rect 36127 22933 36136 22967
rect 36084 22924 36136 22933
rect 4874 22822 4926 22874
rect 4938 22822 4990 22874
rect 5002 22822 5054 22874
rect 5066 22822 5118 22874
rect 5130 22822 5182 22874
rect 35594 22822 35646 22874
rect 35658 22822 35710 22874
rect 35722 22822 35774 22874
rect 35786 22822 35838 22874
rect 35850 22822 35902 22874
rect 2688 22720 2740 22772
rect 3148 22720 3200 22772
rect 3976 22763 4028 22772
rect 3976 22729 3985 22763
rect 3985 22729 4019 22763
rect 4019 22729 4028 22763
rect 3976 22720 4028 22729
rect 4436 22720 4488 22772
rect 2504 22652 2556 22704
rect 2964 22627 3016 22636
rect 2964 22593 2973 22627
rect 2973 22593 3007 22627
rect 3007 22593 3016 22627
rect 2964 22584 3016 22593
rect 4528 22652 4580 22704
rect 4804 22652 4856 22704
rect 5632 22720 5684 22772
rect 9864 22720 9916 22772
rect 11060 22763 11112 22772
rect 11060 22729 11069 22763
rect 11069 22729 11103 22763
rect 11103 22729 11112 22763
rect 11060 22720 11112 22729
rect 12440 22720 12492 22772
rect 12532 22720 12584 22772
rect 3884 22627 3936 22636
rect 3884 22593 3893 22627
rect 3893 22593 3927 22627
rect 3927 22593 3936 22627
rect 3884 22584 3936 22593
rect 2872 22516 2924 22568
rect 3700 22516 3752 22568
rect 4712 22584 4764 22636
rect 5264 22627 5316 22636
rect 5264 22593 5273 22627
rect 5273 22593 5307 22627
rect 5307 22593 5316 22627
rect 5264 22584 5316 22593
rect 7748 22652 7800 22704
rect 6460 22584 6512 22636
rect 8024 22627 8076 22636
rect 8024 22593 8033 22627
rect 8033 22593 8067 22627
rect 8067 22593 8076 22627
rect 8024 22584 8076 22593
rect 8576 22584 8628 22636
rect 5356 22516 5408 22568
rect 7380 22516 7432 22568
rect 11428 22584 11480 22636
rect 3332 22448 3384 22500
rect 4620 22448 4672 22500
rect 8208 22491 8260 22500
rect 8208 22457 8217 22491
rect 8217 22457 8251 22491
rect 8251 22457 8260 22491
rect 8208 22448 8260 22457
rect 11980 22559 12032 22568
rect 11980 22525 11989 22559
rect 11989 22525 12023 22559
rect 12023 22525 12032 22559
rect 11980 22516 12032 22525
rect 12072 22559 12124 22568
rect 12072 22525 12081 22559
rect 12081 22525 12115 22559
rect 12115 22525 12124 22559
rect 12072 22516 12124 22525
rect 10048 22448 10100 22500
rect 11428 22448 11480 22500
rect 11612 22448 11664 22500
rect 12624 22627 12676 22636
rect 12624 22593 12633 22627
rect 12633 22593 12667 22627
rect 12667 22593 12676 22627
rect 12624 22584 12676 22593
rect 15292 22720 15344 22772
rect 15752 22720 15804 22772
rect 18512 22720 18564 22772
rect 22928 22720 22980 22772
rect 23756 22720 23808 22772
rect 25872 22720 25924 22772
rect 26240 22720 26292 22772
rect 27528 22763 27580 22772
rect 27528 22729 27537 22763
rect 27537 22729 27571 22763
rect 27571 22729 27580 22763
rect 27528 22720 27580 22729
rect 27988 22763 28040 22772
rect 27988 22729 27997 22763
rect 27997 22729 28031 22763
rect 28031 22729 28040 22763
rect 27988 22720 28040 22729
rect 29920 22720 29972 22772
rect 32496 22720 32548 22772
rect 34704 22720 34756 22772
rect 35348 22763 35400 22772
rect 35348 22729 35357 22763
rect 35357 22729 35391 22763
rect 35391 22729 35400 22763
rect 35348 22720 35400 22729
rect 35440 22720 35492 22772
rect 13544 22627 13596 22636
rect 13544 22593 13553 22627
rect 13553 22593 13587 22627
rect 13587 22593 13596 22627
rect 13544 22584 13596 22593
rect 14280 22652 14332 22704
rect 14464 22584 14516 22636
rect 14096 22448 14148 22500
rect 15200 22584 15252 22636
rect 16120 22627 16172 22636
rect 16120 22593 16129 22627
rect 16129 22593 16163 22627
rect 16163 22593 16172 22627
rect 16120 22584 16172 22593
rect 16672 22584 16724 22636
rect 16856 22584 16908 22636
rect 17132 22627 17184 22636
rect 17132 22593 17141 22627
rect 17141 22593 17175 22627
rect 17175 22593 17184 22627
rect 17132 22584 17184 22593
rect 14648 22559 14700 22568
rect 14648 22525 14657 22559
rect 14657 22525 14691 22559
rect 14691 22525 14700 22559
rect 14648 22516 14700 22525
rect 15936 22559 15988 22568
rect 15936 22525 15945 22559
rect 15945 22525 15979 22559
rect 15979 22525 15988 22559
rect 15936 22516 15988 22525
rect 16396 22516 16448 22568
rect 16948 22516 17000 22568
rect 20352 22695 20404 22704
rect 20352 22661 20361 22695
rect 20361 22661 20395 22695
rect 20395 22661 20404 22695
rect 20352 22652 20404 22661
rect 17592 22584 17644 22636
rect 20720 22627 20772 22636
rect 20720 22593 20729 22627
rect 20729 22593 20763 22627
rect 20763 22593 20772 22627
rect 20720 22584 20772 22593
rect 21916 22584 21968 22636
rect 22192 22627 22244 22636
rect 22192 22593 22201 22627
rect 22201 22593 22235 22627
rect 22235 22593 22244 22627
rect 22192 22584 22244 22593
rect 22468 22584 22520 22636
rect 22836 22584 22888 22636
rect 22928 22627 22980 22636
rect 22928 22593 22937 22627
rect 22937 22593 22971 22627
rect 22971 22593 22980 22627
rect 22928 22584 22980 22593
rect 23296 22627 23348 22636
rect 23296 22593 23305 22627
rect 23305 22593 23339 22627
rect 23339 22593 23348 22627
rect 23296 22584 23348 22593
rect 23664 22627 23716 22636
rect 23664 22593 23673 22627
rect 23673 22593 23707 22627
rect 23707 22593 23716 22627
rect 23664 22584 23716 22593
rect 24032 22627 24084 22636
rect 24032 22593 24041 22627
rect 24041 22593 24075 22627
rect 24075 22593 24084 22627
rect 24032 22584 24084 22593
rect 18144 22448 18196 22500
rect 4344 22380 4396 22432
rect 4712 22380 4764 22432
rect 5816 22380 5868 22432
rect 7656 22380 7708 22432
rect 10140 22380 10192 22432
rect 14832 22380 14884 22432
rect 15016 22380 15068 22432
rect 24124 22516 24176 22568
rect 25412 22584 25464 22636
rect 26516 22584 26568 22636
rect 26608 22584 26660 22636
rect 27160 22627 27212 22636
rect 27160 22593 27169 22627
rect 27169 22593 27203 22627
rect 27203 22593 27212 22627
rect 27160 22584 27212 22593
rect 25780 22559 25832 22568
rect 25780 22525 25789 22559
rect 25789 22525 25823 22559
rect 25823 22525 25832 22559
rect 25780 22516 25832 22525
rect 26148 22516 26200 22568
rect 26240 22516 26292 22568
rect 27344 22627 27396 22636
rect 27344 22593 27353 22627
rect 27353 22593 27387 22627
rect 27387 22593 27396 22627
rect 27344 22584 27396 22593
rect 27436 22584 27488 22636
rect 30196 22627 30248 22636
rect 30196 22593 30205 22627
rect 30205 22593 30239 22627
rect 30239 22593 30248 22627
rect 30196 22584 30248 22593
rect 32404 22652 32456 22704
rect 23940 22491 23992 22500
rect 23940 22457 23949 22491
rect 23949 22457 23983 22491
rect 23983 22457 23992 22491
rect 23940 22448 23992 22457
rect 31944 22584 31996 22636
rect 32496 22584 32548 22636
rect 35992 22652 36044 22704
rect 32864 22627 32916 22636
rect 32864 22593 32873 22627
rect 32873 22593 32907 22627
rect 32907 22593 32916 22627
rect 32864 22584 32916 22593
rect 31852 22516 31904 22568
rect 32956 22559 33008 22568
rect 32956 22525 32965 22559
rect 32965 22525 32999 22559
rect 32999 22525 33008 22559
rect 32956 22516 33008 22525
rect 24952 22380 25004 22432
rect 25412 22423 25464 22432
rect 25412 22389 25421 22423
rect 25421 22389 25455 22423
rect 25455 22389 25464 22423
rect 25412 22380 25464 22389
rect 31944 22448 31996 22500
rect 33232 22627 33284 22636
rect 33232 22593 33241 22627
rect 33241 22593 33275 22627
rect 33275 22593 33284 22627
rect 33232 22584 33284 22593
rect 33324 22584 33376 22636
rect 34428 22584 34480 22636
rect 34980 22584 35032 22636
rect 35440 22627 35492 22636
rect 35440 22593 35449 22627
rect 35449 22593 35483 22627
rect 35483 22593 35492 22627
rect 35440 22584 35492 22593
rect 37556 22584 37608 22636
rect 37832 22491 37884 22500
rect 37832 22457 37841 22491
rect 37841 22457 37875 22491
rect 37875 22457 37884 22491
rect 37832 22448 37884 22457
rect 28172 22380 28224 22432
rect 29736 22380 29788 22432
rect 30656 22423 30708 22432
rect 30656 22389 30665 22423
rect 30665 22389 30699 22423
rect 30699 22389 30708 22423
rect 30656 22380 30708 22389
rect 32036 22380 32088 22432
rect 32404 22380 32456 22432
rect 32496 22423 32548 22432
rect 32496 22389 32505 22423
rect 32505 22389 32539 22423
rect 32539 22389 32548 22423
rect 32496 22380 32548 22389
rect 34796 22380 34848 22432
rect 36084 22423 36136 22432
rect 36084 22389 36093 22423
rect 36093 22389 36127 22423
rect 36127 22389 36136 22423
rect 36084 22380 36136 22389
rect 36452 22423 36504 22432
rect 36452 22389 36461 22423
rect 36461 22389 36495 22423
rect 36495 22389 36504 22423
rect 36452 22380 36504 22389
rect 37004 22423 37056 22432
rect 37004 22389 37013 22423
rect 37013 22389 37047 22423
rect 37047 22389 37056 22423
rect 37004 22380 37056 22389
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 3608 22176 3660 22228
rect 9680 22176 9732 22228
rect 11980 22176 12032 22228
rect 3056 22108 3108 22160
rect 3424 22108 3476 22160
rect 6184 22108 6236 22160
rect 26240 22176 26292 22228
rect 27160 22176 27212 22228
rect 27712 22176 27764 22228
rect 29276 22176 29328 22228
rect 32864 22176 32916 22228
rect 3792 22040 3844 22092
rect 6276 22040 6328 22092
rect 14556 22151 14608 22160
rect 14556 22117 14565 22151
rect 14565 22117 14599 22151
rect 14599 22117 14608 22151
rect 14556 22108 14608 22117
rect 14648 22108 14700 22160
rect 16028 22108 16080 22160
rect 16304 22108 16356 22160
rect 10048 22083 10100 22092
rect 10048 22049 10057 22083
rect 10057 22049 10091 22083
rect 10091 22049 10100 22083
rect 10048 22040 10100 22049
rect 1952 22015 2004 22024
rect 1952 21981 1961 22015
rect 1961 21981 1995 22015
rect 1995 21981 2004 22015
rect 1952 21972 2004 21981
rect 3792 21947 3844 21956
rect 3792 21913 3801 21947
rect 3801 21913 3835 21947
rect 3835 21913 3844 21947
rect 3792 21904 3844 21913
rect 1768 21879 1820 21888
rect 1768 21845 1777 21879
rect 1777 21845 1811 21879
rect 1811 21845 1820 21879
rect 1768 21836 1820 21845
rect 3884 21836 3936 21888
rect 5724 21972 5776 22024
rect 5816 21972 5868 22024
rect 10416 22015 10468 22024
rect 10416 21981 10425 22015
rect 10425 21981 10459 22015
rect 10459 21981 10468 22015
rect 10416 21972 10468 21981
rect 6184 21904 6236 21956
rect 12072 22040 12124 22092
rect 15476 22040 15528 22092
rect 16764 22108 16816 22160
rect 19340 22151 19392 22160
rect 19340 22117 19349 22151
rect 19349 22117 19383 22151
rect 19383 22117 19392 22151
rect 19340 22108 19392 22117
rect 12808 22015 12860 22024
rect 12808 21981 12817 22015
rect 12817 21981 12851 22015
rect 12851 21981 12860 22015
rect 12808 21972 12860 21981
rect 13544 21972 13596 22024
rect 14556 21972 14608 22024
rect 14832 22015 14884 22024
rect 14832 21981 14841 22015
rect 14841 21981 14875 22015
rect 14875 21981 14884 22015
rect 14832 21972 14884 21981
rect 4344 21879 4396 21888
rect 4344 21845 4353 21879
rect 4353 21845 4387 21879
rect 4387 21845 4396 21879
rect 4344 21836 4396 21845
rect 7748 21836 7800 21888
rect 8208 21879 8260 21888
rect 8208 21845 8217 21879
rect 8217 21845 8251 21879
rect 8251 21845 8260 21879
rect 8208 21836 8260 21845
rect 8484 21836 8536 21888
rect 9772 21879 9824 21888
rect 9772 21845 9781 21879
rect 9781 21845 9815 21879
rect 9815 21845 9824 21879
rect 9772 21836 9824 21845
rect 9864 21879 9916 21888
rect 9864 21845 9873 21879
rect 9873 21845 9907 21879
rect 9907 21845 9916 21879
rect 9864 21836 9916 21845
rect 12440 21947 12492 21956
rect 12440 21913 12449 21947
rect 12449 21913 12483 21947
rect 12483 21913 12492 21947
rect 12440 21904 12492 21913
rect 15200 21972 15252 22024
rect 15752 22015 15804 22024
rect 15752 21981 15761 22015
rect 15761 21981 15795 22015
rect 15795 21981 15804 22015
rect 15752 21972 15804 21981
rect 15844 22015 15896 22024
rect 15844 21981 15853 22015
rect 15853 21981 15887 22015
rect 15887 21981 15896 22015
rect 15844 21972 15896 21981
rect 16396 22015 16448 22024
rect 16396 21981 16405 22015
rect 16405 21981 16439 22015
rect 16439 21981 16448 22015
rect 16396 21972 16448 21981
rect 16488 21972 16540 22024
rect 16764 21972 16816 22024
rect 16948 21972 17000 22024
rect 17040 22015 17092 22024
rect 17040 21981 17049 22015
rect 17049 21981 17083 22015
rect 17083 21981 17092 22015
rect 17040 21972 17092 21981
rect 17868 22040 17920 22092
rect 22376 22108 22428 22160
rect 23112 22108 23164 22160
rect 24032 22040 24084 22092
rect 25320 22083 25372 22092
rect 25320 22049 25329 22083
rect 25329 22049 25363 22083
rect 25363 22049 25372 22083
rect 25320 22040 25372 22049
rect 18052 21972 18104 22024
rect 19248 21972 19300 22024
rect 19708 22015 19760 22024
rect 19708 21981 19717 22015
rect 19717 21981 19751 22015
rect 19751 21981 19760 22015
rect 19708 21972 19760 21981
rect 19800 21972 19852 22024
rect 20076 22015 20128 22024
rect 20076 21981 20085 22015
rect 20085 21981 20119 22015
rect 20119 21981 20128 22015
rect 20076 21972 20128 21981
rect 22008 21972 22060 22024
rect 16212 21904 16264 21956
rect 22652 21972 22704 22024
rect 22744 22015 22796 22024
rect 22744 21981 22753 22015
rect 22753 21981 22787 22015
rect 22787 21981 22796 22015
rect 22744 21972 22796 21981
rect 23756 21972 23808 22024
rect 24584 21972 24636 22024
rect 24768 21972 24820 22024
rect 11612 21836 11664 21888
rect 11704 21879 11756 21888
rect 11704 21845 11713 21879
rect 11713 21845 11747 21879
rect 11747 21845 11756 21879
rect 11704 21836 11756 21845
rect 11796 21879 11848 21888
rect 11796 21845 11805 21879
rect 11805 21845 11839 21879
rect 11839 21845 11848 21879
rect 11796 21836 11848 21845
rect 12164 21836 12216 21888
rect 12624 21879 12676 21888
rect 12624 21845 12633 21879
rect 12633 21845 12667 21879
rect 12667 21845 12676 21879
rect 12624 21836 12676 21845
rect 15476 21836 15528 21888
rect 16028 21836 16080 21888
rect 23112 21904 23164 21956
rect 23296 21904 23348 21956
rect 22376 21836 22428 21888
rect 24676 21836 24728 21888
rect 25780 22015 25832 22026
rect 25780 21981 25789 22015
rect 25789 21981 25823 22015
rect 25823 21981 25832 22015
rect 25780 21974 25832 21981
rect 25136 21904 25188 21956
rect 26240 22015 26292 22024
rect 26240 21981 26243 22015
rect 26243 21981 26292 22015
rect 26240 21972 26292 21981
rect 28264 22108 28316 22160
rect 26608 22040 26660 22092
rect 26516 21904 26568 21956
rect 27712 22015 27764 22024
rect 27712 21981 27721 22015
rect 27721 21981 27755 22015
rect 27755 21981 27764 22015
rect 27712 21972 27764 21981
rect 26056 21836 26108 21888
rect 27528 21836 27580 21888
rect 27620 21879 27672 21888
rect 27620 21845 27629 21879
rect 27629 21845 27663 21879
rect 27663 21845 27672 21879
rect 27620 21836 27672 21845
rect 27896 21836 27948 21888
rect 28356 22015 28408 22024
rect 28356 21981 28365 22015
rect 28365 21981 28399 22015
rect 28399 21981 28408 22015
rect 28356 21972 28408 21981
rect 28172 21947 28224 21956
rect 28172 21913 28181 21947
rect 28181 21913 28215 21947
rect 28215 21913 28224 21947
rect 28172 21904 28224 21913
rect 28264 21947 28316 21956
rect 28264 21913 28273 21947
rect 28273 21913 28307 21947
rect 28307 21913 28316 21947
rect 28264 21904 28316 21913
rect 28816 22015 28868 22024
rect 28816 21981 28825 22015
rect 28825 21981 28859 22015
rect 28859 21981 28868 22015
rect 28816 21972 28868 21981
rect 30012 22040 30064 22092
rect 29828 21972 29880 22024
rect 30564 22040 30616 22092
rect 31208 22083 31260 22092
rect 31208 22049 31217 22083
rect 31217 22049 31251 22083
rect 31251 22049 31260 22083
rect 31208 22040 31260 22049
rect 31484 22040 31536 22092
rect 31116 22015 31168 22024
rect 31116 21981 31125 22015
rect 31125 21981 31159 22015
rect 31159 21981 31168 22015
rect 32404 22108 32456 22160
rect 31116 21972 31168 21981
rect 31852 22015 31904 22024
rect 31852 21981 31861 22015
rect 31861 21981 31895 22015
rect 31895 21981 31904 22015
rect 31852 21972 31904 21981
rect 32036 21972 32088 22024
rect 32864 22083 32916 22092
rect 32864 22049 32873 22083
rect 32873 22049 32907 22083
rect 32907 22049 32916 22083
rect 32864 22040 32916 22049
rect 28540 21879 28592 21888
rect 28540 21845 28549 21879
rect 28549 21845 28583 21879
rect 28583 21845 28592 21879
rect 28540 21836 28592 21845
rect 29828 21836 29880 21888
rect 32220 21836 32272 21888
rect 32680 22015 32732 22024
rect 32680 21981 32689 22015
rect 32689 21981 32723 22015
rect 32723 21981 32732 22015
rect 32680 21972 32732 21981
rect 33140 22083 33192 22092
rect 33140 22049 33149 22083
rect 33149 22049 33183 22083
rect 33183 22049 33192 22083
rect 33140 22040 33192 22049
rect 35164 22040 35216 22092
rect 35256 22083 35308 22092
rect 35256 22049 35265 22083
rect 35265 22049 35299 22083
rect 35299 22049 35308 22083
rect 35256 22040 35308 22049
rect 36268 22176 36320 22228
rect 36084 22040 36136 22092
rect 33508 21972 33560 22024
rect 34796 21972 34848 22024
rect 34428 21904 34480 21956
rect 33324 21836 33376 21888
rect 34704 21879 34756 21888
rect 34704 21845 34713 21879
rect 34713 21845 34747 21879
rect 34747 21845 34756 21879
rect 34704 21836 34756 21845
rect 36452 22040 36504 22092
rect 36912 21972 36964 22024
rect 36360 21836 36412 21888
rect 4874 21734 4926 21786
rect 4938 21734 4990 21786
rect 5002 21734 5054 21786
rect 5066 21734 5118 21786
rect 5130 21734 5182 21786
rect 35594 21734 35646 21786
rect 35658 21734 35710 21786
rect 35722 21734 35774 21786
rect 35786 21734 35838 21786
rect 35850 21734 35902 21786
rect 1768 21632 1820 21684
rect 1952 21632 2004 21684
rect 4344 21632 4396 21684
rect 4712 21632 4764 21684
rect 8852 21632 8904 21684
rect 9588 21632 9640 21684
rect 11152 21632 11204 21684
rect 14924 21675 14976 21684
rect 14924 21641 14933 21675
rect 14933 21641 14967 21675
rect 14967 21641 14976 21675
rect 14924 21632 14976 21641
rect 15108 21632 15160 21684
rect 16304 21632 16356 21684
rect 17316 21675 17368 21684
rect 17316 21641 17325 21675
rect 17325 21641 17359 21675
rect 17359 21641 17368 21675
rect 17316 21632 17368 21641
rect 17868 21632 17920 21684
rect 2780 21496 2832 21548
rect 3608 21539 3660 21548
rect 1400 21471 1452 21480
rect 1400 21437 1409 21471
rect 1409 21437 1443 21471
rect 1443 21437 1452 21471
rect 1400 21428 1452 21437
rect 3608 21505 3617 21539
rect 3617 21505 3651 21539
rect 3651 21505 3660 21539
rect 3608 21496 3660 21505
rect 5172 21607 5224 21616
rect 5172 21573 5181 21607
rect 5181 21573 5215 21607
rect 5215 21573 5224 21607
rect 5172 21564 5224 21573
rect 7288 21564 7340 21616
rect 3056 21292 3108 21344
rect 3976 21428 4028 21480
rect 4896 21496 4948 21548
rect 4528 21428 4580 21480
rect 5724 21539 5776 21548
rect 5724 21505 5733 21539
rect 5733 21505 5767 21539
rect 5767 21505 5776 21539
rect 5724 21496 5776 21505
rect 5816 21539 5868 21548
rect 5816 21505 5825 21539
rect 5825 21505 5859 21539
rect 5859 21505 5868 21539
rect 5816 21496 5868 21505
rect 4620 21360 4672 21412
rect 5264 21428 5316 21480
rect 6184 21496 6236 21548
rect 6828 21471 6880 21480
rect 6828 21437 6837 21471
rect 6837 21437 6871 21471
rect 6871 21437 6880 21471
rect 6828 21428 6880 21437
rect 9404 21539 9456 21548
rect 9404 21505 9413 21539
rect 9413 21505 9447 21539
rect 9447 21505 9456 21539
rect 9404 21496 9456 21505
rect 9588 21496 9640 21548
rect 9680 21539 9732 21548
rect 9680 21505 9689 21539
rect 9689 21505 9723 21539
rect 9723 21505 9732 21539
rect 9680 21496 9732 21505
rect 10048 21539 10100 21548
rect 10048 21505 10057 21539
rect 10057 21505 10091 21539
rect 10091 21505 10100 21539
rect 10048 21496 10100 21505
rect 10232 21496 10284 21548
rect 10324 21539 10376 21548
rect 10324 21505 10333 21539
rect 10333 21505 10367 21539
rect 10367 21505 10376 21539
rect 10324 21496 10376 21505
rect 11888 21539 11940 21548
rect 11888 21505 11897 21539
rect 11897 21505 11931 21539
rect 11931 21505 11940 21539
rect 11888 21496 11940 21505
rect 11980 21471 12032 21480
rect 11980 21437 11989 21471
rect 11989 21437 12023 21471
rect 12023 21437 12032 21471
rect 11980 21428 12032 21437
rect 12164 21471 12216 21480
rect 12164 21437 12173 21471
rect 12173 21437 12207 21471
rect 12207 21437 12216 21471
rect 12164 21428 12216 21437
rect 12808 21428 12860 21480
rect 9956 21360 10008 21412
rect 14004 21428 14056 21480
rect 13912 21360 13964 21412
rect 5356 21292 5408 21344
rect 5448 21335 5500 21344
rect 5448 21301 5457 21335
rect 5457 21301 5491 21335
rect 5491 21301 5500 21335
rect 5448 21292 5500 21301
rect 6644 21292 6696 21344
rect 7932 21292 7984 21344
rect 8208 21292 8260 21344
rect 10968 21292 11020 21344
rect 11612 21292 11664 21344
rect 14648 21428 14700 21480
rect 15292 21539 15344 21548
rect 15292 21505 15301 21539
rect 15301 21505 15335 21539
rect 15335 21505 15344 21539
rect 15292 21496 15344 21505
rect 15476 21539 15528 21548
rect 15476 21505 15484 21539
rect 15484 21505 15518 21539
rect 15518 21505 15528 21539
rect 15476 21496 15528 21505
rect 15660 21496 15712 21548
rect 16488 21496 16540 21548
rect 17132 21496 17184 21548
rect 17592 21496 17644 21548
rect 16948 21428 17000 21480
rect 18144 21564 18196 21616
rect 18880 21607 18932 21616
rect 18880 21573 18889 21607
rect 18889 21573 18923 21607
rect 18923 21573 18932 21607
rect 18880 21564 18932 21573
rect 19340 21564 19392 21616
rect 19800 21564 19852 21616
rect 19248 21496 19300 21548
rect 18144 21471 18196 21480
rect 18144 21437 18153 21471
rect 18153 21437 18187 21471
rect 18187 21437 18196 21471
rect 18144 21428 18196 21437
rect 18972 21428 19024 21480
rect 19708 21428 19760 21480
rect 20076 21564 20128 21616
rect 22192 21632 22244 21684
rect 19984 21496 20036 21548
rect 20352 21539 20404 21548
rect 20352 21505 20361 21539
rect 20361 21505 20395 21539
rect 20395 21505 20404 21539
rect 20352 21496 20404 21505
rect 20996 21496 21048 21548
rect 22928 21496 22980 21548
rect 23112 21539 23164 21548
rect 23112 21505 23121 21539
rect 23121 21505 23155 21539
rect 23155 21505 23164 21539
rect 23112 21496 23164 21505
rect 25504 21632 25556 21684
rect 25688 21632 25740 21684
rect 23572 21564 23624 21616
rect 24768 21564 24820 21616
rect 24860 21539 24912 21548
rect 24860 21505 24869 21539
rect 24869 21505 24903 21539
rect 24903 21505 24912 21539
rect 24860 21496 24912 21505
rect 25320 21564 25372 21616
rect 25504 21496 25556 21548
rect 25780 21564 25832 21616
rect 20260 21428 20312 21480
rect 22192 21428 22244 21480
rect 22744 21428 22796 21480
rect 28172 21632 28224 21684
rect 32588 21675 32640 21684
rect 32588 21641 32597 21675
rect 32597 21641 32631 21675
rect 32631 21641 32640 21675
rect 32588 21632 32640 21641
rect 34704 21632 34756 21684
rect 35164 21632 35216 21684
rect 35348 21632 35400 21684
rect 28448 21564 28500 21616
rect 29736 21607 29788 21616
rect 29736 21573 29745 21607
rect 29745 21573 29779 21607
rect 29779 21573 29788 21607
rect 29736 21564 29788 21573
rect 30104 21564 30156 21616
rect 27712 21539 27764 21548
rect 27712 21505 27721 21539
rect 27721 21505 27755 21539
rect 27755 21505 27764 21539
rect 27712 21496 27764 21505
rect 30564 21496 30616 21548
rect 31116 21496 31168 21548
rect 32220 21496 32272 21548
rect 32680 21539 32732 21548
rect 32680 21505 32689 21539
rect 32689 21505 32723 21539
rect 32723 21505 32732 21539
rect 32680 21496 32732 21505
rect 33324 21539 33376 21548
rect 33324 21505 33333 21539
rect 33333 21505 33367 21539
rect 33367 21505 33376 21539
rect 33324 21496 33376 21505
rect 33508 21539 33560 21548
rect 33508 21505 33517 21539
rect 33517 21505 33551 21539
rect 33551 21505 33560 21539
rect 33508 21496 33560 21505
rect 33600 21496 33652 21548
rect 35624 21564 35676 21616
rect 35532 21496 35584 21548
rect 36268 21539 36320 21548
rect 36268 21505 36277 21539
rect 36277 21505 36311 21539
rect 36311 21505 36320 21539
rect 36268 21496 36320 21505
rect 36360 21539 36412 21548
rect 36360 21505 36369 21539
rect 36369 21505 36403 21539
rect 36403 21505 36412 21539
rect 36360 21496 36412 21505
rect 36452 21496 36504 21548
rect 16764 21360 16816 21412
rect 27436 21360 27488 21412
rect 28816 21360 28868 21412
rect 35256 21428 35308 21480
rect 36176 21428 36228 21480
rect 37280 21428 37332 21480
rect 15384 21292 15436 21344
rect 15476 21292 15528 21344
rect 15660 21292 15712 21344
rect 16028 21292 16080 21344
rect 16120 21292 16172 21344
rect 19800 21292 19852 21344
rect 20076 21292 20128 21344
rect 23112 21335 23164 21344
rect 23112 21301 23121 21335
rect 23121 21301 23155 21335
rect 23155 21301 23164 21335
rect 23112 21292 23164 21301
rect 24860 21292 24912 21344
rect 25780 21292 25832 21344
rect 27160 21292 27212 21344
rect 29644 21292 29696 21344
rect 30932 21335 30984 21344
rect 30932 21301 30941 21335
rect 30941 21301 30975 21335
rect 30975 21301 30984 21335
rect 30932 21292 30984 21301
rect 33232 21292 33284 21344
rect 33508 21292 33560 21344
rect 35716 21292 35768 21344
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 4620 21088 4672 21140
rect 6828 21088 6880 21140
rect 9772 21088 9824 21140
rect 10140 21131 10192 21140
rect 10140 21097 10149 21131
rect 10149 21097 10183 21131
rect 10183 21097 10192 21131
rect 10140 21088 10192 21097
rect 3700 20952 3752 21004
rect 3792 20952 3844 21004
rect 4896 20952 4948 21004
rect 1860 20884 1912 20936
rect 3608 20884 3660 20936
rect 3976 20927 4028 20936
rect 3976 20893 3985 20927
rect 3985 20893 4019 20927
rect 4019 20893 4028 20927
rect 3976 20884 4028 20893
rect 5264 20859 5316 20868
rect 5264 20825 5273 20859
rect 5273 20825 5307 20859
rect 5307 20825 5316 20859
rect 5264 20816 5316 20825
rect 5632 20859 5684 20868
rect 5632 20825 5641 20859
rect 5641 20825 5675 20859
rect 5675 20825 5684 20859
rect 5632 20816 5684 20825
rect 7748 20995 7800 21004
rect 7748 20961 7757 20995
rect 7757 20961 7791 20995
rect 7791 20961 7800 20995
rect 7748 20952 7800 20961
rect 8668 20884 8720 20936
rect 9588 20927 9640 20936
rect 9588 20893 9597 20927
rect 9597 20893 9631 20927
rect 9631 20893 9640 20927
rect 9588 20884 9640 20893
rect 7932 20816 7984 20868
rect 1492 20791 1544 20800
rect 1492 20757 1501 20791
rect 1501 20757 1535 20791
rect 1535 20757 1544 20791
rect 1492 20748 1544 20757
rect 2872 20748 2924 20800
rect 4068 20748 4120 20800
rect 8208 20748 8260 20800
rect 9220 20859 9272 20868
rect 9220 20825 9229 20859
rect 9229 20825 9263 20859
rect 9263 20825 9272 20859
rect 9220 20816 9272 20825
rect 9496 20816 9548 20868
rect 9956 20927 10008 20936
rect 9956 20893 9965 20927
rect 9965 20893 9999 20927
rect 9999 20893 10008 20927
rect 9956 20884 10008 20893
rect 10140 20884 10192 20936
rect 9680 20748 9732 20800
rect 10048 20816 10100 20868
rect 10232 20816 10284 20868
rect 16764 21088 16816 21140
rect 17040 21088 17092 21140
rect 14004 21020 14056 21072
rect 14464 21020 14516 21072
rect 14372 20995 14424 21004
rect 14372 20961 14381 20995
rect 14381 20961 14415 20995
rect 14415 20961 14424 20995
rect 14372 20952 14424 20961
rect 11520 20884 11572 20936
rect 14556 20927 14608 20936
rect 14556 20893 14565 20927
rect 14565 20893 14599 20927
rect 14599 20893 14608 20927
rect 14556 20884 14608 20893
rect 14740 20927 14792 20936
rect 14740 20893 14749 20927
rect 14749 20893 14783 20927
rect 14783 20893 14792 20927
rect 14740 20884 14792 20893
rect 15108 20952 15160 21004
rect 14924 20927 14976 20936
rect 14924 20893 14933 20927
rect 14933 20893 14967 20927
rect 14967 20893 14976 20927
rect 14924 20884 14976 20893
rect 15568 21020 15620 21072
rect 15752 21020 15804 21072
rect 16672 21020 16724 21072
rect 18328 21088 18380 21140
rect 18420 21131 18472 21140
rect 18420 21097 18429 21131
rect 18429 21097 18463 21131
rect 18463 21097 18472 21131
rect 18420 21088 18472 21097
rect 17868 21020 17920 21072
rect 19984 21088 20036 21140
rect 20536 21088 20588 21140
rect 21088 21088 21140 21140
rect 21916 21088 21968 21140
rect 22008 21131 22060 21140
rect 22008 21097 22017 21131
rect 22017 21097 22051 21131
rect 22051 21097 22060 21131
rect 22008 21088 22060 21097
rect 22836 21131 22888 21140
rect 22836 21097 22845 21131
rect 22845 21097 22879 21131
rect 22879 21097 22888 21131
rect 22836 21088 22888 21097
rect 24952 21088 25004 21140
rect 25320 21088 25372 21140
rect 25688 21088 25740 21140
rect 25872 21088 25924 21140
rect 26516 21088 26568 21140
rect 27344 21088 27396 21140
rect 27528 21088 27580 21140
rect 27620 21088 27672 21140
rect 30932 21088 30984 21140
rect 33600 21088 33652 21140
rect 35256 21088 35308 21140
rect 35624 21088 35676 21140
rect 21824 21020 21876 21072
rect 14188 20816 14240 20868
rect 15108 20859 15160 20868
rect 15108 20825 15117 20859
rect 15117 20825 15151 20859
rect 15151 20825 15160 20859
rect 15108 20816 15160 20825
rect 18696 20952 18748 21004
rect 15568 20884 15620 20936
rect 15936 20884 15988 20936
rect 16120 20927 16172 20936
rect 16120 20893 16129 20927
rect 16129 20893 16163 20927
rect 16163 20893 16172 20927
rect 16120 20884 16172 20893
rect 15752 20859 15804 20868
rect 15752 20825 15761 20859
rect 15761 20825 15795 20859
rect 15795 20825 15804 20859
rect 15752 20816 15804 20825
rect 10968 20748 11020 20800
rect 12164 20748 12216 20800
rect 16212 20748 16264 20800
rect 16304 20748 16356 20800
rect 16948 20884 17000 20936
rect 17132 20927 17184 20936
rect 17132 20893 17136 20927
rect 17136 20893 17170 20927
rect 17170 20893 17184 20927
rect 17132 20884 17184 20893
rect 17960 20884 18012 20936
rect 18788 20884 18840 20936
rect 17040 20748 17092 20800
rect 17408 20816 17460 20868
rect 17868 20748 17920 20800
rect 18512 20748 18564 20800
rect 19432 20884 19484 20936
rect 19524 20927 19576 20936
rect 19524 20893 19533 20927
rect 19533 20893 19567 20927
rect 19567 20893 19576 20927
rect 19524 20884 19576 20893
rect 20904 20952 20956 21004
rect 20352 20927 20404 20936
rect 20352 20893 20361 20927
rect 20361 20893 20395 20927
rect 20395 20893 20404 20927
rect 20352 20884 20404 20893
rect 20536 20927 20588 20936
rect 20536 20893 20545 20927
rect 20545 20893 20579 20927
rect 20579 20893 20588 20927
rect 20536 20884 20588 20893
rect 21180 20952 21232 21004
rect 21364 20927 21416 20936
rect 21364 20893 21373 20927
rect 21373 20893 21407 20927
rect 21407 20893 21416 20927
rect 21364 20884 21416 20893
rect 21456 20927 21508 20936
rect 21456 20893 21466 20927
rect 21466 20893 21500 20927
rect 21500 20893 21508 20927
rect 21456 20884 21508 20893
rect 22376 21020 22428 21072
rect 24584 21020 24636 21072
rect 20812 20859 20864 20868
rect 20812 20825 20821 20859
rect 20821 20825 20855 20859
rect 20855 20825 20864 20859
rect 20812 20816 20864 20825
rect 21088 20816 21140 20868
rect 21272 20816 21324 20868
rect 20352 20748 20404 20800
rect 22192 20927 22244 20936
rect 22192 20893 22201 20927
rect 22201 20893 22235 20927
rect 22235 20893 22244 20927
rect 22192 20884 22244 20893
rect 22376 20927 22428 20936
rect 22376 20893 22385 20927
rect 22385 20893 22419 20927
rect 22419 20893 22428 20927
rect 22376 20884 22428 20893
rect 22652 20952 22704 21004
rect 23296 20952 23348 21004
rect 24676 20952 24728 21004
rect 24400 20884 24452 20936
rect 24860 20884 24912 20936
rect 27252 21020 27304 21072
rect 26700 20952 26752 21004
rect 30472 20952 30524 21004
rect 30656 20995 30708 21004
rect 30656 20961 30665 20995
rect 30665 20961 30699 20995
rect 30699 20961 30708 20995
rect 30656 20952 30708 20961
rect 21916 20816 21968 20868
rect 23112 20748 23164 20800
rect 24860 20791 24912 20800
rect 24860 20757 24869 20791
rect 24869 20757 24903 20791
rect 24903 20757 24912 20791
rect 24860 20748 24912 20757
rect 26884 20884 26936 20936
rect 27068 20927 27120 20936
rect 27068 20893 27077 20927
rect 27077 20893 27111 20927
rect 27111 20893 27120 20927
rect 27068 20884 27120 20893
rect 27344 20927 27396 20936
rect 27344 20893 27353 20927
rect 27353 20893 27387 20927
rect 27387 20893 27396 20927
rect 27344 20884 27396 20893
rect 27528 20884 27580 20936
rect 29368 20884 29420 20936
rect 30380 20927 30432 20936
rect 30380 20893 30389 20927
rect 30389 20893 30423 20927
rect 30423 20893 30432 20927
rect 30380 20884 30432 20893
rect 29828 20816 29880 20868
rect 32404 20816 32456 20868
rect 34520 20816 34572 20868
rect 27252 20748 27304 20800
rect 30104 20748 30156 20800
rect 30288 20748 30340 20800
rect 35716 21020 35768 21072
rect 35072 20927 35124 20936
rect 35072 20893 35081 20927
rect 35081 20893 35115 20927
rect 35115 20893 35124 20927
rect 35072 20884 35124 20893
rect 35256 20884 35308 20936
rect 4874 20646 4926 20698
rect 4938 20646 4990 20698
rect 5002 20646 5054 20698
rect 5066 20646 5118 20698
rect 5130 20646 5182 20698
rect 35594 20646 35646 20698
rect 35658 20646 35710 20698
rect 35722 20646 35774 20698
rect 35786 20646 35838 20698
rect 35850 20646 35902 20698
rect 38384 20680 38436 20732
rect 3148 20408 3200 20460
rect 2872 20383 2924 20392
rect 2872 20349 2881 20383
rect 2881 20349 2915 20383
rect 2915 20349 2924 20383
rect 2872 20340 2924 20349
rect 3056 20383 3108 20392
rect 3056 20349 3065 20383
rect 3065 20349 3099 20383
rect 3099 20349 3108 20383
rect 3056 20340 3108 20349
rect 3608 20408 3660 20460
rect 3884 20544 3936 20596
rect 10416 20544 10468 20596
rect 13636 20544 13688 20596
rect 14280 20544 14332 20596
rect 14556 20544 14608 20596
rect 15200 20544 15252 20596
rect 13176 20476 13228 20528
rect 3976 20408 4028 20460
rect 6552 20408 6604 20460
rect 11980 20408 12032 20460
rect 14372 20408 14424 20460
rect 14648 20519 14700 20528
rect 14648 20485 14657 20519
rect 14657 20485 14691 20519
rect 14691 20485 14700 20519
rect 14648 20476 14700 20485
rect 16028 20476 16080 20528
rect 16580 20408 16632 20460
rect 17316 20408 17368 20460
rect 18328 20476 18380 20528
rect 21088 20544 21140 20596
rect 22928 20544 22980 20596
rect 24400 20544 24452 20596
rect 7748 20383 7800 20392
rect 7748 20349 7757 20383
rect 7757 20349 7791 20383
rect 7791 20349 7800 20383
rect 7748 20340 7800 20349
rect 8392 20340 8444 20392
rect 11612 20383 11664 20392
rect 11612 20349 11621 20383
rect 11621 20349 11655 20383
rect 11655 20349 11664 20383
rect 11612 20340 11664 20349
rect 14832 20340 14884 20392
rect 15476 20383 15528 20392
rect 15476 20349 15485 20383
rect 15485 20349 15519 20383
rect 15519 20349 15528 20383
rect 15476 20340 15528 20349
rect 16304 20340 16356 20392
rect 3792 20272 3844 20324
rect 2412 20247 2464 20256
rect 2412 20213 2421 20247
rect 2421 20213 2455 20247
rect 2455 20213 2464 20247
rect 2412 20204 2464 20213
rect 3976 20204 4028 20256
rect 5080 20204 5132 20256
rect 6368 20204 6420 20256
rect 7196 20247 7248 20256
rect 7196 20213 7205 20247
rect 7205 20213 7239 20247
rect 7239 20213 7248 20247
rect 7196 20204 7248 20213
rect 10048 20272 10100 20324
rect 13912 20272 13964 20324
rect 18144 20451 18196 20460
rect 18144 20417 18153 20451
rect 18153 20417 18187 20451
rect 18187 20417 18196 20451
rect 18144 20408 18196 20417
rect 18512 20451 18564 20460
rect 18512 20417 18521 20451
rect 18521 20417 18555 20451
rect 18555 20417 18564 20451
rect 18512 20408 18564 20417
rect 19340 20408 19392 20460
rect 20076 20451 20128 20460
rect 20076 20417 20085 20451
rect 20085 20417 20119 20451
rect 20119 20417 20128 20451
rect 20076 20408 20128 20417
rect 20352 20451 20404 20460
rect 20352 20417 20361 20451
rect 20361 20417 20395 20451
rect 20395 20417 20404 20451
rect 20352 20408 20404 20417
rect 18604 20383 18656 20392
rect 18604 20349 18613 20383
rect 18613 20349 18647 20383
rect 18647 20349 18656 20383
rect 18788 20383 18840 20392
rect 18604 20340 18656 20349
rect 18788 20349 18797 20383
rect 18797 20349 18831 20383
rect 18831 20349 18840 20383
rect 18788 20340 18840 20349
rect 20628 20451 20680 20460
rect 20628 20417 20637 20451
rect 20637 20417 20671 20451
rect 20671 20417 20680 20451
rect 20628 20408 20680 20417
rect 20904 20451 20956 20460
rect 20904 20417 20913 20451
rect 20913 20417 20947 20451
rect 20947 20417 20956 20451
rect 20904 20408 20956 20417
rect 20996 20451 21048 20460
rect 20996 20417 21005 20451
rect 21005 20417 21039 20451
rect 21039 20417 21048 20451
rect 20996 20408 21048 20417
rect 24492 20476 24544 20528
rect 23756 20408 23808 20460
rect 18420 20272 18472 20324
rect 21272 20340 21324 20392
rect 24400 20451 24452 20460
rect 24400 20417 24409 20451
rect 24409 20417 24443 20451
rect 24443 20417 24452 20451
rect 24400 20408 24452 20417
rect 24860 20408 24912 20460
rect 25872 20476 25924 20528
rect 27988 20544 28040 20596
rect 35440 20587 35492 20596
rect 35440 20553 35449 20587
rect 35449 20553 35483 20587
rect 35483 20553 35492 20587
rect 35440 20544 35492 20553
rect 25228 20451 25280 20460
rect 25228 20417 25237 20451
rect 25237 20417 25271 20451
rect 25271 20417 25280 20451
rect 25228 20408 25280 20417
rect 25320 20408 25372 20460
rect 25964 20451 26016 20460
rect 25964 20417 25973 20451
rect 25973 20417 26007 20451
rect 26007 20417 26016 20451
rect 25964 20408 26016 20417
rect 19616 20272 19668 20324
rect 21456 20272 21508 20324
rect 24676 20272 24728 20324
rect 11428 20204 11480 20256
rect 11888 20204 11940 20256
rect 12164 20204 12216 20256
rect 14280 20204 14332 20256
rect 16304 20204 16356 20256
rect 18052 20204 18104 20256
rect 19432 20247 19484 20256
rect 19432 20213 19441 20247
rect 19441 20213 19475 20247
rect 19475 20213 19484 20247
rect 19432 20204 19484 20213
rect 19524 20204 19576 20256
rect 20168 20204 20220 20256
rect 23296 20204 23348 20256
rect 23940 20204 23992 20256
rect 24860 20204 24912 20256
rect 25320 20272 25372 20324
rect 26148 20451 26200 20460
rect 26148 20417 26157 20451
rect 26157 20417 26191 20451
rect 26191 20417 26200 20451
rect 26148 20408 26200 20417
rect 27068 20476 27120 20528
rect 28264 20476 28316 20528
rect 27344 20408 27396 20460
rect 27620 20451 27672 20460
rect 27620 20417 27629 20451
rect 27629 20417 27663 20451
rect 27663 20417 27672 20451
rect 27620 20408 27672 20417
rect 28540 20408 28592 20460
rect 29000 20408 29052 20460
rect 32036 20476 32088 20528
rect 34428 20476 34480 20528
rect 30380 20408 30432 20460
rect 30656 20408 30708 20460
rect 30932 20408 30984 20460
rect 31116 20408 31168 20460
rect 32588 20408 32640 20460
rect 35900 20451 35952 20460
rect 35900 20417 35909 20451
rect 35909 20417 35943 20451
rect 35943 20417 35952 20451
rect 35900 20408 35952 20417
rect 29644 20383 29696 20392
rect 29644 20349 29653 20383
rect 29653 20349 29687 20383
rect 29687 20349 29696 20383
rect 29644 20340 29696 20349
rect 26056 20272 26108 20324
rect 26240 20272 26292 20324
rect 30656 20315 30708 20324
rect 30656 20281 30665 20315
rect 30665 20281 30699 20315
rect 30699 20281 30708 20315
rect 30656 20272 30708 20281
rect 33232 20383 33284 20392
rect 33232 20349 33241 20383
rect 33241 20349 33275 20383
rect 33275 20349 33284 20383
rect 33232 20340 33284 20349
rect 34428 20340 34480 20392
rect 33140 20272 33192 20324
rect 34520 20272 34572 20324
rect 35808 20383 35860 20392
rect 35808 20349 35817 20383
rect 35817 20349 35851 20383
rect 35851 20349 35860 20383
rect 35808 20340 35860 20349
rect 25964 20204 26016 20256
rect 27160 20204 27212 20256
rect 27436 20204 27488 20256
rect 27620 20204 27672 20256
rect 29552 20204 29604 20256
rect 31208 20204 31260 20256
rect 34796 20204 34848 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 2412 20000 2464 20052
rect 2872 20000 2924 20052
rect 2964 19864 3016 19916
rect 3056 19864 3108 19916
rect 3792 19864 3844 19916
rect 7380 20000 7432 20052
rect 7932 20000 7984 20052
rect 10784 20000 10836 20052
rect 11612 20043 11664 20052
rect 11612 20009 11621 20043
rect 11621 20009 11655 20043
rect 11655 20009 11664 20043
rect 11612 20000 11664 20009
rect 12164 20043 12216 20052
rect 12164 20009 12173 20043
rect 12173 20009 12207 20043
rect 12207 20009 12216 20043
rect 12164 20000 12216 20009
rect 13912 20000 13964 20052
rect 15108 20000 15160 20052
rect 15200 20000 15252 20052
rect 15568 20000 15620 20052
rect 3884 19796 3936 19848
rect 4804 19907 4856 19916
rect 4804 19873 4813 19907
rect 4813 19873 4847 19907
rect 4847 19873 4856 19907
rect 4804 19864 4856 19873
rect 5080 19975 5132 19984
rect 5080 19941 5089 19975
rect 5089 19941 5123 19975
rect 5123 19941 5132 19975
rect 5080 19932 5132 19941
rect 5908 19796 5960 19848
rect 6552 19932 6604 19984
rect 1768 19703 1820 19712
rect 1768 19669 1777 19703
rect 1777 19669 1811 19703
rect 1811 19669 1820 19703
rect 1768 19660 1820 19669
rect 3976 19660 4028 19712
rect 4620 19728 4672 19780
rect 4988 19660 5040 19712
rect 5264 19660 5316 19712
rect 6368 19771 6420 19780
rect 6368 19737 6377 19771
rect 6377 19737 6411 19771
rect 6411 19737 6420 19771
rect 6368 19728 6420 19737
rect 7472 19864 7524 19916
rect 9680 19932 9732 19984
rect 11796 19932 11848 19984
rect 8208 19864 8260 19916
rect 6552 19839 6604 19848
rect 6552 19805 6561 19839
rect 6561 19805 6595 19839
rect 6595 19805 6604 19839
rect 6552 19796 6604 19805
rect 6644 19839 6696 19848
rect 6644 19805 6653 19839
rect 6653 19805 6687 19839
rect 6687 19805 6696 19839
rect 6644 19796 6696 19805
rect 9312 19796 9364 19848
rect 9496 19839 9548 19848
rect 9496 19805 9505 19839
rect 9505 19805 9539 19839
rect 9539 19805 9548 19839
rect 9496 19796 9548 19805
rect 9588 19839 9640 19848
rect 9588 19805 9597 19839
rect 9597 19805 9631 19839
rect 9631 19805 9640 19839
rect 9588 19796 9640 19805
rect 9956 19796 10008 19848
rect 10048 19839 10100 19848
rect 10048 19805 10057 19839
rect 10057 19805 10091 19839
rect 10091 19805 10100 19839
rect 10048 19796 10100 19805
rect 10140 19839 10192 19848
rect 10140 19805 10149 19839
rect 10149 19805 10183 19839
rect 10183 19805 10192 19839
rect 10140 19796 10192 19805
rect 12900 19975 12952 19984
rect 12900 19941 12909 19975
rect 12909 19941 12943 19975
rect 12943 19941 12952 19975
rect 12900 19932 12952 19941
rect 14740 19932 14792 19984
rect 15476 19932 15528 19984
rect 16856 20043 16908 20052
rect 16856 20009 16865 20043
rect 16865 20009 16899 20043
rect 16899 20009 16908 20043
rect 16856 20000 16908 20009
rect 17684 20000 17736 20052
rect 20812 20000 20864 20052
rect 22836 20043 22888 20052
rect 22836 20009 22845 20043
rect 22845 20009 22879 20043
rect 22879 20009 22888 20043
rect 22836 20000 22888 20009
rect 23480 20043 23532 20052
rect 23480 20009 23489 20043
rect 23489 20009 23523 20043
rect 23523 20009 23532 20043
rect 23480 20000 23532 20009
rect 23940 20043 23992 20052
rect 23940 20009 23949 20043
rect 23949 20009 23983 20043
rect 23983 20009 23992 20043
rect 23940 20000 23992 20009
rect 26240 20000 26292 20052
rect 26332 20043 26384 20052
rect 26332 20009 26341 20043
rect 26341 20009 26375 20043
rect 26375 20009 26384 20043
rect 26332 20000 26384 20009
rect 26424 20043 26476 20052
rect 26424 20009 26433 20043
rect 26433 20009 26467 20043
rect 26467 20009 26476 20043
rect 26424 20000 26476 20009
rect 30656 20000 30708 20052
rect 32036 20000 32088 20052
rect 32312 20000 32364 20052
rect 16580 19932 16632 19984
rect 18236 19932 18288 19984
rect 24400 19932 24452 19984
rect 24492 19932 24544 19984
rect 24952 19932 25004 19984
rect 25964 19932 26016 19984
rect 11428 19796 11480 19848
rect 11980 19796 12032 19848
rect 6920 19771 6972 19780
rect 6920 19737 6929 19771
rect 6929 19737 6963 19771
rect 6963 19737 6972 19771
rect 6920 19728 6972 19737
rect 8300 19728 8352 19780
rect 8392 19703 8444 19712
rect 8392 19669 8401 19703
rect 8401 19669 8435 19703
rect 8435 19669 8444 19703
rect 8392 19660 8444 19669
rect 8852 19660 8904 19712
rect 12164 19728 12216 19780
rect 12440 19796 12492 19848
rect 14004 19864 14056 19916
rect 12532 19728 12584 19780
rect 13544 19839 13596 19848
rect 13544 19805 13553 19839
rect 13553 19805 13587 19839
rect 13587 19805 13596 19839
rect 13544 19796 13596 19805
rect 13728 19796 13780 19848
rect 14280 19864 14332 19916
rect 13452 19771 13504 19780
rect 13452 19737 13461 19771
rect 13461 19737 13495 19771
rect 13495 19737 13504 19771
rect 13452 19728 13504 19737
rect 14464 19839 14516 19848
rect 14464 19805 14473 19839
rect 14473 19805 14507 19839
rect 14507 19805 14516 19839
rect 14464 19796 14516 19805
rect 15200 19839 15252 19848
rect 15200 19805 15209 19839
rect 15209 19805 15243 19839
rect 15243 19805 15252 19839
rect 15200 19796 15252 19805
rect 16028 19796 16080 19848
rect 11428 19703 11480 19712
rect 11428 19669 11437 19703
rect 11437 19669 11471 19703
rect 11471 19669 11480 19703
rect 11428 19660 11480 19669
rect 11796 19660 11848 19712
rect 13360 19660 13412 19712
rect 13544 19660 13596 19712
rect 15844 19703 15896 19712
rect 15844 19669 15853 19703
rect 15853 19669 15887 19703
rect 15887 19669 15896 19703
rect 15844 19660 15896 19669
rect 16120 19660 16172 19712
rect 16304 19839 16356 19848
rect 16304 19805 16313 19839
rect 16313 19805 16347 19839
rect 16347 19805 16356 19839
rect 16304 19796 16356 19805
rect 16488 19839 16540 19848
rect 16488 19805 16497 19839
rect 16497 19805 16531 19839
rect 16531 19805 16540 19839
rect 16488 19796 16540 19805
rect 17408 19839 17460 19848
rect 17408 19805 17417 19839
rect 17417 19805 17451 19839
rect 17451 19805 17460 19839
rect 17408 19796 17460 19805
rect 17868 19839 17920 19848
rect 17868 19805 17877 19839
rect 17877 19805 17911 19839
rect 17911 19805 17920 19839
rect 17868 19796 17920 19805
rect 16580 19728 16632 19780
rect 20076 19864 20128 19916
rect 18972 19839 19024 19848
rect 18972 19805 18981 19839
rect 18981 19805 19015 19839
rect 19015 19805 19024 19839
rect 19616 19839 19668 19848
rect 18972 19796 19024 19805
rect 19616 19805 19625 19839
rect 19625 19805 19659 19839
rect 19659 19805 19668 19839
rect 19616 19796 19668 19805
rect 18144 19660 18196 19712
rect 19340 19660 19392 19712
rect 19524 19660 19576 19712
rect 19984 19839 20036 19848
rect 19984 19805 19993 19839
rect 19993 19805 20027 19839
rect 20027 19805 20036 19839
rect 19984 19796 20036 19805
rect 20352 19796 20404 19848
rect 20628 19839 20680 19848
rect 20628 19805 20637 19839
rect 20637 19805 20671 19839
rect 20671 19805 20680 19839
rect 20628 19796 20680 19805
rect 21088 19864 21140 19916
rect 23296 19864 23348 19916
rect 23848 19907 23900 19916
rect 23848 19873 23857 19907
rect 23857 19873 23891 19907
rect 23891 19873 23900 19907
rect 23848 19864 23900 19873
rect 19800 19728 19852 19780
rect 20076 19660 20128 19712
rect 21824 19796 21876 19848
rect 22836 19771 22888 19780
rect 22836 19737 22845 19771
rect 22845 19737 22879 19771
rect 22879 19737 22888 19771
rect 22836 19728 22888 19737
rect 23112 19839 23164 19848
rect 23112 19805 23121 19839
rect 23121 19805 23155 19839
rect 23155 19805 23164 19839
rect 23112 19796 23164 19805
rect 23572 19660 23624 19712
rect 24676 19864 24728 19916
rect 24768 19839 24820 19848
rect 24768 19805 24777 19839
rect 24777 19805 24811 19839
rect 24811 19805 24820 19839
rect 24768 19796 24820 19805
rect 24676 19728 24728 19780
rect 25136 19796 25188 19848
rect 25596 19796 25648 19848
rect 25964 19796 26016 19848
rect 27160 19864 27212 19916
rect 25228 19771 25280 19780
rect 25228 19737 25237 19771
rect 25237 19737 25271 19771
rect 25271 19737 25280 19771
rect 25228 19728 25280 19737
rect 25320 19771 25372 19780
rect 25320 19737 25329 19771
rect 25329 19737 25363 19771
rect 25363 19737 25372 19771
rect 25320 19728 25372 19737
rect 26148 19728 26200 19780
rect 24492 19660 24544 19712
rect 26792 19771 26844 19780
rect 26792 19737 26801 19771
rect 26801 19737 26835 19771
rect 26835 19737 26844 19771
rect 26792 19728 26844 19737
rect 27344 19796 27396 19848
rect 28540 19864 28592 19916
rect 28908 19839 28960 19848
rect 28908 19805 28917 19839
rect 28917 19805 28951 19839
rect 28951 19805 28960 19839
rect 28908 19796 28960 19805
rect 29092 19864 29144 19916
rect 29552 19864 29604 19916
rect 29644 19796 29696 19848
rect 29828 19839 29880 19848
rect 29828 19805 29837 19839
rect 29837 19805 29871 19839
rect 29871 19805 29880 19839
rect 29828 19796 29880 19805
rect 27068 19728 27120 19780
rect 27620 19728 27672 19780
rect 29276 19728 29328 19780
rect 29552 19703 29604 19712
rect 29552 19669 29561 19703
rect 29561 19669 29595 19703
rect 29595 19669 29604 19703
rect 29552 19660 29604 19669
rect 29736 19660 29788 19712
rect 30288 19796 30340 19848
rect 30472 19728 30524 19780
rect 31208 19907 31260 19916
rect 31208 19873 31217 19907
rect 31217 19873 31251 19907
rect 31251 19873 31260 19907
rect 31208 19864 31260 19873
rect 31576 19796 31628 19848
rect 33416 19932 33468 19984
rect 33140 19864 33192 19916
rect 33048 19796 33100 19848
rect 35164 19932 35216 19984
rect 35808 20000 35860 20052
rect 36360 19932 36412 19984
rect 35716 19864 35768 19916
rect 36176 19864 36228 19916
rect 36452 19907 36504 19916
rect 36452 19873 36461 19907
rect 36461 19873 36495 19907
rect 36495 19873 36504 19907
rect 36452 19864 36504 19873
rect 34612 19728 34664 19780
rect 34704 19728 34756 19780
rect 35164 19839 35216 19848
rect 35164 19805 35173 19839
rect 35173 19805 35207 19839
rect 35207 19805 35216 19839
rect 35164 19796 35216 19805
rect 35256 19796 35308 19848
rect 35440 19839 35492 19848
rect 35440 19805 35449 19839
rect 35449 19805 35483 19839
rect 35483 19805 35492 19839
rect 35440 19796 35492 19805
rect 35992 19839 36044 19848
rect 35992 19805 36001 19839
rect 36001 19805 36035 19839
rect 36035 19805 36044 19839
rect 35992 19796 36044 19805
rect 30104 19660 30156 19712
rect 33416 19660 33468 19712
rect 34796 19660 34848 19712
rect 36084 19660 36136 19712
rect 4874 19558 4926 19610
rect 4938 19558 4990 19610
rect 5002 19558 5054 19610
rect 5066 19558 5118 19610
rect 5130 19558 5182 19610
rect 35594 19558 35646 19610
rect 35658 19558 35710 19610
rect 35722 19558 35774 19610
rect 35786 19558 35838 19610
rect 35850 19558 35902 19610
rect 1400 19456 1452 19508
rect 3516 19456 3568 19508
rect 5908 19499 5960 19508
rect 5908 19465 5917 19499
rect 5917 19465 5951 19499
rect 5951 19465 5960 19499
rect 5908 19456 5960 19465
rect 6920 19456 6972 19508
rect 7196 19456 7248 19508
rect 8116 19456 8168 19508
rect 9588 19456 9640 19508
rect 1768 19388 1820 19440
rect 2964 19388 3016 19440
rect 4712 19388 4764 19440
rect 4896 19388 4948 19440
rect 3608 19320 3660 19372
rect 8852 19388 8904 19440
rect 3148 19227 3200 19236
rect 3148 19193 3157 19227
rect 3157 19193 3191 19227
rect 3191 19193 3200 19227
rect 3148 19184 3200 19193
rect 3884 19295 3936 19304
rect 3884 19261 3893 19295
rect 3893 19261 3927 19295
rect 3927 19261 3936 19295
rect 3884 19252 3936 19261
rect 4804 19252 4856 19304
rect 4896 19252 4948 19304
rect 8760 19363 8812 19372
rect 8760 19329 8769 19363
rect 8769 19329 8803 19363
rect 8803 19329 8812 19363
rect 8760 19320 8812 19329
rect 9036 19363 9088 19372
rect 9036 19329 9045 19363
rect 9045 19329 9079 19363
rect 9079 19329 9088 19363
rect 9036 19320 9088 19329
rect 9496 19320 9548 19372
rect 11796 19456 11848 19508
rect 9956 19320 10008 19372
rect 10232 19320 10284 19372
rect 8300 19295 8352 19304
rect 8300 19261 8309 19295
rect 8309 19261 8343 19295
rect 8343 19261 8352 19295
rect 8300 19252 8352 19261
rect 9312 19252 9364 19304
rect 11520 19363 11572 19372
rect 11520 19329 11529 19363
rect 11529 19329 11563 19363
rect 11563 19329 11572 19363
rect 11520 19320 11572 19329
rect 11796 19320 11848 19372
rect 13176 19499 13228 19508
rect 13176 19465 13185 19499
rect 13185 19465 13219 19499
rect 13219 19465 13228 19499
rect 13176 19456 13228 19465
rect 14464 19456 14516 19508
rect 14740 19456 14792 19508
rect 15476 19456 15528 19508
rect 15752 19456 15804 19508
rect 15844 19456 15896 19508
rect 19984 19456 20036 19508
rect 22008 19456 22060 19508
rect 22836 19456 22888 19508
rect 22928 19456 22980 19508
rect 25136 19456 25188 19508
rect 28724 19456 28776 19508
rect 29552 19456 29604 19508
rect 29736 19456 29788 19508
rect 29828 19456 29880 19508
rect 30380 19456 30432 19508
rect 12440 19388 12492 19440
rect 14648 19388 14700 19440
rect 12532 19363 12584 19372
rect 12532 19329 12541 19363
rect 12541 19329 12575 19363
rect 12575 19329 12584 19363
rect 12532 19320 12584 19329
rect 13360 19363 13412 19372
rect 13360 19329 13369 19363
rect 13369 19329 13403 19363
rect 13403 19329 13412 19363
rect 13360 19320 13412 19329
rect 14372 19363 14424 19372
rect 14372 19329 14381 19363
rect 14381 19329 14415 19363
rect 14415 19329 14424 19363
rect 14372 19320 14424 19329
rect 14556 19363 14608 19372
rect 14556 19329 14565 19363
rect 14565 19329 14599 19363
rect 14599 19329 14608 19363
rect 14556 19320 14608 19329
rect 16120 19388 16172 19440
rect 20904 19388 20956 19440
rect 23756 19388 23808 19440
rect 24492 19388 24544 19440
rect 11888 19295 11940 19304
rect 11888 19261 11897 19295
rect 11897 19261 11931 19295
rect 11931 19261 11940 19295
rect 11888 19252 11940 19261
rect 12072 19252 12124 19304
rect 14924 19252 14976 19304
rect 16396 19252 16448 19304
rect 12348 19184 12400 19236
rect 14648 19227 14700 19236
rect 14648 19193 14657 19227
rect 14657 19193 14691 19227
rect 14691 19193 14700 19227
rect 14648 19184 14700 19193
rect 3516 19116 3568 19168
rect 11336 19159 11388 19168
rect 11336 19125 11345 19159
rect 11345 19125 11379 19159
rect 11379 19125 11388 19159
rect 11336 19116 11388 19125
rect 11888 19116 11940 19168
rect 12256 19159 12308 19168
rect 12256 19125 12265 19159
rect 12265 19125 12299 19159
rect 12299 19125 12308 19159
rect 12256 19116 12308 19125
rect 13636 19116 13688 19168
rect 16304 19116 16356 19168
rect 17408 19320 17460 19372
rect 19432 19320 19484 19372
rect 19616 19320 19668 19372
rect 18328 19252 18380 19304
rect 19340 19252 19392 19304
rect 22376 19363 22428 19372
rect 22376 19329 22385 19363
rect 22385 19329 22419 19363
rect 22419 19329 22428 19363
rect 22376 19320 22428 19329
rect 22468 19363 22520 19372
rect 22468 19329 22477 19363
rect 22477 19329 22511 19363
rect 22511 19329 22520 19363
rect 22468 19320 22520 19329
rect 22560 19320 22612 19372
rect 23480 19320 23532 19372
rect 23664 19320 23716 19372
rect 27252 19363 27304 19372
rect 27252 19329 27261 19363
rect 27261 19329 27295 19363
rect 27295 19329 27304 19363
rect 27252 19320 27304 19329
rect 27344 19320 27396 19372
rect 27528 19363 27580 19372
rect 27528 19329 27537 19363
rect 27537 19329 27571 19363
rect 27571 19329 27580 19363
rect 27528 19320 27580 19329
rect 23848 19295 23900 19304
rect 23848 19261 23857 19295
rect 23857 19261 23891 19295
rect 23891 19261 23900 19295
rect 23848 19252 23900 19261
rect 17224 19184 17276 19236
rect 25780 19184 25832 19236
rect 27804 19320 27856 19372
rect 28172 19363 28224 19372
rect 28172 19329 28181 19363
rect 28181 19329 28215 19363
rect 28215 19329 28224 19363
rect 28172 19320 28224 19329
rect 28264 19363 28316 19372
rect 28264 19329 28273 19363
rect 28273 19329 28307 19363
rect 28307 19329 28316 19363
rect 28264 19320 28316 19329
rect 29276 19363 29328 19372
rect 29276 19329 29285 19363
rect 29285 19329 29319 19363
rect 29319 19329 29328 19363
rect 29276 19320 29328 19329
rect 29460 19363 29512 19372
rect 29460 19329 29469 19363
rect 29469 19329 29503 19363
rect 29503 19329 29512 19363
rect 29460 19320 29512 19329
rect 33048 19388 33100 19440
rect 33140 19363 33192 19372
rect 33140 19329 33149 19363
rect 33149 19329 33183 19363
rect 33183 19329 33192 19363
rect 33140 19320 33192 19329
rect 30288 19252 30340 19304
rect 30472 19252 30524 19304
rect 31576 19252 31628 19304
rect 18328 19116 18380 19168
rect 19800 19116 19852 19168
rect 21732 19116 21784 19168
rect 24216 19159 24268 19168
rect 24216 19125 24225 19159
rect 24225 19125 24259 19159
rect 24259 19125 24268 19159
rect 24216 19116 24268 19125
rect 26792 19116 26844 19168
rect 29644 19159 29696 19168
rect 29644 19125 29653 19159
rect 29653 19125 29687 19159
rect 29687 19125 29696 19159
rect 29644 19116 29696 19125
rect 33140 19159 33192 19168
rect 33140 19125 33149 19159
rect 33149 19125 33183 19159
rect 33183 19125 33192 19159
rect 34152 19363 34204 19372
rect 34152 19329 34161 19363
rect 34161 19329 34195 19363
rect 34195 19329 34204 19363
rect 34152 19320 34204 19329
rect 34796 19456 34848 19508
rect 36084 19456 36136 19508
rect 34796 19295 34848 19304
rect 34796 19261 34805 19295
rect 34805 19261 34839 19295
rect 34839 19261 34848 19295
rect 34796 19252 34848 19261
rect 34428 19184 34480 19236
rect 33140 19116 33192 19125
rect 35992 19116 36044 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 4804 18912 4856 18964
rect 4068 18776 4120 18828
rect 3148 18708 3200 18760
rect 5264 18708 5316 18760
rect 17224 18912 17276 18964
rect 11152 18844 11204 18896
rect 14004 18844 14056 18896
rect 18052 18912 18104 18964
rect 18236 18912 18288 18964
rect 18420 18912 18472 18964
rect 19708 18912 19760 18964
rect 20720 18912 20772 18964
rect 21088 18912 21140 18964
rect 22100 18912 22152 18964
rect 22468 18912 22520 18964
rect 26792 18912 26844 18964
rect 32864 18912 32916 18964
rect 34428 18912 34480 18964
rect 5908 18776 5960 18828
rect 9220 18776 9272 18828
rect 9864 18776 9916 18828
rect 10876 18819 10928 18828
rect 10876 18785 10885 18819
rect 10885 18785 10919 18819
rect 10919 18785 10928 18819
rect 10876 18776 10928 18785
rect 11336 18776 11388 18828
rect 940 18640 992 18692
rect 1768 18683 1820 18692
rect 1768 18649 1777 18683
rect 1777 18649 1811 18683
rect 1811 18649 1820 18683
rect 1768 18640 1820 18649
rect 6000 18751 6052 18760
rect 6000 18717 6009 18751
rect 6009 18717 6043 18751
rect 6043 18717 6052 18751
rect 6000 18708 6052 18717
rect 1952 18572 2004 18624
rect 5632 18683 5684 18692
rect 5632 18649 5641 18683
rect 5641 18649 5675 18683
rect 5675 18649 5684 18683
rect 5632 18640 5684 18649
rect 5816 18640 5868 18692
rect 8852 18640 8904 18692
rect 11428 18708 11480 18760
rect 11796 18751 11848 18760
rect 11796 18717 11805 18751
rect 11805 18717 11839 18751
rect 11839 18717 11848 18751
rect 11796 18708 11848 18717
rect 11888 18751 11940 18760
rect 11888 18717 11897 18751
rect 11897 18717 11931 18751
rect 11931 18717 11940 18751
rect 11888 18708 11940 18717
rect 12072 18708 12124 18760
rect 15936 18776 15988 18828
rect 18512 18844 18564 18896
rect 21732 18844 21784 18896
rect 25964 18844 26016 18896
rect 15660 18708 15712 18760
rect 17132 18708 17184 18760
rect 4252 18572 4304 18624
rect 6552 18572 6604 18624
rect 10048 18572 10100 18624
rect 10324 18615 10376 18624
rect 10324 18581 10333 18615
rect 10333 18581 10367 18615
rect 10367 18581 10376 18615
rect 10324 18572 10376 18581
rect 13912 18572 13964 18624
rect 17040 18640 17092 18692
rect 17684 18751 17736 18760
rect 17684 18717 17693 18751
rect 17693 18717 17727 18751
rect 17727 18717 17736 18751
rect 17684 18708 17736 18717
rect 19340 18819 19392 18828
rect 19340 18785 19349 18819
rect 19349 18785 19383 18819
rect 19383 18785 19392 18819
rect 19340 18776 19392 18785
rect 18512 18751 18564 18760
rect 18512 18717 18521 18751
rect 18521 18717 18555 18751
rect 18555 18717 18564 18751
rect 18512 18708 18564 18717
rect 18696 18640 18748 18692
rect 18972 18708 19024 18760
rect 19432 18708 19484 18760
rect 19708 18708 19760 18760
rect 19984 18751 20036 18760
rect 19984 18717 19998 18751
rect 19998 18717 20032 18751
rect 20032 18717 20036 18751
rect 19984 18708 20036 18717
rect 20628 18776 20680 18828
rect 20076 18640 20128 18692
rect 21640 18751 21692 18760
rect 21640 18717 21649 18751
rect 21649 18717 21683 18751
rect 21683 18717 21692 18751
rect 21640 18708 21692 18717
rect 21180 18683 21232 18692
rect 21180 18649 21189 18683
rect 21189 18649 21223 18683
rect 21223 18649 21232 18683
rect 21180 18640 21232 18649
rect 23480 18776 23532 18828
rect 22376 18751 22428 18760
rect 22376 18717 22385 18751
rect 22385 18717 22419 18751
rect 22419 18717 22428 18751
rect 22376 18708 22428 18717
rect 27344 18708 27396 18760
rect 24676 18640 24728 18692
rect 25688 18640 25740 18692
rect 30748 18640 30800 18692
rect 31208 18751 31260 18760
rect 31208 18717 31217 18751
rect 31217 18717 31251 18751
rect 31251 18717 31260 18751
rect 31208 18708 31260 18717
rect 31392 18751 31444 18760
rect 31392 18717 31401 18751
rect 31401 18717 31435 18751
rect 31435 18717 31444 18751
rect 31392 18708 31444 18717
rect 33140 18776 33192 18828
rect 32680 18751 32732 18760
rect 32680 18717 32689 18751
rect 32689 18717 32723 18751
rect 32723 18717 32732 18751
rect 32680 18708 32732 18717
rect 32772 18751 32824 18760
rect 32772 18717 32781 18751
rect 32781 18717 32815 18751
rect 32815 18717 32824 18751
rect 32772 18708 32824 18717
rect 33048 18708 33100 18760
rect 33968 18708 34020 18760
rect 35348 18776 35400 18828
rect 36728 18819 36780 18828
rect 36728 18785 36737 18819
rect 36737 18785 36771 18819
rect 36771 18785 36780 18819
rect 36728 18776 36780 18785
rect 36820 18640 36872 18692
rect 14188 18615 14240 18624
rect 14188 18581 14197 18615
rect 14197 18581 14231 18615
rect 14231 18581 14240 18615
rect 14188 18572 14240 18581
rect 16212 18572 16264 18624
rect 18052 18615 18104 18624
rect 18052 18581 18061 18615
rect 18061 18581 18095 18615
rect 18095 18581 18104 18615
rect 18052 18572 18104 18581
rect 18788 18572 18840 18624
rect 20352 18572 20404 18624
rect 20628 18572 20680 18624
rect 22192 18615 22244 18624
rect 22192 18581 22201 18615
rect 22201 18581 22235 18615
rect 22235 18581 22244 18615
rect 22192 18572 22244 18581
rect 25136 18572 25188 18624
rect 25964 18572 26016 18624
rect 28356 18572 28408 18624
rect 30932 18572 30984 18624
rect 31208 18615 31260 18624
rect 31208 18581 31217 18615
rect 31217 18581 31251 18615
rect 31251 18581 31260 18615
rect 31208 18572 31260 18581
rect 32312 18572 32364 18624
rect 33048 18572 33100 18624
rect 33140 18572 33192 18624
rect 34796 18615 34848 18624
rect 34796 18581 34811 18615
rect 34811 18581 34845 18615
rect 34845 18581 34848 18615
rect 34796 18572 34848 18581
rect 34980 18572 35032 18624
rect 35164 18572 35216 18624
rect 37096 18615 37148 18624
rect 37096 18581 37105 18615
rect 37105 18581 37139 18615
rect 37139 18581 37148 18615
rect 37096 18572 37148 18581
rect 4874 18470 4926 18522
rect 4938 18470 4990 18522
rect 5002 18470 5054 18522
rect 5066 18470 5118 18522
rect 5130 18470 5182 18522
rect 35594 18470 35646 18522
rect 35658 18470 35710 18522
rect 35722 18470 35774 18522
rect 35786 18470 35838 18522
rect 35850 18470 35902 18522
rect 4252 18368 4304 18420
rect 8300 18300 8352 18352
rect 10232 18300 10284 18352
rect 1676 18207 1728 18216
rect 1676 18173 1685 18207
rect 1685 18173 1719 18207
rect 1719 18173 1728 18207
rect 1676 18164 1728 18173
rect 6552 18232 6604 18284
rect 4068 18164 4120 18216
rect 5908 18207 5960 18216
rect 5908 18173 5917 18207
rect 5917 18173 5951 18207
rect 5951 18173 5960 18207
rect 5908 18164 5960 18173
rect 3424 18096 3476 18148
rect 3700 18096 3752 18148
rect 6644 18164 6696 18216
rect 2044 18071 2096 18080
rect 2044 18037 2053 18071
rect 2053 18037 2087 18071
rect 2087 18037 2096 18071
rect 2044 18028 2096 18037
rect 2504 18071 2556 18080
rect 2504 18037 2513 18071
rect 2513 18037 2547 18071
rect 2547 18037 2556 18071
rect 2504 18028 2556 18037
rect 2964 18028 3016 18080
rect 3516 18028 3568 18080
rect 6184 18028 6236 18080
rect 7932 18164 7984 18216
rect 9036 18164 9088 18216
rect 13820 18368 13872 18420
rect 13912 18411 13964 18420
rect 13912 18377 13921 18411
rect 13921 18377 13955 18411
rect 13955 18377 13964 18411
rect 13912 18368 13964 18377
rect 14188 18368 14240 18420
rect 15384 18411 15436 18420
rect 15384 18377 15393 18411
rect 15393 18377 15427 18411
rect 15427 18377 15436 18411
rect 15384 18368 15436 18377
rect 18512 18368 18564 18420
rect 12256 18300 12308 18352
rect 11336 18232 11388 18284
rect 11428 18164 11480 18216
rect 12072 18164 12124 18216
rect 11152 18096 11204 18148
rect 12532 18275 12584 18284
rect 12532 18241 12541 18275
rect 12541 18241 12575 18275
rect 12575 18241 12584 18275
rect 12532 18232 12584 18241
rect 13820 18232 13872 18284
rect 14280 18275 14332 18284
rect 14280 18241 14289 18275
rect 14289 18241 14323 18275
rect 14323 18241 14332 18275
rect 14280 18232 14332 18241
rect 15108 18300 15160 18352
rect 19708 18368 19760 18420
rect 20168 18368 20220 18420
rect 30748 18368 30800 18420
rect 16120 18232 16172 18284
rect 16488 18232 16540 18284
rect 16764 18275 16816 18284
rect 16764 18241 16773 18275
rect 16773 18241 16807 18275
rect 16807 18241 16816 18275
rect 16764 18232 16816 18241
rect 16948 18232 17000 18284
rect 18236 18232 18288 18284
rect 18880 18275 18932 18284
rect 18880 18241 18889 18275
rect 18889 18241 18923 18275
rect 18923 18241 18932 18275
rect 18880 18232 18932 18241
rect 22652 18300 22704 18352
rect 25228 18343 25280 18352
rect 25228 18309 25237 18343
rect 25237 18309 25271 18343
rect 25271 18309 25280 18343
rect 25228 18300 25280 18309
rect 27620 18300 27672 18352
rect 15384 18164 15436 18216
rect 15752 18164 15804 18216
rect 15936 18164 15988 18216
rect 19800 18232 19852 18284
rect 19984 18232 20036 18284
rect 20536 18232 20588 18284
rect 22376 18232 22428 18284
rect 22468 18275 22520 18284
rect 22468 18241 22477 18275
rect 22477 18241 22511 18275
rect 22511 18241 22520 18275
rect 22468 18232 22520 18241
rect 22560 18232 22612 18284
rect 23572 18232 23624 18284
rect 24952 18232 25004 18284
rect 25044 18275 25096 18284
rect 25044 18241 25053 18275
rect 25053 18241 25087 18275
rect 25087 18241 25096 18275
rect 25044 18232 25096 18241
rect 23664 18164 23716 18216
rect 19432 18139 19484 18148
rect 19432 18105 19441 18139
rect 19441 18105 19475 18139
rect 19475 18105 19484 18139
rect 19432 18096 19484 18105
rect 8944 18028 8996 18080
rect 10508 18028 10560 18080
rect 11060 18028 11112 18080
rect 11520 18028 11572 18080
rect 12072 18028 12124 18080
rect 12716 18028 12768 18080
rect 14188 18028 14240 18080
rect 17960 18028 18012 18080
rect 18512 18028 18564 18080
rect 18604 18028 18656 18080
rect 19984 18028 20036 18080
rect 20260 18028 20312 18080
rect 20352 18028 20404 18080
rect 20444 18028 20496 18080
rect 21548 18028 21600 18080
rect 23848 18096 23900 18148
rect 25596 18232 25648 18284
rect 25964 18232 26016 18284
rect 27988 18275 28040 18284
rect 27988 18241 27997 18275
rect 27997 18241 28031 18275
rect 28031 18241 28040 18275
rect 27988 18232 28040 18241
rect 28632 18232 28684 18284
rect 29368 18232 29420 18284
rect 29552 18275 29604 18284
rect 29552 18241 29561 18275
rect 29561 18241 29595 18275
rect 29595 18241 29604 18275
rect 29552 18232 29604 18241
rect 25780 18207 25832 18216
rect 25780 18173 25789 18207
rect 25789 18173 25823 18207
rect 25823 18173 25832 18207
rect 25780 18164 25832 18173
rect 26240 18139 26292 18148
rect 26240 18105 26249 18139
rect 26249 18105 26283 18139
rect 26283 18105 26292 18139
rect 26240 18096 26292 18105
rect 28448 18096 28500 18148
rect 30288 18232 30340 18284
rect 30380 18275 30432 18284
rect 30380 18241 30389 18275
rect 30389 18241 30423 18275
rect 30423 18241 30432 18275
rect 30380 18232 30432 18241
rect 30840 18300 30892 18352
rect 31208 18368 31260 18420
rect 34152 18368 34204 18420
rect 34796 18368 34848 18420
rect 37096 18368 37148 18420
rect 31300 18232 31352 18284
rect 32680 18300 32732 18352
rect 33140 18343 33192 18352
rect 33140 18309 33149 18343
rect 33149 18309 33183 18343
rect 33183 18309 33192 18343
rect 33140 18300 33192 18309
rect 32772 18232 32824 18284
rect 30472 18207 30524 18216
rect 30472 18173 30481 18207
rect 30481 18173 30515 18207
rect 30515 18173 30524 18207
rect 30472 18164 30524 18173
rect 31116 18164 31168 18216
rect 31944 18164 31996 18216
rect 32496 18207 32548 18216
rect 32496 18173 32505 18207
rect 32505 18173 32539 18207
rect 32539 18173 32548 18207
rect 32496 18164 32548 18173
rect 32588 18207 32640 18216
rect 32588 18173 32597 18207
rect 32597 18173 32631 18207
rect 32631 18173 32640 18207
rect 32588 18164 32640 18173
rect 26516 18028 26568 18080
rect 27896 18028 27948 18080
rect 29460 18028 29512 18080
rect 31484 18096 31536 18148
rect 34980 18275 35032 18284
rect 34980 18241 34989 18275
rect 34989 18241 35023 18275
rect 35023 18241 35032 18275
rect 34980 18232 35032 18241
rect 35440 18300 35492 18352
rect 35164 18275 35216 18284
rect 35164 18241 35173 18275
rect 35173 18241 35207 18275
rect 35207 18241 35216 18275
rect 35164 18232 35216 18241
rect 37280 18300 37332 18352
rect 32036 18028 32088 18080
rect 33968 18028 34020 18080
rect 37556 18028 37608 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 38384 17960 38436 18012
rect 1768 17824 1820 17876
rect 2136 17824 2188 17876
rect 1676 17688 1728 17740
rect 1952 17620 2004 17672
rect 2044 17620 2096 17672
rect 5632 17824 5684 17876
rect 6920 17824 6972 17876
rect 7656 17824 7708 17876
rect 7932 17824 7984 17876
rect 8300 17756 8352 17808
rect 3516 17688 3568 17740
rect 9772 17824 9824 17876
rect 11428 17824 11480 17876
rect 12440 17867 12492 17876
rect 12440 17833 12449 17867
rect 12449 17833 12483 17867
rect 12483 17833 12492 17867
rect 12440 17824 12492 17833
rect 12532 17824 12584 17876
rect 13360 17824 13412 17876
rect 15292 17867 15344 17876
rect 15292 17833 15301 17867
rect 15301 17833 15335 17867
rect 15335 17833 15344 17867
rect 15292 17824 15344 17833
rect 17684 17867 17736 17876
rect 17684 17833 17693 17867
rect 17693 17833 17727 17867
rect 17727 17833 17736 17867
rect 17684 17824 17736 17833
rect 1952 17527 2004 17536
rect 1952 17493 1961 17527
rect 1961 17493 1995 17527
rect 1995 17493 2004 17527
rect 1952 17484 2004 17493
rect 3424 17663 3476 17672
rect 3424 17629 3433 17663
rect 3433 17629 3467 17663
rect 3467 17629 3476 17663
rect 3424 17620 3476 17629
rect 3700 17620 3752 17672
rect 4252 17595 4304 17604
rect 4252 17561 4261 17595
rect 4261 17561 4295 17595
rect 4295 17561 4304 17595
rect 4252 17552 4304 17561
rect 4712 17552 4764 17604
rect 12716 17756 12768 17808
rect 12900 17756 12952 17808
rect 14188 17756 14240 17808
rect 9036 17688 9088 17740
rect 6368 17595 6420 17604
rect 6368 17561 6377 17595
rect 6377 17561 6411 17595
rect 6411 17561 6420 17595
rect 6368 17552 6420 17561
rect 6920 17552 6972 17604
rect 10048 17731 10100 17740
rect 10048 17697 10057 17731
rect 10057 17697 10091 17731
rect 10091 17697 10100 17731
rect 10048 17688 10100 17697
rect 11152 17688 11204 17740
rect 10324 17620 10376 17672
rect 10508 17620 10560 17672
rect 11060 17663 11112 17672
rect 11060 17629 11069 17663
rect 11069 17629 11103 17663
rect 11103 17629 11112 17663
rect 11060 17620 11112 17629
rect 11704 17688 11756 17740
rect 11612 17620 11664 17672
rect 12256 17688 12308 17740
rect 10876 17552 10928 17604
rect 11704 17595 11756 17604
rect 11704 17561 11713 17595
rect 11713 17561 11747 17595
rect 11747 17561 11756 17595
rect 11704 17552 11756 17561
rect 11980 17552 12032 17604
rect 5724 17527 5776 17536
rect 5724 17493 5733 17527
rect 5733 17493 5767 17527
rect 5767 17493 5776 17527
rect 5724 17484 5776 17493
rect 6184 17484 6236 17536
rect 7748 17484 7800 17536
rect 9588 17484 9640 17536
rect 12348 17620 12400 17672
rect 12716 17663 12768 17672
rect 12716 17629 12725 17663
rect 12725 17629 12759 17663
rect 12759 17629 12768 17663
rect 12716 17620 12768 17629
rect 14096 17688 14148 17740
rect 14832 17688 14884 17740
rect 16212 17688 16264 17740
rect 20812 17824 20864 17876
rect 21640 17824 21692 17876
rect 22100 17824 22152 17876
rect 13728 17484 13780 17536
rect 14004 17484 14056 17536
rect 14188 17620 14240 17672
rect 15844 17663 15896 17672
rect 15844 17629 15853 17663
rect 15853 17629 15887 17663
rect 15887 17629 15896 17663
rect 15844 17620 15896 17629
rect 16028 17620 16080 17672
rect 16396 17663 16448 17672
rect 16396 17629 16405 17663
rect 16405 17629 16439 17663
rect 16439 17629 16448 17663
rect 16396 17620 16448 17629
rect 16488 17663 16540 17672
rect 16488 17629 16497 17663
rect 16497 17629 16531 17663
rect 16531 17629 16540 17663
rect 16488 17620 16540 17629
rect 16580 17620 16632 17672
rect 17224 17620 17276 17672
rect 17316 17620 17368 17672
rect 14372 17552 14424 17604
rect 16212 17552 16264 17604
rect 17040 17552 17092 17604
rect 17960 17620 18012 17672
rect 18052 17663 18104 17672
rect 18052 17629 18061 17663
rect 18061 17629 18095 17663
rect 18095 17629 18104 17663
rect 18052 17620 18104 17629
rect 18144 17663 18196 17672
rect 18144 17629 18153 17663
rect 18153 17629 18187 17663
rect 18187 17629 18196 17663
rect 18144 17620 18196 17629
rect 18604 17756 18656 17808
rect 19156 17756 19208 17808
rect 18696 17688 18748 17740
rect 20260 17688 20312 17740
rect 20628 17688 20680 17740
rect 18788 17663 18840 17672
rect 18788 17629 18797 17663
rect 18797 17629 18831 17663
rect 18831 17629 18840 17663
rect 18788 17620 18840 17629
rect 19524 17620 19576 17672
rect 20076 17620 20128 17672
rect 20168 17620 20220 17672
rect 21180 17620 21232 17672
rect 14280 17484 14332 17536
rect 16396 17484 16448 17536
rect 16488 17484 16540 17536
rect 17500 17484 17552 17536
rect 19248 17552 19300 17604
rect 19800 17552 19852 17604
rect 22652 17824 22704 17876
rect 23204 17824 23256 17876
rect 26240 17824 26292 17876
rect 26884 17824 26936 17876
rect 22468 17663 22520 17672
rect 22468 17629 22477 17663
rect 22477 17629 22511 17663
rect 22511 17629 22520 17663
rect 22468 17620 22520 17629
rect 23480 17731 23532 17740
rect 23480 17697 23489 17731
rect 23489 17697 23523 17731
rect 23523 17697 23532 17731
rect 23480 17688 23532 17697
rect 23756 17620 23808 17672
rect 24676 17731 24728 17740
rect 24676 17697 24685 17731
rect 24685 17697 24719 17731
rect 24719 17697 24728 17731
rect 24676 17688 24728 17697
rect 24768 17620 24820 17672
rect 27988 17824 28040 17876
rect 31208 17824 31260 17876
rect 31392 17824 31444 17876
rect 32496 17824 32548 17876
rect 27712 17731 27764 17740
rect 27712 17697 27721 17731
rect 27721 17697 27755 17731
rect 27755 17697 27764 17731
rect 27712 17688 27764 17697
rect 32312 17756 32364 17808
rect 32404 17756 32456 17808
rect 27436 17620 27488 17672
rect 27896 17663 27948 17672
rect 27896 17629 27905 17663
rect 27905 17629 27939 17663
rect 27939 17629 27948 17663
rect 27896 17620 27948 17629
rect 28172 17620 28224 17672
rect 28356 17663 28408 17672
rect 28356 17629 28365 17663
rect 28365 17629 28399 17663
rect 28399 17629 28408 17663
rect 28356 17620 28408 17629
rect 18604 17527 18656 17536
rect 18604 17493 18613 17527
rect 18613 17493 18647 17527
rect 18647 17493 18656 17527
rect 18604 17484 18656 17493
rect 18880 17527 18932 17536
rect 18880 17493 18889 17527
rect 18889 17493 18923 17527
rect 18923 17493 18932 17527
rect 18880 17484 18932 17493
rect 18972 17484 19024 17536
rect 23664 17484 23716 17536
rect 28264 17552 28316 17604
rect 28632 17620 28684 17672
rect 29736 17663 29788 17672
rect 29736 17629 29745 17663
rect 29745 17629 29779 17663
rect 29779 17629 29788 17663
rect 29736 17620 29788 17629
rect 30012 17688 30064 17740
rect 30288 17663 30340 17672
rect 30288 17629 30297 17663
rect 30297 17629 30331 17663
rect 30331 17629 30340 17663
rect 30288 17620 30340 17629
rect 32588 17688 32640 17740
rect 31300 17620 31352 17672
rect 34060 17799 34112 17808
rect 34060 17765 34069 17799
rect 34069 17765 34103 17799
rect 34103 17765 34112 17799
rect 34060 17756 34112 17765
rect 32956 17620 33008 17672
rect 33968 17620 34020 17672
rect 29184 17484 29236 17536
rect 30196 17527 30248 17536
rect 30196 17493 30205 17527
rect 30205 17493 30239 17527
rect 30239 17493 30248 17527
rect 30196 17484 30248 17493
rect 31944 17552 31996 17604
rect 32496 17484 32548 17536
rect 33784 17484 33836 17536
rect 4874 17382 4926 17434
rect 4938 17382 4990 17434
rect 5002 17382 5054 17434
rect 5066 17382 5118 17434
rect 5130 17382 5182 17434
rect 35594 17382 35646 17434
rect 35658 17382 35710 17434
rect 35722 17382 35774 17434
rect 35786 17382 35838 17434
rect 35850 17382 35902 17434
rect 3424 17323 3476 17332
rect 3424 17289 3433 17323
rect 3433 17289 3467 17323
rect 3467 17289 3476 17323
rect 3424 17280 3476 17289
rect 4252 17323 4304 17332
rect 4252 17289 4261 17323
rect 4261 17289 4295 17323
rect 4295 17289 4304 17323
rect 4252 17280 4304 17289
rect 3240 17187 3292 17196
rect 3240 17153 3249 17187
rect 3249 17153 3283 17187
rect 3283 17153 3292 17187
rect 3240 17144 3292 17153
rect 3792 17144 3844 17196
rect 5724 17280 5776 17332
rect 6368 17280 6420 17332
rect 4804 17212 4856 17264
rect 5264 17144 5316 17196
rect 3056 17076 3108 17128
rect 3792 16940 3844 16992
rect 4068 16940 4120 16992
rect 7656 17280 7708 17332
rect 8484 17144 8536 17196
rect 9220 17280 9272 17332
rect 10140 17280 10192 17332
rect 10876 17280 10928 17332
rect 11612 17280 11664 17332
rect 11980 17323 12032 17332
rect 11980 17289 11989 17323
rect 11989 17289 12023 17323
rect 12023 17289 12032 17323
rect 11980 17280 12032 17289
rect 12348 17323 12400 17332
rect 9496 17212 9548 17264
rect 9680 17212 9732 17264
rect 9036 17144 9088 17196
rect 7656 17076 7708 17128
rect 10324 17187 10376 17196
rect 10324 17153 10333 17187
rect 10333 17153 10367 17187
rect 10367 17153 10376 17187
rect 10324 17144 10376 17153
rect 10416 17187 10468 17196
rect 10416 17153 10425 17187
rect 10425 17153 10459 17187
rect 10459 17153 10468 17187
rect 10416 17144 10468 17153
rect 12348 17289 12357 17323
rect 12357 17289 12391 17323
rect 12391 17289 12400 17323
rect 12348 17280 12400 17289
rect 12440 17280 12492 17332
rect 12716 17280 12768 17332
rect 13820 17280 13872 17332
rect 14004 17323 14056 17332
rect 14004 17289 14013 17323
rect 14013 17289 14047 17323
rect 14047 17289 14056 17323
rect 14004 17280 14056 17289
rect 15752 17280 15804 17332
rect 16212 17280 16264 17332
rect 16580 17280 16632 17332
rect 11796 17144 11848 17196
rect 11152 17076 11204 17128
rect 12072 17076 12124 17128
rect 12532 17144 12584 17196
rect 13544 17144 13596 17196
rect 7932 17008 7984 17060
rect 18972 17212 19024 17264
rect 19156 17212 19208 17264
rect 15752 17144 15804 17196
rect 16856 17187 16908 17196
rect 16856 17153 16865 17187
rect 16865 17153 16899 17187
rect 16899 17153 16908 17187
rect 16856 17144 16908 17153
rect 17316 17144 17368 17196
rect 18052 17144 18104 17196
rect 18420 17144 18472 17196
rect 14464 17119 14516 17128
rect 14464 17085 14473 17119
rect 14473 17085 14507 17119
rect 14507 17085 14516 17119
rect 14464 17076 14516 17085
rect 14188 17051 14240 17060
rect 14188 17017 14197 17051
rect 14197 17017 14231 17051
rect 14231 17017 14240 17051
rect 17500 17076 17552 17128
rect 18788 17076 18840 17128
rect 14188 17008 14240 17017
rect 15844 17008 15896 17060
rect 16396 17008 16448 17060
rect 6092 16983 6144 16992
rect 6092 16949 6101 16983
rect 6101 16949 6135 16983
rect 6135 16949 6144 16983
rect 6092 16940 6144 16949
rect 9588 16940 9640 16992
rect 11796 16940 11848 16992
rect 16672 16983 16724 16992
rect 16672 16949 16681 16983
rect 16681 16949 16715 16983
rect 16715 16949 16724 16983
rect 16672 16940 16724 16949
rect 17684 16940 17736 16992
rect 18328 16940 18380 16992
rect 19800 17212 19852 17264
rect 21088 17280 21140 17332
rect 20168 17212 20220 17264
rect 19708 17187 19760 17196
rect 19708 17153 19718 17187
rect 19718 17153 19752 17187
rect 19752 17153 19760 17187
rect 19708 17144 19760 17153
rect 20168 17076 20220 17128
rect 20352 17119 20404 17128
rect 20352 17085 20361 17119
rect 20361 17085 20395 17119
rect 20395 17085 20404 17119
rect 20352 17076 20404 17085
rect 20444 17076 20496 17128
rect 20812 17187 20864 17196
rect 20812 17153 20821 17187
rect 20821 17153 20855 17187
rect 20855 17153 20864 17187
rect 20812 17144 20864 17153
rect 23112 17280 23164 17332
rect 28264 17280 28316 17332
rect 28356 17323 28408 17332
rect 28356 17289 28365 17323
rect 28365 17289 28399 17323
rect 28399 17289 28408 17323
rect 28356 17280 28408 17289
rect 20720 17008 20772 17060
rect 22560 17144 22612 17196
rect 27804 17144 27856 17196
rect 28632 17212 28684 17264
rect 23296 17076 23348 17128
rect 29184 17323 29236 17332
rect 29184 17289 29193 17323
rect 29193 17289 29227 17323
rect 29227 17289 29236 17323
rect 29184 17280 29236 17289
rect 30196 17280 30248 17332
rect 31944 17280 31996 17332
rect 32404 17280 32456 17332
rect 32864 17280 32916 17332
rect 33048 17280 33100 17332
rect 33968 17323 34020 17332
rect 33968 17289 33993 17323
rect 33993 17289 34020 17323
rect 33968 17280 34020 17289
rect 32496 17212 32548 17264
rect 33784 17255 33836 17264
rect 33784 17221 33793 17255
rect 33793 17221 33827 17255
rect 33827 17221 33836 17255
rect 33784 17212 33836 17221
rect 29184 17187 29236 17196
rect 29184 17153 29193 17187
rect 29193 17153 29227 17187
rect 29227 17153 29236 17187
rect 29184 17144 29236 17153
rect 29644 17144 29696 17196
rect 32128 17144 32180 17196
rect 23480 17008 23532 17060
rect 29368 17008 29420 17060
rect 32312 17119 32364 17128
rect 32312 17085 32321 17119
rect 32321 17085 32355 17119
rect 32355 17085 32364 17119
rect 32312 17076 32364 17085
rect 32404 17119 32456 17128
rect 32404 17085 32413 17119
rect 32413 17085 32447 17119
rect 32447 17085 32456 17119
rect 32404 17076 32456 17085
rect 32496 17119 32548 17128
rect 32496 17085 32505 17119
rect 32505 17085 32539 17119
rect 32539 17085 32548 17119
rect 32496 17076 32548 17085
rect 34520 17212 34572 17264
rect 34060 17076 34112 17128
rect 34520 17119 34572 17128
rect 34520 17085 34529 17119
rect 34529 17085 34563 17119
rect 34563 17085 34572 17119
rect 34520 17076 34572 17085
rect 31852 16940 31904 16992
rect 32956 16940 33008 16992
rect 34520 16940 34572 16992
rect 34704 16940 34756 16992
rect 34796 16983 34848 16992
rect 34796 16949 34805 16983
rect 34805 16949 34839 16983
rect 34839 16949 34848 16983
rect 34796 16940 34848 16949
rect 35348 16940 35400 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 3608 16736 3660 16788
rect 3056 16600 3108 16652
rect 4436 16643 4488 16652
rect 4436 16609 4445 16643
rect 4445 16609 4479 16643
rect 4479 16609 4488 16643
rect 4436 16600 4488 16609
rect 2136 16532 2188 16584
rect 1768 16439 1820 16448
rect 1768 16405 1777 16439
rect 1777 16405 1811 16439
rect 1811 16405 1820 16439
rect 1768 16396 1820 16405
rect 1952 16396 2004 16448
rect 3976 16575 4028 16584
rect 3976 16541 3985 16575
rect 3985 16541 4019 16575
rect 4019 16541 4028 16575
rect 3976 16532 4028 16541
rect 4160 16575 4212 16584
rect 4160 16541 4169 16575
rect 4169 16541 4203 16575
rect 4203 16541 4212 16575
rect 4160 16532 4212 16541
rect 3148 16396 3200 16448
rect 4252 16464 4304 16516
rect 6092 16736 6144 16788
rect 8484 16668 8536 16720
rect 6184 16600 6236 16652
rect 5908 16464 5960 16516
rect 9036 16668 9088 16720
rect 12992 16736 13044 16788
rect 16028 16736 16080 16788
rect 16580 16736 16632 16788
rect 16672 16779 16724 16788
rect 16672 16745 16681 16779
rect 16681 16745 16715 16779
rect 16715 16745 16724 16779
rect 16672 16736 16724 16745
rect 22468 16736 22520 16788
rect 27804 16736 27856 16788
rect 29184 16736 29236 16788
rect 31208 16779 31260 16788
rect 31208 16745 31217 16779
rect 31217 16745 31251 16779
rect 31251 16745 31260 16779
rect 31208 16736 31260 16745
rect 31852 16736 31904 16788
rect 8576 16575 8628 16584
rect 8576 16541 8585 16575
rect 8585 16541 8619 16575
rect 8619 16541 8628 16575
rect 8576 16532 8628 16541
rect 15660 16600 15712 16652
rect 16396 16600 16448 16652
rect 8944 16532 8996 16584
rect 14188 16575 14240 16584
rect 14188 16541 14197 16575
rect 14197 16541 14231 16575
rect 14231 16541 14240 16575
rect 14188 16532 14240 16541
rect 9404 16507 9456 16516
rect 9404 16473 9413 16507
rect 9413 16473 9447 16507
rect 9447 16473 9456 16507
rect 9404 16464 9456 16473
rect 9680 16464 9732 16516
rect 11244 16464 11296 16516
rect 13084 16464 13136 16516
rect 11060 16396 11112 16448
rect 12256 16396 12308 16448
rect 14464 16396 14516 16448
rect 16304 16396 16356 16448
rect 16672 16532 16724 16584
rect 16580 16464 16632 16516
rect 17592 16532 17644 16584
rect 20720 16668 20772 16720
rect 22284 16668 22336 16720
rect 23112 16668 23164 16720
rect 30288 16668 30340 16720
rect 32128 16779 32180 16788
rect 32128 16745 32137 16779
rect 32137 16745 32171 16779
rect 32171 16745 32180 16779
rect 32128 16736 32180 16745
rect 35256 16736 35308 16788
rect 35440 16779 35492 16788
rect 35440 16745 35449 16779
rect 35449 16745 35483 16779
rect 35483 16745 35492 16779
rect 35440 16736 35492 16745
rect 18236 16600 18288 16652
rect 20168 16600 20220 16652
rect 20536 16600 20588 16652
rect 20628 16600 20680 16652
rect 17408 16464 17460 16516
rect 18604 16575 18656 16584
rect 18604 16541 18613 16575
rect 18613 16541 18647 16575
rect 18647 16541 18656 16575
rect 18604 16532 18656 16541
rect 18788 16532 18840 16584
rect 20076 16532 20128 16584
rect 20352 16575 20404 16584
rect 20352 16541 20362 16575
rect 20362 16541 20396 16575
rect 20396 16541 20404 16575
rect 20352 16532 20404 16541
rect 18696 16464 18748 16516
rect 19064 16507 19116 16516
rect 19064 16473 19073 16507
rect 19073 16473 19107 16507
rect 19107 16473 19116 16507
rect 19064 16464 19116 16473
rect 20812 16532 20864 16584
rect 20996 16575 21048 16584
rect 20996 16541 21005 16575
rect 21005 16541 21039 16575
rect 21039 16541 21048 16575
rect 20996 16532 21048 16541
rect 23204 16643 23256 16652
rect 23204 16609 23213 16643
rect 23213 16609 23247 16643
rect 23247 16609 23256 16643
rect 23204 16600 23256 16609
rect 23848 16600 23900 16652
rect 24860 16600 24912 16652
rect 22284 16575 22336 16584
rect 22284 16541 22293 16575
rect 22293 16541 22327 16575
rect 22327 16541 22336 16575
rect 22284 16532 22336 16541
rect 23296 16532 23348 16584
rect 23388 16575 23440 16584
rect 23388 16541 23421 16575
rect 23421 16541 23440 16575
rect 23388 16532 23440 16541
rect 25228 16575 25280 16584
rect 25228 16541 25237 16575
rect 25237 16541 25271 16575
rect 25271 16541 25280 16575
rect 25228 16532 25280 16541
rect 26240 16600 26292 16652
rect 26056 16575 26108 16584
rect 16948 16396 17000 16448
rect 17684 16396 17736 16448
rect 18052 16396 18104 16448
rect 18144 16396 18196 16448
rect 18512 16396 18564 16448
rect 22468 16464 22520 16516
rect 23204 16464 23256 16516
rect 23756 16507 23808 16516
rect 23756 16473 23765 16507
rect 23765 16473 23799 16507
rect 23799 16473 23808 16507
rect 23756 16464 23808 16473
rect 26056 16541 26065 16575
rect 26065 16541 26099 16575
rect 26099 16541 26108 16575
rect 26056 16532 26108 16541
rect 31760 16600 31812 16652
rect 30196 16575 30248 16584
rect 30196 16541 30205 16575
rect 30205 16541 30239 16575
rect 30239 16541 30248 16575
rect 30196 16532 30248 16541
rect 30288 16532 30340 16584
rect 30656 16532 30708 16584
rect 31116 16532 31168 16584
rect 31484 16532 31536 16584
rect 34704 16600 34756 16652
rect 25964 16464 26016 16516
rect 29368 16464 29420 16516
rect 32772 16464 32824 16516
rect 20904 16439 20956 16448
rect 20904 16405 20913 16439
rect 20913 16405 20947 16439
rect 20947 16405 20956 16439
rect 20904 16396 20956 16405
rect 22652 16396 22704 16448
rect 24952 16396 25004 16448
rect 25136 16396 25188 16448
rect 26424 16439 26476 16448
rect 26424 16405 26433 16439
rect 26433 16405 26467 16439
rect 26467 16405 26476 16439
rect 26424 16396 26476 16405
rect 27160 16396 27212 16448
rect 30656 16396 30708 16448
rect 30748 16439 30800 16448
rect 30748 16405 30757 16439
rect 30757 16405 30791 16439
rect 30791 16405 30800 16439
rect 30748 16396 30800 16405
rect 35072 16532 35124 16584
rect 34796 16464 34848 16516
rect 35164 16439 35216 16448
rect 35164 16405 35189 16439
rect 35189 16405 35216 16439
rect 35164 16396 35216 16405
rect 4874 16294 4926 16346
rect 4938 16294 4990 16346
rect 5002 16294 5054 16346
rect 5066 16294 5118 16346
rect 5130 16294 5182 16346
rect 35594 16294 35646 16346
rect 35658 16294 35710 16346
rect 35722 16294 35774 16346
rect 35786 16294 35838 16346
rect 35850 16294 35902 16346
rect 1400 16192 1452 16244
rect 2964 16192 3016 16244
rect 3608 16192 3660 16244
rect 4620 16192 4672 16244
rect 5264 16192 5316 16244
rect 9404 16192 9456 16244
rect 1952 16124 2004 16176
rect 4804 16124 4856 16176
rect 4712 16056 4764 16108
rect 1400 16031 1452 16040
rect 1400 15997 1409 16031
rect 1409 15997 1443 16031
rect 1443 15997 1452 16031
rect 1400 15988 1452 15997
rect 2136 15988 2188 16040
rect 5632 16031 5684 16040
rect 5632 15997 5641 16031
rect 5641 15997 5675 16031
rect 5675 15997 5684 16031
rect 5632 15988 5684 15997
rect 5908 15988 5960 16040
rect 11244 16192 11296 16244
rect 14096 16192 14148 16244
rect 16672 16192 16724 16244
rect 18236 16192 18288 16244
rect 11060 16124 11112 16176
rect 12624 16124 12676 16176
rect 12256 16099 12308 16108
rect 12256 16065 12265 16099
rect 12265 16065 12299 16099
rect 12299 16065 12308 16099
rect 12256 16056 12308 16065
rect 12348 16099 12400 16108
rect 12348 16065 12357 16099
rect 12357 16065 12391 16099
rect 12391 16065 12400 16099
rect 12348 16056 12400 16065
rect 14464 16099 14516 16108
rect 14464 16065 14473 16099
rect 14473 16065 14507 16099
rect 14507 16065 14516 16099
rect 14464 16056 14516 16065
rect 14740 16099 14792 16108
rect 14740 16065 14749 16099
rect 14749 16065 14783 16099
rect 14783 16065 14792 16099
rect 14740 16056 14792 16065
rect 14832 16056 14884 16108
rect 10324 16031 10376 16040
rect 10324 15997 10333 16031
rect 10333 15997 10367 16031
rect 10367 15997 10376 16031
rect 10324 15988 10376 15997
rect 12164 15988 12216 16040
rect 12532 16031 12584 16040
rect 12532 15997 12541 16031
rect 12541 15997 12575 16031
rect 12575 15997 12584 16031
rect 12532 15988 12584 15997
rect 16764 16124 16816 16176
rect 17316 16124 17368 16176
rect 16396 16056 16448 16108
rect 3148 15895 3200 15904
rect 3148 15861 3157 15895
rect 3157 15861 3191 15895
rect 3191 15861 3200 15895
rect 3148 15852 3200 15861
rect 3884 15852 3936 15904
rect 16764 15920 16816 15972
rect 17500 15988 17552 16040
rect 17868 16124 17920 16176
rect 19064 16192 19116 16244
rect 20352 16167 20404 16176
rect 20352 16133 20361 16167
rect 20361 16133 20395 16167
rect 20395 16133 20404 16167
rect 20352 16124 20404 16133
rect 20720 16235 20772 16244
rect 20720 16201 20729 16235
rect 20729 16201 20763 16235
rect 20763 16201 20772 16235
rect 20720 16192 20772 16201
rect 22284 16192 22336 16244
rect 17592 15920 17644 15972
rect 18052 16056 18104 16108
rect 18144 16099 18196 16108
rect 18144 16065 18153 16099
rect 18153 16065 18187 16099
rect 18187 16065 18196 16099
rect 18144 16056 18196 16065
rect 17868 15963 17920 15972
rect 17868 15929 17877 15963
rect 17877 15929 17911 15963
rect 17911 15929 17920 15963
rect 17868 15920 17920 15929
rect 14188 15852 14240 15904
rect 14740 15852 14792 15904
rect 16672 15895 16724 15904
rect 16672 15861 16681 15895
rect 16681 15861 16715 15895
rect 16715 15861 16724 15895
rect 16672 15852 16724 15861
rect 18880 16056 18932 16108
rect 19708 16056 19760 16108
rect 20444 16056 20496 16108
rect 23020 16167 23072 16176
rect 23020 16133 23029 16167
rect 23029 16133 23063 16167
rect 23063 16133 23072 16167
rect 23020 16124 23072 16133
rect 25136 16124 25188 16176
rect 20904 16056 20956 16108
rect 21548 16056 21600 16108
rect 22008 16056 22060 16108
rect 20536 15988 20588 16040
rect 20996 16031 21048 16040
rect 20996 15997 21005 16031
rect 21005 15997 21039 16031
rect 21039 15997 21048 16031
rect 20996 15988 21048 15997
rect 20352 15920 20404 15972
rect 18604 15895 18656 15904
rect 18604 15861 18613 15895
rect 18613 15861 18647 15895
rect 18647 15861 18656 15895
rect 18604 15852 18656 15861
rect 18880 15895 18932 15904
rect 18880 15861 18889 15895
rect 18889 15861 18923 15895
rect 18923 15861 18932 15895
rect 18880 15852 18932 15861
rect 20168 15852 20220 15904
rect 20720 15852 20772 15904
rect 22928 15852 22980 15904
rect 23296 16056 23348 16108
rect 24676 16099 24728 16108
rect 24676 16065 24685 16099
rect 24685 16065 24719 16099
rect 24719 16065 24728 16099
rect 24676 16056 24728 16065
rect 24860 16056 24912 16108
rect 25228 15920 25280 15972
rect 26424 16056 26476 16108
rect 27252 16124 27304 16176
rect 27344 16099 27396 16108
rect 27344 16065 27353 16099
rect 27353 16065 27387 16099
rect 27387 16065 27396 16099
rect 27344 16056 27396 16065
rect 30196 16192 30248 16244
rect 30748 16192 30800 16244
rect 34796 16192 34848 16244
rect 35072 16192 35124 16244
rect 35440 16192 35492 16244
rect 29552 16099 29604 16108
rect 29552 16065 29561 16099
rect 29561 16065 29595 16099
rect 29595 16065 29604 16099
rect 29552 16056 29604 16065
rect 29644 16056 29696 16108
rect 30288 16124 30340 16176
rect 31116 16124 31168 16176
rect 29184 15988 29236 16040
rect 27344 15920 27396 15972
rect 32220 15988 32272 16040
rect 35164 16099 35216 16108
rect 35164 16065 35173 16099
rect 35173 16065 35207 16099
rect 35207 16065 35216 16099
rect 35164 16056 35216 16065
rect 35256 15988 35308 16040
rect 24032 15852 24084 15904
rect 25044 15852 25096 15904
rect 27160 15852 27212 15904
rect 30012 15852 30064 15904
rect 30196 15852 30248 15904
rect 30380 15852 30432 15904
rect 35072 15920 35124 15972
rect 31392 15895 31444 15904
rect 31392 15861 31401 15895
rect 31401 15861 31435 15895
rect 31435 15861 31444 15895
rect 31392 15852 31444 15861
rect 31760 15852 31812 15904
rect 32496 15852 32548 15904
rect 35348 15852 35400 15904
rect 37832 15895 37884 15904
rect 37832 15861 37841 15895
rect 37841 15861 37875 15895
rect 37875 15861 37884 15895
rect 37832 15852 37884 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 940 15648 992 15700
rect 3976 15648 4028 15700
rect 4712 15648 4764 15700
rect 5632 15648 5684 15700
rect 7932 15691 7984 15700
rect 7932 15657 7941 15691
rect 7941 15657 7975 15691
rect 7975 15657 7984 15691
rect 7932 15648 7984 15657
rect 9496 15648 9548 15700
rect 10232 15691 10284 15700
rect 10232 15657 10241 15691
rect 10241 15657 10275 15691
rect 10275 15657 10284 15691
rect 10232 15648 10284 15657
rect 4620 15580 4672 15632
rect 1768 15487 1820 15496
rect 1768 15453 1777 15487
rect 1777 15453 1811 15487
rect 1811 15453 1820 15487
rect 1768 15444 1820 15453
rect 3884 15444 3936 15496
rect 3976 15487 4028 15496
rect 3976 15453 3985 15487
rect 3985 15453 4019 15487
rect 4019 15453 4028 15487
rect 3976 15444 4028 15453
rect 4160 15487 4212 15496
rect 4160 15453 4169 15487
rect 4169 15453 4203 15487
rect 4203 15453 4212 15487
rect 4160 15444 4212 15453
rect 6184 15555 6236 15564
rect 6184 15521 6193 15555
rect 6193 15521 6227 15555
rect 6227 15521 6236 15555
rect 6184 15512 6236 15521
rect 4804 15444 4856 15496
rect 7840 15444 7892 15496
rect 11244 15512 11296 15564
rect 12532 15648 12584 15700
rect 14188 15648 14240 15700
rect 15476 15648 15528 15700
rect 17776 15648 17828 15700
rect 11152 15444 11204 15496
rect 11428 15487 11480 15496
rect 11428 15453 11437 15487
rect 11437 15453 11471 15487
rect 11471 15453 11480 15487
rect 11428 15444 11480 15453
rect 6368 15376 6420 15428
rect 6460 15419 6512 15428
rect 6460 15385 6469 15419
rect 6469 15385 6503 15419
rect 6503 15385 6512 15419
rect 6460 15376 6512 15385
rect 6920 15376 6972 15428
rect 5356 15308 5408 15360
rect 11888 15487 11940 15496
rect 11888 15453 11897 15487
rect 11897 15453 11931 15487
rect 11931 15453 11940 15487
rect 11888 15444 11940 15453
rect 14096 15444 14148 15496
rect 14648 15444 14700 15496
rect 15752 15487 15804 15496
rect 15752 15453 15761 15487
rect 15761 15453 15795 15487
rect 15795 15453 15804 15487
rect 15752 15444 15804 15453
rect 15844 15487 15896 15496
rect 15844 15453 15853 15487
rect 15853 15453 15887 15487
rect 15887 15453 15896 15487
rect 15844 15444 15896 15453
rect 15936 15487 15988 15496
rect 15936 15453 15945 15487
rect 15945 15453 15979 15487
rect 15979 15453 15988 15487
rect 15936 15444 15988 15453
rect 16396 15512 16448 15564
rect 16488 15512 16540 15564
rect 19064 15580 19116 15632
rect 18604 15512 18656 15564
rect 21088 15648 21140 15700
rect 24492 15648 24544 15700
rect 19248 15580 19300 15632
rect 11612 15376 11664 15428
rect 12440 15376 12492 15428
rect 13820 15376 13872 15428
rect 14740 15376 14792 15428
rect 15660 15376 15712 15428
rect 18236 15487 18288 15496
rect 18236 15453 18245 15487
rect 18245 15453 18279 15487
rect 18279 15453 18288 15487
rect 18236 15444 18288 15453
rect 20628 15555 20680 15564
rect 20628 15521 20637 15555
rect 20637 15521 20671 15555
rect 20671 15521 20680 15555
rect 20628 15512 20680 15521
rect 22652 15512 22704 15564
rect 22744 15512 22796 15564
rect 18696 15376 18748 15428
rect 18788 15308 18840 15360
rect 19616 15376 19668 15428
rect 20076 15376 20128 15428
rect 20536 15376 20588 15428
rect 22008 15444 22060 15496
rect 23020 15444 23072 15496
rect 23572 15376 23624 15428
rect 24492 15487 24544 15496
rect 24492 15453 24501 15487
rect 24501 15453 24535 15487
rect 24535 15453 24544 15487
rect 24492 15444 24544 15453
rect 24676 15444 24728 15496
rect 25228 15487 25280 15496
rect 25228 15453 25237 15487
rect 25237 15453 25271 15487
rect 25271 15453 25280 15487
rect 25228 15444 25280 15453
rect 27344 15648 27396 15700
rect 30748 15648 30800 15700
rect 31392 15648 31444 15700
rect 32220 15648 32272 15700
rect 32496 15648 32548 15700
rect 32864 15648 32916 15700
rect 34704 15648 34756 15700
rect 35348 15648 35400 15700
rect 29184 15512 29236 15564
rect 29552 15512 29604 15564
rect 25504 15444 25556 15496
rect 25964 15487 26016 15496
rect 25964 15453 25973 15487
rect 25973 15453 26007 15487
rect 26007 15453 26016 15487
rect 25964 15444 26016 15453
rect 26056 15444 26108 15496
rect 26240 15444 26292 15496
rect 27160 15444 27212 15496
rect 27620 15487 27672 15496
rect 27620 15453 27629 15487
rect 27629 15453 27663 15487
rect 27663 15453 27672 15487
rect 27620 15444 27672 15453
rect 29644 15487 29696 15496
rect 25320 15376 25372 15428
rect 29644 15453 29653 15487
rect 29653 15453 29687 15487
rect 29687 15453 29696 15487
rect 29644 15444 29696 15453
rect 34520 15512 34572 15564
rect 32864 15444 32916 15496
rect 33416 15487 33468 15496
rect 33416 15453 33425 15487
rect 33425 15453 33459 15487
rect 33459 15453 33468 15487
rect 33416 15444 33468 15453
rect 34612 15444 34664 15496
rect 34796 15555 34848 15564
rect 34796 15521 34805 15555
rect 34805 15521 34839 15555
rect 34839 15521 34848 15555
rect 34796 15512 34848 15521
rect 35348 15512 35400 15564
rect 19156 15308 19208 15360
rect 22928 15308 22980 15360
rect 24676 15308 24728 15360
rect 25504 15308 25556 15360
rect 25688 15308 25740 15360
rect 26700 15308 26752 15360
rect 27344 15308 27396 15360
rect 30748 15376 30800 15428
rect 32220 15376 32272 15428
rect 28356 15351 28408 15360
rect 28356 15317 28365 15351
rect 28365 15317 28399 15351
rect 28399 15317 28408 15351
rect 28356 15308 28408 15317
rect 30472 15308 30524 15360
rect 32588 15351 32640 15360
rect 32588 15317 32597 15351
rect 32597 15317 32631 15351
rect 32631 15317 32640 15351
rect 32588 15308 32640 15317
rect 4874 15206 4926 15258
rect 4938 15206 4990 15258
rect 5002 15206 5054 15258
rect 5066 15206 5118 15258
rect 5130 15206 5182 15258
rect 35594 15206 35646 15258
rect 35658 15206 35710 15258
rect 35722 15206 35774 15258
rect 35786 15206 35838 15258
rect 35850 15206 35902 15258
rect 5356 15104 5408 15156
rect 6460 15104 6512 15156
rect 7932 15104 7984 15156
rect 3240 14968 3292 15020
rect 4160 15036 4212 15088
rect 3976 14968 4028 15020
rect 3148 14943 3200 14952
rect 3148 14909 3157 14943
rect 3157 14909 3191 14943
rect 3191 14909 3200 14943
rect 3148 14900 3200 14909
rect 4252 14943 4304 14952
rect 4252 14909 4261 14943
rect 4261 14909 4295 14943
rect 4295 14909 4304 14943
rect 4252 14900 4304 14909
rect 4068 14832 4120 14884
rect 2504 14807 2556 14816
rect 2504 14773 2513 14807
rect 2513 14773 2547 14807
rect 2547 14773 2556 14807
rect 2504 14764 2556 14773
rect 3608 14807 3660 14816
rect 3608 14773 3617 14807
rect 3617 14773 3651 14807
rect 3651 14773 3660 14807
rect 3608 14764 3660 14773
rect 3884 14764 3936 14816
rect 4620 15036 4672 15088
rect 4712 15011 4764 15020
rect 4712 14977 4721 15011
rect 4721 14977 4755 15011
rect 4755 14977 4764 15011
rect 4712 14968 4764 14977
rect 8208 15104 8260 15156
rect 8576 15104 8628 15156
rect 8760 15104 8812 15156
rect 9220 15104 9272 15156
rect 12440 15104 12492 15156
rect 8392 15011 8444 15020
rect 8392 14977 8401 15011
rect 8401 14977 8435 15011
rect 8435 14977 8444 15011
rect 8392 14968 8444 14977
rect 8944 14968 8996 15020
rect 9588 15036 9640 15088
rect 11060 15036 11112 15088
rect 12072 15036 12124 15088
rect 12900 15036 12952 15088
rect 7656 14943 7708 14952
rect 7656 14909 7665 14943
rect 7665 14909 7699 14943
rect 7699 14909 7708 14943
rect 7656 14900 7708 14909
rect 9404 14900 9456 14952
rect 9036 14875 9088 14884
rect 9036 14841 9045 14875
rect 9045 14841 9079 14875
rect 9079 14841 9088 14875
rect 9036 14832 9088 14841
rect 12992 15011 13044 15020
rect 12992 14977 13001 15011
rect 13001 14977 13035 15011
rect 13035 14977 13044 15011
rect 12992 14968 13044 14977
rect 13360 15011 13412 15020
rect 13360 14977 13369 15011
rect 13369 14977 13403 15011
rect 13403 14977 13412 15011
rect 13360 14968 13412 14977
rect 14096 15011 14148 15020
rect 14096 14977 14105 15011
rect 14105 14977 14139 15011
rect 14139 14977 14148 15011
rect 14096 14968 14148 14977
rect 15568 15104 15620 15156
rect 16396 15104 16448 15156
rect 16488 15104 16540 15156
rect 12532 14900 12584 14952
rect 12256 14832 12308 14884
rect 14372 14968 14424 15020
rect 14464 14832 14516 14884
rect 14832 15011 14884 15020
rect 14832 14977 14841 15011
rect 14841 14977 14875 15011
rect 14875 14977 14884 15011
rect 14832 14968 14884 14977
rect 14648 14900 14700 14952
rect 14740 14832 14792 14884
rect 15384 15011 15436 15020
rect 15384 14977 15393 15011
rect 15393 14977 15427 15011
rect 15427 14977 15436 15011
rect 15384 14968 15436 14977
rect 16120 15036 16172 15088
rect 16212 15011 16264 15020
rect 16212 14977 16221 15011
rect 16221 14977 16255 15011
rect 16255 14977 16264 15011
rect 16212 14968 16264 14977
rect 19064 15104 19116 15156
rect 20168 15147 20220 15156
rect 20168 15113 20177 15147
rect 20177 15113 20211 15147
rect 20211 15113 20220 15147
rect 20168 15104 20220 15113
rect 26056 15104 26108 15156
rect 27344 15104 27396 15156
rect 27712 15104 27764 15156
rect 17868 15036 17920 15088
rect 24216 15036 24268 15088
rect 17040 15011 17092 15020
rect 17040 14977 17049 15011
rect 17049 14977 17083 15011
rect 17083 14977 17092 15011
rect 17040 14968 17092 14977
rect 16304 14900 16356 14952
rect 17592 15011 17644 15020
rect 17592 14977 17601 15011
rect 17601 14977 17635 15011
rect 17635 14977 17644 15011
rect 17592 14968 17644 14977
rect 17684 15011 17736 15020
rect 17684 14977 17693 15011
rect 17693 14977 17727 15011
rect 17727 14977 17736 15011
rect 17684 14968 17736 14977
rect 18236 15011 18288 15020
rect 18236 14977 18245 15011
rect 18245 14977 18279 15011
rect 18279 14977 18288 15011
rect 18236 14968 18288 14977
rect 18604 14968 18656 15020
rect 19064 14968 19116 15020
rect 19616 15011 19668 15020
rect 19616 14977 19625 15011
rect 19625 14977 19659 15011
rect 19659 14977 19668 15011
rect 19616 14968 19668 14977
rect 20076 15011 20128 15020
rect 20076 14977 20085 15011
rect 20085 14977 20119 15011
rect 20119 14977 20128 15011
rect 20076 14968 20128 14977
rect 18696 14943 18748 14952
rect 18696 14909 18705 14943
rect 18705 14909 18739 14943
rect 18739 14909 18748 14943
rect 18696 14900 18748 14909
rect 19432 14900 19484 14952
rect 20996 14968 21048 15020
rect 21916 14968 21968 15020
rect 25688 15011 25740 15020
rect 25688 14977 25697 15011
rect 25697 14977 25731 15011
rect 25731 14977 25740 15011
rect 25688 14968 25740 14977
rect 21824 14943 21876 14952
rect 21824 14909 21833 14943
rect 21833 14909 21867 14943
rect 21867 14909 21876 14943
rect 21824 14900 21876 14909
rect 23296 14900 23348 14952
rect 25596 14900 25648 14952
rect 26424 14968 26476 15020
rect 27160 14968 27212 15020
rect 32588 15104 32640 15156
rect 34796 15104 34848 15156
rect 27988 15036 28040 15088
rect 27896 15011 27948 15020
rect 27896 14977 27905 15011
rect 27905 14977 27939 15011
rect 27939 14977 27948 15011
rect 27896 14968 27948 14977
rect 26148 14900 26200 14952
rect 28816 15011 28868 15020
rect 28816 14977 28825 15011
rect 28825 14977 28859 15011
rect 28859 14977 28868 15011
rect 28816 14968 28868 14977
rect 30472 14968 30524 15020
rect 30748 15011 30800 15020
rect 30748 14977 30757 15011
rect 30757 14977 30791 15011
rect 30791 14977 30800 15011
rect 30748 14968 30800 14977
rect 30840 15011 30892 15020
rect 30840 14977 30849 15011
rect 30849 14977 30883 15011
rect 30883 14977 30892 15011
rect 30840 14968 30892 14977
rect 8668 14807 8720 14816
rect 8668 14773 8677 14807
rect 8677 14773 8711 14807
rect 8711 14773 8720 14807
rect 8668 14764 8720 14773
rect 8944 14764 8996 14816
rect 9772 14807 9824 14816
rect 9772 14773 9781 14807
rect 9781 14773 9815 14807
rect 9815 14773 9824 14807
rect 9772 14764 9824 14773
rect 10232 14764 10284 14816
rect 13544 14807 13596 14816
rect 13544 14773 13553 14807
rect 13553 14773 13587 14807
rect 13587 14773 13596 14807
rect 21272 14832 21324 14884
rect 23664 14832 23716 14884
rect 24768 14832 24820 14884
rect 13544 14764 13596 14773
rect 16396 14807 16448 14816
rect 16396 14773 16405 14807
rect 16405 14773 16439 14807
rect 16439 14773 16448 14807
rect 16396 14764 16448 14773
rect 16580 14764 16632 14816
rect 17684 14764 17736 14816
rect 18788 14764 18840 14816
rect 19248 14764 19300 14816
rect 20536 14807 20588 14816
rect 20536 14773 20545 14807
rect 20545 14773 20579 14807
rect 20579 14773 20588 14807
rect 20536 14764 20588 14773
rect 20812 14764 20864 14816
rect 22192 14764 22244 14816
rect 25596 14807 25648 14816
rect 25596 14773 25605 14807
rect 25605 14773 25639 14807
rect 25639 14773 25648 14807
rect 25596 14764 25648 14773
rect 26332 14764 26384 14816
rect 28724 14900 28776 14952
rect 28540 14832 28592 14884
rect 28816 14832 28868 14884
rect 29460 14900 29512 14952
rect 30380 14900 30432 14952
rect 31116 15011 31168 15020
rect 31116 14977 31125 15011
rect 31125 14977 31159 15011
rect 31159 14977 31168 15011
rect 31116 14968 31168 14977
rect 33048 15011 33100 15020
rect 33048 14977 33057 15011
rect 33057 14977 33091 15011
rect 33091 14977 33100 15011
rect 33048 14968 33100 14977
rect 31668 14900 31720 14952
rect 32956 14943 33008 14952
rect 32956 14909 32965 14943
rect 32965 14909 32999 14943
rect 32999 14909 33008 14943
rect 32956 14900 33008 14909
rect 31208 14764 31260 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 3240 14560 3292 14612
rect 3608 14560 3660 14612
rect 4068 14603 4120 14612
rect 4068 14569 4077 14603
rect 4077 14569 4111 14603
rect 4111 14569 4120 14603
rect 4068 14560 4120 14569
rect 7380 14603 7432 14612
rect 7380 14569 7389 14603
rect 7389 14569 7423 14603
rect 7423 14569 7432 14603
rect 7380 14560 7432 14569
rect 8668 14560 8720 14612
rect 8852 14560 8904 14612
rect 14096 14560 14148 14612
rect 14832 14560 14884 14612
rect 15568 14560 15620 14612
rect 15936 14560 15988 14612
rect 16580 14603 16632 14612
rect 16580 14569 16589 14603
rect 16589 14569 16623 14603
rect 16623 14569 16632 14603
rect 16580 14560 16632 14569
rect 17040 14603 17092 14612
rect 17040 14569 17049 14603
rect 17049 14569 17083 14603
rect 17083 14569 17092 14603
rect 17040 14560 17092 14569
rect 17408 14603 17460 14612
rect 17408 14569 17417 14603
rect 17417 14569 17451 14603
rect 17451 14569 17460 14603
rect 17408 14560 17460 14569
rect 22928 14560 22980 14612
rect 1400 14399 1452 14408
rect 1400 14365 1409 14399
rect 1409 14365 1443 14399
rect 1443 14365 1452 14399
rect 1400 14356 1452 14365
rect 2780 14356 2832 14408
rect 9128 14492 9180 14544
rect 3700 14424 3752 14476
rect 4620 14356 4672 14408
rect 5632 14399 5684 14408
rect 5632 14365 5641 14399
rect 5641 14365 5675 14399
rect 5675 14365 5684 14399
rect 5632 14356 5684 14365
rect 9036 14356 9088 14408
rect 10232 14424 10284 14476
rect 12072 14424 12124 14476
rect 12532 14424 12584 14476
rect 14372 14424 14424 14476
rect 1676 14331 1728 14340
rect 1676 14297 1685 14331
rect 1685 14297 1719 14331
rect 1719 14297 1728 14331
rect 1676 14288 1728 14297
rect 5908 14331 5960 14340
rect 5908 14297 5917 14331
rect 5917 14297 5951 14331
rect 5951 14297 5960 14331
rect 5908 14288 5960 14297
rect 6920 14288 6972 14340
rect 8760 14288 8812 14340
rect 9864 14399 9916 14408
rect 9864 14365 9873 14399
rect 9873 14365 9907 14399
rect 9907 14365 9916 14399
rect 9864 14356 9916 14365
rect 11152 14356 11204 14408
rect 11704 14356 11756 14408
rect 14464 14356 14516 14408
rect 14832 14356 14884 14408
rect 15292 14399 15344 14408
rect 15292 14365 15301 14399
rect 15301 14365 15335 14399
rect 15335 14365 15344 14399
rect 15292 14356 15344 14365
rect 16396 14424 16448 14476
rect 16488 14356 16540 14408
rect 16672 14356 16724 14408
rect 9588 14331 9640 14340
rect 9588 14297 9597 14331
rect 9597 14297 9631 14331
rect 9631 14297 9640 14331
rect 9588 14288 9640 14297
rect 8668 14220 8720 14272
rect 15568 14288 15620 14340
rect 16948 14288 17000 14340
rect 14004 14220 14056 14272
rect 16120 14220 16172 14272
rect 17316 14399 17368 14408
rect 17316 14365 17325 14399
rect 17325 14365 17359 14399
rect 17359 14365 17368 14399
rect 17316 14356 17368 14365
rect 20536 14492 20588 14544
rect 20628 14492 20680 14544
rect 18052 14424 18104 14476
rect 19524 14288 19576 14340
rect 20444 14288 20496 14340
rect 20904 14356 20956 14408
rect 21088 14356 21140 14408
rect 23940 14492 23992 14544
rect 28356 14560 28408 14612
rect 31760 14560 31812 14612
rect 32956 14560 33008 14612
rect 29184 14492 29236 14544
rect 31300 14492 31352 14544
rect 21916 14424 21968 14476
rect 23296 14467 23348 14476
rect 23296 14433 23305 14467
rect 23305 14433 23339 14467
rect 23339 14433 23348 14467
rect 23296 14424 23348 14433
rect 30840 14424 30892 14476
rect 21824 14288 21876 14340
rect 23204 14288 23256 14340
rect 24124 14356 24176 14408
rect 24492 14356 24544 14408
rect 26240 14288 26292 14340
rect 27160 14288 27212 14340
rect 30472 14288 30524 14340
rect 30748 14288 30800 14340
rect 31208 14399 31260 14408
rect 31208 14365 31217 14399
rect 31217 14365 31251 14399
rect 31251 14365 31260 14399
rect 31208 14356 31260 14365
rect 31392 14399 31444 14408
rect 31392 14365 31401 14399
rect 31401 14365 31435 14399
rect 31435 14365 31444 14399
rect 31392 14356 31444 14365
rect 31668 14424 31720 14476
rect 33784 14424 33836 14476
rect 31760 14399 31812 14408
rect 31760 14365 31769 14399
rect 31769 14365 31803 14399
rect 31803 14365 31812 14399
rect 31760 14356 31812 14365
rect 34060 14356 34112 14408
rect 19432 14220 19484 14272
rect 23848 14220 23900 14272
rect 26424 14220 26476 14272
rect 30288 14220 30340 14272
rect 30380 14220 30432 14272
rect 32128 14220 32180 14272
rect 4874 14118 4926 14170
rect 4938 14118 4990 14170
rect 5002 14118 5054 14170
rect 5066 14118 5118 14170
rect 5130 14118 5182 14170
rect 35594 14118 35646 14170
rect 35658 14118 35710 14170
rect 35722 14118 35774 14170
rect 35786 14118 35838 14170
rect 35850 14118 35902 14170
rect 1676 14016 1728 14068
rect 2504 14016 2556 14068
rect 5908 14016 5960 14068
rect 8668 14059 8720 14068
rect 8668 14025 8677 14059
rect 8677 14025 8711 14059
rect 8711 14025 8720 14059
rect 8668 14016 8720 14025
rect 16764 14016 16816 14068
rect 17868 14059 17920 14068
rect 17868 14025 17877 14059
rect 17877 14025 17911 14059
rect 17911 14025 17920 14059
rect 17868 14016 17920 14025
rect 21088 14016 21140 14068
rect 7380 13948 7432 14000
rect 1492 13855 1544 13864
rect 1492 13821 1501 13855
rect 1501 13821 1535 13855
rect 1535 13821 1544 13855
rect 1492 13812 1544 13821
rect 8392 13923 8444 13932
rect 8392 13889 8401 13923
rect 8401 13889 8435 13923
rect 8435 13889 8444 13923
rect 8392 13880 8444 13889
rect 8576 13948 8628 14000
rect 10140 13948 10192 14000
rect 12992 13948 13044 14000
rect 13268 13948 13320 14000
rect 9956 13880 10008 13932
rect 12440 13880 12492 13932
rect 13360 13880 13412 13932
rect 15108 13948 15160 14000
rect 15200 13880 15252 13932
rect 17500 13948 17552 14000
rect 20536 13948 20588 14000
rect 17316 13880 17368 13932
rect 19708 13923 19760 13932
rect 19708 13889 19717 13923
rect 19717 13889 19751 13923
rect 19751 13889 19760 13923
rect 19708 13880 19760 13889
rect 6000 13812 6052 13864
rect 7656 13812 7708 13864
rect 15568 13855 15620 13864
rect 15568 13821 15577 13855
rect 15577 13821 15611 13855
rect 15611 13821 15620 13855
rect 15568 13812 15620 13821
rect 10968 13744 11020 13796
rect 18420 13744 18472 13796
rect 18972 13744 19024 13796
rect 7104 13676 7156 13728
rect 15660 13676 15712 13728
rect 17408 13719 17460 13728
rect 17408 13685 17417 13719
rect 17417 13685 17451 13719
rect 17451 13685 17460 13719
rect 17408 13676 17460 13685
rect 17868 13676 17920 13728
rect 19616 13676 19668 13728
rect 20444 13880 20496 13932
rect 20720 13880 20772 13932
rect 22560 13948 22612 14000
rect 22100 13923 22152 13932
rect 22100 13889 22109 13923
rect 22109 13889 22143 13923
rect 22143 13889 22152 13923
rect 22100 13880 22152 13889
rect 24124 13923 24176 13932
rect 24124 13889 24133 13923
rect 24133 13889 24167 13923
rect 24167 13889 24176 13923
rect 24124 13880 24176 13889
rect 24492 13923 24544 13932
rect 24492 13889 24501 13923
rect 24501 13889 24535 13923
rect 24535 13889 24544 13923
rect 24492 13880 24544 13889
rect 20904 13744 20956 13796
rect 21364 13744 21416 13796
rect 22468 13855 22520 13864
rect 22468 13821 22477 13855
rect 22477 13821 22511 13855
rect 22511 13821 22520 13855
rect 22468 13812 22520 13821
rect 22928 13812 22980 13864
rect 23112 13855 23164 13864
rect 23112 13821 23121 13855
rect 23121 13821 23155 13855
rect 23155 13821 23164 13855
rect 23112 13812 23164 13821
rect 23204 13855 23256 13864
rect 23204 13821 23213 13855
rect 23213 13821 23247 13855
rect 23247 13821 23256 13855
rect 23204 13812 23256 13821
rect 22744 13744 22796 13796
rect 23388 13812 23440 13864
rect 23664 13855 23716 13864
rect 23664 13821 23673 13855
rect 23673 13821 23707 13855
rect 23707 13821 23716 13855
rect 23664 13812 23716 13821
rect 24308 13812 24360 13864
rect 24216 13744 24268 13796
rect 24768 13923 24820 13932
rect 24768 13889 24777 13923
rect 24777 13889 24811 13923
rect 24811 13889 24820 13923
rect 24768 13880 24820 13889
rect 25044 13923 25096 13932
rect 25044 13889 25053 13923
rect 25053 13889 25087 13923
rect 25087 13889 25096 13923
rect 25044 13880 25096 13889
rect 25780 13880 25832 13932
rect 26332 14016 26384 14068
rect 26056 13923 26108 13932
rect 26056 13889 26065 13923
rect 26065 13889 26099 13923
rect 26099 13889 26108 13923
rect 26056 13880 26108 13889
rect 26148 13880 26200 13932
rect 27252 14016 27304 14068
rect 28540 14016 28592 14068
rect 29276 14016 29328 14068
rect 30196 14016 30248 14068
rect 25044 13744 25096 13796
rect 23112 13676 23164 13728
rect 25964 13744 26016 13796
rect 26424 13812 26476 13864
rect 26700 13880 26752 13932
rect 27804 13948 27856 14000
rect 31484 14016 31536 14068
rect 32864 14059 32916 14068
rect 32864 14025 32873 14059
rect 32873 14025 32907 14059
rect 32907 14025 32916 14059
rect 32864 14016 32916 14025
rect 27620 13880 27672 13932
rect 28816 13923 28868 13932
rect 28816 13889 28825 13923
rect 28825 13889 28859 13923
rect 28859 13889 28868 13923
rect 28816 13880 28868 13889
rect 29000 13812 29052 13864
rect 29184 13880 29236 13932
rect 30380 13923 30432 13932
rect 30380 13889 30389 13923
rect 30389 13889 30423 13923
rect 30423 13889 30432 13923
rect 30380 13880 30432 13889
rect 30472 13923 30524 13932
rect 30472 13889 30481 13923
rect 30481 13889 30515 13923
rect 30515 13889 30524 13923
rect 30472 13880 30524 13889
rect 30564 13855 30616 13864
rect 30564 13821 30573 13855
rect 30573 13821 30607 13855
rect 30607 13821 30616 13855
rect 30564 13812 30616 13821
rect 32404 13812 32456 13864
rect 26056 13676 26108 13728
rect 26240 13676 26292 13728
rect 26976 13676 27028 13728
rect 27344 13676 27396 13728
rect 28540 13719 28592 13728
rect 28540 13685 28549 13719
rect 28549 13685 28583 13719
rect 28583 13685 28592 13719
rect 28540 13676 28592 13685
rect 32588 13744 32640 13796
rect 32956 13923 33008 13932
rect 32956 13889 32965 13923
rect 32965 13889 32999 13923
rect 32999 13889 33008 13923
rect 32956 13880 33008 13889
rect 33232 13923 33284 13932
rect 33232 13889 33241 13923
rect 33241 13889 33275 13923
rect 33275 13889 33284 13923
rect 33232 13880 33284 13889
rect 29368 13676 29420 13728
rect 30196 13676 30248 13728
rect 30472 13676 30524 13728
rect 31852 13719 31904 13728
rect 31852 13685 31861 13719
rect 31861 13685 31895 13719
rect 31895 13685 31904 13719
rect 31852 13676 31904 13685
rect 33140 13676 33192 13728
rect 33508 13676 33560 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 9036 13472 9088 13524
rect 10324 13472 10376 13524
rect 10416 13472 10468 13524
rect 1400 13336 1452 13388
rect 5632 13336 5684 13388
rect 6276 13336 6328 13388
rect 2964 13268 3016 13320
rect 3792 13268 3844 13320
rect 3976 13200 4028 13252
rect 4620 13243 4672 13252
rect 4620 13209 4629 13243
rect 4629 13209 4663 13243
rect 4663 13209 4672 13243
rect 4620 13200 4672 13209
rect 2780 13132 2832 13184
rect 6920 13336 6972 13388
rect 7104 13379 7156 13388
rect 7104 13345 7113 13379
rect 7113 13345 7147 13379
rect 7147 13345 7156 13379
rect 7104 13336 7156 13345
rect 9588 13336 9640 13388
rect 9220 13268 9272 13320
rect 9956 13243 10008 13252
rect 9956 13209 9965 13243
rect 9965 13209 9999 13243
rect 9999 13209 10008 13243
rect 9956 13200 10008 13209
rect 10140 13311 10192 13320
rect 10140 13277 10149 13311
rect 10149 13277 10183 13311
rect 10183 13277 10192 13311
rect 10140 13268 10192 13277
rect 11244 13472 11296 13524
rect 15292 13472 15344 13524
rect 16856 13472 16908 13524
rect 17868 13515 17920 13524
rect 17868 13481 17877 13515
rect 17877 13481 17911 13515
rect 17911 13481 17920 13515
rect 17868 13472 17920 13481
rect 18420 13515 18472 13524
rect 18420 13481 18429 13515
rect 18429 13481 18463 13515
rect 18463 13481 18472 13515
rect 18420 13472 18472 13481
rect 11888 13336 11940 13388
rect 12532 13336 12584 13388
rect 13084 13268 13136 13320
rect 16764 13404 16816 13456
rect 17592 13404 17644 13456
rect 19708 13515 19760 13524
rect 19708 13481 19717 13515
rect 19717 13481 19751 13515
rect 19751 13481 19760 13515
rect 19708 13472 19760 13481
rect 19248 13404 19300 13456
rect 19340 13404 19392 13456
rect 16948 13336 17000 13388
rect 15108 13268 15160 13320
rect 16028 13268 16080 13320
rect 18420 13336 18472 13388
rect 20904 13472 20956 13524
rect 11152 13200 11204 13252
rect 6552 13175 6604 13184
rect 6552 13141 6561 13175
rect 6561 13141 6595 13175
rect 6595 13141 6604 13175
rect 6552 13132 6604 13141
rect 8024 13132 8076 13184
rect 8576 13175 8628 13184
rect 8576 13141 8585 13175
rect 8585 13141 8619 13175
rect 8619 13141 8628 13175
rect 8576 13132 8628 13141
rect 9404 13132 9456 13184
rect 9588 13175 9640 13184
rect 9588 13141 9597 13175
rect 9597 13141 9631 13175
rect 9631 13141 9640 13175
rect 9588 13132 9640 13141
rect 11704 13200 11756 13252
rect 12716 13175 12768 13184
rect 12716 13141 12725 13175
rect 12725 13141 12759 13175
rect 12759 13141 12768 13175
rect 12716 13132 12768 13141
rect 13360 13132 13412 13184
rect 15200 13243 15252 13252
rect 15200 13209 15209 13243
rect 15209 13209 15243 13243
rect 15243 13209 15252 13243
rect 15200 13200 15252 13209
rect 16672 13243 16724 13252
rect 16672 13209 16681 13243
rect 16681 13209 16715 13243
rect 16715 13209 16724 13243
rect 16672 13200 16724 13209
rect 13544 13132 13596 13184
rect 13636 13175 13688 13184
rect 13636 13141 13645 13175
rect 13645 13141 13679 13175
rect 13679 13141 13688 13175
rect 13636 13132 13688 13141
rect 15476 13132 15528 13184
rect 20444 13404 20496 13456
rect 16856 13243 16908 13252
rect 16856 13209 16865 13243
rect 16865 13209 16899 13243
rect 16899 13209 16908 13243
rect 16856 13200 16908 13209
rect 18236 13243 18288 13252
rect 18236 13209 18245 13243
rect 18245 13209 18279 13243
rect 18279 13209 18288 13243
rect 18236 13200 18288 13209
rect 19524 13268 19576 13320
rect 19984 13311 20036 13320
rect 19984 13277 19993 13311
rect 19993 13277 20027 13311
rect 20027 13277 20036 13311
rect 19984 13268 20036 13277
rect 20076 13311 20128 13320
rect 20076 13277 20085 13311
rect 20085 13277 20119 13311
rect 20119 13277 20128 13311
rect 20076 13268 20128 13277
rect 20628 13336 20680 13388
rect 22744 13404 22796 13456
rect 23112 13404 23164 13456
rect 18880 13243 18932 13252
rect 18420 13175 18472 13184
rect 18420 13141 18445 13175
rect 18445 13141 18472 13175
rect 18420 13132 18472 13141
rect 18696 13175 18748 13184
rect 18696 13141 18705 13175
rect 18705 13141 18739 13175
rect 18739 13141 18748 13175
rect 18696 13132 18748 13141
rect 18880 13209 18907 13243
rect 18907 13209 18932 13243
rect 18880 13200 18932 13209
rect 18972 13200 19024 13252
rect 20536 13268 20588 13320
rect 21088 13311 21140 13320
rect 21088 13277 21097 13311
rect 21097 13277 21131 13311
rect 21131 13277 21140 13311
rect 21088 13268 21140 13277
rect 21364 13311 21416 13320
rect 21364 13277 21373 13311
rect 21373 13277 21407 13311
rect 21407 13277 21416 13311
rect 21364 13268 21416 13277
rect 21732 13311 21784 13320
rect 21732 13277 21741 13311
rect 21741 13277 21775 13311
rect 21775 13277 21784 13311
rect 21732 13268 21784 13277
rect 21916 13268 21968 13320
rect 23204 13311 23256 13320
rect 23204 13277 23213 13311
rect 23213 13277 23247 13311
rect 23247 13277 23256 13311
rect 23204 13268 23256 13277
rect 24124 13268 24176 13320
rect 25780 13336 25832 13388
rect 24492 13200 24544 13252
rect 19248 13132 19300 13184
rect 21088 13132 21140 13184
rect 21180 13132 21232 13184
rect 21548 13175 21600 13184
rect 21548 13141 21557 13175
rect 21557 13141 21591 13175
rect 21591 13141 21600 13175
rect 21548 13132 21600 13141
rect 22744 13132 22796 13184
rect 22928 13132 22980 13184
rect 23112 13132 23164 13184
rect 25596 13268 25648 13320
rect 25872 13311 25924 13320
rect 25872 13277 25881 13311
rect 25881 13277 25915 13311
rect 25915 13277 25924 13311
rect 25872 13268 25924 13277
rect 26056 13336 26108 13388
rect 26240 13379 26292 13388
rect 26240 13345 26249 13379
rect 26249 13345 26283 13379
rect 26283 13345 26292 13379
rect 26240 13336 26292 13345
rect 27068 13404 27120 13456
rect 27804 13472 27856 13524
rect 27896 13472 27948 13524
rect 28172 13472 28224 13524
rect 28448 13472 28500 13524
rect 29000 13472 29052 13524
rect 29184 13515 29236 13524
rect 29184 13481 29193 13515
rect 29193 13481 29227 13515
rect 29227 13481 29236 13515
rect 29184 13472 29236 13481
rect 32404 13472 32456 13524
rect 33232 13515 33284 13524
rect 33232 13481 33241 13515
rect 33241 13481 33275 13515
rect 33275 13481 33284 13515
rect 33232 13472 33284 13481
rect 33416 13472 33468 13524
rect 28264 13447 28316 13456
rect 28264 13413 28273 13447
rect 28273 13413 28307 13447
rect 28307 13413 28316 13447
rect 28264 13404 28316 13413
rect 30288 13404 30340 13456
rect 26148 13311 26200 13320
rect 26148 13277 26157 13311
rect 26157 13277 26191 13311
rect 26191 13277 26200 13311
rect 26148 13268 26200 13277
rect 26516 13311 26568 13320
rect 26516 13277 26525 13311
rect 26525 13277 26559 13311
rect 26559 13277 26568 13311
rect 26516 13268 26568 13277
rect 26792 13311 26844 13320
rect 26792 13277 26801 13311
rect 26801 13277 26835 13311
rect 26835 13277 26844 13311
rect 26792 13268 26844 13277
rect 27344 13336 27396 13388
rect 26884 13200 26936 13252
rect 24860 13132 24912 13184
rect 26240 13132 26292 13184
rect 26700 13132 26752 13184
rect 27436 13268 27488 13320
rect 28356 13268 28408 13320
rect 28540 13311 28592 13320
rect 28540 13277 28549 13311
rect 28549 13277 28583 13311
rect 28583 13277 28592 13311
rect 28540 13268 28592 13277
rect 29276 13311 29328 13320
rect 29276 13277 29285 13311
rect 29285 13277 29319 13311
rect 29319 13277 29328 13311
rect 29276 13268 29328 13277
rect 29368 13268 29420 13320
rect 31208 13268 31260 13320
rect 32864 13311 32916 13320
rect 32864 13277 32873 13311
rect 32873 13277 32907 13311
rect 32907 13277 32916 13311
rect 32864 13268 32916 13277
rect 33140 13268 33192 13320
rect 32404 13200 32456 13252
rect 32588 13243 32640 13252
rect 32588 13209 32597 13243
rect 32597 13209 32631 13243
rect 32631 13209 32640 13243
rect 32588 13200 32640 13209
rect 33048 13200 33100 13252
rect 33508 13311 33560 13320
rect 33508 13277 33517 13311
rect 33517 13277 33551 13311
rect 33551 13277 33560 13311
rect 33508 13268 33560 13277
rect 33876 13311 33928 13320
rect 33876 13277 33885 13311
rect 33885 13277 33919 13311
rect 33919 13277 33928 13311
rect 33876 13268 33928 13277
rect 29644 13175 29696 13184
rect 29644 13141 29653 13175
rect 29653 13141 29687 13175
rect 29687 13141 29696 13175
rect 29644 13132 29696 13141
rect 4874 13030 4926 13082
rect 4938 13030 4990 13082
rect 5002 13030 5054 13082
rect 5066 13030 5118 13082
rect 5130 13030 5182 13082
rect 35594 13030 35646 13082
rect 35658 13030 35710 13082
rect 35722 13030 35774 13082
rect 35786 13030 35838 13082
rect 35850 13030 35902 13082
rect 3976 12928 4028 12980
rect 4620 12928 4672 12980
rect 6552 12928 6604 12980
rect 1400 12835 1452 12844
rect 1400 12801 1409 12835
rect 1409 12801 1443 12835
rect 1443 12801 1452 12835
rect 1400 12792 1452 12801
rect 2780 12792 2832 12844
rect 3976 12835 4028 12844
rect 3976 12801 3985 12835
rect 3985 12801 4019 12835
rect 4019 12801 4028 12835
rect 3976 12792 4028 12801
rect 4436 12835 4488 12844
rect 4436 12801 4445 12835
rect 4445 12801 4479 12835
rect 4479 12801 4488 12835
rect 4436 12792 4488 12801
rect 1676 12767 1728 12776
rect 1676 12733 1685 12767
rect 1685 12733 1719 12767
rect 1719 12733 1728 12767
rect 1676 12724 1728 12733
rect 3884 12724 3936 12776
rect 3792 12656 3844 12708
rect 4712 12792 4764 12844
rect 5816 12792 5868 12844
rect 6920 12860 6972 12912
rect 6368 12835 6420 12844
rect 6368 12801 6377 12835
rect 6377 12801 6411 12835
rect 6411 12801 6420 12835
rect 6368 12792 6420 12801
rect 8024 12928 8076 12980
rect 9864 12928 9916 12980
rect 10416 12928 10468 12980
rect 8576 12903 8628 12912
rect 8576 12869 8585 12903
rect 8585 12869 8619 12903
rect 8619 12869 8628 12903
rect 8576 12860 8628 12869
rect 9680 12792 9732 12844
rect 10232 12792 10284 12844
rect 9588 12656 9640 12708
rect 11888 12860 11940 12912
rect 13636 12928 13688 12980
rect 12256 12767 12308 12776
rect 12256 12733 12265 12767
rect 12265 12733 12299 12767
rect 12299 12733 12308 12767
rect 12256 12724 12308 12733
rect 12716 12792 12768 12844
rect 13544 12860 13596 12912
rect 15200 12928 15252 12980
rect 14832 12860 14884 12912
rect 19432 12928 19484 12980
rect 20076 12928 20128 12980
rect 21180 12928 21232 12980
rect 21732 12928 21784 12980
rect 15292 12792 15344 12844
rect 15844 12792 15896 12844
rect 16856 12835 16908 12844
rect 16856 12801 16865 12835
rect 16865 12801 16899 12835
rect 16899 12801 16908 12835
rect 16856 12792 16908 12801
rect 19524 12903 19576 12912
rect 19524 12869 19533 12903
rect 19533 12869 19567 12903
rect 19567 12869 19576 12903
rect 19524 12860 19576 12869
rect 18420 12792 18472 12844
rect 22744 12928 22796 12980
rect 23112 12860 23164 12912
rect 24400 12860 24452 12912
rect 21088 12835 21140 12844
rect 21088 12801 21119 12835
rect 21119 12801 21140 12835
rect 21088 12792 21140 12801
rect 21456 12835 21508 12844
rect 21456 12801 21465 12835
rect 21465 12801 21499 12835
rect 21499 12801 21508 12835
rect 21456 12792 21508 12801
rect 22100 12792 22152 12844
rect 22468 12792 22520 12844
rect 20260 12656 20312 12708
rect 3056 12588 3108 12640
rect 10140 12631 10192 12640
rect 10140 12597 10149 12631
rect 10149 12597 10183 12631
rect 10183 12597 10192 12631
rect 10140 12588 10192 12597
rect 14648 12588 14700 12640
rect 15108 12631 15160 12640
rect 15108 12597 15117 12631
rect 15117 12597 15151 12631
rect 15151 12597 15160 12631
rect 15108 12588 15160 12597
rect 19616 12588 19668 12640
rect 19984 12631 20036 12640
rect 19984 12597 19993 12631
rect 19993 12597 20027 12631
rect 20027 12597 20036 12631
rect 19984 12588 20036 12597
rect 21364 12588 21416 12640
rect 23204 12724 23256 12776
rect 24308 12792 24360 12844
rect 25872 12928 25924 12980
rect 26148 12860 26200 12912
rect 24400 12767 24452 12776
rect 24400 12733 24409 12767
rect 24409 12733 24443 12767
rect 24443 12733 24452 12767
rect 24400 12724 24452 12733
rect 24492 12767 24544 12776
rect 24492 12733 24501 12767
rect 24501 12733 24535 12767
rect 24535 12733 24544 12767
rect 24492 12724 24544 12733
rect 23756 12588 23808 12640
rect 24860 12724 24912 12776
rect 24768 12656 24820 12708
rect 25596 12792 25648 12844
rect 26332 12792 26384 12844
rect 26700 12928 26752 12980
rect 26976 12928 27028 12980
rect 29644 12928 29696 12980
rect 31208 12971 31260 12980
rect 31208 12937 31217 12971
rect 31217 12937 31251 12971
rect 31251 12937 31260 12971
rect 31208 12928 31260 12937
rect 31852 12971 31904 12980
rect 31852 12937 31861 12971
rect 31861 12937 31895 12971
rect 31895 12937 31904 12971
rect 31852 12928 31904 12937
rect 32864 12971 32916 12980
rect 32864 12937 32873 12971
rect 32873 12937 32907 12971
rect 32907 12937 32916 12971
rect 32864 12928 32916 12937
rect 33140 12928 33192 12980
rect 25228 12767 25280 12776
rect 25228 12733 25237 12767
rect 25237 12733 25271 12767
rect 25271 12733 25280 12767
rect 25228 12724 25280 12733
rect 30380 12792 30432 12844
rect 28448 12724 28500 12776
rect 25136 12631 25188 12640
rect 25136 12597 25145 12631
rect 25145 12597 25179 12631
rect 25179 12597 25188 12631
rect 25136 12588 25188 12597
rect 26240 12656 26292 12708
rect 29000 12656 29052 12708
rect 29092 12656 29144 12708
rect 29920 12656 29972 12708
rect 26884 12588 26936 12640
rect 27160 12588 27212 12640
rect 30012 12588 30064 12640
rect 30288 12724 30340 12776
rect 31300 12792 31352 12844
rect 31392 12835 31444 12844
rect 31392 12801 31401 12835
rect 31401 12801 31435 12835
rect 31435 12801 31444 12835
rect 31392 12792 31444 12801
rect 32404 12792 32456 12844
rect 33876 12792 33928 12844
rect 32496 12724 32548 12776
rect 33324 12724 33376 12776
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 1676 12384 1728 12436
rect 3792 12427 3844 12436
rect 3792 12393 3801 12427
rect 3801 12393 3835 12427
rect 3835 12393 3844 12427
rect 3792 12384 3844 12393
rect 4068 12384 4120 12436
rect 4620 12384 4672 12436
rect 5816 12384 5868 12436
rect 8852 12384 8904 12436
rect 10232 12384 10284 12436
rect 11152 12384 11204 12436
rect 16856 12427 16908 12436
rect 16856 12393 16865 12427
rect 16865 12393 16899 12427
rect 16899 12393 16908 12427
rect 16856 12384 16908 12393
rect 21916 12384 21968 12436
rect 3056 12291 3108 12300
rect 3056 12257 3065 12291
rect 3065 12257 3099 12291
rect 3099 12257 3108 12291
rect 3056 12248 3108 12257
rect 3240 12291 3292 12300
rect 3240 12257 3249 12291
rect 3249 12257 3283 12291
rect 3283 12257 3292 12291
rect 3240 12248 3292 12257
rect 4068 12248 4120 12300
rect 6276 12248 6328 12300
rect 7104 12291 7156 12300
rect 7104 12257 7113 12291
rect 7113 12257 7147 12291
rect 7147 12257 7156 12291
rect 7104 12248 7156 12257
rect 3148 12112 3200 12164
rect 3424 12044 3476 12096
rect 8024 12180 8076 12232
rect 12532 12248 12584 12300
rect 15752 12248 15804 12300
rect 22836 12316 22888 12368
rect 8300 12180 8352 12232
rect 8760 12180 8812 12232
rect 9404 12180 9456 12232
rect 10048 12180 10100 12232
rect 10232 12180 10284 12232
rect 12256 12180 12308 12232
rect 14832 12180 14884 12232
rect 15108 12223 15160 12232
rect 15108 12189 15117 12223
rect 15117 12189 15151 12223
rect 15151 12189 15160 12223
rect 15108 12180 15160 12189
rect 16488 12180 16540 12232
rect 7840 12044 7892 12096
rect 15292 12044 15344 12096
rect 17684 12112 17736 12164
rect 18420 12291 18472 12300
rect 18420 12257 18429 12291
rect 18429 12257 18463 12291
rect 18463 12257 18472 12291
rect 18420 12248 18472 12257
rect 18328 12180 18380 12232
rect 18880 12248 18932 12300
rect 20812 12248 20864 12300
rect 20904 12248 20956 12300
rect 21548 12248 21600 12300
rect 18788 12180 18840 12232
rect 19340 12223 19392 12232
rect 19340 12189 19349 12223
rect 19349 12189 19383 12223
rect 19383 12189 19392 12223
rect 19340 12180 19392 12189
rect 21456 12180 21508 12232
rect 23020 12291 23072 12300
rect 23020 12257 23029 12291
rect 23029 12257 23063 12291
rect 23063 12257 23072 12291
rect 23020 12248 23072 12257
rect 23204 12291 23256 12300
rect 23204 12257 23213 12291
rect 23213 12257 23247 12291
rect 23247 12257 23256 12291
rect 23204 12248 23256 12257
rect 20076 12112 20128 12164
rect 22100 12112 22152 12164
rect 17592 12044 17644 12096
rect 19524 12087 19576 12096
rect 19524 12053 19533 12087
rect 19533 12053 19567 12087
rect 19567 12053 19576 12087
rect 19524 12044 19576 12053
rect 22192 12044 22244 12096
rect 24216 12384 24268 12436
rect 24400 12384 24452 12436
rect 25136 12384 25188 12436
rect 25228 12427 25280 12436
rect 25228 12393 25237 12427
rect 25237 12393 25271 12427
rect 25271 12393 25280 12427
rect 25228 12384 25280 12393
rect 26792 12384 26844 12436
rect 29736 12384 29788 12436
rect 31760 12384 31812 12436
rect 32772 12384 32824 12436
rect 26516 12316 26568 12368
rect 27804 12316 27856 12368
rect 32680 12316 32732 12368
rect 24768 12248 24820 12300
rect 26148 12248 26200 12300
rect 28908 12248 28960 12300
rect 25044 12180 25096 12232
rect 26424 12223 26476 12232
rect 26424 12189 26433 12223
rect 26433 12189 26467 12223
rect 26467 12189 26476 12223
rect 26424 12180 26476 12189
rect 26792 12180 26844 12232
rect 30012 12223 30064 12232
rect 30012 12189 30021 12223
rect 30021 12189 30055 12223
rect 30055 12189 30064 12223
rect 30012 12180 30064 12189
rect 30288 12223 30340 12232
rect 30288 12189 30297 12223
rect 30297 12189 30331 12223
rect 30331 12189 30340 12223
rect 30288 12180 30340 12189
rect 32312 12248 32364 12300
rect 26056 12044 26108 12096
rect 26608 12044 26660 12096
rect 28172 12044 28224 12096
rect 28908 12044 28960 12096
rect 32036 12180 32088 12232
rect 32956 12180 33008 12232
rect 33600 12180 33652 12232
rect 30380 12044 30432 12096
rect 30472 12087 30524 12096
rect 30472 12053 30481 12087
rect 30481 12053 30515 12087
rect 30515 12053 30524 12087
rect 30472 12044 30524 12053
rect 32588 12044 32640 12096
rect 4874 11942 4926 11994
rect 4938 11942 4990 11994
rect 5002 11942 5054 11994
rect 5066 11942 5118 11994
rect 5130 11942 5182 11994
rect 35594 11942 35646 11994
rect 35658 11942 35710 11994
rect 35722 11942 35774 11994
rect 35786 11942 35838 11994
rect 35850 11942 35902 11994
rect 8208 11840 8260 11892
rect 8760 11840 8812 11892
rect 9312 11840 9364 11892
rect 940 11704 992 11756
rect 9312 11704 9364 11756
rect 11060 11772 11112 11824
rect 13544 11840 13596 11892
rect 15292 11840 15344 11892
rect 12992 11772 13044 11824
rect 14464 11772 14516 11824
rect 20352 11840 20404 11892
rect 24216 11840 24268 11892
rect 26792 11840 26844 11892
rect 27620 11840 27672 11892
rect 29092 11840 29144 11892
rect 15844 11772 15896 11824
rect 10784 11747 10836 11756
rect 10784 11713 10793 11747
rect 10793 11713 10827 11747
rect 10827 11713 10836 11747
rect 10784 11704 10836 11713
rect 11888 11704 11940 11756
rect 11980 11747 12032 11756
rect 11980 11713 11989 11747
rect 11989 11713 12023 11747
rect 12023 11713 12032 11747
rect 11980 11704 12032 11713
rect 14832 11704 14884 11756
rect 10324 11636 10376 11688
rect 10876 11679 10928 11688
rect 10876 11645 10885 11679
rect 10885 11645 10919 11679
rect 10919 11645 10928 11679
rect 10876 11636 10928 11645
rect 12256 11679 12308 11688
rect 12256 11645 12265 11679
rect 12265 11645 12299 11679
rect 12299 11645 12308 11679
rect 12256 11636 12308 11645
rect 12900 11636 12952 11688
rect 14740 11636 14792 11688
rect 9496 11568 9548 11620
rect 5448 11500 5500 11552
rect 8300 11500 8352 11552
rect 10324 11543 10376 11552
rect 10324 11509 10333 11543
rect 10333 11509 10367 11543
rect 10367 11509 10376 11543
rect 10324 11500 10376 11509
rect 19156 11772 19208 11824
rect 20260 11772 20312 11824
rect 23480 11747 23532 11756
rect 23480 11713 23489 11747
rect 23489 11713 23523 11747
rect 23523 11713 23532 11747
rect 23480 11704 23532 11713
rect 23756 11747 23808 11756
rect 23756 11713 23765 11747
rect 23765 11713 23799 11747
rect 23799 11713 23808 11747
rect 23756 11704 23808 11713
rect 24216 11747 24268 11756
rect 24216 11713 24225 11747
rect 24225 11713 24259 11747
rect 24259 11713 24268 11747
rect 24216 11704 24268 11713
rect 24400 11704 24452 11756
rect 17592 11568 17644 11620
rect 18696 11611 18748 11620
rect 18696 11577 18705 11611
rect 18705 11577 18739 11611
rect 18739 11577 18748 11611
rect 18696 11568 18748 11577
rect 15568 11543 15620 11552
rect 15568 11509 15577 11543
rect 15577 11509 15611 11543
rect 15611 11509 15620 11543
rect 15568 11500 15620 11509
rect 18144 11500 18196 11552
rect 19248 11500 19300 11552
rect 23572 11636 23624 11688
rect 24584 11747 24636 11756
rect 24584 11713 24593 11747
rect 24593 11713 24627 11747
rect 24627 11713 24636 11747
rect 24584 11704 24636 11713
rect 24768 11747 24820 11756
rect 24768 11713 24777 11747
rect 24777 11713 24811 11747
rect 24811 11713 24820 11747
rect 24768 11704 24820 11713
rect 25320 11772 25372 11824
rect 25044 11747 25096 11756
rect 25044 11713 25053 11747
rect 25053 11713 25087 11747
rect 25087 11713 25096 11747
rect 25044 11704 25096 11713
rect 26608 11704 26660 11756
rect 26424 11636 26476 11688
rect 26976 11636 27028 11688
rect 27344 11747 27396 11756
rect 27344 11713 27353 11747
rect 27353 11713 27387 11747
rect 27387 11713 27396 11747
rect 27344 11704 27396 11713
rect 27804 11772 27856 11824
rect 27988 11772 28040 11824
rect 30104 11840 30156 11892
rect 30472 11840 30524 11892
rect 33048 11840 33100 11892
rect 28816 11704 28868 11756
rect 29000 11704 29052 11756
rect 27528 11611 27580 11620
rect 27528 11577 27537 11611
rect 27537 11577 27571 11611
rect 27571 11577 27580 11611
rect 27528 11568 27580 11577
rect 30380 11772 30432 11824
rect 29736 11704 29788 11756
rect 32588 11747 32640 11756
rect 32588 11713 32597 11747
rect 32597 11713 32631 11747
rect 32631 11713 32640 11747
rect 32588 11704 32640 11713
rect 32680 11747 32732 11756
rect 32680 11713 32689 11747
rect 32689 11713 32723 11747
rect 32723 11713 32732 11747
rect 32680 11704 32732 11713
rect 29828 11679 29880 11688
rect 29828 11645 29837 11679
rect 29837 11645 29871 11679
rect 29871 11645 29880 11679
rect 29828 11636 29880 11645
rect 30656 11679 30708 11688
rect 30656 11645 30665 11679
rect 30665 11645 30699 11679
rect 30699 11645 30708 11679
rect 30656 11636 30708 11645
rect 32220 11636 32272 11688
rect 23388 11500 23440 11552
rect 26056 11500 26108 11552
rect 26700 11500 26752 11552
rect 34612 11568 34664 11620
rect 27712 11543 27764 11552
rect 27712 11509 27721 11543
rect 27721 11509 27755 11543
rect 27755 11509 27764 11543
rect 27712 11500 27764 11509
rect 29092 11500 29144 11552
rect 30380 11500 30432 11552
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 3148 11339 3200 11348
rect 3148 11305 3157 11339
rect 3157 11305 3191 11339
rect 3191 11305 3200 11339
rect 3148 11296 3200 11305
rect 3424 11296 3476 11348
rect 5724 11339 5776 11348
rect 5724 11305 5733 11339
rect 5733 11305 5767 11339
rect 5767 11305 5776 11339
rect 5724 11296 5776 11305
rect 7840 11296 7892 11348
rect 9036 11296 9088 11348
rect 3884 11228 3936 11280
rect 4068 11160 4120 11212
rect 5540 11160 5592 11212
rect 5908 11135 5960 11144
rect 5908 11101 5917 11135
rect 5917 11101 5951 11135
rect 5951 11101 5960 11135
rect 5908 11092 5960 11101
rect 6092 11135 6144 11144
rect 6092 11101 6101 11135
rect 6101 11101 6135 11135
rect 6135 11101 6144 11135
rect 6092 11092 6144 11101
rect 1676 11067 1728 11076
rect 1676 11033 1685 11067
rect 1685 11033 1719 11067
rect 1719 11033 1728 11067
rect 1676 11024 1728 11033
rect 2964 11024 3016 11076
rect 3884 11024 3936 11076
rect 5816 11024 5868 11076
rect 7472 11135 7524 11144
rect 7472 11101 7481 11135
rect 7481 11101 7515 11135
rect 7515 11101 7524 11135
rect 7472 11092 7524 11101
rect 9312 11271 9364 11280
rect 9312 11237 9321 11271
rect 9321 11237 9355 11271
rect 9355 11237 9364 11271
rect 9312 11228 9364 11237
rect 9496 11228 9548 11280
rect 8208 11160 8260 11212
rect 8852 11160 8904 11212
rect 8576 11135 8628 11144
rect 8576 11101 8585 11135
rect 8585 11101 8619 11135
rect 8619 11101 8628 11135
rect 8576 11092 8628 11101
rect 9036 11092 9088 11144
rect 9404 11135 9456 11144
rect 9404 11101 9413 11135
rect 9413 11101 9447 11135
rect 9447 11101 9456 11135
rect 9404 11092 9456 11101
rect 10324 11296 10376 11348
rect 11980 11296 12032 11348
rect 14464 11296 14516 11348
rect 9864 11160 9916 11212
rect 10784 11160 10836 11212
rect 12532 11160 12584 11212
rect 11704 11092 11756 11144
rect 12440 11092 12492 11144
rect 13360 11092 13412 11144
rect 7840 11024 7892 11076
rect 8116 11024 8168 11076
rect 12900 11067 12952 11076
rect 12900 11033 12909 11067
rect 12909 11033 12943 11067
rect 12943 11033 12952 11067
rect 12900 11024 12952 11033
rect 14648 11203 14700 11212
rect 14648 11169 14657 11203
rect 14657 11169 14691 11203
rect 14691 11169 14700 11203
rect 14648 11160 14700 11169
rect 14832 11160 14884 11212
rect 15568 11135 15620 11144
rect 15568 11101 15577 11135
rect 15577 11101 15611 11135
rect 15611 11101 15620 11135
rect 15568 11092 15620 11101
rect 16120 11296 16172 11348
rect 17592 11339 17644 11348
rect 17592 11305 17601 11339
rect 17601 11305 17635 11339
rect 17635 11305 17644 11339
rect 17592 11296 17644 11305
rect 22100 11296 22152 11348
rect 23388 11296 23440 11348
rect 23480 11296 23532 11348
rect 26516 11296 26568 11348
rect 27344 11296 27396 11348
rect 27620 11296 27672 11348
rect 29184 11296 29236 11348
rect 30104 11296 30156 11348
rect 30380 11296 30432 11348
rect 30472 11296 30524 11348
rect 30656 11296 30708 11348
rect 32128 11339 32180 11348
rect 32128 11305 32137 11339
rect 32137 11305 32171 11339
rect 32171 11305 32180 11339
rect 32128 11296 32180 11305
rect 34612 11296 34664 11348
rect 19248 11228 19300 11280
rect 19892 11228 19944 11280
rect 22284 11228 22336 11280
rect 22468 11228 22520 11280
rect 18328 11092 18380 11144
rect 19524 11092 19576 11144
rect 20536 11160 20588 11212
rect 18512 11024 18564 11076
rect 20076 11135 20128 11144
rect 20076 11101 20085 11135
rect 20085 11101 20119 11135
rect 20119 11101 20128 11135
rect 20076 11092 20128 11101
rect 20996 11024 21048 11076
rect 22192 11135 22244 11144
rect 22192 11101 22201 11135
rect 22201 11101 22235 11135
rect 22235 11101 22244 11135
rect 22192 11092 22244 11101
rect 23388 11092 23440 11144
rect 23572 11228 23624 11280
rect 24584 11228 24636 11280
rect 25044 11160 25096 11212
rect 24308 11092 24360 11144
rect 26148 11092 26200 11144
rect 26424 11135 26476 11144
rect 26424 11101 26433 11135
rect 26433 11101 26467 11135
rect 26467 11101 26476 11135
rect 26424 11092 26476 11101
rect 26516 11092 26568 11144
rect 3792 10999 3844 11008
rect 3792 10965 3801 10999
rect 3801 10965 3835 10999
rect 3835 10965 3844 10999
rect 3792 10956 3844 10965
rect 4252 10999 4304 11008
rect 4252 10965 4261 10999
rect 4261 10965 4295 10999
rect 4295 10965 4304 10999
rect 4252 10956 4304 10965
rect 7564 10956 7616 11008
rect 14096 10956 14148 11008
rect 15108 10956 15160 11008
rect 15752 10956 15804 11008
rect 16488 10956 16540 11008
rect 20168 10956 20220 11008
rect 22100 11024 22152 11076
rect 24216 11024 24268 11076
rect 27068 11135 27120 11144
rect 27068 11101 27077 11135
rect 27077 11101 27111 11135
rect 27111 11101 27120 11135
rect 27068 11092 27120 11101
rect 27712 11228 27764 11280
rect 27160 11024 27212 11076
rect 27804 11092 27856 11144
rect 27896 11135 27948 11144
rect 27896 11101 27905 11135
rect 27905 11101 27939 11135
rect 27939 11101 27948 11135
rect 27896 11092 27948 11101
rect 31760 11228 31812 11280
rect 29092 11135 29144 11144
rect 29092 11101 29101 11135
rect 29101 11101 29135 11135
rect 29135 11101 29144 11135
rect 29092 11092 29144 11101
rect 30012 11024 30064 11076
rect 30288 11135 30340 11144
rect 30288 11101 30297 11135
rect 30297 11101 30331 11135
rect 30331 11101 30340 11135
rect 30288 11092 30340 11101
rect 31852 11135 31904 11144
rect 31852 11101 31861 11135
rect 31861 11101 31895 11135
rect 31895 11101 31904 11135
rect 31852 11092 31904 11101
rect 32312 11135 32364 11144
rect 32312 11101 32321 11135
rect 32321 11101 32355 11135
rect 32355 11101 32364 11135
rect 32312 11092 32364 11101
rect 32496 11092 32548 11144
rect 32772 11135 32824 11144
rect 32772 11101 32781 11135
rect 32781 11101 32815 11135
rect 32815 11101 32824 11135
rect 32772 11092 32824 11101
rect 33048 11135 33100 11144
rect 33048 11101 33057 11135
rect 33057 11101 33091 11135
rect 33091 11101 33100 11135
rect 33048 11092 33100 11101
rect 21824 10956 21876 11008
rect 23388 10999 23440 11008
rect 23388 10965 23397 10999
rect 23397 10965 23431 10999
rect 23431 10965 23440 10999
rect 23388 10956 23440 10965
rect 26056 10956 26108 11008
rect 26792 10999 26844 11008
rect 26792 10965 26801 10999
rect 26801 10965 26835 10999
rect 26835 10965 26844 10999
rect 26792 10956 26844 10965
rect 27620 10999 27672 11008
rect 27620 10965 27629 10999
rect 27629 10965 27663 10999
rect 27663 10965 27672 10999
rect 27620 10956 27672 10965
rect 37924 11067 37976 11076
rect 37924 11033 37933 11067
rect 37933 11033 37967 11067
rect 37967 11033 37976 11067
rect 37924 11024 37976 11033
rect 30656 10956 30708 11008
rect 32864 10956 32916 11008
rect 4874 10854 4926 10906
rect 4938 10854 4990 10906
rect 5002 10854 5054 10906
rect 5066 10854 5118 10906
rect 5130 10854 5182 10906
rect 35594 10854 35646 10906
rect 35658 10854 35710 10906
rect 35722 10854 35774 10906
rect 35786 10854 35838 10906
rect 35850 10854 35902 10906
rect 1676 10752 1728 10804
rect 3792 10752 3844 10804
rect 3884 10752 3936 10804
rect 3148 10616 3200 10668
rect 3424 10591 3476 10600
rect 3424 10557 3433 10591
rect 3433 10557 3467 10591
rect 3467 10557 3476 10591
rect 3424 10548 3476 10557
rect 4252 10684 4304 10736
rect 6092 10752 6144 10804
rect 8944 10752 8996 10804
rect 9404 10752 9456 10804
rect 5724 10616 5776 10668
rect 6184 10659 6236 10668
rect 6184 10625 6193 10659
rect 6193 10625 6227 10659
rect 6227 10625 6236 10659
rect 6184 10616 6236 10625
rect 6736 10659 6788 10668
rect 6736 10625 6745 10659
rect 6745 10625 6779 10659
rect 6779 10625 6788 10659
rect 6736 10616 6788 10625
rect 4068 10591 4120 10600
rect 4068 10557 4077 10591
rect 4077 10557 4111 10591
rect 4111 10557 4120 10591
rect 4068 10548 4120 10557
rect 4712 10548 4764 10600
rect 5540 10548 5592 10600
rect 5816 10548 5868 10600
rect 13820 10684 13872 10736
rect 7196 10659 7248 10668
rect 7196 10625 7205 10659
rect 7205 10625 7239 10659
rect 7239 10625 7248 10659
rect 7196 10616 7248 10625
rect 8852 10659 8904 10668
rect 8852 10625 8861 10659
rect 8861 10625 8895 10659
rect 8895 10625 8904 10659
rect 8852 10616 8904 10625
rect 10784 10616 10836 10668
rect 11520 10616 11572 10668
rect 12256 10616 12308 10668
rect 15108 10752 15160 10804
rect 19156 10795 19208 10804
rect 19156 10761 19165 10795
rect 19165 10761 19199 10795
rect 19199 10761 19208 10795
rect 19156 10752 19208 10761
rect 14096 10684 14148 10736
rect 16120 10684 16172 10736
rect 20720 10752 20772 10804
rect 22376 10752 22428 10804
rect 27620 10752 27672 10804
rect 28724 10752 28776 10804
rect 32128 10752 32180 10804
rect 32312 10752 32364 10804
rect 15292 10616 15344 10668
rect 10232 10548 10284 10600
rect 11244 10591 11296 10600
rect 11244 10557 11253 10591
rect 11253 10557 11287 10591
rect 11287 10557 11296 10591
rect 11244 10548 11296 10557
rect 16948 10616 17000 10668
rect 3240 10412 3292 10464
rect 5816 10412 5868 10464
rect 6368 10455 6420 10464
rect 6368 10421 6377 10455
rect 6377 10421 6411 10455
rect 6411 10421 6420 10455
rect 6368 10412 6420 10421
rect 7932 10412 7984 10464
rect 8208 10412 8260 10464
rect 8300 10412 8352 10464
rect 13820 10412 13872 10464
rect 17132 10659 17184 10668
rect 17132 10625 17141 10659
rect 17141 10625 17175 10659
rect 17175 10625 17184 10659
rect 17132 10616 17184 10625
rect 17500 10523 17552 10532
rect 17500 10489 17509 10523
rect 17509 10489 17543 10523
rect 17543 10489 17552 10523
rect 17500 10480 17552 10489
rect 18328 10659 18380 10668
rect 18328 10625 18337 10659
rect 18337 10625 18371 10659
rect 18371 10625 18380 10659
rect 18328 10616 18380 10625
rect 18512 10616 18564 10668
rect 20996 10727 21048 10736
rect 20996 10693 21021 10727
rect 21021 10693 21048 10727
rect 20996 10684 21048 10693
rect 22008 10684 22060 10736
rect 22836 10684 22888 10736
rect 23112 10727 23164 10736
rect 23112 10693 23121 10727
rect 23121 10693 23155 10727
rect 23155 10693 23164 10727
rect 23112 10684 23164 10693
rect 23388 10684 23440 10736
rect 21180 10548 21232 10600
rect 21640 10591 21692 10600
rect 21640 10557 21649 10591
rect 21649 10557 21683 10591
rect 21683 10557 21692 10591
rect 21640 10548 21692 10557
rect 22652 10616 22704 10668
rect 22744 10616 22796 10668
rect 22928 10659 22980 10668
rect 22928 10625 22937 10659
rect 22937 10625 22971 10659
rect 22971 10625 22980 10659
rect 22928 10616 22980 10625
rect 22192 10480 22244 10532
rect 22376 10480 22428 10532
rect 18052 10455 18104 10464
rect 18052 10421 18061 10455
rect 18061 10421 18095 10455
rect 18095 10421 18104 10455
rect 18052 10412 18104 10421
rect 20168 10455 20220 10464
rect 20168 10421 20177 10455
rect 20177 10421 20211 10455
rect 20211 10421 20220 10455
rect 20168 10412 20220 10421
rect 21088 10412 21140 10464
rect 21456 10412 21508 10464
rect 21548 10412 21600 10464
rect 22008 10412 22060 10464
rect 23112 10548 23164 10600
rect 24400 10616 24452 10668
rect 26792 10616 26844 10668
rect 29092 10684 29144 10736
rect 27252 10659 27304 10668
rect 27252 10625 27261 10659
rect 27261 10625 27295 10659
rect 27295 10625 27304 10659
rect 27252 10616 27304 10625
rect 27528 10616 27580 10668
rect 28172 10659 28224 10668
rect 28172 10625 28181 10659
rect 28181 10625 28215 10659
rect 28215 10625 28224 10659
rect 28172 10616 28224 10625
rect 28264 10616 28316 10668
rect 23664 10548 23716 10600
rect 24492 10548 24544 10600
rect 30196 10616 30248 10668
rect 31300 10684 31352 10736
rect 32588 10752 32640 10804
rect 32680 10752 32732 10804
rect 35348 10752 35400 10804
rect 31852 10616 31904 10668
rect 32220 10616 32272 10668
rect 33232 10684 33284 10736
rect 33600 10684 33652 10736
rect 32772 10616 32824 10668
rect 33508 10659 33560 10668
rect 33508 10625 33517 10659
rect 33517 10625 33551 10659
rect 33551 10625 33560 10659
rect 33508 10616 33560 10625
rect 23572 10480 23624 10532
rect 26424 10480 26476 10532
rect 22744 10455 22796 10464
rect 22744 10421 22753 10455
rect 22753 10421 22787 10455
rect 22787 10421 22796 10455
rect 22744 10412 22796 10421
rect 23480 10412 23532 10464
rect 23848 10412 23900 10464
rect 26608 10412 26660 10464
rect 27620 10455 27672 10464
rect 27620 10421 27629 10455
rect 27629 10421 27663 10455
rect 27663 10421 27672 10455
rect 27620 10412 27672 10421
rect 28540 10480 28592 10532
rect 28724 10523 28776 10532
rect 28724 10489 28733 10523
rect 28733 10489 28767 10523
rect 28767 10489 28776 10523
rect 28724 10480 28776 10489
rect 29000 10548 29052 10600
rect 32496 10591 32548 10600
rect 32496 10557 32505 10591
rect 32505 10557 32539 10591
rect 32539 10557 32548 10591
rect 32496 10548 32548 10557
rect 30288 10412 30340 10464
rect 32956 10412 33008 10464
rect 34428 10616 34480 10668
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 4712 10208 4764 10260
rect 6184 10251 6236 10260
rect 6184 10217 6193 10251
rect 6193 10217 6227 10251
rect 6227 10217 6236 10251
rect 6184 10208 6236 10217
rect 6368 10208 6420 10260
rect 7564 10251 7616 10260
rect 7564 10217 7573 10251
rect 7573 10217 7607 10251
rect 7607 10217 7616 10251
rect 7564 10208 7616 10217
rect 9956 10208 10008 10260
rect 10508 10208 10560 10260
rect 13084 10208 13136 10260
rect 14464 10208 14516 10260
rect 17132 10208 17184 10260
rect 7472 10140 7524 10192
rect 8392 10140 8444 10192
rect 5816 10115 5868 10124
rect 5816 10081 5825 10115
rect 5825 10081 5859 10115
rect 5859 10081 5868 10115
rect 5816 10072 5868 10081
rect 5908 10072 5960 10124
rect 3148 10004 3200 10056
rect 3056 9936 3108 9988
rect 3148 9911 3200 9920
rect 3148 9877 3157 9911
rect 3157 9877 3191 9911
rect 3191 9877 3200 9911
rect 3148 9868 3200 9877
rect 6092 10004 6144 10056
rect 8208 10072 8260 10124
rect 8668 10072 8720 10124
rect 9772 10072 9824 10124
rect 7932 10004 7984 10056
rect 8024 10004 8076 10056
rect 8944 10004 8996 10056
rect 13176 10072 13228 10124
rect 13268 10072 13320 10124
rect 5632 9868 5684 9920
rect 5816 9868 5868 9920
rect 8484 9936 8536 9988
rect 11428 10047 11480 10056
rect 11428 10013 11437 10047
rect 11437 10013 11471 10047
rect 11471 10013 11480 10047
rect 11428 10004 11480 10013
rect 11520 10004 11572 10056
rect 13452 10004 13504 10056
rect 16672 10004 16724 10056
rect 9496 9911 9548 9920
rect 9496 9877 9505 9911
rect 9505 9877 9539 9911
rect 9539 9877 9548 9911
rect 9496 9868 9548 9877
rect 12992 9936 13044 9988
rect 18144 10072 18196 10124
rect 22008 10208 22060 10260
rect 22376 10251 22428 10260
rect 22376 10217 22385 10251
rect 22385 10217 22419 10251
rect 22419 10217 22428 10251
rect 22376 10208 22428 10217
rect 22560 10208 22612 10260
rect 22652 10251 22704 10260
rect 22652 10217 22661 10251
rect 22661 10217 22695 10251
rect 22695 10217 22704 10251
rect 22652 10208 22704 10217
rect 22744 10208 22796 10260
rect 27252 10208 27304 10260
rect 27896 10208 27948 10260
rect 28448 10208 28500 10260
rect 30564 10208 30616 10260
rect 32772 10208 32824 10260
rect 33508 10251 33560 10260
rect 33508 10217 33517 10251
rect 33517 10217 33551 10251
rect 33551 10217 33560 10251
rect 33508 10208 33560 10217
rect 18052 10047 18104 10056
rect 18052 10013 18061 10047
rect 18061 10013 18095 10047
rect 18095 10013 18104 10047
rect 18052 10004 18104 10013
rect 18236 10047 18288 10056
rect 18236 10013 18245 10047
rect 18245 10013 18279 10047
rect 18279 10013 18288 10047
rect 18236 10004 18288 10013
rect 18420 10047 18472 10056
rect 18420 10013 18429 10047
rect 18429 10013 18463 10047
rect 18463 10013 18472 10047
rect 18420 10004 18472 10013
rect 18512 10004 18564 10056
rect 20168 10004 20220 10056
rect 20536 10047 20588 10056
rect 20536 10013 20545 10047
rect 20545 10013 20579 10047
rect 20579 10013 20588 10047
rect 20536 10004 20588 10013
rect 20628 10004 20680 10056
rect 21180 10004 21232 10056
rect 21456 10004 21508 10056
rect 22192 10140 22244 10192
rect 25964 10140 26016 10192
rect 29092 10140 29144 10192
rect 30386 10140 30438 10192
rect 21916 10047 21968 10056
rect 21916 10013 21925 10047
rect 21925 10013 21959 10047
rect 21959 10013 21968 10047
rect 21916 10004 21968 10013
rect 22284 10047 22336 10056
rect 22284 10013 22293 10047
rect 22293 10013 22327 10047
rect 22327 10013 22336 10047
rect 22284 10004 22336 10013
rect 18696 9911 18748 9920
rect 18696 9877 18705 9911
rect 18705 9877 18739 9911
rect 18739 9877 18748 9911
rect 18696 9868 18748 9877
rect 20076 9868 20128 9920
rect 20904 9936 20956 9988
rect 24400 10072 24452 10124
rect 25044 10072 25096 10124
rect 27620 10072 27672 10124
rect 23940 10004 23992 10056
rect 26240 10004 26292 10056
rect 28264 10004 28316 10056
rect 28724 10047 28776 10056
rect 28724 10013 28733 10047
rect 28733 10013 28767 10047
rect 28767 10013 28776 10047
rect 28724 10004 28776 10013
rect 28816 10004 28868 10056
rect 30288 10047 30340 10056
rect 30288 10013 30297 10047
rect 30297 10013 30331 10047
rect 30331 10013 30340 10047
rect 30288 10004 30340 10013
rect 32956 10072 33008 10124
rect 30656 10047 30708 10056
rect 30656 10013 30665 10047
rect 30665 10013 30699 10047
rect 30699 10013 30708 10047
rect 30656 10004 30708 10013
rect 32864 10004 32916 10056
rect 23756 9936 23808 9988
rect 29000 9936 29052 9988
rect 33968 10047 34020 10056
rect 33968 10013 33977 10047
rect 33977 10013 34011 10047
rect 34011 10013 34020 10047
rect 33968 10004 34020 10013
rect 34060 10004 34112 10056
rect 21824 9911 21876 9920
rect 21824 9877 21833 9911
rect 21833 9877 21867 9911
rect 21867 9877 21876 9911
rect 21824 9868 21876 9877
rect 22100 9868 22152 9920
rect 26148 9868 26200 9920
rect 27896 9868 27948 9920
rect 30840 9911 30892 9920
rect 30840 9877 30849 9911
rect 30849 9877 30883 9911
rect 30883 9877 30892 9911
rect 30840 9868 30892 9877
rect 4874 9766 4926 9818
rect 4938 9766 4990 9818
rect 5002 9766 5054 9818
rect 5066 9766 5118 9818
rect 5130 9766 5182 9818
rect 35594 9766 35646 9818
rect 35658 9766 35710 9818
rect 35722 9766 35774 9818
rect 35786 9766 35838 9818
rect 35850 9766 35902 9818
rect 3148 9664 3200 9716
rect 3240 9571 3292 9580
rect 3240 9537 3249 9571
rect 3249 9537 3283 9571
rect 3283 9537 3292 9571
rect 3240 9528 3292 9537
rect 3332 9571 3384 9580
rect 3332 9537 3341 9571
rect 3341 9537 3375 9571
rect 3375 9537 3384 9571
rect 3332 9528 3384 9537
rect 6000 9596 6052 9648
rect 3700 9528 3752 9580
rect 4620 9528 4672 9580
rect 6644 9571 6696 9580
rect 6644 9537 6653 9571
rect 6653 9537 6687 9571
rect 6687 9537 6696 9571
rect 6644 9528 6696 9537
rect 6736 9571 6788 9580
rect 6736 9537 6745 9571
rect 6745 9537 6779 9571
rect 6779 9537 6788 9571
rect 6736 9528 6788 9537
rect 6828 9571 6880 9580
rect 6828 9537 6837 9571
rect 6837 9537 6871 9571
rect 6871 9537 6880 9571
rect 6828 9528 6880 9537
rect 8208 9596 8260 9648
rect 11428 9664 11480 9716
rect 13176 9664 13228 9716
rect 15292 9664 15344 9716
rect 7840 9528 7892 9580
rect 8116 9528 8168 9580
rect 8484 9571 8536 9580
rect 8484 9537 8493 9571
rect 8493 9537 8527 9571
rect 8527 9537 8536 9571
rect 8484 9528 8536 9537
rect 8944 9528 8996 9580
rect 9312 9596 9364 9648
rect 16028 9707 16080 9716
rect 16028 9673 16037 9707
rect 16037 9673 16071 9707
rect 16071 9673 16080 9707
rect 16028 9664 16080 9673
rect 18696 9664 18748 9716
rect 9956 9528 10008 9580
rect 7472 9435 7524 9444
rect 7472 9401 7481 9435
rect 7481 9401 7515 9435
rect 7515 9401 7524 9435
rect 7472 9392 7524 9401
rect 8208 9392 8260 9444
rect 10508 9528 10560 9580
rect 2964 9367 3016 9376
rect 2964 9333 2973 9367
rect 2973 9333 3007 9367
rect 3007 9333 3016 9367
rect 2964 9324 3016 9333
rect 6736 9324 6788 9376
rect 10048 9367 10100 9376
rect 10048 9333 10057 9367
rect 10057 9333 10091 9367
rect 10091 9333 10100 9367
rect 10048 9324 10100 9333
rect 11612 9528 11664 9580
rect 10876 9503 10928 9512
rect 10876 9469 10885 9503
rect 10885 9469 10919 9503
rect 10919 9469 10928 9503
rect 10876 9460 10928 9469
rect 13268 9528 13320 9580
rect 12532 9460 12584 9512
rect 15568 9571 15620 9580
rect 15568 9537 15577 9571
rect 15577 9537 15611 9571
rect 15611 9537 15620 9571
rect 15568 9528 15620 9537
rect 15936 9528 15988 9580
rect 16672 9528 16724 9580
rect 16948 9528 17000 9580
rect 10508 9324 10560 9376
rect 13084 9367 13136 9376
rect 13084 9333 13093 9367
rect 13093 9333 13127 9367
rect 13127 9333 13136 9367
rect 13084 9324 13136 9333
rect 13452 9324 13504 9376
rect 13728 9392 13780 9444
rect 15844 9392 15896 9444
rect 15936 9435 15988 9444
rect 15936 9401 15945 9435
rect 15945 9401 15979 9435
rect 15979 9401 15988 9435
rect 15936 9392 15988 9401
rect 17132 9503 17184 9512
rect 17132 9469 17141 9503
rect 17141 9469 17175 9503
rect 17175 9469 17184 9503
rect 17132 9460 17184 9469
rect 18052 9528 18104 9580
rect 18512 9528 18564 9580
rect 19984 9596 20036 9648
rect 21088 9596 21140 9648
rect 21640 9596 21692 9648
rect 22376 9664 22428 9716
rect 23940 9664 23992 9716
rect 24032 9664 24084 9716
rect 28816 9664 28868 9716
rect 20168 9528 20220 9580
rect 20260 9528 20312 9580
rect 20536 9528 20588 9580
rect 18236 9503 18288 9512
rect 18236 9469 18245 9503
rect 18245 9469 18279 9503
rect 18279 9469 18288 9503
rect 18236 9460 18288 9469
rect 18880 9503 18932 9512
rect 18880 9469 18889 9503
rect 18889 9469 18923 9503
rect 18923 9469 18932 9503
rect 18880 9460 18932 9469
rect 19432 9503 19484 9512
rect 19432 9469 19441 9503
rect 19441 9469 19475 9503
rect 19475 9469 19484 9503
rect 19432 9460 19484 9469
rect 22744 9571 22796 9580
rect 22744 9537 22753 9571
rect 22753 9537 22787 9571
rect 22787 9537 22796 9571
rect 22744 9528 22796 9537
rect 22928 9528 22980 9580
rect 23388 9528 23440 9580
rect 24216 9528 24268 9580
rect 20076 9392 20128 9444
rect 23020 9392 23072 9444
rect 23296 9460 23348 9512
rect 24400 9571 24452 9580
rect 24400 9537 24409 9571
rect 24409 9537 24443 9571
rect 24443 9537 24452 9571
rect 24400 9528 24452 9537
rect 26148 9571 26200 9580
rect 26148 9537 26157 9571
rect 26157 9537 26191 9571
rect 26191 9537 26200 9571
rect 26148 9528 26200 9537
rect 24216 9392 24268 9444
rect 24768 9392 24820 9444
rect 13912 9324 13964 9376
rect 18512 9324 18564 9376
rect 19616 9367 19668 9376
rect 19616 9333 19625 9367
rect 19625 9333 19659 9367
rect 19659 9333 19668 9367
rect 19616 9324 19668 9333
rect 24308 9367 24360 9376
rect 24308 9333 24317 9367
rect 24317 9333 24351 9367
rect 24351 9333 24360 9367
rect 24308 9324 24360 9333
rect 24584 9324 24636 9376
rect 26976 9571 27028 9580
rect 26976 9537 26985 9571
rect 26985 9537 27019 9571
rect 27019 9537 27028 9571
rect 26976 9528 27028 9537
rect 27160 9571 27212 9580
rect 27160 9537 27169 9571
rect 27169 9537 27203 9571
rect 27203 9537 27212 9571
rect 27160 9528 27212 9537
rect 27344 9528 27396 9580
rect 27436 9571 27488 9580
rect 27436 9537 27445 9571
rect 27445 9537 27479 9571
rect 27479 9537 27488 9571
rect 27436 9528 27488 9537
rect 27528 9528 27580 9580
rect 27712 9528 27764 9580
rect 29460 9634 29512 9686
rect 30380 9664 30432 9716
rect 33140 9664 33192 9716
rect 33968 9664 34020 9716
rect 29460 9528 29512 9580
rect 29552 9528 29604 9580
rect 30012 9596 30064 9648
rect 27436 9392 27488 9444
rect 28724 9460 28776 9512
rect 30104 9392 30156 9444
rect 30748 9571 30800 9580
rect 30748 9537 30757 9571
rect 30757 9537 30791 9571
rect 30791 9537 30800 9571
rect 30748 9528 30800 9537
rect 30840 9528 30892 9580
rect 31392 9528 31444 9580
rect 30932 9392 30984 9444
rect 26516 9367 26568 9376
rect 26516 9333 26525 9367
rect 26525 9333 26559 9367
rect 26559 9333 26568 9367
rect 26516 9324 26568 9333
rect 27528 9324 27580 9376
rect 28080 9324 28132 9376
rect 29736 9324 29788 9376
rect 33048 9639 33100 9648
rect 33048 9605 33057 9639
rect 33057 9605 33091 9639
rect 33091 9605 33100 9639
rect 33048 9596 33100 9605
rect 32772 9528 32824 9580
rect 32036 9392 32088 9444
rect 31576 9324 31628 9376
rect 31668 9324 31720 9376
rect 33232 9324 33284 9376
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 2964 9120 3016 9172
rect 6736 9120 6788 9172
rect 6920 9120 6972 9172
rect 3332 9052 3384 9104
rect 11612 9120 11664 9172
rect 13084 9120 13136 9172
rect 13820 9120 13872 9172
rect 13912 9120 13964 9172
rect 3056 8916 3108 8968
rect 4160 8959 4212 8968
rect 4160 8925 4169 8959
rect 4169 8925 4203 8959
rect 4203 8925 4212 8959
rect 4160 8916 4212 8925
rect 5632 8984 5684 9036
rect 4528 8959 4580 8968
rect 4528 8925 4537 8959
rect 4537 8925 4571 8959
rect 4571 8925 4580 8959
rect 4528 8916 4580 8925
rect 940 8848 992 8900
rect 7196 8916 7248 8968
rect 4712 8848 4764 8900
rect 6000 8891 6052 8900
rect 6000 8857 6009 8891
rect 6009 8857 6043 8891
rect 6043 8857 6052 8891
rect 6000 8848 6052 8857
rect 6828 8848 6880 8900
rect 3884 8823 3936 8832
rect 3884 8789 3893 8823
rect 3893 8789 3927 8823
rect 3927 8789 3936 8823
rect 3884 8780 3936 8789
rect 8024 8823 8076 8832
rect 8024 8789 8033 8823
rect 8033 8789 8067 8823
rect 8067 8789 8076 8823
rect 8024 8780 8076 8789
rect 8484 8823 8536 8832
rect 8484 8789 8493 8823
rect 8493 8789 8527 8823
rect 8527 8789 8536 8823
rect 8484 8780 8536 8789
rect 8668 8780 8720 8832
rect 9772 9027 9824 9036
rect 9772 8993 9781 9027
rect 9781 8993 9815 9027
rect 9815 8993 9824 9027
rect 9772 8984 9824 8993
rect 10048 9027 10100 9036
rect 10048 8993 10057 9027
rect 10057 8993 10091 9027
rect 10091 8993 10100 9027
rect 10048 8984 10100 8993
rect 10508 8984 10560 9036
rect 11704 8916 11756 8968
rect 12716 8959 12768 8968
rect 12716 8925 12725 8959
rect 12725 8925 12759 8959
rect 12759 8925 12768 8959
rect 12716 8916 12768 8925
rect 13360 8959 13412 8968
rect 13360 8925 13369 8959
rect 13369 8925 13403 8959
rect 13403 8925 13412 8959
rect 13360 8916 13412 8925
rect 13544 8984 13596 9036
rect 13728 8984 13780 9036
rect 14464 9052 14516 9104
rect 18236 9120 18288 9172
rect 13912 8916 13964 8968
rect 15384 9027 15436 9036
rect 15384 8993 15393 9027
rect 15393 8993 15427 9027
rect 15427 8993 15436 9027
rect 15384 8984 15436 8993
rect 17592 8984 17644 9036
rect 20812 9120 20864 9172
rect 21088 9120 21140 9172
rect 22100 9120 22152 9172
rect 18512 9052 18564 9104
rect 22284 9052 22336 9104
rect 22744 9052 22796 9104
rect 11060 8780 11112 8832
rect 12992 8823 13044 8832
rect 12992 8789 13001 8823
rect 13001 8789 13035 8823
rect 13035 8789 13044 8823
rect 12992 8780 13044 8789
rect 13452 8823 13504 8832
rect 13452 8789 13461 8823
rect 13461 8789 13495 8823
rect 13495 8789 13504 8823
rect 13452 8780 13504 8789
rect 13912 8780 13964 8832
rect 15016 8916 15068 8968
rect 15292 8959 15344 8968
rect 15292 8925 15301 8959
rect 15301 8925 15335 8959
rect 15335 8925 15344 8959
rect 15292 8916 15344 8925
rect 14740 8823 14792 8832
rect 14740 8789 14749 8823
rect 14749 8789 14783 8823
rect 14783 8789 14792 8823
rect 14740 8780 14792 8789
rect 14924 8823 14976 8832
rect 14924 8789 14933 8823
rect 14933 8789 14967 8823
rect 14967 8789 14976 8823
rect 14924 8780 14976 8789
rect 22192 9027 22244 9036
rect 22192 8993 22201 9027
rect 22201 8993 22235 9027
rect 22235 8993 22244 9027
rect 22192 8984 22244 8993
rect 15752 8959 15804 8968
rect 15752 8925 15761 8959
rect 15761 8925 15795 8959
rect 15795 8925 15804 8959
rect 15752 8916 15804 8925
rect 16028 8891 16080 8900
rect 16028 8857 16037 8891
rect 16037 8857 16071 8891
rect 16071 8857 16080 8891
rect 16028 8848 16080 8857
rect 16764 8848 16816 8900
rect 18144 8916 18196 8968
rect 19524 8916 19576 8968
rect 19708 8780 19760 8832
rect 19984 8959 20036 8968
rect 19984 8925 19993 8959
rect 19993 8925 20027 8959
rect 20027 8925 20036 8959
rect 19984 8916 20036 8925
rect 20076 8916 20128 8968
rect 22376 8916 22428 8968
rect 22560 8959 22612 8968
rect 22560 8925 22569 8959
rect 22569 8925 22603 8959
rect 22603 8925 22612 8959
rect 22560 8916 22612 8925
rect 19892 8891 19944 8900
rect 19892 8857 19901 8891
rect 19901 8857 19935 8891
rect 19935 8857 19944 8891
rect 19892 8848 19944 8857
rect 20260 8891 20312 8900
rect 20260 8857 20269 8891
rect 20269 8857 20303 8891
rect 20303 8857 20312 8891
rect 20260 8848 20312 8857
rect 22284 8891 22336 8900
rect 22284 8857 22293 8891
rect 22293 8857 22327 8891
rect 22327 8857 22336 8891
rect 22284 8848 22336 8857
rect 22928 9052 22980 9104
rect 23112 9052 23164 9104
rect 23572 9052 23624 9104
rect 23020 8959 23072 8968
rect 23020 8925 23030 8959
rect 23030 8925 23064 8959
rect 23064 8925 23072 8959
rect 23020 8916 23072 8925
rect 23388 8959 23440 8968
rect 23388 8925 23402 8959
rect 23402 8925 23436 8959
rect 23436 8925 23440 8959
rect 23388 8916 23440 8925
rect 23296 8891 23348 8900
rect 23296 8857 23305 8891
rect 23305 8857 23339 8891
rect 23339 8857 23348 8891
rect 23296 8848 23348 8857
rect 23572 8823 23624 8832
rect 23572 8789 23581 8823
rect 23581 8789 23615 8823
rect 23615 8789 23624 8823
rect 23572 8780 23624 8789
rect 24216 8984 24268 9036
rect 24676 9052 24728 9104
rect 26332 9120 26384 9172
rect 25320 9027 25372 9036
rect 25320 8993 25329 9027
rect 25329 8993 25363 9027
rect 25363 8993 25372 9027
rect 25320 8984 25372 8993
rect 24860 8959 24912 8968
rect 24860 8925 24893 8959
rect 24893 8925 24912 8959
rect 24860 8916 24912 8925
rect 25044 8916 25096 8968
rect 24584 8848 24636 8900
rect 25964 8916 26016 8968
rect 26976 9052 27028 9104
rect 27068 9052 27120 9104
rect 26516 8916 26568 8968
rect 26884 8984 26936 9036
rect 28080 8984 28132 9036
rect 25136 8780 25188 8832
rect 25412 8848 25464 8900
rect 26332 8780 26384 8832
rect 26516 8823 26568 8832
rect 26516 8789 26525 8823
rect 26525 8789 26559 8823
rect 26559 8789 26568 8823
rect 26516 8780 26568 8789
rect 26884 8848 26936 8900
rect 27252 8916 27304 8968
rect 27620 8959 27672 8968
rect 27620 8925 27629 8959
rect 27629 8925 27663 8959
rect 27663 8925 27672 8959
rect 27620 8916 27672 8925
rect 27712 8848 27764 8900
rect 28448 8959 28500 8968
rect 28448 8925 28457 8959
rect 28457 8925 28491 8959
rect 28491 8925 28500 8959
rect 28448 8916 28500 8925
rect 29184 9052 29236 9104
rect 29276 8984 29328 9036
rect 29644 9120 29696 9172
rect 29736 9163 29788 9172
rect 29736 9129 29745 9163
rect 29745 9129 29779 9163
rect 29779 9129 29788 9163
rect 29736 9120 29788 9129
rect 27160 8780 27212 8832
rect 29276 8848 29328 8900
rect 28816 8823 28868 8832
rect 28816 8789 28825 8823
rect 28825 8789 28859 8823
rect 28859 8789 28868 8823
rect 28816 8780 28868 8789
rect 28908 8780 28960 8832
rect 29000 8823 29052 8832
rect 29000 8789 29009 8823
rect 29009 8789 29043 8823
rect 29043 8789 29052 8823
rect 29000 8780 29052 8789
rect 29092 8780 29144 8832
rect 30196 8959 30248 8968
rect 30196 8925 30205 8959
rect 30205 8925 30239 8959
rect 30239 8925 30248 8959
rect 30196 8916 30248 8925
rect 30380 8891 30432 8900
rect 30380 8857 30389 8891
rect 30389 8857 30423 8891
rect 30423 8857 30432 8891
rect 30380 8848 30432 8857
rect 30748 9120 30800 9172
rect 31576 9120 31628 9172
rect 33140 9120 33192 9172
rect 33324 9120 33376 9172
rect 32036 8984 32088 9036
rect 31760 8916 31812 8968
rect 31852 8959 31904 8968
rect 31852 8925 31861 8959
rect 31861 8925 31895 8959
rect 31895 8925 31904 8959
rect 31852 8916 31904 8925
rect 30840 8780 30892 8832
rect 31944 8823 31996 8832
rect 31944 8789 31953 8823
rect 31953 8789 31987 8823
rect 31987 8789 31996 8823
rect 31944 8780 31996 8789
rect 32772 8916 32824 8968
rect 32864 8848 32916 8900
rect 33048 8959 33100 8968
rect 33048 8925 33057 8959
rect 33057 8925 33091 8959
rect 33091 8925 33100 8959
rect 33048 8916 33100 8925
rect 33140 8916 33192 8968
rect 33508 8959 33560 8968
rect 33508 8925 33517 8959
rect 33517 8925 33551 8959
rect 33551 8925 33560 8959
rect 33508 8916 33560 8925
rect 38292 8916 38344 8968
rect 35992 8848 36044 8900
rect 36820 8848 36872 8900
rect 33232 8780 33284 8832
rect 4874 8678 4926 8730
rect 4938 8678 4990 8730
rect 5002 8678 5054 8730
rect 5066 8678 5118 8730
rect 5130 8678 5182 8730
rect 35594 8678 35646 8730
rect 35658 8678 35710 8730
rect 35722 8678 35774 8730
rect 35786 8678 35838 8730
rect 35850 8678 35902 8730
rect 6000 8508 6052 8560
rect 7104 8576 7156 8628
rect 9220 8576 9272 8628
rect 9404 8576 9456 8628
rect 9864 8576 9916 8628
rect 10140 8576 10192 8628
rect 4712 8440 4764 8492
rect 4068 8304 4120 8356
rect 5540 8415 5592 8424
rect 5540 8381 5549 8415
rect 5549 8381 5583 8415
rect 5583 8381 5592 8415
rect 5540 8372 5592 8381
rect 5632 8372 5684 8424
rect 5724 8415 5776 8424
rect 5724 8381 5733 8415
rect 5733 8381 5767 8415
rect 5767 8381 5776 8415
rect 5724 8372 5776 8381
rect 6276 8440 6328 8492
rect 9588 8508 9640 8560
rect 12716 8576 12768 8628
rect 12992 8576 13044 8628
rect 8668 8440 8720 8492
rect 11152 8440 11204 8492
rect 11796 8440 11848 8492
rect 12624 8551 12676 8560
rect 12624 8517 12633 8551
rect 12633 8517 12667 8551
rect 12667 8517 12676 8551
rect 12624 8508 12676 8517
rect 13452 8576 13504 8628
rect 18420 8576 18472 8628
rect 22376 8576 22428 8628
rect 23572 8576 23624 8628
rect 24308 8576 24360 8628
rect 12348 8483 12400 8492
rect 12348 8449 12357 8483
rect 12357 8449 12391 8483
rect 12391 8449 12400 8483
rect 12348 8440 12400 8449
rect 12532 8483 12584 8492
rect 12532 8449 12541 8483
rect 12541 8449 12575 8483
rect 12575 8449 12584 8483
rect 12532 8440 12584 8449
rect 12992 8483 13044 8492
rect 12992 8449 13001 8483
rect 13001 8449 13035 8483
rect 13035 8449 13044 8483
rect 12992 8440 13044 8449
rect 15016 8508 15068 8560
rect 16764 8440 16816 8492
rect 17132 8440 17184 8492
rect 17408 8483 17460 8492
rect 17408 8449 17417 8483
rect 17417 8449 17451 8483
rect 17451 8449 17460 8483
rect 17408 8440 17460 8449
rect 5908 8347 5960 8356
rect 5908 8313 5917 8347
rect 5917 8313 5951 8347
rect 5951 8313 5960 8347
rect 5908 8304 5960 8313
rect 6460 8304 6512 8356
rect 8484 8304 8536 8356
rect 10416 8372 10468 8424
rect 10600 8372 10652 8424
rect 12256 8372 12308 8424
rect 14924 8372 14976 8424
rect 19524 8551 19576 8560
rect 19524 8517 19533 8551
rect 19533 8517 19567 8551
rect 19567 8517 19576 8551
rect 19524 8508 19576 8517
rect 19892 8508 19944 8560
rect 19984 8508 20036 8560
rect 21456 8508 21508 8560
rect 18972 8483 19024 8492
rect 18972 8449 18981 8483
rect 18981 8449 19015 8483
rect 19015 8449 19024 8483
rect 18972 8440 19024 8449
rect 19156 8440 19208 8492
rect 20812 8440 20864 8492
rect 21824 8440 21876 8492
rect 22008 8440 22060 8492
rect 25320 8508 25372 8560
rect 28908 8576 28960 8628
rect 26884 8508 26936 8560
rect 23572 8440 23624 8492
rect 24216 8440 24268 8492
rect 21548 8372 21600 8424
rect 25412 8440 25464 8492
rect 26516 8440 26568 8492
rect 29000 8508 29052 8560
rect 30196 8576 30248 8628
rect 31392 8576 31444 8628
rect 32036 8576 32088 8628
rect 32772 8576 32824 8628
rect 33508 8576 33560 8628
rect 27344 8483 27396 8492
rect 27344 8449 27353 8483
rect 27353 8449 27387 8483
rect 27387 8449 27396 8483
rect 27344 8440 27396 8449
rect 27436 8440 27488 8492
rect 27620 8440 27672 8492
rect 30012 8508 30064 8560
rect 31944 8508 31996 8560
rect 31668 8440 31720 8492
rect 16948 8304 17000 8356
rect 2964 8236 3016 8288
rect 4620 8236 4672 8288
rect 6276 8236 6328 8288
rect 6828 8236 6880 8288
rect 8668 8236 8720 8288
rect 17224 8347 17276 8356
rect 17224 8313 17233 8347
rect 17233 8313 17267 8347
rect 17267 8313 17276 8347
rect 17224 8304 17276 8313
rect 27804 8304 27856 8356
rect 29276 8372 29328 8424
rect 31024 8372 31076 8424
rect 35992 8508 36044 8560
rect 33048 8440 33100 8492
rect 33232 8415 33284 8424
rect 33232 8381 33241 8415
rect 33241 8381 33275 8415
rect 33275 8381 33284 8415
rect 33232 8372 33284 8381
rect 32588 8304 32640 8356
rect 19524 8279 19576 8288
rect 19524 8245 19533 8279
rect 19533 8245 19567 8279
rect 19567 8245 19576 8279
rect 19524 8236 19576 8245
rect 20904 8236 20956 8288
rect 21916 8236 21968 8288
rect 22376 8236 22428 8288
rect 23020 8279 23072 8288
rect 23020 8245 23029 8279
rect 23029 8245 23063 8279
rect 23063 8245 23072 8279
rect 23020 8236 23072 8245
rect 25320 8279 25372 8288
rect 25320 8245 25329 8279
rect 25329 8245 25363 8279
rect 25363 8245 25372 8279
rect 25320 8236 25372 8245
rect 29000 8279 29052 8288
rect 29000 8245 29009 8279
rect 29009 8245 29043 8279
rect 29043 8245 29052 8279
rect 29000 8236 29052 8245
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 5540 8032 5592 8084
rect 5816 8032 5868 8084
rect 6368 8032 6420 8084
rect 5724 7828 5776 7880
rect 5908 7828 5960 7880
rect 8668 8075 8720 8084
rect 8668 8041 8677 8075
rect 8677 8041 8711 8075
rect 8711 8041 8720 8075
rect 8668 8032 8720 8041
rect 8852 8032 8904 8084
rect 9864 8032 9916 8084
rect 12532 8032 12584 8084
rect 12992 8032 13044 8084
rect 13728 8075 13780 8084
rect 13728 8041 13737 8075
rect 13737 8041 13771 8075
rect 13771 8041 13780 8075
rect 13728 8032 13780 8041
rect 23572 8032 23624 8084
rect 26240 8032 26292 8084
rect 29368 8032 29420 8084
rect 29460 8032 29512 8084
rect 22652 7964 22704 8016
rect 22744 7964 22796 8016
rect 6920 7939 6972 7948
rect 6920 7905 6929 7939
rect 6929 7905 6963 7939
rect 6963 7905 6972 7939
rect 6920 7896 6972 7905
rect 9404 7896 9456 7948
rect 8300 7828 8352 7880
rect 8852 7828 8904 7880
rect 9220 7828 9272 7880
rect 10600 7896 10652 7948
rect 12256 7896 12308 7948
rect 10876 7828 10928 7880
rect 13544 7896 13596 7948
rect 14004 7896 14056 7948
rect 15936 7939 15988 7948
rect 15936 7905 15945 7939
rect 15945 7905 15979 7939
rect 15979 7905 15988 7939
rect 15936 7896 15988 7905
rect 12900 7828 12952 7880
rect 19524 7896 19576 7948
rect 17592 7871 17644 7880
rect 7196 7803 7248 7812
rect 7196 7769 7205 7803
rect 7205 7769 7239 7803
rect 7239 7769 7248 7803
rect 7196 7760 7248 7769
rect 12348 7803 12400 7812
rect 12348 7769 12357 7803
rect 12357 7769 12391 7803
rect 12391 7769 12400 7803
rect 12348 7760 12400 7769
rect 12532 7760 12584 7812
rect 13544 7760 13596 7812
rect 17592 7837 17601 7871
rect 17601 7837 17635 7871
rect 17635 7837 17644 7871
rect 17592 7828 17644 7837
rect 17776 7871 17828 7880
rect 17776 7837 17785 7871
rect 17785 7837 17819 7871
rect 17819 7837 17828 7871
rect 17776 7828 17828 7837
rect 19708 7871 19760 7880
rect 19708 7837 19717 7871
rect 19717 7837 19751 7871
rect 19751 7837 19760 7871
rect 19708 7828 19760 7837
rect 20628 7896 20680 7948
rect 16856 7760 16908 7812
rect 21456 7828 21508 7880
rect 22284 7896 22336 7948
rect 22376 7939 22428 7948
rect 22376 7905 22385 7939
rect 22385 7905 22419 7939
rect 22419 7905 22428 7939
rect 22376 7896 22428 7905
rect 21824 7871 21876 7880
rect 21824 7837 21833 7871
rect 21833 7837 21867 7871
rect 21867 7837 21876 7871
rect 21824 7828 21876 7837
rect 23020 7896 23072 7948
rect 28540 7896 28592 7948
rect 28724 7896 28776 7948
rect 6092 7735 6144 7744
rect 6092 7701 6101 7735
rect 6101 7701 6135 7735
rect 6135 7701 6144 7735
rect 6092 7692 6144 7701
rect 6552 7735 6604 7744
rect 6552 7701 6561 7735
rect 6561 7701 6595 7735
rect 6595 7701 6604 7735
rect 6552 7692 6604 7701
rect 9680 7692 9732 7744
rect 9772 7735 9824 7744
rect 9772 7701 9781 7735
rect 9781 7701 9815 7735
rect 9815 7701 9824 7735
rect 9772 7692 9824 7701
rect 15384 7735 15436 7744
rect 15384 7701 15393 7735
rect 15393 7701 15427 7735
rect 15427 7701 15436 7735
rect 15384 7692 15436 7701
rect 17316 7735 17368 7744
rect 17316 7701 17325 7735
rect 17325 7701 17359 7735
rect 17359 7701 17368 7735
rect 17316 7692 17368 7701
rect 20536 7692 20588 7744
rect 22652 7871 22704 7880
rect 22652 7837 22661 7871
rect 22661 7837 22695 7871
rect 22695 7837 22704 7871
rect 22652 7828 22704 7837
rect 30012 7871 30064 7880
rect 30012 7837 30021 7871
rect 30021 7837 30055 7871
rect 30055 7837 30064 7871
rect 30012 7828 30064 7837
rect 30472 7896 30524 7948
rect 31484 8032 31536 8084
rect 31760 8032 31812 8084
rect 33048 7964 33100 8016
rect 30380 7871 30432 7880
rect 30380 7837 30389 7871
rect 30389 7837 30423 7871
rect 30423 7837 30432 7871
rect 30380 7828 30432 7837
rect 30564 7871 30616 7880
rect 30564 7837 30573 7871
rect 30573 7837 30607 7871
rect 30607 7837 30616 7871
rect 30564 7828 30616 7837
rect 30840 7828 30892 7880
rect 31024 7828 31076 7880
rect 22376 7760 22428 7812
rect 22744 7803 22796 7812
rect 22744 7769 22753 7803
rect 22753 7769 22787 7803
rect 22787 7769 22796 7803
rect 22744 7760 22796 7769
rect 23112 7803 23164 7812
rect 23112 7769 23121 7803
rect 23121 7769 23155 7803
rect 23155 7769 23164 7803
rect 23112 7760 23164 7769
rect 30748 7760 30800 7812
rect 22100 7692 22152 7744
rect 22284 7735 22336 7744
rect 22284 7701 22293 7735
rect 22293 7701 22327 7735
rect 22327 7701 22336 7735
rect 22284 7692 22336 7701
rect 22468 7692 22520 7744
rect 23204 7692 23256 7744
rect 24032 7692 24084 7744
rect 24308 7692 24360 7744
rect 31116 7692 31168 7744
rect 31208 7735 31260 7744
rect 31208 7701 31217 7735
rect 31217 7701 31251 7735
rect 31251 7701 31260 7735
rect 31208 7692 31260 7701
rect 31668 7803 31720 7812
rect 31668 7769 31677 7803
rect 31677 7769 31711 7803
rect 31711 7769 31720 7803
rect 31668 7760 31720 7769
rect 4874 7590 4926 7642
rect 4938 7590 4990 7642
rect 5002 7590 5054 7642
rect 5066 7590 5118 7642
rect 5130 7590 5182 7642
rect 35594 7590 35646 7642
rect 35658 7590 35710 7642
rect 35722 7590 35774 7642
rect 35786 7590 35838 7642
rect 35850 7590 35902 7642
rect 1492 7395 1544 7404
rect 1492 7361 1501 7395
rect 1501 7361 1535 7395
rect 1535 7361 1544 7395
rect 1492 7352 1544 7361
rect 4620 7488 4672 7540
rect 6092 7488 6144 7540
rect 6552 7488 6604 7540
rect 7196 7488 7248 7540
rect 8024 7488 8076 7540
rect 2964 7420 3016 7472
rect 3976 7352 4028 7404
rect 5448 7352 5500 7404
rect 6000 7352 6052 7404
rect 4712 7284 4764 7336
rect 5632 7284 5684 7336
rect 9772 7488 9824 7540
rect 9864 7488 9916 7540
rect 13636 7488 13688 7540
rect 15384 7488 15436 7540
rect 19156 7488 19208 7540
rect 21088 7488 21140 7540
rect 22284 7488 22336 7540
rect 22376 7531 22428 7540
rect 22376 7497 22385 7531
rect 22385 7497 22419 7531
rect 22419 7497 22428 7531
rect 22376 7488 22428 7497
rect 11796 7463 11848 7472
rect 11796 7429 11805 7463
rect 11805 7429 11839 7463
rect 11839 7429 11848 7463
rect 11796 7420 11848 7429
rect 12072 7420 12124 7472
rect 9404 7395 9456 7404
rect 9404 7361 9413 7395
rect 9413 7361 9447 7395
rect 9447 7361 9456 7395
rect 9404 7352 9456 7361
rect 12808 7352 12860 7404
rect 14188 7352 14240 7404
rect 6828 7327 6880 7336
rect 6828 7293 6837 7327
rect 6837 7293 6871 7327
rect 6871 7293 6880 7327
rect 6828 7284 6880 7293
rect 11888 7284 11940 7336
rect 12256 7284 12308 7336
rect 14464 7352 14516 7404
rect 15292 7420 15344 7472
rect 17776 7395 17828 7404
rect 17776 7361 17785 7395
rect 17785 7361 17819 7395
rect 17819 7361 17828 7395
rect 17776 7352 17828 7361
rect 18512 7420 18564 7472
rect 15292 7284 15344 7336
rect 14924 7216 14976 7268
rect 15476 7216 15528 7268
rect 18696 7284 18748 7336
rect 19708 7352 19760 7404
rect 20628 7352 20680 7404
rect 4804 7148 4856 7200
rect 11152 7191 11204 7200
rect 11152 7157 11161 7191
rect 11161 7157 11195 7191
rect 11195 7157 11204 7191
rect 11152 7148 11204 7157
rect 12900 7148 12952 7200
rect 15568 7148 15620 7200
rect 17868 7191 17920 7200
rect 17868 7157 17877 7191
rect 17877 7157 17911 7191
rect 17911 7157 17920 7191
rect 17868 7148 17920 7157
rect 18052 7148 18104 7200
rect 20536 7148 20588 7200
rect 22100 7395 22152 7404
rect 22100 7361 22109 7395
rect 22109 7361 22143 7395
rect 22143 7361 22152 7395
rect 22100 7352 22152 7361
rect 22192 7395 22244 7404
rect 22192 7361 22201 7395
rect 22201 7361 22235 7395
rect 22235 7361 22244 7395
rect 22192 7352 22244 7361
rect 22928 7463 22980 7472
rect 22928 7429 22937 7463
rect 22937 7429 22971 7463
rect 22971 7429 22980 7463
rect 22928 7420 22980 7429
rect 23112 7488 23164 7540
rect 26424 7488 26476 7540
rect 26608 7531 26660 7540
rect 26608 7497 26617 7531
rect 26617 7497 26651 7531
rect 26651 7497 26660 7531
rect 26608 7488 26660 7497
rect 27436 7488 27488 7540
rect 27620 7488 27672 7540
rect 27712 7488 27764 7540
rect 21272 7284 21324 7336
rect 23572 7352 23624 7404
rect 24032 7395 24084 7404
rect 24032 7361 24041 7395
rect 24041 7361 24075 7395
rect 24075 7361 24084 7395
rect 24032 7352 24084 7361
rect 24492 7395 24544 7404
rect 24492 7361 24501 7395
rect 24501 7361 24535 7395
rect 24535 7361 24544 7395
rect 24492 7352 24544 7361
rect 24584 7352 24636 7404
rect 22008 7216 22060 7268
rect 23296 7216 23348 7268
rect 25320 7420 25372 7472
rect 26240 7420 26292 7472
rect 26332 7420 26384 7472
rect 30012 7488 30064 7540
rect 31208 7488 31260 7540
rect 25228 7352 25280 7404
rect 25412 7284 25464 7336
rect 25964 7284 26016 7336
rect 21364 7148 21416 7200
rect 21916 7191 21968 7200
rect 21916 7157 21925 7191
rect 21925 7157 21959 7191
rect 21959 7157 21968 7191
rect 21916 7148 21968 7157
rect 24768 7148 24820 7200
rect 24860 7191 24912 7200
rect 24860 7157 24869 7191
rect 24869 7157 24903 7191
rect 24903 7157 24912 7191
rect 24860 7148 24912 7157
rect 25044 7148 25096 7200
rect 25136 7191 25188 7200
rect 25136 7157 25145 7191
rect 25145 7157 25179 7191
rect 25179 7157 25188 7191
rect 25136 7148 25188 7157
rect 28540 7352 28592 7404
rect 28632 7327 28684 7336
rect 28632 7293 28641 7327
rect 28641 7293 28675 7327
rect 28675 7293 28684 7327
rect 28632 7284 28684 7293
rect 28080 7216 28132 7268
rect 29184 7352 29236 7404
rect 29460 7352 29512 7404
rect 31576 7420 31628 7472
rect 30656 7352 30708 7404
rect 31392 7395 31444 7404
rect 31392 7361 31401 7395
rect 31401 7361 31435 7395
rect 31435 7361 31444 7395
rect 31392 7352 31444 7361
rect 31760 7395 31812 7404
rect 31760 7361 31769 7395
rect 31769 7361 31803 7395
rect 31803 7361 31812 7395
rect 31760 7352 31812 7361
rect 30380 7284 30432 7336
rect 31300 7327 31352 7336
rect 31300 7293 31309 7327
rect 31309 7293 31343 7327
rect 31343 7293 31352 7327
rect 31300 7284 31352 7293
rect 34060 7216 34112 7268
rect 30564 7148 30616 7200
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 3976 6944 4028 6996
rect 4620 6808 4672 6860
rect 6000 6987 6052 6996
rect 6000 6953 6009 6987
rect 6009 6953 6043 6987
rect 6043 6953 6052 6987
rect 6000 6944 6052 6953
rect 12348 6987 12400 6996
rect 12348 6953 12357 6987
rect 12357 6953 12391 6987
rect 12391 6953 12400 6987
rect 12348 6944 12400 6953
rect 13544 6944 13596 6996
rect 15568 6944 15620 6996
rect 17776 6944 17828 6996
rect 18052 6987 18104 6996
rect 18052 6953 18061 6987
rect 18061 6953 18095 6987
rect 18095 6953 18104 6987
rect 18052 6944 18104 6953
rect 21272 6944 21324 6996
rect 23204 6944 23256 6996
rect 23848 6944 23900 6996
rect 25412 6987 25464 6996
rect 25412 6953 25421 6987
rect 25421 6953 25455 6987
rect 25455 6953 25464 6987
rect 25412 6944 25464 6953
rect 11152 6876 11204 6928
rect 17316 6876 17368 6928
rect 4528 6715 4580 6724
rect 4528 6681 4537 6715
rect 4537 6681 4571 6715
rect 4571 6681 4580 6715
rect 4528 6672 4580 6681
rect 13728 6808 13780 6860
rect 15752 6808 15804 6860
rect 17868 6851 17920 6860
rect 17868 6817 17877 6851
rect 17877 6817 17911 6851
rect 17911 6817 17920 6851
rect 17868 6808 17920 6817
rect 8208 6740 8260 6792
rect 9496 6740 9548 6792
rect 10692 6740 10744 6792
rect 12808 6740 12860 6792
rect 12900 6783 12952 6792
rect 12900 6749 12909 6783
rect 12909 6749 12943 6783
rect 12943 6749 12952 6783
rect 12900 6740 12952 6749
rect 15200 6783 15252 6792
rect 15200 6749 15209 6783
rect 15209 6749 15243 6783
rect 15243 6749 15252 6783
rect 15200 6740 15252 6749
rect 6460 6672 6512 6724
rect 16764 6672 16816 6724
rect 18236 6740 18288 6792
rect 19984 6851 20036 6860
rect 19984 6817 19993 6851
rect 19993 6817 20027 6851
rect 20027 6817 20036 6851
rect 19984 6808 20036 6817
rect 30380 6944 30432 6996
rect 30840 6944 30892 6996
rect 31300 6944 31352 6996
rect 31392 6944 31444 6996
rect 31944 6944 31996 6996
rect 18512 6783 18564 6792
rect 18512 6749 18521 6783
rect 18521 6749 18555 6783
rect 18555 6749 18564 6783
rect 18512 6740 18564 6749
rect 18972 6740 19024 6792
rect 20628 6740 20680 6792
rect 21272 6783 21324 6792
rect 21272 6749 21281 6783
rect 21281 6749 21315 6783
rect 21315 6749 21324 6783
rect 21272 6740 21324 6749
rect 21364 6740 21416 6792
rect 22100 6672 22152 6724
rect 24860 6851 24912 6860
rect 24860 6817 24869 6851
rect 24869 6817 24903 6851
rect 24903 6817 24912 6851
rect 24860 6808 24912 6817
rect 24952 6783 25004 6792
rect 24952 6749 24961 6783
rect 24961 6749 24995 6783
rect 24995 6749 25004 6783
rect 24952 6740 25004 6749
rect 26056 6740 26108 6792
rect 26608 6808 26660 6860
rect 26240 6783 26292 6792
rect 26240 6749 26249 6783
rect 26249 6749 26283 6783
rect 26283 6749 26292 6783
rect 26240 6740 26292 6749
rect 27804 6808 27856 6860
rect 25504 6672 25556 6724
rect 8300 6604 8352 6656
rect 9036 6647 9088 6656
rect 9036 6613 9045 6647
rect 9045 6613 9079 6647
rect 9079 6613 9088 6647
rect 9036 6604 9088 6613
rect 14556 6647 14608 6656
rect 14556 6613 14565 6647
rect 14565 6613 14599 6647
rect 14599 6613 14608 6647
rect 14556 6604 14608 6613
rect 22376 6604 22428 6656
rect 23572 6604 23624 6656
rect 23848 6604 23900 6656
rect 25320 6647 25372 6656
rect 25320 6613 25329 6647
rect 25329 6613 25363 6647
rect 25363 6613 25372 6647
rect 25320 6604 25372 6613
rect 26976 6783 27028 6792
rect 26976 6749 26985 6783
rect 26985 6749 27019 6783
rect 27019 6749 27028 6783
rect 26976 6740 27028 6749
rect 27436 6740 27488 6792
rect 28448 6808 28500 6860
rect 28540 6851 28592 6860
rect 28540 6817 28549 6851
rect 28549 6817 28583 6851
rect 28583 6817 28592 6851
rect 28540 6808 28592 6817
rect 28632 6808 28684 6860
rect 30564 6808 30616 6860
rect 26700 6604 26752 6656
rect 27988 6783 28040 6792
rect 27988 6749 28002 6783
rect 28002 6749 28036 6783
rect 28036 6749 28040 6783
rect 27988 6740 28040 6749
rect 28172 6740 28224 6792
rect 28264 6783 28316 6792
rect 28264 6749 28273 6783
rect 28273 6749 28307 6783
rect 28307 6749 28316 6783
rect 28264 6740 28316 6749
rect 28080 6672 28132 6724
rect 28816 6740 28868 6792
rect 30012 6740 30064 6792
rect 30472 6740 30524 6792
rect 30748 6783 30800 6792
rect 30748 6749 30757 6783
rect 30757 6749 30791 6783
rect 30791 6749 30800 6783
rect 30748 6740 30800 6749
rect 32496 6876 32548 6928
rect 31760 6783 31812 6792
rect 31760 6749 31769 6783
rect 31769 6749 31803 6783
rect 31803 6749 31812 6783
rect 31760 6740 31812 6749
rect 31852 6783 31904 6792
rect 31852 6749 31861 6783
rect 31861 6749 31895 6783
rect 31895 6749 31904 6783
rect 31852 6740 31904 6749
rect 32864 6808 32916 6860
rect 32128 6783 32180 6792
rect 32128 6749 32137 6783
rect 32137 6749 32171 6783
rect 32171 6749 32180 6783
rect 32128 6740 32180 6749
rect 32220 6740 32272 6792
rect 28448 6672 28500 6724
rect 32588 6783 32640 6792
rect 32588 6749 32597 6783
rect 32597 6749 32631 6783
rect 32631 6749 32640 6783
rect 32588 6740 32640 6749
rect 33048 6740 33100 6792
rect 34428 6672 34480 6724
rect 28356 6604 28408 6656
rect 32680 6604 32732 6656
rect 4874 6502 4926 6554
rect 4938 6502 4990 6554
rect 5002 6502 5054 6554
rect 5066 6502 5118 6554
rect 5130 6502 5182 6554
rect 35594 6502 35646 6554
rect 35658 6502 35710 6554
rect 35722 6502 35774 6554
rect 35786 6502 35838 6554
rect 35850 6502 35902 6554
rect 4528 6400 4580 6452
rect 4804 6400 4856 6452
rect 9496 6400 9548 6452
rect 8852 6332 8904 6384
rect 9404 6332 9456 6384
rect 11060 6332 11112 6384
rect 8208 6264 8260 6316
rect 7472 6196 7524 6248
rect 9312 6239 9364 6248
rect 9312 6205 9321 6239
rect 9321 6205 9355 6239
rect 9355 6205 9364 6239
rect 9312 6196 9364 6205
rect 10232 6264 10284 6316
rect 9772 6196 9824 6248
rect 13544 6264 13596 6316
rect 14464 6400 14516 6452
rect 15476 6400 15528 6452
rect 17868 6400 17920 6452
rect 18696 6443 18748 6452
rect 18696 6409 18705 6443
rect 18705 6409 18739 6443
rect 18739 6409 18748 6443
rect 18696 6400 18748 6409
rect 19616 6400 19668 6452
rect 19800 6400 19852 6452
rect 19984 6400 20036 6452
rect 15384 6332 15436 6384
rect 15200 6264 15252 6316
rect 15292 6264 15344 6316
rect 18144 6264 18196 6316
rect 18512 6332 18564 6384
rect 12348 6128 12400 6180
rect 18144 6171 18196 6180
rect 18144 6137 18153 6171
rect 18153 6137 18187 6171
rect 18187 6137 18196 6171
rect 18144 6128 18196 6137
rect 7380 6103 7432 6112
rect 7380 6069 7389 6103
rect 7389 6069 7423 6103
rect 7423 6069 7432 6103
rect 7380 6060 7432 6069
rect 8208 6103 8260 6112
rect 8208 6069 8217 6103
rect 8217 6069 8251 6103
rect 8251 6069 8260 6103
rect 8208 6060 8260 6069
rect 8852 6060 8904 6112
rect 9496 6060 9548 6112
rect 12532 6060 12584 6112
rect 16488 6060 16540 6112
rect 18972 6264 19024 6316
rect 22744 6400 22796 6452
rect 22928 6332 22980 6384
rect 23480 6375 23532 6384
rect 23480 6341 23489 6375
rect 23489 6341 23523 6375
rect 23523 6341 23532 6375
rect 23480 6332 23532 6341
rect 24952 6400 25004 6452
rect 25228 6400 25280 6452
rect 27988 6443 28040 6452
rect 27988 6409 27997 6443
rect 27997 6409 28031 6443
rect 28031 6409 28040 6443
rect 27988 6400 28040 6409
rect 28172 6443 28224 6452
rect 28172 6409 28181 6443
rect 28181 6409 28215 6443
rect 28215 6409 28224 6443
rect 28172 6400 28224 6409
rect 31024 6400 31076 6452
rect 25320 6332 25372 6384
rect 32496 6400 32548 6452
rect 32588 6400 32640 6452
rect 22652 6264 22704 6316
rect 23112 6264 23164 6316
rect 23572 6307 23624 6316
rect 23572 6273 23581 6307
rect 23581 6273 23615 6307
rect 23615 6273 23624 6307
rect 23572 6264 23624 6273
rect 24308 6307 24360 6316
rect 24308 6273 24317 6307
rect 24317 6273 24351 6307
rect 24351 6273 24360 6307
rect 24308 6264 24360 6273
rect 24768 6264 24820 6316
rect 26056 6264 26108 6316
rect 27804 6307 27856 6316
rect 19524 6060 19576 6112
rect 23020 6103 23072 6112
rect 23020 6069 23029 6103
rect 23029 6069 23063 6103
rect 23063 6069 23072 6103
rect 23020 6060 23072 6069
rect 23296 6128 23348 6180
rect 27804 6273 27813 6307
rect 27813 6273 27847 6307
rect 27847 6273 27856 6307
rect 27804 6264 27856 6273
rect 27528 6239 27580 6248
rect 27528 6205 27537 6239
rect 27537 6205 27571 6239
rect 27571 6205 27580 6239
rect 27528 6196 27580 6205
rect 27712 6196 27764 6248
rect 32220 6264 32272 6316
rect 32680 6264 32732 6316
rect 32772 6171 32824 6180
rect 32772 6137 32781 6171
rect 32781 6137 32815 6171
rect 32815 6137 32824 6171
rect 32772 6128 32824 6137
rect 27620 6103 27672 6112
rect 27620 6069 27629 6103
rect 27629 6069 27663 6103
rect 27663 6069 27672 6103
rect 27620 6060 27672 6069
rect 32036 6060 32088 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 8208 5856 8260 5908
rect 4620 5720 4672 5772
rect 6920 5763 6972 5772
rect 6920 5729 6929 5763
rect 6929 5729 6963 5763
rect 6963 5729 6972 5763
rect 6920 5720 6972 5729
rect 9312 5856 9364 5908
rect 9680 5788 9732 5840
rect 6460 5652 6512 5704
rect 8300 5652 8352 5704
rect 9404 5695 9456 5704
rect 9404 5661 9413 5695
rect 9413 5661 9447 5695
rect 9447 5661 9456 5695
rect 9404 5652 9456 5661
rect 9496 5695 9548 5704
rect 9496 5661 9506 5695
rect 9506 5661 9540 5695
rect 9540 5661 9548 5695
rect 9496 5652 9548 5661
rect 9772 5695 9824 5704
rect 9772 5661 9781 5695
rect 9781 5661 9815 5695
rect 9815 5661 9824 5695
rect 9772 5652 9824 5661
rect 10784 5856 10836 5908
rect 14096 5856 14148 5908
rect 15292 5856 15344 5908
rect 16304 5856 16356 5908
rect 18144 5856 18196 5908
rect 22560 5856 22612 5908
rect 27804 5856 27856 5908
rect 28632 5856 28684 5908
rect 30472 5899 30524 5908
rect 30472 5865 30481 5899
rect 30481 5865 30515 5899
rect 30515 5865 30524 5899
rect 30472 5856 30524 5865
rect 32036 5899 32088 5908
rect 32036 5865 32045 5899
rect 32045 5865 32079 5899
rect 32079 5865 32088 5899
rect 32036 5856 32088 5865
rect 32220 5899 32272 5908
rect 32220 5865 32229 5899
rect 32229 5865 32263 5899
rect 32263 5865 32272 5899
rect 32220 5856 32272 5865
rect 10692 5788 10744 5840
rect 12440 5720 12492 5772
rect 14924 5763 14976 5772
rect 5632 5584 5684 5636
rect 8208 5516 8260 5568
rect 9864 5516 9916 5568
rect 10048 5559 10100 5568
rect 10048 5525 10057 5559
rect 10057 5525 10091 5559
rect 10091 5525 10100 5559
rect 10048 5516 10100 5525
rect 10692 5652 10744 5704
rect 10416 5627 10468 5636
rect 10416 5593 10425 5627
rect 10425 5593 10459 5627
rect 10459 5593 10468 5627
rect 10416 5584 10468 5593
rect 12440 5584 12492 5636
rect 12992 5652 13044 5704
rect 14924 5729 14933 5763
rect 14933 5729 14967 5763
rect 14967 5729 14976 5763
rect 14924 5720 14976 5729
rect 14556 5652 14608 5704
rect 15200 5652 15252 5704
rect 15752 5720 15804 5772
rect 17132 5695 17184 5704
rect 17132 5661 17141 5695
rect 17141 5661 17175 5695
rect 17175 5661 17184 5695
rect 17132 5652 17184 5661
rect 23204 5788 23256 5840
rect 27528 5788 27580 5840
rect 29368 5788 29420 5840
rect 19340 5720 19392 5772
rect 19524 5720 19576 5772
rect 19800 5720 19852 5772
rect 20076 5695 20128 5704
rect 20076 5661 20085 5695
rect 20085 5661 20119 5695
rect 20119 5661 20128 5695
rect 20076 5652 20128 5661
rect 20444 5695 20496 5704
rect 20444 5661 20453 5695
rect 20453 5661 20487 5695
rect 20487 5661 20496 5695
rect 20444 5652 20496 5661
rect 20536 5652 20588 5704
rect 24216 5720 24268 5772
rect 14188 5584 14240 5636
rect 10692 5516 10744 5568
rect 11704 5516 11756 5568
rect 13636 5516 13688 5568
rect 15936 5584 15988 5636
rect 16120 5584 16172 5636
rect 22652 5652 22704 5704
rect 22928 5695 22980 5704
rect 22928 5661 22937 5695
rect 22937 5661 22971 5695
rect 22971 5661 22980 5695
rect 22928 5652 22980 5661
rect 23112 5695 23164 5704
rect 23112 5661 23121 5695
rect 23121 5661 23155 5695
rect 23155 5661 23164 5695
rect 23112 5652 23164 5661
rect 23296 5652 23348 5704
rect 23572 5695 23624 5704
rect 23572 5661 23581 5695
rect 23581 5661 23615 5695
rect 23615 5661 23624 5695
rect 23572 5652 23624 5661
rect 23664 5695 23716 5704
rect 23664 5661 23673 5695
rect 23673 5661 23707 5695
rect 23707 5661 23716 5695
rect 23664 5652 23716 5661
rect 24768 5652 24820 5704
rect 29184 5720 29236 5772
rect 30012 5652 30064 5704
rect 31760 5652 31812 5704
rect 32128 5695 32180 5704
rect 32128 5661 32137 5695
rect 32137 5661 32171 5695
rect 32171 5661 32180 5695
rect 32128 5652 32180 5661
rect 14372 5559 14424 5568
rect 14372 5525 14381 5559
rect 14381 5525 14415 5559
rect 14415 5525 14424 5559
rect 14372 5516 14424 5525
rect 15384 5516 15436 5568
rect 19616 5516 19668 5568
rect 20996 5516 21048 5568
rect 30196 5584 30248 5636
rect 30288 5627 30340 5636
rect 30288 5593 30297 5627
rect 30297 5593 30331 5627
rect 30331 5593 30340 5627
rect 30288 5584 30340 5593
rect 22928 5516 22980 5568
rect 23756 5516 23808 5568
rect 24400 5559 24452 5568
rect 24400 5525 24409 5559
rect 24409 5525 24443 5559
rect 24443 5525 24452 5559
rect 24400 5516 24452 5525
rect 29460 5516 29512 5568
rect 31944 5584 31996 5636
rect 4874 5414 4926 5466
rect 4938 5414 4990 5466
rect 5002 5414 5054 5466
rect 5066 5414 5118 5466
rect 5130 5414 5182 5466
rect 35594 5414 35646 5466
rect 35658 5414 35710 5466
rect 35722 5414 35774 5466
rect 35786 5414 35838 5466
rect 35850 5414 35902 5466
rect 5632 5312 5684 5364
rect 7380 5312 7432 5364
rect 8852 5355 8904 5364
rect 8852 5321 8861 5355
rect 8861 5321 8895 5355
rect 8895 5321 8904 5355
rect 8852 5312 8904 5321
rect 8208 5219 8260 5228
rect 8208 5185 8217 5219
rect 8217 5185 8251 5219
rect 8251 5185 8260 5219
rect 8208 5176 8260 5185
rect 9036 5176 9088 5228
rect 9864 5312 9916 5364
rect 9864 5176 9916 5228
rect 10416 5244 10468 5296
rect 10048 5176 10100 5228
rect 11888 5312 11940 5364
rect 12164 5312 12216 5364
rect 11704 5244 11756 5296
rect 12900 5176 12952 5228
rect 15200 5355 15252 5364
rect 15200 5321 15209 5355
rect 15209 5321 15243 5355
rect 15243 5321 15252 5355
rect 15200 5312 15252 5321
rect 17132 5312 17184 5364
rect 20168 5312 20220 5364
rect 20444 5312 20496 5364
rect 23572 5312 23624 5364
rect 23664 5355 23716 5364
rect 23664 5321 23673 5355
rect 23673 5321 23707 5355
rect 23707 5321 23716 5355
rect 23664 5312 23716 5321
rect 27620 5312 27672 5364
rect 13636 5244 13688 5296
rect 9680 5108 9732 5160
rect 12992 5108 13044 5160
rect 16120 5244 16172 5296
rect 19340 5287 19392 5296
rect 19340 5253 19349 5287
rect 19349 5253 19383 5287
rect 19383 5253 19392 5287
rect 19340 5244 19392 5253
rect 19524 5287 19576 5296
rect 19524 5253 19533 5287
rect 19533 5253 19567 5287
rect 19567 5253 19576 5287
rect 19524 5244 19576 5253
rect 20996 5244 21048 5296
rect 20904 5219 20956 5228
rect 20904 5185 20913 5219
rect 20913 5185 20947 5219
rect 20947 5185 20956 5219
rect 20904 5176 20956 5185
rect 22652 5176 22704 5228
rect 23020 5219 23072 5228
rect 23020 5185 23029 5219
rect 23029 5185 23063 5219
rect 23063 5185 23072 5219
rect 23020 5176 23072 5185
rect 23112 5176 23164 5228
rect 23204 5219 23256 5228
rect 23204 5185 23213 5219
rect 23213 5185 23247 5219
rect 23247 5185 23256 5219
rect 23204 5176 23256 5185
rect 15384 5108 15436 5160
rect 15844 5151 15896 5160
rect 15844 5117 15853 5151
rect 15853 5117 15887 5151
rect 15887 5117 15896 5151
rect 15844 5108 15896 5117
rect 16672 5151 16724 5160
rect 16672 5117 16681 5151
rect 16681 5117 16715 5151
rect 16715 5117 16724 5151
rect 16672 5108 16724 5117
rect 22376 5151 22428 5160
rect 22376 5117 22385 5151
rect 22385 5117 22419 5151
rect 22419 5117 22428 5151
rect 22376 5108 22428 5117
rect 23296 5040 23348 5092
rect 24860 5176 24912 5228
rect 25504 5176 25556 5228
rect 26240 5176 26292 5228
rect 27620 5219 27672 5228
rect 27620 5185 27629 5219
rect 27629 5185 27663 5219
rect 27663 5185 27672 5219
rect 27620 5176 27672 5185
rect 27712 5219 27764 5228
rect 27712 5185 27721 5219
rect 27721 5185 27755 5219
rect 27755 5185 27764 5219
rect 27712 5176 27764 5185
rect 27804 5176 27856 5228
rect 28448 5244 28500 5296
rect 29736 5312 29788 5364
rect 30288 5312 30340 5364
rect 32128 5312 32180 5364
rect 29368 5244 29420 5296
rect 24400 5108 24452 5160
rect 26976 5108 27028 5160
rect 28264 5108 28316 5160
rect 29460 5176 29512 5228
rect 30380 5244 30432 5296
rect 26056 5040 26108 5092
rect 29184 5040 29236 5092
rect 9128 5015 9180 5024
rect 9128 4981 9137 5015
rect 9137 4981 9171 5015
rect 9171 4981 9180 5015
rect 9128 4972 9180 4981
rect 11152 5015 11204 5024
rect 11152 4981 11161 5015
rect 11161 4981 11195 5015
rect 11195 4981 11204 5015
rect 11152 4972 11204 4981
rect 16396 5015 16448 5024
rect 16396 4981 16405 5015
rect 16405 4981 16439 5015
rect 16439 4981 16448 5015
rect 16396 4972 16448 4981
rect 19892 5015 19944 5024
rect 19892 4981 19901 5015
rect 19901 4981 19935 5015
rect 19935 4981 19944 5015
rect 19892 4972 19944 4981
rect 23388 4972 23440 5024
rect 24400 4972 24452 5024
rect 29828 5176 29880 5228
rect 30104 5176 30156 5228
rect 29828 5083 29880 5092
rect 29828 5049 29837 5083
rect 29837 5049 29871 5083
rect 29871 5049 29880 5083
rect 29828 5040 29880 5049
rect 30012 4972 30064 5024
rect 30288 5015 30340 5024
rect 30288 4981 30297 5015
rect 30297 4981 30331 5015
rect 30331 4981 30340 5015
rect 30288 4972 30340 4981
rect 30656 5083 30708 5092
rect 30656 5049 30665 5083
rect 30665 5049 30699 5083
rect 30699 5049 30708 5083
rect 30656 5040 30708 5049
rect 31760 5176 31812 5228
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 9864 4811 9916 4820
rect 9864 4777 9873 4811
rect 9873 4777 9907 4811
rect 9907 4777 9916 4811
rect 9864 4768 9916 4777
rect 11152 4768 11204 4820
rect 12440 4811 12492 4820
rect 12440 4777 12449 4811
rect 12449 4777 12483 4811
rect 12483 4777 12492 4811
rect 12440 4768 12492 4777
rect 15844 4768 15896 4820
rect 16396 4768 16448 4820
rect 16672 4768 16724 4820
rect 19432 4768 19484 4820
rect 20168 4811 20220 4820
rect 20168 4777 20177 4811
rect 20177 4777 20211 4811
rect 20211 4777 20220 4811
rect 20168 4768 20220 4777
rect 20904 4768 20956 4820
rect 23388 4768 23440 4820
rect 23572 4768 23624 4820
rect 24400 4811 24452 4820
rect 24400 4777 24409 4811
rect 24409 4777 24443 4811
rect 24443 4777 24452 4811
rect 24400 4768 24452 4777
rect 12164 4632 12216 4684
rect 19892 4700 19944 4752
rect 25504 4768 25556 4820
rect 26056 4811 26108 4820
rect 26056 4777 26065 4811
rect 26065 4777 26099 4811
rect 26099 4777 26108 4811
rect 26056 4768 26108 4777
rect 27620 4768 27672 4820
rect 29184 4768 29236 4820
rect 30012 4811 30064 4820
rect 30012 4777 30021 4811
rect 30021 4777 30055 4811
rect 30055 4777 30064 4811
rect 30012 4768 30064 4777
rect 30288 4768 30340 4820
rect 3884 4564 3936 4616
rect 9772 4564 9824 4616
rect 10232 4607 10284 4616
rect 10232 4573 10241 4607
rect 10241 4573 10275 4607
rect 10275 4573 10284 4607
rect 10232 4564 10284 4573
rect 15936 4564 15988 4616
rect 16304 4607 16356 4616
rect 16304 4573 16313 4607
rect 16313 4573 16347 4607
rect 16347 4573 16356 4607
rect 16304 4564 16356 4573
rect 16488 4564 16540 4616
rect 20812 4564 20864 4616
rect 22928 4632 22980 4684
rect 24676 4700 24728 4752
rect 23756 4632 23808 4684
rect 24584 4675 24636 4684
rect 24584 4641 24593 4675
rect 24593 4641 24627 4675
rect 24627 4641 24636 4675
rect 24584 4632 24636 4641
rect 24860 4700 24912 4752
rect 27804 4700 27856 4752
rect 29368 4700 29420 4752
rect 940 4496 992 4548
rect 12900 4496 12952 4548
rect 14464 4539 14516 4548
rect 14464 4505 14473 4539
rect 14473 4505 14507 4539
rect 14507 4505 14516 4539
rect 14464 4496 14516 4505
rect 16764 4428 16816 4480
rect 20076 4496 20128 4548
rect 20536 4496 20588 4548
rect 22652 4496 22704 4548
rect 23204 4428 23256 4480
rect 23480 4539 23532 4548
rect 23480 4505 23489 4539
rect 23489 4505 23523 4539
rect 23523 4505 23532 4539
rect 23480 4496 23532 4505
rect 24584 4496 24636 4548
rect 24952 4564 25004 4616
rect 25412 4632 25464 4684
rect 26976 4632 27028 4684
rect 23388 4428 23440 4480
rect 25044 4428 25096 4480
rect 26332 4607 26384 4616
rect 26332 4573 26341 4607
rect 26341 4573 26375 4607
rect 26375 4573 26384 4607
rect 27988 4675 28040 4684
rect 27988 4641 27997 4675
rect 27997 4641 28031 4675
rect 28031 4641 28040 4675
rect 27988 4632 28040 4641
rect 28080 4632 28132 4684
rect 26332 4564 26384 4573
rect 30196 4607 30248 4616
rect 30196 4573 30205 4607
rect 30205 4573 30239 4607
rect 30239 4573 30248 4607
rect 30196 4564 30248 4573
rect 30380 4564 30432 4616
rect 27712 4428 27764 4480
rect 31944 4428 31996 4480
rect 4874 4326 4926 4378
rect 4938 4326 4990 4378
rect 5002 4326 5054 4378
rect 5066 4326 5118 4378
rect 5130 4326 5182 4378
rect 35594 4326 35646 4378
rect 35658 4326 35710 4378
rect 35722 4326 35774 4378
rect 35786 4326 35838 4378
rect 35850 4326 35902 4378
rect 9128 4224 9180 4276
rect 9680 4224 9732 4276
rect 14464 4224 14516 4276
rect 20996 4224 21048 4276
rect 8392 4156 8444 4208
rect 22652 4156 22704 4208
rect 23480 4156 23532 4208
rect 25044 4156 25096 4208
rect 26332 4224 26384 4276
rect 27988 4224 28040 4276
rect 6920 4088 6972 4140
rect 14372 4131 14424 4140
rect 14372 4097 14381 4131
rect 14381 4097 14415 4131
rect 14415 4097 14424 4131
rect 14372 4088 14424 4097
rect 25504 4088 25556 4140
rect 29828 4156 29880 4208
rect 30656 4156 30708 4208
rect 30104 4088 30156 4140
rect 25412 3952 25464 4004
rect 25504 3884 25556 3936
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 4874 3238 4926 3290
rect 4938 3238 4990 3290
rect 5002 3238 5054 3290
rect 5066 3238 5118 3290
rect 5130 3238 5182 3290
rect 35594 3238 35646 3290
rect 35658 3238 35710 3290
rect 35722 3238 35774 3290
rect 35786 3238 35838 3290
rect 35850 3238 35902 3290
rect 17224 3136 17276 3188
rect 1952 3043 2004 3052
rect 1952 3009 1961 3043
rect 1961 3009 1995 3043
rect 1995 3009 2004 3043
rect 1952 3000 2004 3009
rect 2412 3043 2464 3052
rect 2412 3009 2421 3043
rect 2421 3009 2455 3043
rect 2455 3009 2464 3043
rect 2412 3000 2464 3009
rect 12532 3043 12584 3052
rect 12532 3009 12541 3043
rect 12541 3009 12575 3043
rect 12575 3009 12584 3043
rect 12532 3000 12584 3009
rect 13176 3043 13228 3052
rect 13176 3009 13185 3043
rect 13185 3009 13219 3043
rect 13219 3009 13228 3043
rect 13176 3000 13228 3009
rect 15108 3043 15160 3052
rect 15108 3009 15117 3043
rect 15117 3009 15151 3043
rect 15151 3009 15160 3043
rect 15108 3000 15160 3009
rect 37556 3111 37608 3120
rect 37556 3077 37565 3111
rect 37565 3077 37599 3111
rect 37599 3077 37608 3111
rect 37556 3068 37608 3077
rect 25596 3000 25648 3052
rect 1768 2839 1820 2848
rect 1768 2805 1777 2839
rect 1777 2805 1811 2839
rect 1811 2805 1820 2839
rect 1768 2796 1820 2805
rect 2228 2839 2280 2848
rect 2228 2805 2237 2839
rect 2237 2805 2271 2839
rect 2271 2805 2280 2839
rect 2228 2796 2280 2805
rect 8392 2796 8444 2848
rect 12992 2839 13044 2848
rect 12992 2805 13001 2839
rect 13001 2805 13035 2839
rect 13035 2805 13044 2839
rect 12992 2796 13044 2805
rect 14924 2839 14976 2848
rect 14924 2805 14933 2839
rect 14933 2805 14967 2839
rect 14967 2805 14976 2839
rect 14924 2796 14976 2805
rect 17408 2839 17460 2848
rect 17408 2805 17417 2839
rect 17417 2805 17451 2839
rect 17451 2805 17460 2839
rect 17408 2796 17460 2805
rect 19800 2839 19852 2848
rect 19800 2805 19809 2839
rect 19809 2805 19843 2839
rect 19843 2805 19852 2839
rect 19800 2796 19852 2805
rect 37188 2796 37240 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 8760 2592 8812 2644
rect 10140 2592 10192 2644
rect 8944 2456 8996 2508
rect 1768 2431 1820 2440
rect 1768 2397 1777 2431
rect 1777 2397 1811 2431
rect 1811 2397 1820 2431
rect 1768 2388 1820 2397
rect 2228 2388 2280 2440
rect 5448 2388 5500 2440
rect 8392 2388 8444 2440
rect 8484 2431 8536 2440
rect 8484 2397 8493 2431
rect 8493 2397 8527 2431
rect 8527 2397 8536 2431
rect 8484 2388 8536 2397
rect 12992 2388 13044 2440
rect 14924 2388 14976 2440
rect 17408 2388 17460 2440
rect 19800 2431 19852 2440
rect 19800 2397 19809 2431
rect 19809 2397 19843 2431
rect 19843 2397 19852 2431
rect 19800 2388 19852 2397
rect 37464 2431 37516 2440
rect 37464 2397 37473 2431
rect 37473 2397 37507 2431
rect 37507 2397 37516 2431
rect 37464 2388 37516 2397
rect 20 2320 72 2372
rect 2044 2363 2096 2372
rect 2044 2329 2053 2363
rect 2053 2329 2087 2363
rect 2087 2329 2096 2363
rect 2044 2320 2096 2329
rect 3976 2363 4028 2372
rect 3976 2329 3985 2363
rect 3985 2329 4019 2363
rect 4019 2329 4028 2363
rect 3976 2320 4028 2329
rect 6552 2363 6604 2372
rect 6552 2329 6561 2363
rect 6561 2329 6595 2363
rect 6595 2329 6604 2363
rect 6552 2320 6604 2329
rect 10968 2320 11020 2372
rect 14648 2320 14700 2372
rect 12900 2252 12952 2304
rect 15016 2252 15068 2304
rect 17408 2252 17460 2304
rect 19432 2363 19484 2372
rect 19432 2329 19441 2363
rect 19441 2329 19475 2363
rect 19475 2329 19484 2363
rect 19432 2320 19484 2329
rect 26424 2252 26476 2304
rect 4874 2150 4926 2202
rect 4938 2150 4990 2202
rect 5002 2150 5054 2202
rect 5066 2150 5118 2202
rect 5130 2150 5182 2202
rect 35594 2150 35646 2202
rect 35658 2150 35710 2202
rect 35722 2150 35774 2202
rect 35786 2150 35838 2202
rect 35850 2150 35902 2202
<< metal2 >>
rect 18 40762 74 41562
rect 1950 40762 2006 41562
rect 4526 40762 4582 41562
rect 6458 40762 6514 41562
rect 9034 40762 9090 41562
rect 10966 40762 11022 41562
rect 12898 40882 12954 41562
rect 12898 40854 13216 40882
rect 12898 40762 12954 40854
rect 32 39098 60 40762
rect 4540 39098 4568 40762
rect 4874 39196 5182 39205
rect 4874 39194 4880 39196
rect 4936 39194 4960 39196
rect 5016 39194 5040 39196
rect 5096 39194 5120 39196
rect 5176 39194 5182 39196
rect 4936 39142 4938 39194
rect 5118 39142 5120 39194
rect 4874 39140 4880 39142
rect 4936 39140 4960 39142
rect 5016 39140 5040 39142
rect 5096 39140 5120 39142
rect 5176 39140 5182 39142
rect 4874 39131 5182 39140
rect 9048 39098 9076 40762
rect 10980 39114 11008 40762
rect 10980 39098 11100 39114
rect 13188 39098 13216 40854
rect 15474 40762 15530 41562
rect 17406 40762 17462 41562
rect 19982 40882 20038 41562
rect 19982 40854 20116 40882
rect 19982 40762 20038 40854
rect 20 39092 72 39098
rect 20 39034 72 39040
rect 4528 39092 4580 39098
rect 4528 39034 4580 39040
rect 9036 39092 9088 39098
rect 10980 39092 11112 39098
rect 10980 39086 11060 39092
rect 9036 39034 9088 39040
rect 11060 39034 11112 39040
rect 13176 39092 13228 39098
rect 13176 39034 13228 39040
rect 15488 39030 15516 40762
rect 17420 39098 17448 40762
rect 17408 39092 17460 39098
rect 17408 39034 17460 39040
rect 12348 39024 12400 39030
rect 12348 38966 12400 38972
rect 15476 39024 15528 39030
rect 15476 38966 15528 38972
rect 1768 38956 1820 38962
rect 1768 38898 1820 38904
rect 5080 38956 5132 38962
rect 5080 38898 5132 38904
rect 9220 38956 9272 38962
rect 9220 38898 9272 38904
rect 12072 38956 12124 38962
rect 12072 38898 12124 38904
rect 940 37188 992 37194
rect 940 37130 992 37136
rect 952 36825 980 37130
rect 938 36816 994 36825
rect 938 36751 994 36760
rect 1780 35894 1808 38898
rect 4214 38652 4522 38661
rect 4214 38650 4220 38652
rect 4276 38650 4300 38652
rect 4356 38650 4380 38652
rect 4436 38650 4460 38652
rect 4516 38650 4522 38652
rect 4276 38598 4278 38650
rect 4458 38598 4460 38650
rect 4214 38596 4220 38598
rect 4276 38596 4300 38598
rect 4356 38596 4380 38598
rect 4436 38596 4460 38598
rect 4516 38596 4522 38598
rect 4214 38587 4522 38596
rect 5092 38554 5120 38898
rect 9232 38554 9260 38898
rect 5080 38548 5132 38554
rect 5080 38490 5132 38496
rect 9220 38548 9272 38554
rect 9220 38490 9272 38496
rect 5170 38448 5226 38457
rect 5170 38383 5226 38392
rect 5184 38350 5212 38383
rect 5172 38344 5224 38350
rect 5172 38286 5224 38292
rect 8576 38344 8628 38350
rect 8576 38286 8628 38292
rect 9036 38344 9088 38350
rect 9036 38286 9088 38292
rect 4874 38108 5182 38117
rect 4874 38106 4880 38108
rect 4936 38106 4960 38108
rect 5016 38106 5040 38108
rect 5096 38106 5120 38108
rect 5176 38106 5182 38108
rect 4936 38054 4938 38106
rect 5118 38054 5120 38106
rect 4874 38052 4880 38054
rect 4936 38052 4960 38054
rect 5016 38052 5040 38054
rect 5096 38052 5120 38054
rect 5176 38052 5182 38054
rect 4874 38043 5182 38052
rect 4214 37564 4522 37573
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37499 4522 37508
rect 8392 37324 8444 37330
rect 8392 37266 8444 37272
rect 8300 37256 8352 37262
rect 8300 37198 8352 37204
rect 6920 37188 6972 37194
rect 6920 37130 6972 37136
rect 4874 37020 5182 37029
rect 4874 37018 4880 37020
rect 4936 37018 4960 37020
rect 5016 37018 5040 37020
rect 5096 37018 5120 37020
rect 5176 37018 5182 37020
rect 4936 36966 4938 37018
rect 5118 36966 5120 37018
rect 4874 36964 4880 36966
rect 4936 36964 4960 36966
rect 5016 36964 5040 36966
rect 5096 36964 5120 36966
rect 5176 36964 5182 36966
rect 4874 36955 5182 36964
rect 4214 36476 4522 36485
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36411 4522 36420
rect 4712 36168 4764 36174
rect 4712 36110 4764 36116
rect 1780 35866 2176 35894
rect 1768 25900 1820 25906
rect 1768 25842 1820 25848
rect 940 25696 992 25702
rect 940 25638 992 25644
rect 952 25265 980 25638
rect 1400 25288 1452 25294
rect 938 25256 994 25265
rect 1400 25230 1452 25236
rect 938 25191 994 25200
rect 1412 24750 1440 25230
rect 1400 24744 1452 24750
rect 1400 24686 1452 24692
rect 1676 24744 1728 24750
rect 1676 24686 1728 24692
rect 1412 24342 1440 24686
rect 1688 24410 1716 24686
rect 1676 24404 1728 24410
rect 1676 24346 1728 24352
rect 1400 24336 1452 24342
rect 1400 24278 1452 24284
rect 1412 21486 1440 24278
rect 1780 23322 1808 25842
rect 1860 25832 1912 25838
rect 1860 25774 1912 25780
rect 1872 25294 1900 25774
rect 1860 25288 1912 25294
rect 1860 25230 1912 25236
rect 1952 23860 2004 23866
rect 1952 23802 2004 23808
rect 1768 23316 1820 23322
rect 1768 23258 1820 23264
rect 1964 23118 1992 23802
rect 1952 23112 2004 23118
rect 1952 23054 2004 23060
rect 1860 22976 1912 22982
rect 1860 22918 1912 22924
rect 1768 21888 1820 21894
rect 1768 21830 1820 21836
rect 1780 21690 1808 21830
rect 1768 21684 1820 21690
rect 1768 21626 1820 21632
rect 1400 21480 1452 21486
rect 1400 21422 1452 21428
rect 1412 19514 1440 21422
rect 1872 20942 1900 22918
rect 1952 22024 2004 22030
rect 1952 21966 2004 21972
rect 1964 21690 1992 21966
rect 1952 21684 2004 21690
rect 1952 21626 2004 21632
rect 1860 20936 1912 20942
rect 1860 20878 1912 20884
rect 1492 20800 1544 20806
rect 1492 20742 1544 20748
rect 1504 20641 1532 20742
rect 1490 20632 1546 20641
rect 1490 20567 1546 20576
rect 1768 19712 1820 19718
rect 1768 19654 1820 19660
rect 1400 19508 1452 19514
rect 1400 19450 1452 19456
rect 1780 19446 1808 19654
rect 1768 19440 1820 19446
rect 1768 19382 1820 19388
rect 940 18692 992 18698
rect 940 18634 992 18640
rect 1768 18692 1820 18698
rect 1768 18634 1820 18640
rect 952 18465 980 18634
rect 938 18456 994 18465
rect 938 18391 994 18400
rect 1676 18216 1728 18222
rect 1676 18158 1728 18164
rect 1688 17746 1716 18158
rect 1780 17882 1808 18634
rect 1952 18624 2004 18630
rect 1952 18566 2004 18572
rect 1768 17876 1820 17882
rect 1768 17818 1820 17824
rect 1676 17740 1728 17746
rect 1676 17682 1728 17688
rect 1964 17678 1992 18566
rect 2044 18080 2096 18086
rect 2044 18022 2096 18028
rect 2056 17678 2084 18022
rect 2148 17882 2176 35866
rect 4214 35388 4522 35397
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35323 4522 35332
rect 4214 34300 4522 34309
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34235 4522 34244
rect 4724 33998 4752 36110
rect 6276 36100 6328 36106
rect 6276 36042 6328 36048
rect 4874 35932 5182 35941
rect 4874 35930 4880 35932
rect 4936 35930 4960 35932
rect 5016 35930 5040 35932
rect 5096 35930 5120 35932
rect 5176 35930 5182 35932
rect 4936 35878 4938 35930
rect 5118 35878 5120 35930
rect 4874 35876 4880 35878
rect 4936 35876 4960 35878
rect 5016 35876 5040 35878
rect 5096 35876 5120 35878
rect 5176 35876 5182 35878
rect 4874 35867 5182 35876
rect 6288 35834 6316 36042
rect 6644 36032 6696 36038
rect 6644 35974 6696 35980
rect 6276 35828 6328 35834
rect 6276 35770 6328 35776
rect 4874 34844 5182 34853
rect 4874 34842 4880 34844
rect 4936 34842 4960 34844
rect 5016 34842 5040 34844
rect 5096 34842 5120 34844
rect 5176 34842 5182 34844
rect 4936 34790 4938 34842
rect 5118 34790 5120 34842
rect 4874 34788 4880 34790
rect 4936 34788 4960 34790
rect 5016 34788 5040 34790
rect 5096 34788 5120 34790
rect 5176 34788 5182 34790
rect 4874 34779 5182 34788
rect 5632 34604 5684 34610
rect 5632 34546 5684 34552
rect 5356 34400 5408 34406
rect 5356 34342 5408 34348
rect 5368 34066 5396 34342
rect 5356 34060 5408 34066
rect 5356 34002 5408 34008
rect 4712 33992 4764 33998
rect 4764 33952 4844 33980
rect 4712 33934 4764 33940
rect 4214 33212 4522 33221
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33147 4522 33156
rect 4620 32972 4672 32978
rect 4620 32914 4672 32920
rect 4214 32124 4522 32133
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32059 4522 32068
rect 4632 32026 4660 32914
rect 4712 32836 4764 32842
rect 4712 32778 4764 32784
rect 4724 32570 4752 32778
rect 4712 32564 4764 32570
rect 4712 32506 4764 32512
rect 4620 32020 4672 32026
rect 4620 31962 4672 31968
rect 4214 31036 4522 31045
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30971 4522 30980
rect 4632 30598 4660 31962
rect 4816 30734 4844 33952
rect 4874 33756 5182 33765
rect 4874 33754 4880 33756
rect 4936 33754 4960 33756
rect 5016 33754 5040 33756
rect 5096 33754 5120 33756
rect 5176 33754 5182 33756
rect 4936 33702 4938 33754
rect 5118 33702 5120 33754
rect 4874 33700 4880 33702
rect 4936 33700 4960 33702
rect 5016 33700 5040 33702
rect 5096 33700 5120 33702
rect 5176 33700 5182 33702
rect 4874 33691 5182 33700
rect 5644 33658 5672 34546
rect 6656 33998 6684 35974
rect 6932 35222 6960 37130
rect 8312 36922 8340 37198
rect 8300 36916 8352 36922
rect 8300 36858 8352 36864
rect 8404 36854 8432 37266
rect 8392 36848 8444 36854
rect 8392 36790 8444 36796
rect 7656 36576 7708 36582
rect 7656 36518 7708 36524
rect 7668 36106 7696 36518
rect 7656 36100 7708 36106
rect 7656 36042 7708 36048
rect 7748 36032 7800 36038
rect 7748 35974 7800 35980
rect 7760 35834 7788 35974
rect 7748 35828 7800 35834
rect 7748 35770 7800 35776
rect 8208 35828 8260 35834
rect 8208 35770 8260 35776
rect 7840 35624 7892 35630
rect 7840 35566 7892 35572
rect 8116 35624 8168 35630
rect 8116 35566 8168 35572
rect 6920 35216 6972 35222
rect 6920 35158 6972 35164
rect 6736 34196 6788 34202
rect 6736 34138 6788 34144
rect 6368 33992 6420 33998
rect 6368 33934 6420 33940
rect 6644 33992 6696 33998
rect 6644 33934 6696 33940
rect 5632 33652 5684 33658
rect 5632 33594 5684 33600
rect 5908 33448 5960 33454
rect 5908 33390 5960 33396
rect 5920 32910 5948 33390
rect 5908 32904 5960 32910
rect 5908 32846 5960 32852
rect 6380 32842 6408 33934
rect 6748 33658 6776 34138
rect 6932 34066 6960 35158
rect 7196 35012 7248 35018
rect 7196 34954 7248 34960
rect 7208 34746 7236 34954
rect 7196 34740 7248 34746
rect 7196 34682 7248 34688
rect 6920 34060 6972 34066
rect 6920 34002 6972 34008
rect 7564 33992 7616 33998
rect 7564 33934 7616 33940
rect 7196 33856 7248 33862
rect 7196 33798 7248 33804
rect 7208 33658 7236 33798
rect 6736 33652 6788 33658
rect 6736 33594 6788 33600
rect 7196 33652 7248 33658
rect 7196 33594 7248 33600
rect 7288 33448 7340 33454
rect 7288 33390 7340 33396
rect 7012 33312 7064 33318
rect 7012 33254 7064 33260
rect 6736 32972 6788 32978
rect 6736 32914 6788 32920
rect 6828 32972 6880 32978
rect 6828 32914 6880 32920
rect 6644 32904 6696 32910
rect 6644 32846 6696 32852
rect 6368 32836 6420 32842
rect 6368 32778 6420 32784
rect 6276 32768 6328 32774
rect 6276 32710 6328 32716
rect 4874 32668 5182 32677
rect 4874 32666 4880 32668
rect 4936 32666 4960 32668
rect 5016 32666 5040 32668
rect 5096 32666 5120 32668
rect 5176 32666 5182 32668
rect 4936 32614 4938 32666
rect 5118 32614 5120 32666
rect 4874 32612 4880 32614
rect 4936 32612 4960 32614
rect 5016 32612 5040 32614
rect 5096 32612 5120 32614
rect 5176 32612 5182 32614
rect 4874 32603 5182 32612
rect 6288 32570 6316 32710
rect 6276 32564 6328 32570
rect 6276 32506 6328 32512
rect 5724 32292 5776 32298
rect 5724 32234 5776 32240
rect 5736 31770 5764 32234
rect 5816 31816 5868 31822
rect 5736 31764 5816 31770
rect 5736 31758 5868 31764
rect 5736 31742 5856 31758
rect 4874 31580 5182 31589
rect 4874 31578 4880 31580
rect 4936 31578 4960 31580
rect 5016 31578 5040 31580
rect 5096 31578 5120 31580
rect 5176 31578 5182 31580
rect 4936 31526 4938 31578
rect 5118 31526 5120 31578
rect 4874 31524 4880 31526
rect 4936 31524 4960 31526
rect 5016 31524 5040 31526
rect 5096 31524 5120 31526
rect 5176 31524 5182 31526
rect 4874 31515 5182 31524
rect 4804 30728 4856 30734
rect 4804 30670 4856 30676
rect 5632 30728 5684 30734
rect 5632 30670 5684 30676
rect 4252 30592 4304 30598
rect 4252 30534 4304 30540
rect 4620 30592 4672 30598
rect 4620 30534 4672 30540
rect 4264 30190 4292 30534
rect 4252 30184 4304 30190
rect 4252 30126 4304 30132
rect 4214 29948 4522 29957
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29883 4522 29892
rect 4632 29578 4660 30534
rect 4874 30492 5182 30501
rect 4874 30490 4880 30492
rect 4936 30490 4960 30492
rect 5016 30490 5040 30492
rect 5096 30490 5120 30492
rect 5176 30490 5182 30492
rect 4936 30438 4938 30490
rect 5118 30438 5120 30490
rect 4874 30436 4880 30438
rect 4936 30436 4960 30438
rect 5016 30436 5040 30438
rect 5096 30436 5120 30438
rect 5176 30436 5182 30438
rect 4874 30427 5182 30436
rect 5264 30320 5316 30326
rect 5264 30262 5316 30268
rect 5276 30054 5304 30262
rect 5264 30048 5316 30054
rect 5264 29990 5316 29996
rect 4620 29572 4672 29578
rect 4620 29514 4672 29520
rect 4068 29504 4120 29510
rect 4068 29446 4120 29452
rect 4080 29306 4108 29446
rect 4068 29300 4120 29306
rect 4068 29242 4120 29248
rect 4214 28860 4522 28869
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28795 4522 28804
rect 4252 28416 4304 28422
rect 4252 28358 4304 28364
rect 4264 28218 4292 28358
rect 4252 28212 4304 28218
rect 4252 28154 4304 28160
rect 4214 27772 4522 27781
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27707 4522 27716
rect 4066 27296 4122 27305
rect 4066 27231 4122 27240
rect 3884 26240 3936 26246
rect 3884 26182 3936 26188
rect 3896 25974 3924 26182
rect 3884 25968 3936 25974
rect 3884 25910 3936 25916
rect 3056 25900 3108 25906
rect 3056 25842 3108 25848
rect 3240 25900 3292 25906
rect 3240 25842 3292 25848
rect 2872 25696 2924 25702
rect 2872 25638 2924 25644
rect 2884 25362 2912 25638
rect 2872 25356 2924 25362
rect 2872 25298 2924 25304
rect 2964 25152 3016 25158
rect 2964 25094 3016 25100
rect 2976 24818 3004 25094
rect 2964 24812 3016 24818
rect 2964 24754 3016 24760
rect 2688 24608 2740 24614
rect 2688 24550 2740 24556
rect 2700 24070 2728 24550
rect 2504 24064 2556 24070
rect 2504 24006 2556 24012
rect 2688 24064 2740 24070
rect 2688 24006 2740 24012
rect 2780 24064 2832 24070
rect 2780 24006 2832 24012
rect 2516 23118 2544 24006
rect 2792 23322 2820 24006
rect 2780 23316 2832 23322
rect 2780 23258 2832 23264
rect 2504 23112 2556 23118
rect 2504 23054 2556 23060
rect 2688 23112 2740 23118
rect 2976 23100 3004 24754
rect 3068 24410 3096 25842
rect 3252 25294 3280 25842
rect 3608 25832 3660 25838
rect 3608 25774 3660 25780
rect 3620 25498 3648 25774
rect 3608 25492 3660 25498
rect 3608 25434 3660 25440
rect 3240 25288 3292 25294
rect 3240 25230 3292 25236
rect 3976 24608 4028 24614
rect 3976 24550 4028 24556
rect 3056 24404 3108 24410
rect 3056 24346 3108 24352
rect 3988 24290 4016 24550
rect 4080 24410 4108 27231
rect 4214 26684 4522 26693
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26619 4522 26628
rect 4528 26376 4580 26382
rect 4632 26364 4660 29514
rect 4874 29404 5182 29413
rect 4874 29402 4880 29404
rect 4936 29402 4960 29404
rect 5016 29402 5040 29404
rect 5096 29402 5120 29404
rect 5176 29402 5182 29404
rect 4936 29350 4938 29402
rect 5118 29350 5120 29402
rect 4874 29348 4880 29350
rect 4936 29348 4960 29350
rect 5016 29348 5040 29350
rect 5096 29348 5120 29350
rect 5176 29348 5182 29350
rect 4874 29339 5182 29348
rect 5276 29170 5304 29990
rect 5448 29504 5500 29510
rect 5448 29446 5500 29452
rect 5264 29164 5316 29170
rect 5264 29106 5316 29112
rect 4712 28960 4764 28966
rect 4712 28902 4764 28908
rect 5356 28960 5408 28966
rect 5356 28902 5408 28908
rect 4724 28762 4752 28902
rect 4712 28756 4764 28762
rect 4712 28698 4764 28704
rect 4874 28316 5182 28325
rect 4874 28314 4880 28316
rect 4936 28314 4960 28316
rect 5016 28314 5040 28316
rect 5096 28314 5120 28316
rect 5176 28314 5182 28316
rect 4936 28262 4938 28314
rect 5118 28262 5120 28314
rect 4874 28260 4880 28262
rect 4936 28260 4960 28262
rect 5016 28260 5040 28262
rect 5096 28260 5120 28262
rect 5176 28260 5182 28262
rect 4874 28251 5182 28260
rect 5368 28064 5396 28902
rect 5460 28558 5488 29446
rect 5644 29073 5672 30670
rect 5736 30054 5764 31742
rect 6184 30660 6236 30666
rect 6184 30602 6236 30608
rect 6196 30394 6224 30602
rect 6380 30598 6408 32778
rect 6552 32224 6604 32230
rect 6552 32166 6604 32172
rect 6564 31822 6592 32166
rect 6656 31822 6684 32846
rect 6748 32570 6776 32914
rect 6736 32564 6788 32570
rect 6736 32506 6788 32512
rect 6552 31816 6604 31822
rect 6552 31758 6604 31764
rect 6644 31816 6696 31822
rect 6644 31758 6696 31764
rect 6368 30592 6420 30598
rect 6368 30534 6420 30540
rect 6184 30388 6236 30394
rect 6184 30330 6236 30336
rect 6840 30054 6868 32914
rect 7024 30818 7052 33254
rect 7300 33114 7328 33390
rect 7288 33108 7340 33114
rect 7288 33050 7340 33056
rect 7576 32042 7604 33934
rect 7852 33318 7880 35566
rect 8128 35170 8156 35566
rect 7944 35154 8156 35170
rect 7932 35148 8156 35154
rect 7984 35142 8156 35148
rect 7932 35090 7984 35096
rect 8128 34524 8156 35142
rect 8220 34678 8248 35770
rect 8300 35624 8352 35630
rect 8300 35566 8352 35572
rect 8312 35086 8340 35566
rect 8300 35080 8352 35086
rect 8300 35022 8352 35028
rect 8208 34672 8260 34678
rect 8208 34614 8260 34620
rect 8208 34536 8260 34542
rect 8128 34496 8208 34524
rect 8208 34478 8260 34484
rect 7840 33312 7892 33318
rect 7840 33254 7892 33260
rect 8220 32910 8248 34478
rect 8312 33590 8340 35022
rect 8484 34944 8536 34950
rect 8404 34892 8484 34898
rect 8404 34886 8536 34892
rect 8404 34870 8524 34886
rect 8404 34610 8432 34870
rect 8392 34604 8444 34610
rect 8392 34546 8444 34552
rect 8404 34066 8432 34546
rect 8392 34060 8444 34066
rect 8392 34002 8444 34008
rect 8300 33584 8352 33590
rect 8300 33526 8352 33532
rect 8208 32904 8260 32910
rect 8208 32846 8260 32852
rect 7208 32026 7604 32042
rect 7196 32020 7604 32026
rect 7248 32014 7604 32020
rect 7196 31962 7248 31968
rect 7472 31952 7524 31958
rect 7472 31894 7524 31900
rect 7484 31822 7512 31894
rect 7472 31816 7524 31822
rect 7472 31758 7524 31764
rect 7024 30802 7420 30818
rect 7024 30796 7432 30802
rect 7024 30790 7380 30796
rect 5724 30048 5776 30054
rect 5724 29990 5776 29996
rect 6828 30048 6880 30054
rect 6828 29990 6880 29996
rect 6840 29714 6868 29990
rect 6828 29708 6880 29714
rect 6828 29650 6880 29656
rect 6828 29572 6880 29578
rect 6828 29514 6880 29520
rect 5908 29504 5960 29510
rect 5908 29446 5960 29452
rect 5920 29306 5948 29446
rect 5908 29300 5960 29306
rect 5908 29242 5960 29248
rect 6840 29102 6868 29514
rect 6828 29096 6880 29102
rect 5630 29064 5686 29073
rect 6828 29038 6880 29044
rect 5630 28999 5686 29008
rect 5644 28558 5672 28999
rect 6552 28960 6604 28966
rect 6552 28902 6604 28908
rect 6564 28626 6592 28902
rect 6552 28620 6604 28626
rect 6552 28562 6604 28568
rect 5448 28552 5500 28558
rect 5448 28494 5500 28500
rect 5632 28552 5684 28558
rect 5632 28494 5684 28500
rect 6840 28150 6868 29038
rect 6828 28144 6880 28150
rect 6828 28086 6880 28092
rect 5448 28076 5500 28082
rect 5368 28036 5448 28064
rect 5500 28036 5580 28064
rect 5448 28018 5500 28024
rect 4712 28008 4764 28014
rect 4712 27950 4764 27956
rect 4724 27674 4752 27950
rect 4712 27668 4764 27674
rect 4712 27610 4764 27616
rect 4874 27228 5182 27237
rect 4874 27226 4880 27228
rect 4936 27226 4960 27228
rect 5016 27226 5040 27228
rect 5096 27226 5120 27228
rect 5176 27226 5182 27228
rect 4936 27174 4938 27226
rect 5118 27174 5120 27226
rect 4874 27172 4880 27174
rect 4936 27172 4960 27174
rect 5016 27172 5040 27174
rect 5096 27172 5120 27174
rect 5176 27172 5182 27174
rect 4874 27163 5182 27172
rect 4580 26336 4660 26364
rect 4528 26318 4580 26324
rect 5552 26314 5580 28036
rect 7024 28014 7052 30790
rect 7380 30738 7432 30744
rect 7484 30258 7512 31758
rect 7472 30252 7524 30258
rect 7472 30194 7524 30200
rect 7484 29306 7512 30194
rect 7576 29306 7604 32014
rect 7656 31816 7708 31822
rect 8116 31816 8168 31822
rect 7708 31776 7972 31804
rect 7656 31758 7708 31764
rect 7840 31680 7892 31686
rect 7840 31622 7892 31628
rect 7852 31278 7880 31622
rect 7840 31272 7892 31278
rect 7840 31214 7892 31220
rect 7840 30932 7892 30938
rect 7840 30874 7892 30880
rect 7748 30592 7800 30598
rect 7748 30534 7800 30540
rect 7760 30258 7788 30534
rect 7852 30394 7880 30874
rect 7840 30388 7892 30394
rect 7840 30330 7892 30336
rect 7944 30258 7972 31776
rect 8116 31758 8168 31764
rect 7748 30252 7800 30258
rect 7748 30194 7800 30200
rect 7932 30252 7984 30258
rect 7932 30194 7984 30200
rect 7944 30054 7972 30194
rect 7932 30048 7984 30054
rect 7932 29990 7984 29996
rect 7472 29300 7524 29306
rect 7472 29242 7524 29248
rect 7564 29300 7616 29306
rect 7564 29242 7616 29248
rect 7196 28484 7248 28490
rect 7196 28426 7248 28432
rect 7012 28008 7064 28014
rect 7012 27950 7064 27956
rect 6368 27872 6420 27878
rect 6368 27814 6420 27820
rect 6380 27470 6408 27814
rect 6368 27464 6420 27470
rect 6368 27406 6420 27412
rect 6828 27328 6880 27334
rect 6828 27270 6880 27276
rect 6840 27130 6868 27270
rect 7024 27130 7052 27950
rect 7208 27878 7236 28426
rect 7196 27872 7248 27878
rect 7196 27814 7248 27820
rect 6828 27124 6880 27130
rect 6828 27066 6880 27072
rect 7012 27124 7064 27130
rect 7012 27066 7064 27072
rect 7208 27062 7236 27814
rect 7196 27056 7248 27062
rect 7196 26998 7248 27004
rect 6920 26920 6972 26926
rect 6920 26862 6972 26868
rect 6932 26586 6960 26862
rect 6920 26580 6972 26586
rect 6920 26522 6972 26528
rect 7208 26314 7236 26998
rect 5356 26308 5408 26314
rect 5356 26250 5408 26256
rect 5540 26308 5592 26314
rect 5540 26250 5592 26256
rect 7196 26308 7248 26314
rect 7196 26250 7248 26256
rect 4874 26140 5182 26149
rect 4874 26138 4880 26140
rect 4936 26138 4960 26140
rect 5016 26138 5040 26140
rect 5096 26138 5120 26140
rect 5176 26138 5182 26140
rect 4936 26086 4938 26138
rect 5118 26086 5120 26138
rect 4874 26084 4880 26086
rect 4936 26084 4960 26086
rect 5016 26084 5040 26086
rect 5096 26084 5120 26086
rect 5176 26084 5182 26086
rect 4874 26075 5182 26084
rect 5368 26042 5396 26250
rect 6000 26240 6052 26246
rect 6000 26182 6052 26188
rect 6920 26240 6972 26246
rect 6920 26182 6972 26188
rect 5356 26036 5408 26042
rect 5356 25978 5408 25984
rect 4712 25696 4764 25702
rect 4712 25638 4764 25644
rect 4214 25596 4522 25605
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25531 4522 25540
rect 4344 25288 4396 25294
rect 4344 25230 4396 25236
rect 4356 24954 4384 25230
rect 4620 25152 4672 25158
rect 4620 25094 4672 25100
rect 4344 24948 4396 24954
rect 4344 24890 4396 24896
rect 4214 24508 4522 24517
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24443 4522 24452
rect 4068 24404 4120 24410
rect 4068 24346 4120 24352
rect 3988 24274 4108 24290
rect 3988 24268 4120 24274
rect 3988 24262 4068 24268
rect 4068 24210 4120 24216
rect 4080 23662 4108 24210
rect 4632 24206 4660 25094
rect 4724 24954 4752 25638
rect 4874 25052 5182 25061
rect 4874 25050 4880 25052
rect 4936 25050 4960 25052
rect 5016 25050 5040 25052
rect 5096 25050 5120 25052
rect 5176 25050 5182 25052
rect 4936 24998 4938 25050
rect 5118 24998 5120 25050
rect 4874 24996 4880 24998
rect 4936 24996 4960 24998
rect 5016 24996 5040 24998
rect 5096 24996 5120 24998
rect 5176 24996 5182 24998
rect 4874 24987 5182 24996
rect 4712 24948 4764 24954
rect 4712 24890 4764 24896
rect 5816 24948 5868 24954
rect 5816 24890 5868 24896
rect 4804 24744 4856 24750
rect 4804 24686 4856 24692
rect 4620 24200 4672 24206
rect 4672 24160 4752 24188
rect 4620 24142 4672 24148
rect 4620 24064 4672 24070
rect 4620 24006 4672 24012
rect 4068 23656 4120 23662
rect 4068 23598 4120 23604
rect 2688 23054 2740 23060
rect 2792 23072 3004 23100
rect 3056 23112 3108 23118
rect 2516 22710 2544 23054
rect 2700 22778 2728 23054
rect 2688 22772 2740 22778
rect 2688 22714 2740 22720
rect 2504 22704 2556 22710
rect 2504 22646 2556 22652
rect 2792 21554 2820 23072
rect 3056 23054 3108 23060
rect 3148 23112 3200 23118
rect 3148 23054 3200 23060
rect 3608 23112 3660 23118
rect 3660 23072 3832 23100
rect 3608 23054 3660 23060
rect 2872 22976 2924 22982
rect 2872 22918 2924 22924
rect 2884 22574 2912 22918
rect 2962 22672 3018 22681
rect 2962 22607 2964 22616
rect 3016 22607 3018 22616
rect 2964 22578 3016 22584
rect 2872 22568 2924 22574
rect 2872 22510 2924 22516
rect 2780 21548 2832 21554
rect 2780 21490 2832 21496
rect 2884 20806 2912 22510
rect 3068 22166 3096 23054
rect 3160 22778 3188 23054
rect 3332 23044 3384 23050
rect 3332 22986 3384 22992
rect 3148 22772 3200 22778
rect 3148 22714 3200 22720
rect 3344 22506 3372 22986
rect 3700 22568 3752 22574
rect 3700 22510 3752 22516
rect 3332 22500 3384 22506
rect 3332 22442 3384 22448
rect 3608 22228 3660 22234
rect 3608 22170 3660 22176
rect 3056 22160 3108 22166
rect 3056 22102 3108 22108
rect 3424 22160 3476 22166
rect 3424 22102 3476 22108
rect 3056 21344 3108 21350
rect 3056 21286 3108 21292
rect 2872 20800 2924 20806
rect 2872 20742 2924 20748
rect 3068 20398 3096 21286
rect 3148 20460 3200 20466
rect 3148 20402 3200 20408
rect 2872 20392 2924 20398
rect 2872 20334 2924 20340
rect 3056 20392 3108 20398
rect 3056 20334 3108 20340
rect 2412 20256 2464 20262
rect 2412 20198 2464 20204
rect 2424 20058 2452 20198
rect 2884 20058 2912 20334
rect 2412 20052 2464 20058
rect 2412 19994 2464 20000
rect 2872 20052 2924 20058
rect 2872 19994 2924 20000
rect 3068 19922 3096 20334
rect 2964 19916 3016 19922
rect 2964 19858 3016 19864
rect 3056 19916 3108 19922
rect 3056 19858 3108 19864
rect 2976 19446 3004 19858
rect 2964 19440 3016 19446
rect 2964 19382 3016 19388
rect 2504 18080 2556 18086
rect 2504 18022 2556 18028
rect 2964 18080 3016 18086
rect 2964 18022 3016 18028
rect 2136 17876 2188 17882
rect 2136 17818 2188 17824
rect 1952 17672 2004 17678
rect 1952 17614 2004 17620
rect 2044 17672 2096 17678
rect 2044 17614 2096 17620
rect 1952 17536 2004 17542
rect 1952 17478 2004 17484
rect 1964 16574 1992 17478
rect 1872 16546 1992 16574
rect 2136 16584 2188 16590
rect 1768 16448 1820 16454
rect 1768 16390 1820 16396
rect 1400 16244 1452 16250
rect 1400 16186 1452 16192
rect 1412 16046 1440 16186
rect 1400 16040 1452 16046
rect 1400 15982 1452 15988
rect 938 15736 994 15745
rect 938 15671 940 15680
rect 992 15671 994 15680
rect 940 15642 992 15648
rect 1412 14414 1440 15982
rect 1780 15502 1808 16390
rect 1768 15496 1820 15502
rect 1768 15438 1820 15444
rect 1400 14408 1452 14414
rect 1400 14350 1452 14356
rect 1412 13394 1440 14350
rect 1676 14340 1728 14346
rect 1676 14282 1728 14288
rect 1688 14074 1716 14282
rect 1676 14068 1728 14074
rect 1676 14010 1728 14016
rect 1492 13864 1544 13870
rect 1492 13806 1544 13812
rect 1504 13705 1532 13806
rect 1490 13696 1546 13705
rect 1490 13631 1546 13640
rect 1400 13388 1452 13394
rect 1400 13330 1452 13336
rect 1412 12850 1440 13330
rect 1400 12844 1452 12850
rect 1400 12786 1452 12792
rect 1676 12776 1728 12782
rect 1676 12718 1728 12724
rect 1688 12442 1716 12718
rect 1676 12436 1728 12442
rect 1676 12378 1728 12384
rect 940 11756 992 11762
rect 940 11698 992 11704
rect 952 11665 980 11698
rect 938 11656 994 11665
rect 938 11591 994 11600
rect 1676 11076 1728 11082
rect 1676 11018 1728 11024
rect 1688 10810 1716 11018
rect 1676 10804 1728 10810
rect 1676 10746 1728 10752
rect 938 8936 994 8945
rect 938 8871 940 8880
rect 992 8871 994 8880
rect 940 8842 992 8848
rect 1492 7404 1544 7410
rect 1492 7346 1544 7352
rect 1504 6905 1532 7346
rect 1872 6914 1900 16546
rect 2516 16574 2544 18022
rect 2136 16526 2188 16532
rect 2424 16546 2544 16574
rect 1952 16448 2004 16454
rect 1952 16390 2004 16396
rect 1964 16182 1992 16390
rect 1952 16176 2004 16182
rect 1952 16118 2004 16124
rect 2148 16046 2176 16526
rect 2136 16040 2188 16046
rect 2136 15982 2188 15988
rect 1490 6896 1546 6905
rect 1872 6886 1992 6914
rect 1490 6831 1546 6840
rect 940 4548 992 4554
rect 940 4490 992 4496
rect 952 4185 980 4490
rect 938 4176 994 4185
rect 938 4111 994 4120
rect 1964 3058 1992 6886
rect 2424 3058 2452 16546
rect 2976 16250 3004 18022
rect 3068 17134 3096 19858
rect 3160 19242 3188 20402
rect 3148 19236 3200 19242
rect 3148 19178 3200 19184
rect 3160 18766 3188 19178
rect 3148 18760 3200 18766
rect 3148 18702 3200 18708
rect 3436 18154 3464 22102
rect 3620 21554 3648 22170
rect 3712 21944 3740 22510
rect 3804 22098 3832 23072
rect 3976 22976 4028 22982
rect 3976 22918 4028 22924
rect 3988 22778 4016 22918
rect 3976 22772 4028 22778
rect 3976 22714 4028 22720
rect 4080 22658 4108 23598
rect 4214 23420 4522 23429
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23355 4522 23364
rect 4632 23322 4660 24006
rect 4620 23316 4672 23322
rect 4620 23258 4672 23264
rect 4436 23112 4488 23118
rect 4436 23054 4488 23060
rect 4344 23044 4396 23050
rect 4344 22986 4396 22992
rect 3884 22636 3936 22642
rect 3884 22578 3936 22584
rect 3988 22630 4108 22658
rect 3792 22092 3844 22098
rect 3792 22034 3844 22040
rect 3792 21956 3844 21962
rect 3712 21916 3792 21944
rect 3792 21898 3844 21904
rect 3608 21548 3660 21554
rect 3608 21490 3660 21496
rect 3620 20942 3648 21490
rect 3804 21010 3832 21898
rect 3896 21894 3924 22578
rect 3884 21888 3936 21894
rect 3884 21830 3936 21836
rect 3700 21004 3752 21010
rect 3700 20946 3752 20952
rect 3792 21004 3844 21010
rect 3792 20946 3844 20952
rect 3608 20936 3660 20942
rect 3608 20878 3660 20884
rect 3712 20754 3740 20946
rect 3620 20726 3740 20754
rect 3620 20466 3648 20726
rect 3896 20602 3924 21830
rect 3988 21486 4016 22630
rect 4356 22438 4384 22986
rect 4448 22778 4476 23054
rect 4528 23044 4580 23050
rect 4528 22986 4580 22992
rect 4620 23044 4672 23050
rect 4620 22986 4672 22992
rect 4436 22772 4488 22778
rect 4436 22714 4488 22720
rect 4540 22710 4568 22986
rect 4528 22704 4580 22710
rect 4528 22646 4580 22652
rect 4632 22506 4660 22986
rect 4724 22642 4752 24160
rect 4816 23322 4844 24686
rect 5632 24608 5684 24614
rect 5632 24550 5684 24556
rect 5644 24274 5672 24550
rect 5632 24268 5684 24274
rect 5632 24210 5684 24216
rect 4874 23964 5182 23973
rect 4874 23962 4880 23964
rect 4936 23962 4960 23964
rect 5016 23962 5040 23964
rect 5096 23962 5120 23964
rect 5176 23962 5182 23964
rect 4936 23910 4938 23962
rect 5118 23910 5120 23962
rect 4874 23908 4880 23910
rect 4936 23908 4960 23910
rect 5016 23908 5040 23910
rect 5096 23908 5120 23910
rect 5176 23908 5182 23910
rect 4874 23899 5182 23908
rect 5632 23724 5684 23730
rect 5632 23666 5684 23672
rect 5264 23520 5316 23526
rect 5264 23462 5316 23468
rect 4804 23316 4856 23322
rect 4804 23258 4856 23264
rect 4896 23112 4948 23118
rect 4894 23080 4896 23089
rect 4948 23080 4950 23089
rect 5276 23050 5304 23462
rect 5644 23322 5672 23666
rect 5632 23316 5684 23322
rect 5632 23258 5684 23264
rect 5356 23112 5408 23118
rect 5356 23054 5408 23060
rect 4894 23015 4950 23024
rect 5264 23044 5316 23050
rect 5264 22986 5316 22992
rect 4874 22876 5182 22885
rect 4874 22874 4880 22876
rect 4936 22874 4960 22876
rect 5016 22874 5040 22876
rect 5096 22874 5120 22876
rect 5176 22874 5182 22876
rect 4936 22822 4938 22874
rect 5118 22822 5120 22874
rect 4874 22820 4880 22822
rect 4936 22820 4960 22822
rect 5016 22820 5040 22822
rect 5096 22820 5120 22822
rect 5176 22820 5182 22822
rect 4874 22811 5182 22820
rect 4804 22704 4856 22710
rect 4804 22646 4856 22652
rect 4712 22636 4764 22642
rect 4712 22578 4764 22584
rect 4620 22500 4672 22506
rect 4620 22442 4672 22448
rect 4344 22432 4396 22438
rect 4344 22374 4396 22380
rect 4214 22332 4522 22341
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22267 4522 22276
rect 4344 21888 4396 21894
rect 4344 21830 4396 21836
rect 4356 21690 4384 21830
rect 4344 21684 4396 21690
rect 4344 21626 4396 21632
rect 4632 21570 4660 22442
rect 4712 22432 4764 22438
rect 4712 22374 4764 22380
rect 4724 21690 4752 22374
rect 4712 21684 4764 21690
rect 4712 21626 4764 21632
rect 4540 21542 4660 21570
rect 4540 21486 4568 21542
rect 3976 21480 4028 21486
rect 3976 21422 4028 21428
rect 4528 21480 4580 21486
rect 4528 21422 4580 21428
rect 4620 21412 4672 21418
rect 4620 21354 4672 21360
rect 4214 21244 4522 21253
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21179 4522 21188
rect 4632 21146 4660 21354
rect 4620 21140 4672 21146
rect 4620 21082 4672 21088
rect 3976 20936 4028 20942
rect 3976 20878 4028 20884
rect 3884 20596 3936 20602
rect 3884 20538 3936 20544
rect 3988 20466 4016 20878
rect 4068 20800 4120 20806
rect 4068 20742 4120 20748
rect 3608 20460 3660 20466
rect 3608 20402 3660 20408
rect 3976 20460 4028 20466
rect 3976 20402 4028 20408
rect 3516 19508 3568 19514
rect 3516 19450 3568 19456
rect 3528 19174 3556 19450
rect 3620 19378 3648 20402
rect 3792 20324 3844 20330
rect 3792 20266 3844 20272
rect 3804 19922 3832 20266
rect 3976 20256 4028 20262
rect 3976 20198 4028 20204
rect 3792 19916 3844 19922
rect 3792 19858 3844 19864
rect 3884 19848 3936 19854
rect 3884 19790 3936 19796
rect 3608 19372 3660 19378
rect 3608 19314 3660 19320
rect 3516 19168 3568 19174
rect 3516 19110 3568 19116
rect 3424 18148 3476 18154
rect 3424 18090 3476 18096
rect 3528 18086 3556 19110
rect 3516 18080 3568 18086
rect 3516 18022 3568 18028
rect 3528 17746 3556 18022
rect 3516 17740 3568 17746
rect 3516 17682 3568 17688
rect 3424 17672 3476 17678
rect 3424 17614 3476 17620
rect 3436 17338 3464 17614
rect 3424 17332 3476 17338
rect 3424 17274 3476 17280
rect 3240 17196 3292 17202
rect 3240 17138 3292 17144
rect 3056 17128 3108 17134
rect 3056 17070 3108 17076
rect 3068 16658 3096 17070
rect 3056 16652 3108 16658
rect 3056 16594 3108 16600
rect 2964 16244 3016 16250
rect 2964 16186 3016 16192
rect 3068 14940 3096 16594
rect 3148 16448 3200 16454
rect 3148 16390 3200 16396
rect 3160 15910 3188 16390
rect 3148 15904 3200 15910
rect 3148 15846 3200 15852
rect 3252 15026 3280 17138
rect 3620 16794 3648 19314
rect 3896 19310 3924 19790
rect 3988 19718 4016 20198
rect 3976 19712 4028 19718
rect 3976 19654 4028 19660
rect 3884 19304 3936 19310
rect 3884 19246 3936 19252
rect 4080 18834 4108 20742
rect 4214 20156 4522 20165
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20091 4522 20100
rect 4620 19780 4672 19786
rect 4724 19768 4752 21626
rect 4816 19922 4844 22646
rect 5264 22636 5316 22642
rect 5264 22578 5316 22584
rect 4874 21788 5182 21797
rect 4874 21786 4880 21788
rect 4936 21786 4960 21788
rect 5016 21786 5040 21788
rect 5096 21786 5120 21788
rect 5176 21786 5182 21788
rect 4936 21734 4938 21786
rect 5118 21734 5120 21786
rect 4874 21732 4880 21734
rect 4936 21732 4960 21734
rect 5016 21732 5040 21734
rect 5096 21732 5120 21734
rect 5176 21732 5182 21734
rect 4874 21723 5182 21732
rect 5172 21616 5224 21622
rect 5276 21570 5304 22578
rect 5368 22574 5396 23054
rect 5644 22778 5672 23258
rect 5828 23254 5856 24890
rect 5908 24812 5960 24818
rect 5908 24754 5960 24760
rect 5920 23866 5948 24754
rect 6012 24138 6040 26182
rect 6932 26042 6960 26182
rect 6920 26036 6972 26042
rect 6920 25978 6972 25984
rect 7288 25152 7340 25158
rect 7288 25094 7340 25100
rect 7300 24750 7328 25094
rect 7288 24744 7340 24750
rect 7288 24686 7340 24692
rect 7288 24608 7340 24614
rect 7288 24550 7340 24556
rect 6644 24336 6696 24342
rect 6644 24278 6696 24284
rect 6000 24132 6052 24138
rect 6000 24074 6052 24080
rect 5908 23860 5960 23866
rect 5908 23802 5960 23808
rect 6012 23594 6040 24074
rect 6656 23730 6684 24278
rect 6644 23724 6696 23730
rect 6644 23666 6696 23672
rect 7012 23724 7064 23730
rect 7012 23666 7064 23672
rect 6000 23588 6052 23594
rect 6000 23530 6052 23536
rect 6460 23316 6512 23322
rect 6460 23258 6512 23264
rect 5816 23248 5868 23254
rect 5816 23190 5868 23196
rect 5816 23112 5868 23118
rect 5816 23054 5868 23060
rect 5724 22976 5776 22982
rect 5724 22918 5776 22924
rect 5632 22772 5684 22778
rect 5632 22714 5684 22720
rect 5356 22568 5408 22574
rect 5356 22510 5408 22516
rect 5224 21564 5304 21570
rect 5172 21558 5304 21564
rect 4896 21548 4948 21554
rect 5184 21542 5304 21558
rect 4896 21490 4948 21496
rect 4908 21010 4936 21490
rect 5264 21480 5316 21486
rect 5264 21422 5316 21428
rect 4896 21004 4948 21010
rect 4896 20946 4948 20952
rect 5276 20874 5304 21422
rect 5368 21350 5396 22510
rect 5736 22030 5764 22918
rect 5828 22438 5856 23054
rect 6472 22642 6500 23258
rect 6656 23186 6684 23666
rect 7024 23322 7052 23666
rect 7300 23594 7328 24550
rect 7288 23588 7340 23594
rect 7288 23530 7340 23536
rect 7012 23316 7064 23322
rect 7012 23258 7064 23264
rect 6644 23180 6696 23186
rect 6644 23122 6696 23128
rect 6460 22636 6512 22642
rect 6460 22578 6512 22584
rect 5816 22432 5868 22438
rect 5816 22374 5868 22380
rect 6184 22160 6236 22166
rect 6184 22102 6236 22108
rect 5724 22024 5776 22030
rect 5724 21966 5776 21972
rect 5816 22024 5868 22030
rect 5816 21966 5868 21972
rect 5828 21554 5856 21966
rect 6196 21962 6224 22102
rect 6276 22092 6328 22098
rect 6276 22034 6328 22040
rect 6184 21956 6236 21962
rect 6184 21898 6236 21904
rect 6196 21554 6224 21898
rect 5724 21548 5776 21554
rect 5724 21490 5776 21496
rect 5816 21548 5868 21554
rect 5816 21490 5868 21496
rect 6184 21548 6236 21554
rect 6184 21490 6236 21496
rect 5356 21344 5408 21350
rect 5356 21286 5408 21292
rect 5448 21344 5500 21350
rect 5448 21286 5500 21292
rect 5264 20868 5316 20874
rect 5264 20810 5316 20816
rect 4874 20700 5182 20709
rect 4874 20698 4880 20700
rect 4936 20698 4960 20700
rect 5016 20698 5040 20700
rect 5096 20698 5120 20700
rect 5176 20698 5182 20700
rect 4936 20646 4938 20698
rect 5118 20646 5120 20698
rect 4874 20644 4880 20646
rect 4936 20644 4960 20646
rect 5016 20644 5040 20646
rect 5096 20644 5120 20646
rect 5176 20644 5182 20646
rect 4874 20635 5182 20644
rect 5080 20256 5132 20262
rect 5080 20198 5132 20204
rect 5092 19990 5120 20198
rect 5080 19984 5132 19990
rect 5080 19926 5132 19932
rect 4804 19916 4856 19922
rect 4804 19858 4856 19864
rect 5368 19825 5396 21286
rect 4672 19740 4752 19768
rect 4986 19816 5042 19825
rect 4986 19751 5042 19760
rect 5354 19816 5410 19825
rect 5354 19751 5410 19760
rect 4620 19722 4672 19728
rect 4214 19068 4522 19077
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 19003 4522 19012
rect 4068 18828 4120 18834
rect 4068 18770 4120 18776
rect 4080 18222 4108 18770
rect 4252 18624 4304 18630
rect 4252 18566 4304 18572
rect 4264 18426 4292 18566
rect 4252 18420 4304 18426
rect 4252 18362 4304 18368
rect 4068 18216 4120 18222
rect 4068 18158 4120 18164
rect 3700 18148 3752 18154
rect 3700 18090 3752 18096
rect 3712 17678 3740 18090
rect 3700 17672 3752 17678
rect 3700 17614 3752 17620
rect 3608 16788 3660 16794
rect 3608 16730 3660 16736
rect 3620 16250 3648 16730
rect 3608 16244 3660 16250
rect 3608 16186 3660 16192
rect 3240 15020 3292 15026
rect 3240 14962 3292 14968
rect 3148 14952 3200 14958
rect 3068 14912 3148 14940
rect 3148 14894 3200 14900
rect 2504 14816 2556 14822
rect 2504 14758 2556 14764
rect 2516 14074 2544 14758
rect 2780 14408 2832 14414
rect 2780 14350 2832 14356
rect 2504 14068 2556 14074
rect 2504 14010 2556 14016
rect 2792 13190 2820 14350
rect 2964 13320 3016 13326
rect 2964 13262 3016 13268
rect 2780 13184 2832 13190
rect 2780 13126 2832 13132
rect 2792 12850 2820 13126
rect 2780 12844 2832 12850
rect 2780 12786 2832 12792
rect 2792 11506 2820 12786
rect 2976 11642 3004 13262
rect 3056 12640 3108 12646
rect 3056 12582 3108 12588
rect 3068 12306 3096 12582
rect 3160 12434 3188 14894
rect 3252 14618 3280 14962
rect 3608 14816 3660 14822
rect 3608 14758 3660 14764
rect 3620 14618 3648 14758
rect 3240 14612 3292 14618
rect 3240 14554 3292 14560
rect 3608 14612 3660 14618
rect 3608 14554 3660 14560
rect 3712 14482 3740 17614
rect 3792 17196 3844 17202
rect 3792 17138 3844 17144
rect 3804 16998 3832 17138
rect 4080 16998 4108 18158
rect 4214 17980 4522 17989
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17915 4522 17924
rect 4252 17604 4304 17610
rect 4252 17546 4304 17552
rect 4264 17338 4292 17546
rect 4252 17332 4304 17338
rect 4252 17274 4304 17280
rect 3792 16992 3844 16998
rect 3792 16934 3844 16940
rect 4068 16992 4120 16998
rect 4068 16934 4120 16940
rect 3700 14476 3752 14482
rect 3700 14418 3752 14424
rect 3160 12406 3280 12434
rect 3252 12306 3280 12406
rect 3056 12300 3108 12306
rect 3056 12242 3108 12248
rect 3240 12300 3292 12306
rect 3240 12242 3292 12248
rect 3148 12164 3200 12170
rect 3148 12106 3200 12112
rect 2976 11614 3096 11642
rect 2792 11478 3004 11506
rect 2976 11082 3004 11478
rect 2964 11076 3016 11082
rect 2964 11018 3016 11024
rect 3068 9994 3096 11614
rect 3160 11354 3188 12106
rect 3148 11348 3200 11354
rect 3148 11290 3200 11296
rect 3160 10674 3188 11290
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 3160 10062 3188 10610
rect 3252 10470 3280 12242
rect 3424 12096 3476 12102
rect 3424 12038 3476 12044
rect 3436 11354 3464 12038
rect 3424 11348 3476 11354
rect 3424 11290 3476 11296
rect 3436 10606 3464 11290
rect 3424 10600 3476 10606
rect 3424 10542 3476 10548
rect 3240 10464 3292 10470
rect 3240 10406 3292 10412
rect 3148 10056 3200 10062
rect 3148 9998 3200 10004
rect 3056 9988 3108 9994
rect 3056 9930 3108 9936
rect 2964 9376 3016 9382
rect 2964 9318 3016 9324
rect 2976 9178 3004 9318
rect 2964 9172 3016 9178
rect 2964 9114 3016 9120
rect 3068 8974 3096 9930
rect 3148 9920 3200 9926
rect 3148 9862 3200 9868
rect 3160 9722 3188 9862
rect 3148 9716 3200 9722
rect 3148 9658 3200 9664
rect 3238 9616 3294 9625
rect 3712 9586 3740 14418
rect 3804 13326 3832 16934
rect 4214 16892 4522 16901
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16827 4522 16836
rect 4434 16688 4490 16697
rect 4434 16623 4436 16632
rect 4488 16623 4490 16632
rect 4436 16594 4488 16600
rect 3976 16584 4028 16590
rect 4160 16584 4212 16590
rect 3976 16526 4028 16532
rect 4080 16544 4160 16572
rect 3884 15904 3936 15910
rect 3884 15846 3936 15852
rect 3896 15502 3924 15846
rect 3988 15706 4016 16526
rect 3976 15700 4028 15706
rect 3976 15642 4028 15648
rect 4080 15586 4108 16544
rect 4160 16526 4212 16532
rect 4252 16516 4304 16522
rect 4632 16504 4660 19722
rect 5000 19718 5028 19751
rect 4988 19712 5040 19718
rect 4988 19654 5040 19660
rect 5264 19712 5316 19718
rect 5264 19654 5316 19660
rect 4874 19612 5182 19621
rect 4874 19610 4880 19612
rect 4936 19610 4960 19612
rect 5016 19610 5040 19612
rect 5096 19610 5120 19612
rect 5176 19610 5182 19612
rect 4936 19558 4938 19610
rect 5118 19558 5120 19610
rect 4874 19556 4880 19558
rect 4936 19556 4960 19558
rect 5016 19556 5040 19558
rect 5096 19556 5120 19558
rect 5176 19556 5182 19558
rect 4874 19547 5182 19556
rect 4712 19440 4764 19446
rect 4712 19382 4764 19388
rect 4896 19440 4948 19446
rect 4896 19382 4948 19388
rect 4724 17610 4752 19382
rect 4908 19310 4936 19382
rect 4804 19304 4856 19310
rect 4804 19246 4856 19252
rect 4896 19304 4948 19310
rect 4896 19246 4948 19252
rect 4816 18970 4844 19246
rect 4804 18964 4856 18970
rect 4804 18906 4856 18912
rect 5276 18766 5304 19654
rect 5264 18760 5316 18766
rect 5264 18702 5316 18708
rect 4874 18524 5182 18533
rect 4874 18522 4880 18524
rect 4936 18522 4960 18524
rect 5016 18522 5040 18524
rect 5096 18522 5120 18524
rect 5176 18522 5182 18524
rect 4936 18470 4938 18522
rect 5118 18470 5120 18522
rect 4874 18468 4880 18470
rect 4936 18468 4960 18470
rect 5016 18468 5040 18470
rect 5096 18468 5120 18470
rect 5176 18468 5182 18470
rect 4874 18459 5182 18468
rect 4712 17604 4764 17610
rect 4712 17546 4764 17552
rect 4304 16476 4660 16504
rect 4252 16458 4304 16464
rect 4620 16244 4672 16250
rect 4620 16186 4672 16192
rect 4214 15804 4522 15813
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15739 4522 15748
rect 4632 15638 4660 16186
rect 4724 16114 4752 17546
rect 4874 17436 5182 17445
rect 4874 17434 4880 17436
rect 4936 17434 4960 17436
rect 5016 17434 5040 17436
rect 5096 17434 5120 17436
rect 5176 17434 5182 17436
rect 4936 17382 4938 17434
rect 5118 17382 5120 17434
rect 4874 17380 4880 17382
rect 4936 17380 4960 17382
rect 5016 17380 5040 17382
rect 5096 17380 5120 17382
rect 5176 17380 5182 17382
rect 4874 17371 5182 17380
rect 4804 17264 4856 17270
rect 4804 17206 4856 17212
rect 4816 16182 4844 17206
rect 5264 17196 5316 17202
rect 5264 17138 5316 17144
rect 4874 16348 5182 16357
rect 4874 16346 4880 16348
rect 4936 16346 4960 16348
rect 5016 16346 5040 16348
rect 5096 16346 5120 16348
rect 5176 16346 5182 16348
rect 4936 16294 4938 16346
rect 5118 16294 5120 16346
rect 4874 16292 4880 16294
rect 4936 16292 4960 16294
rect 5016 16292 5040 16294
rect 5096 16292 5120 16294
rect 5176 16292 5182 16294
rect 4874 16283 5182 16292
rect 5276 16250 5304 17138
rect 5264 16244 5316 16250
rect 5264 16186 5316 16192
rect 4804 16176 4856 16182
rect 4804 16118 4856 16124
rect 4712 16108 4764 16114
rect 4712 16050 4764 16056
rect 4724 15706 4752 16050
rect 4712 15700 4764 15706
rect 4712 15642 4764 15648
rect 4620 15632 4672 15638
rect 4080 15558 4292 15586
rect 4620 15574 4672 15580
rect 3884 15496 3936 15502
rect 3884 15438 3936 15444
rect 3976 15496 4028 15502
rect 3976 15438 4028 15444
rect 4160 15496 4212 15502
rect 4160 15438 4212 15444
rect 3988 15026 4016 15438
rect 4172 15094 4200 15438
rect 4160 15088 4212 15094
rect 4160 15030 4212 15036
rect 3976 15020 4028 15026
rect 3976 14962 4028 14968
rect 4264 14958 4292 15558
rect 4632 15094 4660 15574
rect 4816 15502 4844 16118
rect 4804 15496 4856 15502
rect 4804 15438 4856 15444
rect 5356 15360 5408 15366
rect 5356 15302 5408 15308
rect 4874 15260 5182 15269
rect 4874 15258 4880 15260
rect 4936 15258 4960 15260
rect 5016 15258 5040 15260
rect 5096 15258 5120 15260
rect 5176 15258 5182 15260
rect 4936 15206 4938 15258
rect 5118 15206 5120 15258
rect 4874 15204 4880 15206
rect 4936 15204 4960 15206
rect 5016 15204 5040 15206
rect 5096 15204 5120 15206
rect 5176 15204 5182 15206
rect 4874 15195 5182 15204
rect 5368 15162 5396 15302
rect 5356 15156 5408 15162
rect 5356 15098 5408 15104
rect 4620 15088 4672 15094
rect 4620 15030 4672 15036
rect 4252 14952 4304 14958
rect 4252 14894 4304 14900
rect 4068 14884 4120 14890
rect 4068 14826 4120 14832
rect 3884 14816 3936 14822
rect 3884 14758 3936 14764
rect 3792 13320 3844 13326
rect 3792 13262 3844 13268
rect 3896 12782 3924 14758
rect 4080 14618 4108 14826
rect 4214 14716 4522 14725
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14651 4522 14660
rect 4068 14612 4120 14618
rect 4068 14554 4120 14560
rect 4632 14414 4660 15030
rect 4712 15020 4764 15026
rect 4712 14962 4764 14968
rect 4620 14408 4672 14414
rect 4620 14350 4672 14356
rect 4214 13628 4522 13637
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13563 4522 13572
rect 3976 13252 4028 13258
rect 3976 13194 4028 13200
rect 4620 13252 4672 13258
rect 4620 13194 4672 13200
rect 3988 13002 4016 13194
rect 3988 12986 4108 13002
rect 4632 12986 4660 13194
rect 3976 12980 4108 12986
rect 4028 12974 4108 12980
rect 3976 12922 4028 12928
rect 3976 12844 4028 12850
rect 3976 12786 4028 12792
rect 3884 12776 3936 12782
rect 3884 12718 3936 12724
rect 3792 12708 3844 12714
rect 3792 12650 3844 12656
rect 3804 12442 3832 12650
rect 3792 12436 3844 12442
rect 3792 12378 3844 12384
rect 3896 11286 3924 12718
rect 3988 12322 4016 12786
rect 4080 12442 4108 12974
rect 4620 12980 4672 12986
rect 4620 12922 4672 12928
rect 4724 12850 4752 14962
rect 4874 14172 5182 14181
rect 4874 14170 4880 14172
rect 4936 14170 4960 14172
rect 5016 14170 5040 14172
rect 5096 14170 5120 14172
rect 5176 14170 5182 14172
rect 4936 14118 4938 14170
rect 5118 14118 5120 14170
rect 4874 14116 4880 14118
rect 4936 14116 4960 14118
rect 5016 14116 5040 14118
rect 5096 14116 5120 14118
rect 5176 14116 5182 14118
rect 4874 14107 5182 14116
rect 4874 13084 5182 13093
rect 4874 13082 4880 13084
rect 4936 13082 4960 13084
rect 5016 13082 5040 13084
rect 5096 13082 5120 13084
rect 5176 13082 5182 13084
rect 4936 13030 4938 13082
rect 5118 13030 5120 13082
rect 4874 13028 4880 13030
rect 4936 13028 4960 13030
rect 5016 13028 5040 13030
rect 5096 13028 5120 13030
rect 5176 13028 5182 13030
rect 4874 13019 5182 13028
rect 4436 12844 4488 12850
rect 4712 12844 4764 12850
rect 4488 12804 4660 12832
rect 4436 12786 4488 12792
rect 4214 12540 4522 12549
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12475 4522 12484
rect 4632 12442 4660 12804
rect 4712 12786 4764 12792
rect 4068 12436 4120 12442
rect 4068 12378 4120 12384
rect 4620 12436 4672 12442
rect 5460 12434 5488 21286
rect 5736 21185 5764 21490
rect 5722 21176 5778 21185
rect 5722 21111 5778 21120
rect 5630 20904 5686 20913
rect 5630 20839 5632 20848
rect 5684 20839 5686 20848
rect 5632 20810 5684 20816
rect 5828 18698 5856 21490
rect 5908 19848 5960 19854
rect 5908 19790 5960 19796
rect 5920 19514 5948 19790
rect 5908 19508 5960 19514
rect 5908 19450 5960 19456
rect 5920 18834 5948 19450
rect 5998 18864 6054 18873
rect 5908 18828 5960 18834
rect 5998 18799 6054 18808
rect 5908 18770 5960 18776
rect 6012 18766 6040 18799
rect 6000 18760 6052 18766
rect 6000 18702 6052 18708
rect 5632 18692 5684 18698
rect 5632 18634 5684 18640
rect 5816 18692 5868 18698
rect 5816 18634 5868 18640
rect 5644 17882 5672 18634
rect 5908 18216 5960 18222
rect 5908 18158 5960 18164
rect 5632 17876 5684 17882
rect 5632 17818 5684 17824
rect 5724 17536 5776 17542
rect 5724 17478 5776 17484
rect 5736 17338 5764 17478
rect 5724 17332 5776 17338
rect 5724 17274 5776 17280
rect 5920 16522 5948 18158
rect 6184 18080 6236 18086
rect 6184 18022 6236 18028
rect 6196 17542 6224 18022
rect 6184 17536 6236 17542
rect 6184 17478 6236 17484
rect 6092 16992 6144 16998
rect 6092 16934 6144 16940
rect 6104 16794 6132 16934
rect 6092 16788 6144 16794
rect 6092 16730 6144 16736
rect 6196 16658 6224 17478
rect 6184 16652 6236 16658
rect 6184 16594 6236 16600
rect 5908 16516 5960 16522
rect 5908 16458 5960 16464
rect 5920 16046 5948 16458
rect 5632 16040 5684 16046
rect 5632 15982 5684 15988
rect 5908 16040 5960 16046
rect 5908 15982 5960 15988
rect 5644 15706 5672 15982
rect 5632 15700 5684 15706
rect 5632 15642 5684 15648
rect 6196 15570 6224 16594
rect 6184 15564 6236 15570
rect 6184 15506 6236 15512
rect 5632 14408 5684 14414
rect 5632 14350 5684 14356
rect 5644 13394 5672 14350
rect 5908 14340 5960 14346
rect 5908 14282 5960 14288
rect 5920 14074 5948 14282
rect 5908 14068 5960 14074
rect 5908 14010 5960 14016
rect 6000 13864 6052 13870
rect 6000 13806 6052 13812
rect 5632 13388 5684 13394
rect 5632 13330 5684 13336
rect 5816 12844 5868 12850
rect 5816 12786 5868 12792
rect 5828 12442 5856 12786
rect 4620 12378 4672 12384
rect 5368 12406 5488 12434
rect 5816 12436 5868 12442
rect 3988 12306 4108 12322
rect 3988 12300 4120 12306
rect 3988 12294 4068 12300
rect 4068 12242 4120 12248
rect 4874 11996 5182 12005
rect 4874 11994 4880 11996
rect 4936 11994 4960 11996
rect 5016 11994 5040 11996
rect 5096 11994 5120 11996
rect 5176 11994 5182 11996
rect 4936 11942 4938 11994
rect 5118 11942 5120 11994
rect 4874 11940 4880 11942
rect 4936 11940 4960 11942
rect 5016 11940 5040 11942
rect 5096 11940 5120 11942
rect 5176 11940 5182 11942
rect 4874 11931 5182 11940
rect 4214 11452 4522 11461
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11387 4522 11396
rect 3884 11280 3936 11286
rect 3884 11222 3936 11228
rect 4068 11212 4120 11218
rect 4068 11154 4120 11160
rect 3884 11076 3936 11082
rect 3884 11018 3936 11024
rect 3792 11008 3844 11014
rect 3792 10950 3844 10956
rect 3804 10810 3832 10950
rect 3896 10810 3924 11018
rect 3792 10804 3844 10810
rect 3792 10746 3844 10752
rect 3884 10804 3936 10810
rect 3884 10746 3936 10752
rect 4080 10606 4108 11154
rect 4252 11008 4304 11014
rect 4252 10950 4304 10956
rect 4264 10742 4292 10950
rect 4874 10908 5182 10917
rect 4874 10906 4880 10908
rect 4936 10906 4960 10908
rect 5016 10906 5040 10908
rect 5096 10906 5120 10908
rect 5176 10906 5182 10908
rect 4936 10854 4938 10906
rect 5118 10854 5120 10906
rect 4874 10852 4880 10854
rect 4936 10852 4960 10854
rect 5016 10852 5040 10854
rect 5096 10852 5120 10854
rect 5176 10852 5182 10854
rect 4874 10843 5182 10852
rect 4252 10736 4304 10742
rect 4252 10678 4304 10684
rect 4068 10600 4120 10606
rect 4068 10542 4120 10548
rect 4712 10600 4764 10606
rect 4712 10542 4764 10548
rect 3238 9551 3240 9560
rect 3292 9551 3294 9560
rect 3332 9580 3384 9586
rect 3240 9522 3292 9528
rect 3332 9522 3384 9528
rect 3700 9580 3752 9586
rect 3700 9522 3752 9528
rect 3344 9110 3372 9522
rect 3332 9104 3384 9110
rect 3332 9046 3384 9052
rect 3056 8968 3108 8974
rect 3056 8910 3108 8916
rect 3884 8832 3936 8838
rect 3884 8774 3936 8780
rect 2964 8288 3016 8294
rect 2964 8230 3016 8236
rect 2976 7478 3004 8230
rect 2964 7472 3016 7478
rect 2964 7414 3016 7420
rect 3896 4622 3924 8774
rect 4080 8362 4108 10542
rect 4214 10364 4522 10373
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10299 4522 10308
rect 4724 10266 4752 10542
rect 4712 10260 4764 10266
rect 4712 10202 4764 10208
rect 4874 9820 5182 9829
rect 4874 9818 4880 9820
rect 4936 9818 4960 9820
rect 5016 9818 5040 9820
rect 5096 9818 5120 9820
rect 5176 9818 5182 9820
rect 4936 9766 4938 9818
rect 5118 9766 5120 9818
rect 4874 9764 4880 9766
rect 4936 9764 4960 9766
rect 5016 9764 5040 9766
rect 5096 9764 5120 9766
rect 5176 9764 5182 9766
rect 4874 9755 5182 9764
rect 4620 9580 4672 9586
rect 4620 9522 4672 9528
rect 4214 9276 4522 9285
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9211 4522 9220
rect 4158 9072 4214 9081
rect 4158 9007 4214 9016
rect 4172 8974 4200 9007
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 4528 8968 4580 8974
rect 4632 8956 4660 9522
rect 4580 8928 4660 8956
rect 4528 8910 4580 8916
rect 4712 8900 4764 8906
rect 4712 8842 4764 8848
rect 4724 8498 4752 8842
rect 4874 8732 5182 8741
rect 4874 8730 4880 8732
rect 4936 8730 4960 8732
rect 5016 8730 5040 8732
rect 5096 8730 5120 8732
rect 5176 8730 5182 8732
rect 4936 8678 4938 8730
rect 5118 8678 5120 8730
rect 4874 8676 4880 8678
rect 4936 8676 4960 8678
rect 5016 8676 5040 8678
rect 5096 8676 5120 8678
rect 5176 8676 5182 8678
rect 4874 8667 5182 8676
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 4068 8356 4120 8362
rect 4068 8298 4120 8304
rect 4620 8288 4672 8294
rect 4620 8230 4672 8236
rect 4214 8188 4522 8197
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8123 4522 8132
rect 4632 7546 4660 8230
rect 4620 7540 4672 7546
rect 4620 7482 4672 7488
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 3988 7002 4016 7346
rect 4214 7100 4522 7109
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7035 4522 7044
rect 3976 6996 4028 7002
rect 3976 6938 4028 6944
rect 4632 6866 4660 7482
rect 4724 7342 4752 8434
rect 4874 7644 5182 7653
rect 4874 7642 4880 7644
rect 4936 7642 4960 7644
rect 5016 7642 5040 7644
rect 5096 7642 5120 7644
rect 5176 7642 5182 7644
rect 4936 7590 4938 7642
rect 5118 7590 5120 7642
rect 4874 7588 4880 7590
rect 4936 7588 4960 7590
rect 5016 7588 5040 7590
rect 5096 7588 5120 7590
rect 5176 7588 5182 7590
rect 4874 7579 5182 7588
rect 4712 7336 4764 7342
rect 4712 7278 4764 7284
rect 4804 7200 4856 7206
rect 4804 7142 4856 7148
rect 4620 6860 4672 6866
rect 4620 6802 4672 6808
rect 4528 6724 4580 6730
rect 4528 6666 4580 6672
rect 4540 6458 4568 6666
rect 4528 6452 4580 6458
rect 4528 6394 4580 6400
rect 4214 6012 4522 6021
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5947 4522 5956
rect 4632 5778 4660 6802
rect 4816 6458 4844 7142
rect 4874 6556 5182 6565
rect 4874 6554 4880 6556
rect 4936 6554 4960 6556
rect 5016 6554 5040 6556
rect 5096 6554 5120 6556
rect 5176 6554 5182 6556
rect 4936 6502 4938 6554
rect 5118 6502 5120 6554
rect 4874 6500 4880 6502
rect 4936 6500 4960 6502
rect 5016 6500 5040 6502
rect 5096 6500 5120 6502
rect 5176 6500 5182 6502
rect 4874 6491 5182 6500
rect 4804 6452 4856 6458
rect 4804 6394 4856 6400
rect 4620 5772 4672 5778
rect 4620 5714 4672 5720
rect 4874 5468 5182 5477
rect 4874 5466 4880 5468
rect 4936 5466 4960 5468
rect 5016 5466 5040 5468
rect 5096 5466 5120 5468
rect 5176 5466 5182 5468
rect 4936 5414 4938 5466
rect 5118 5414 5120 5466
rect 4874 5412 4880 5414
rect 4936 5412 4960 5414
rect 5016 5412 5040 5414
rect 5096 5412 5120 5414
rect 5176 5412 5182 5414
rect 4874 5403 5182 5412
rect 4214 4924 4522 4933
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4859 4522 4868
rect 3884 4616 3936 4622
rect 3884 4558 3936 4564
rect 4874 4380 5182 4389
rect 4874 4378 4880 4380
rect 4936 4378 4960 4380
rect 5016 4378 5040 4380
rect 5096 4378 5120 4380
rect 5176 4378 5182 4380
rect 4936 4326 4938 4378
rect 5118 4326 5120 4378
rect 4874 4324 4880 4326
rect 4936 4324 4960 4326
rect 5016 4324 5040 4326
rect 5096 4324 5120 4326
rect 5176 4324 5182 4326
rect 4874 4315 5182 4324
rect 4214 3836 4522 3845
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3771 4522 3780
rect 4874 3292 5182 3301
rect 4874 3290 4880 3292
rect 4936 3290 4960 3292
rect 5016 3290 5040 3292
rect 5096 3290 5120 3292
rect 5176 3290 5182 3292
rect 4936 3238 4938 3290
rect 5118 3238 5120 3290
rect 4874 3236 4880 3238
rect 4936 3236 4960 3238
rect 5016 3236 5040 3238
rect 5096 3236 5120 3238
rect 5176 3236 5182 3238
rect 4874 3227 5182 3236
rect 1952 3052 2004 3058
rect 1952 2994 2004 3000
rect 2412 3052 2464 3058
rect 2412 2994 2464 3000
rect 1768 2848 1820 2854
rect 1768 2790 1820 2796
rect 2228 2848 2280 2854
rect 2228 2790 2280 2796
rect 1780 2446 1808 2790
rect 2240 2446 2268 2790
rect 5368 2774 5396 12406
rect 5816 12378 5868 12384
rect 5448 11552 5500 11558
rect 5448 11494 5500 11500
rect 5460 7410 5488 11494
rect 5724 11348 5776 11354
rect 5724 11290 5776 11296
rect 5540 11212 5592 11218
rect 5540 11154 5592 11160
rect 5552 10606 5580 11154
rect 5736 10674 5764 11290
rect 5908 11144 5960 11150
rect 5908 11086 5960 11092
rect 5816 11076 5868 11082
rect 5816 11018 5868 11024
rect 5724 10668 5776 10674
rect 5724 10610 5776 10616
rect 5828 10606 5856 11018
rect 5540 10600 5592 10606
rect 5540 10542 5592 10548
rect 5816 10600 5868 10606
rect 5816 10542 5868 10548
rect 5552 10010 5580 10542
rect 5816 10464 5868 10470
rect 5816 10406 5868 10412
rect 5828 10130 5856 10406
rect 5920 10130 5948 11086
rect 5816 10124 5868 10130
rect 5816 10066 5868 10072
rect 5908 10124 5960 10130
rect 5908 10066 5960 10072
rect 5552 9982 5764 10010
rect 5632 9920 5684 9926
rect 5632 9862 5684 9868
rect 5644 9042 5672 9862
rect 5632 9036 5684 9042
rect 5632 8978 5684 8984
rect 5644 8430 5672 8978
rect 5736 8430 5764 9982
rect 5828 9926 5856 10066
rect 5816 9920 5868 9926
rect 5816 9862 5868 9868
rect 5920 8480 5948 10066
rect 6012 9654 6040 13806
rect 6288 13394 6316 22034
rect 7300 21622 7328 23530
rect 7484 23526 7512 29242
rect 7576 27538 7604 29242
rect 7944 29238 7972 29990
rect 7932 29232 7984 29238
rect 7932 29174 7984 29180
rect 8024 28756 8076 28762
rect 8024 28698 8076 28704
rect 8036 28218 8064 28698
rect 8128 28490 8156 31758
rect 8220 28506 8248 32846
rect 8312 32298 8340 33526
rect 8484 32904 8536 32910
rect 8484 32846 8536 32852
rect 8392 32836 8444 32842
rect 8392 32778 8444 32784
rect 8300 32292 8352 32298
rect 8300 32234 8352 32240
rect 8300 31680 8352 31686
rect 8300 31622 8352 31628
rect 8312 31482 8340 31622
rect 8300 31476 8352 31482
rect 8300 31418 8352 31424
rect 8404 30326 8432 32778
rect 8496 31958 8524 32846
rect 8588 32842 8616 38286
rect 9048 36242 9076 38286
rect 9588 38276 9640 38282
rect 9588 38218 9640 38224
rect 10232 38276 10284 38282
rect 10232 38218 10284 38224
rect 9128 38208 9180 38214
rect 9128 38150 9180 38156
rect 9140 36718 9168 38150
rect 9600 38010 9628 38218
rect 9588 38004 9640 38010
rect 9588 37946 9640 37952
rect 10244 37262 10272 38218
rect 11244 38208 11296 38214
rect 11244 38150 11296 38156
rect 11336 38208 11388 38214
rect 11336 38150 11388 38156
rect 11256 37874 11284 38150
rect 11348 38010 11376 38150
rect 12084 38010 12112 38898
rect 12360 38010 12388 38966
rect 20088 38962 20116 40854
rect 21914 40762 21970 41562
rect 24490 40762 24546 41562
rect 26422 40762 26478 41562
rect 28354 40762 28410 41562
rect 30930 40762 30986 41562
rect 32862 40882 32918 41562
rect 32862 40854 33088 40882
rect 32862 40762 32918 40854
rect 21928 39098 21956 40762
rect 26436 39098 26464 40762
rect 21916 39092 21968 39098
rect 21916 39034 21968 39040
rect 26424 39092 26476 39098
rect 26424 39034 26476 39040
rect 30944 39030 30972 40762
rect 33060 39794 33088 40854
rect 35438 40762 35494 41562
rect 37370 40762 37426 41562
rect 39302 40762 39358 41562
rect 33060 39766 33180 39794
rect 33152 39098 33180 39766
rect 35452 39098 35480 40762
rect 35594 39196 35902 39205
rect 35594 39194 35600 39196
rect 35656 39194 35680 39196
rect 35736 39194 35760 39196
rect 35816 39194 35840 39196
rect 35896 39194 35902 39196
rect 35656 39142 35658 39194
rect 35838 39142 35840 39194
rect 35594 39140 35600 39142
rect 35656 39140 35680 39142
rect 35736 39140 35760 39142
rect 35816 39140 35840 39142
rect 35896 39140 35902 39142
rect 35594 39131 35902 39140
rect 33140 39092 33192 39098
rect 33140 39034 33192 39040
rect 35440 39092 35492 39098
rect 35440 39034 35492 39040
rect 30932 39024 30984 39030
rect 30932 38966 30984 38972
rect 37384 38962 37412 40762
rect 12532 38956 12584 38962
rect 12532 38898 12584 38904
rect 17960 38956 18012 38962
rect 17960 38898 18012 38904
rect 19432 38956 19484 38962
rect 19432 38898 19484 38904
rect 20076 38956 20128 38962
rect 20076 38898 20128 38904
rect 22376 38956 22428 38962
rect 22376 38898 22428 38904
rect 27068 38956 27120 38962
rect 27068 38898 27120 38904
rect 27712 38956 27764 38962
rect 27712 38898 27764 38904
rect 33048 38956 33100 38962
rect 33048 38898 33100 38904
rect 35624 38956 35676 38962
rect 35624 38898 35676 38904
rect 37372 38956 37424 38962
rect 37372 38898 37424 38904
rect 11336 38004 11388 38010
rect 11336 37946 11388 37952
rect 11888 38004 11940 38010
rect 11888 37946 11940 37952
rect 12072 38004 12124 38010
rect 12072 37946 12124 37952
rect 12348 38004 12400 38010
rect 12348 37946 12400 37952
rect 11244 37868 11296 37874
rect 11244 37810 11296 37816
rect 10784 37800 10836 37806
rect 10784 37742 10836 37748
rect 10600 37664 10652 37670
rect 10600 37606 10652 37612
rect 10232 37256 10284 37262
rect 10232 37198 10284 37204
rect 9128 36712 9180 36718
rect 9128 36654 9180 36660
rect 9864 36712 9916 36718
rect 9864 36654 9916 36660
rect 9036 36236 9088 36242
rect 9036 36178 9088 36184
rect 9048 35834 9076 36178
rect 9036 35828 9088 35834
rect 9036 35770 9088 35776
rect 9048 33998 9076 35770
rect 9140 35698 9168 36654
rect 9772 36168 9824 36174
rect 9772 36110 9824 36116
rect 9220 36032 9272 36038
rect 9220 35974 9272 35980
rect 9588 36032 9640 36038
rect 9588 35974 9640 35980
rect 9128 35692 9180 35698
rect 9128 35634 9180 35640
rect 9232 35630 9260 35974
rect 9600 35766 9628 35974
rect 9588 35760 9640 35766
rect 9588 35702 9640 35708
rect 9220 35624 9272 35630
rect 9220 35566 9272 35572
rect 9784 35290 9812 36110
rect 9772 35284 9824 35290
rect 9772 35226 9824 35232
rect 9680 35148 9732 35154
rect 9680 35090 9732 35096
rect 9496 34468 9548 34474
rect 9496 34410 9548 34416
rect 9036 33992 9088 33998
rect 9036 33934 9088 33940
rect 8668 33856 8720 33862
rect 8668 33798 8720 33804
rect 8944 33856 8996 33862
rect 8944 33798 8996 33804
rect 8680 33658 8708 33798
rect 8668 33652 8720 33658
rect 8668 33594 8720 33600
rect 8956 33114 8984 33798
rect 8944 33108 8996 33114
rect 8944 33050 8996 33056
rect 8576 32836 8628 32842
rect 8576 32778 8628 32784
rect 8852 32768 8904 32774
rect 8852 32710 8904 32716
rect 8484 31952 8536 31958
rect 8484 31894 8536 31900
rect 8864 31822 8892 32710
rect 9048 31822 9076 33934
rect 9404 33856 9456 33862
rect 9404 33798 9456 33804
rect 9416 33658 9444 33798
rect 9404 33652 9456 33658
rect 9404 33594 9456 33600
rect 8484 31816 8536 31822
rect 8484 31758 8536 31764
rect 8852 31816 8904 31822
rect 8852 31758 8904 31764
rect 9036 31816 9088 31822
rect 9036 31758 9088 31764
rect 8496 30938 8524 31758
rect 8576 31408 8628 31414
rect 8576 31350 8628 31356
rect 8484 30932 8536 30938
rect 8484 30874 8536 30880
rect 8588 30802 8616 31350
rect 8576 30796 8628 30802
rect 8576 30738 8628 30744
rect 8392 30320 8444 30326
rect 8392 30262 8444 30268
rect 8576 30252 8628 30258
rect 8576 30194 8628 30200
rect 8300 29640 8352 29646
rect 8300 29582 8352 29588
rect 8312 29102 8340 29582
rect 8392 29504 8444 29510
rect 8392 29446 8444 29452
rect 8404 29345 8432 29446
rect 8390 29336 8446 29345
rect 8390 29271 8446 29280
rect 8300 29096 8352 29102
rect 8300 29038 8352 29044
rect 8300 28960 8352 28966
rect 8300 28902 8352 28908
rect 8312 28694 8340 28902
rect 8300 28688 8352 28694
rect 8300 28630 8352 28636
rect 8116 28484 8168 28490
rect 8220 28478 8340 28506
rect 8116 28426 8168 28432
rect 8208 28416 8260 28422
rect 8208 28358 8260 28364
rect 8220 28218 8248 28358
rect 8024 28212 8076 28218
rect 8024 28154 8076 28160
rect 8208 28212 8260 28218
rect 8208 28154 8260 28160
rect 8312 28098 8340 28478
rect 8128 28070 8340 28098
rect 7564 27532 7616 27538
rect 7564 27474 7616 27480
rect 7576 25294 7604 27474
rect 7656 26784 7708 26790
rect 7656 26726 7708 26732
rect 7668 26518 7696 26726
rect 7656 26512 7708 26518
rect 7656 26454 7708 26460
rect 7564 25288 7616 25294
rect 7564 25230 7616 25236
rect 7932 24744 7984 24750
rect 7932 24686 7984 24692
rect 7944 24410 7972 24686
rect 7840 24404 7892 24410
rect 7840 24346 7892 24352
rect 7932 24404 7984 24410
rect 7932 24346 7984 24352
rect 7472 23520 7524 23526
rect 7472 23462 7524 23468
rect 7656 23316 7708 23322
rect 7656 23258 7708 23264
rect 7380 23044 7432 23050
rect 7380 22986 7432 22992
rect 7472 23044 7524 23050
rect 7472 22986 7524 22992
rect 7392 22574 7420 22986
rect 7380 22568 7432 22574
rect 7380 22510 7432 22516
rect 7288 21616 7340 21622
rect 7288 21558 7340 21564
rect 6828 21480 6880 21486
rect 6828 21422 6880 21428
rect 6644 21344 6696 21350
rect 6644 21286 6696 21292
rect 6552 20460 6604 20466
rect 6552 20402 6604 20408
rect 6368 20256 6420 20262
rect 6368 20198 6420 20204
rect 6380 19786 6408 20198
rect 6564 19990 6592 20402
rect 6552 19984 6604 19990
rect 6552 19926 6604 19932
rect 6656 19854 6684 21286
rect 6840 21146 6868 21422
rect 6828 21140 6880 21146
rect 6828 21082 6880 21088
rect 7196 20256 7248 20262
rect 7196 20198 7248 20204
rect 6552 19848 6604 19854
rect 6550 19816 6552 19825
rect 6644 19848 6696 19854
rect 6604 19816 6606 19825
rect 6368 19780 6420 19786
rect 6644 19790 6696 19796
rect 6550 19751 6606 19760
rect 6368 19722 6420 19728
rect 6564 18630 6592 19751
rect 6552 18624 6604 18630
rect 6552 18566 6604 18572
rect 6564 18290 6592 18566
rect 6552 18284 6604 18290
rect 6552 18226 6604 18232
rect 6656 18222 6684 19790
rect 6920 19780 6972 19786
rect 6920 19722 6972 19728
rect 6932 19514 6960 19722
rect 7208 19514 7236 20198
rect 7380 20052 7432 20058
rect 7380 19994 7432 20000
rect 6920 19508 6972 19514
rect 6920 19450 6972 19456
rect 7196 19508 7248 19514
rect 7196 19450 7248 19456
rect 6644 18216 6696 18222
rect 6644 18158 6696 18164
rect 6920 17876 6972 17882
rect 6920 17818 6972 17824
rect 6932 17610 6960 17818
rect 6368 17604 6420 17610
rect 6368 17546 6420 17552
rect 6920 17604 6972 17610
rect 6920 17546 6972 17552
rect 6380 17338 6408 17546
rect 6368 17332 6420 17338
rect 6368 17274 6420 17280
rect 6932 15434 6960 17546
rect 6368 15428 6420 15434
rect 6368 15370 6420 15376
rect 6460 15428 6512 15434
rect 6460 15370 6512 15376
rect 6920 15428 6972 15434
rect 6920 15370 6972 15376
rect 6276 13388 6328 13394
rect 6276 13330 6328 13336
rect 6288 12306 6316 13330
rect 6380 12850 6408 15370
rect 6472 15162 6500 15370
rect 6460 15156 6512 15162
rect 6460 15098 6512 15104
rect 6932 14346 6960 15370
rect 7392 14618 7420 19994
rect 7484 19922 7512 22986
rect 7668 22438 7696 23258
rect 7748 22704 7800 22710
rect 7748 22646 7800 22652
rect 7656 22432 7708 22438
rect 7656 22374 7708 22380
rect 7472 19916 7524 19922
rect 7472 19858 7524 19864
rect 7668 17882 7696 22374
rect 7760 21894 7788 22646
rect 7748 21888 7800 21894
rect 7748 21830 7800 21836
rect 7748 21004 7800 21010
rect 7748 20946 7800 20952
rect 7760 20398 7788 20946
rect 7748 20392 7800 20398
rect 7748 20334 7800 20340
rect 7656 17876 7708 17882
rect 7656 17818 7708 17824
rect 7668 17338 7696 17818
rect 7760 17542 7788 20334
rect 7748 17536 7800 17542
rect 7748 17478 7800 17484
rect 7656 17332 7708 17338
rect 7656 17274 7708 17280
rect 7760 17218 7788 17478
rect 7668 17190 7788 17218
rect 7668 17134 7696 17190
rect 7656 17128 7708 17134
rect 7656 17070 7708 17076
rect 7668 14958 7696 17070
rect 7852 15502 7880 24346
rect 8024 23248 8076 23254
rect 8024 23190 8076 23196
rect 7930 23080 7986 23089
rect 8036 23050 8064 23190
rect 7930 23015 7986 23024
rect 8024 23044 8076 23050
rect 7944 22094 7972 23015
rect 8024 22986 8076 22992
rect 8036 22642 8064 22986
rect 8024 22636 8076 22642
rect 8024 22578 8076 22584
rect 7944 22066 8064 22094
rect 7932 21344 7984 21350
rect 7932 21286 7984 21292
rect 7944 20874 7972 21286
rect 7932 20868 7984 20874
rect 7932 20810 7984 20816
rect 7932 20052 7984 20058
rect 7932 19994 7984 20000
rect 7944 19825 7972 19994
rect 7930 19816 7986 19825
rect 7930 19751 7986 19760
rect 7932 18216 7984 18222
rect 7932 18158 7984 18164
rect 7944 17882 7972 18158
rect 7932 17876 7984 17882
rect 7932 17818 7984 17824
rect 7932 17060 7984 17066
rect 7932 17002 7984 17008
rect 7944 16697 7972 17002
rect 7930 16688 7986 16697
rect 7930 16623 7986 16632
rect 7944 15706 7972 16623
rect 7932 15700 7984 15706
rect 7932 15642 7984 15648
rect 7840 15496 7892 15502
rect 7840 15438 7892 15444
rect 7944 15162 7972 15642
rect 7932 15156 7984 15162
rect 7932 15098 7984 15104
rect 7656 14952 7708 14958
rect 7656 14894 7708 14900
rect 7380 14612 7432 14618
rect 7380 14554 7432 14560
rect 6920 14340 6972 14346
rect 6920 14282 6972 14288
rect 6932 13394 6960 14282
rect 7392 14006 7420 14554
rect 7380 14000 7432 14006
rect 7380 13942 7432 13948
rect 7668 13870 7696 14894
rect 7656 13864 7708 13870
rect 7656 13806 7708 13812
rect 7104 13728 7156 13734
rect 7104 13670 7156 13676
rect 7116 13394 7144 13670
rect 6920 13388 6972 13394
rect 6920 13330 6972 13336
rect 7104 13388 7156 13394
rect 7104 13330 7156 13336
rect 6552 13184 6604 13190
rect 6552 13126 6604 13132
rect 6564 12986 6592 13126
rect 6552 12980 6604 12986
rect 6552 12922 6604 12928
rect 6932 12918 6960 13330
rect 6920 12912 6972 12918
rect 6920 12854 6972 12860
rect 6368 12844 6420 12850
rect 6368 12786 6420 12792
rect 7116 12306 7144 13330
rect 8036 13190 8064 22066
rect 8128 19514 8156 28070
rect 8300 28008 8352 28014
rect 8300 27950 8352 27956
rect 8312 27674 8340 27950
rect 8300 27668 8352 27674
rect 8300 27610 8352 27616
rect 8588 26858 8616 30194
rect 8576 26852 8628 26858
rect 8576 26794 8628 26800
rect 8392 26784 8444 26790
rect 8392 26726 8444 26732
rect 8404 26518 8432 26726
rect 8392 26512 8444 26518
rect 8392 26454 8444 26460
rect 8588 26450 8616 26794
rect 8576 26444 8628 26450
rect 8576 26386 8628 26392
rect 8484 26308 8536 26314
rect 8484 26250 8536 26256
rect 8206 22536 8262 22545
rect 8206 22471 8208 22480
rect 8260 22471 8262 22480
rect 8208 22442 8260 22448
rect 8496 21894 8524 26250
rect 8588 22642 8616 26386
rect 8668 26240 8720 26246
rect 8668 26182 8720 26188
rect 8680 25838 8708 26182
rect 8668 25832 8720 25838
rect 8668 25774 8720 25780
rect 8668 25288 8720 25294
rect 8668 25230 8720 25236
rect 8680 24274 8708 25230
rect 8668 24268 8720 24274
rect 8668 24210 8720 24216
rect 8576 22636 8628 22642
rect 8576 22578 8628 22584
rect 8208 21888 8260 21894
rect 8208 21830 8260 21836
rect 8484 21888 8536 21894
rect 8484 21830 8536 21836
rect 8220 21350 8248 21830
rect 8864 21690 8892 31758
rect 9048 29510 9076 31758
rect 9404 31272 9456 31278
rect 9404 31214 9456 31220
rect 9416 30802 9444 31214
rect 9508 30802 9536 34410
rect 9588 33924 9640 33930
rect 9588 33866 9640 33872
rect 9600 33454 9628 33866
rect 9588 33448 9640 33454
rect 9588 33390 9640 33396
rect 9692 32978 9720 35090
rect 9876 34474 9904 36654
rect 10244 36106 10272 37198
rect 10612 36786 10640 37606
rect 10692 37120 10744 37126
rect 10692 37062 10744 37068
rect 10704 36922 10732 37062
rect 10692 36916 10744 36922
rect 10692 36858 10744 36864
rect 10600 36780 10652 36786
rect 10600 36722 10652 36728
rect 10612 36258 10640 36722
rect 10704 36378 10732 36858
rect 10692 36372 10744 36378
rect 10692 36314 10744 36320
rect 10612 36230 10732 36258
rect 10232 36100 10284 36106
rect 10232 36042 10284 36048
rect 10244 35766 10272 36042
rect 10232 35760 10284 35766
rect 10232 35702 10284 35708
rect 9864 34468 9916 34474
rect 9864 34410 9916 34416
rect 9864 33992 9916 33998
rect 9864 33934 9916 33940
rect 9876 33114 9904 33934
rect 10244 33590 10272 35702
rect 10232 33584 10284 33590
rect 10232 33526 10284 33532
rect 9864 33108 9916 33114
rect 9864 33050 9916 33056
rect 9680 32972 9732 32978
rect 9680 32914 9732 32920
rect 9692 31210 9720 32914
rect 10244 31754 10272 33526
rect 10704 31754 10732 36230
rect 10796 35154 10824 37742
rect 11256 36174 11284 37810
rect 11900 37806 11928 37946
rect 11888 37800 11940 37806
rect 11888 37742 11940 37748
rect 12440 37664 12492 37670
rect 12440 37606 12492 37612
rect 11244 36168 11296 36174
rect 11520 36168 11572 36174
rect 11244 36110 11296 36116
rect 11518 36136 11520 36145
rect 11796 36168 11848 36174
rect 11572 36136 11574 36145
rect 11256 35562 11284 36110
rect 11428 36100 11480 36106
rect 11796 36110 11848 36116
rect 11518 36071 11574 36080
rect 11704 36100 11756 36106
rect 11428 36042 11480 36048
rect 11704 36042 11756 36048
rect 11336 36032 11388 36038
rect 11336 35974 11388 35980
rect 11060 35556 11112 35562
rect 11060 35498 11112 35504
rect 11244 35556 11296 35562
rect 11244 35498 11296 35504
rect 10784 35148 10836 35154
rect 10784 35090 10836 35096
rect 10968 32836 11020 32842
rect 10968 32778 11020 32784
rect 9772 31748 9824 31754
rect 9772 31690 9824 31696
rect 10232 31748 10284 31754
rect 10232 31690 10284 31696
rect 10612 31726 10732 31754
rect 9784 31482 9812 31690
rect 9772 31476 9824 31482
rect 9772 31418 9824 31424
rect 9680 31204 9732 31210
rect 9680 31146 9732 31152
rect 9404 30796 9456 30802
rect 9404 30738 9456 30744
rect 9496 30796 9548 30802
rect 9496 30738 9548 30744
rect 9508 30258 9536 30738
rect 9588 30388 9640 30394
rect 9588 30330 9640 30336
rect 9496 30252 9548 30258
rect 9496 30194 9548 30200
rect 9508 30122 9536 30194
rect 9496 30116 9548 30122
rect 9496 30058 9548 30064
rect 9404 30048 9456 30054
rect 9404 29990 9456 29996
rect 9036 29504 9088 29510
rect 9036 29446 9088 29452
rect 9128 29096 9180 29102
rect 9128 29038 9180 29044
rect 8944 25832 8996 25838
rect 8944 25774 8996 25780
rect 8956 25498 8984 25774
rect 8944 25492 8996 25498
rect 8944 25434 8996 25440
rect 9140 24290 9168 29038
rect 9220 24608 9272 24614
rect 9220 24550 9272 24556
rect 9232 24410 9260 24550
rect 9220 24404 9272 24410
rect 9220 24346 9272 24352
rect 9140 24262 9260 24290
rect 9128 24200 9180 24206
rect 9128 24142 9180 24148
rect 9036 24064 9088 24070
rect 9036 24006 9088 24012
rect 9048 23798 9076 24006
rect 9036 23792 9088 23798
rect 9036 23734 9088 23740
rect 9140 23186 9168 24142
rect 9128 23180 9180 23186
rect 9128 23122 9180 23128
rect 8944 22976 8996 22982
rect 8944 22918 8996 22924
rect 8852 21684 8904 21690
rect 8852 21626 8904 21632
rect 8208 21344 8260 21350
rect 8208 21286 8260 21292
rect 8220 20806 8248 21286
rect 8668 20936 8720 20942
rect 8668 20878 8720 20884
rect 8208 20800 8260 20806
rect 8208 20742 8260 20748
rect 8392 20392 8444 20398
rect 8392 20334 8444 20340
rect 8208 19916 8260 19922
rect 8208 19858 8260 19864
rect 8116 19508 8168 19514
rect 8116 19450 8168 19456
rect 8220 15162 8248 19858
rect 8300 19780 8352 19786
rect 8300 19722 8352 19728
rect 8312 19310 8340 19722
rect 8404 19718 8432 20334
rect 8392 19712 8444 19718
rect 8390 19680 8392 19689
rect 8444 19680 8446 19689
rect 8390 19615 8446 19624
rect 8300 19304 8352 19310
rect 8300 19246 8352 19252
rect 8312 18358 8340 19246
rect 8300 18352 8352 18358
rect 8300 18294 8352 18300
rect 8312 17814 8340 18294
rect 8300 17808 8352 17814
rect 8300 17750 8352 17756
rect 8484 17196 8536 17202
rect 8484 17138 8536 17144
rect 8496 16726 8524 17138
rect 8484 16720 8536 16726
rect 8484 16662 8536 16668
rect 8208 15156 8260 15162
rect 8208 15098 8260 15104
rect 8024 13184 8076 13190
rect 8024 13126 8076 13132
rect 8036 12986 8064 13126
rect 8024 12980 8076 12986
rect 8024 12922 8076 12928
rect 6276 12300 6328 12306
rect 6276 12242 6328 12248
rect 7104 12300 7156 12306
rect 7104 12242 7156 12248
rect 6092 11144 6144 11150
rect 6092 11086 6144 11092
rect 6104 10810 6132 11086
rect 6092 10804 6144 10810
rect 6092 10746 6144 10752
rect 6104 10062 6132 10746
rect 6184 10668 6236 10674
rect 6184 10610 6236 10616
rect 6736 10668 6788 10674
rect 6736 10610 6788 10616
rect 6196 10266 6224 10610
rect 6748 10554 6776 10610
rect 6748 10526 6960 10554
rect 6368 10464 6420 10470
rect 6368 10406 6420 10412
rect 6380 10266 6408 10406
rect 6184 10260 6236 10266
rect 6184 10202 6236 10208
rect 6368 10260 6420 10266
rect 6368 10202 6420 10208
rect 6092 10056 6144 10062
rect 6092 9998 6144 10004
rect 6000 9648 6052 9654
rect 6000 9590 6052 9596
rect 6644 9580 6696 9586
rect 6644 9522 6696 9528
rect 6736 9580 6788 9586
rect 6736 9522 6788 9528
rect 6828 9580 6880 9586
rect 6828 9522 6880 9528
rect 6656 9489 6684 9522
rect 6642 9480 6698 9489
rect 6642 9415 6698 9424
rect 6748 9382 6776 9522
rect 6736 9376 6788 9382
rect 6736 9318 6788 9324
rect 6748 9178 6776 9318
rect 6736 9172 6788 9178
rect 6736 9114 6788 9120
rect 6840 8906 6868 9522
rect 6932 9178 6960 10526
rect 6920 9172 6972 9178
rect 6920 9114 6972 9120
rect 6000 8900 6052 8906
rect 6000 8842 6052 8848
rect 6828 8900 6880 8906
rect 6828 8842 6880 8848
rect 6012 8566 6040 8842
rect 7116 8634 7144 12242
rect 8024 12232 8076 12238
rect 8024 12174 8076 12180
rect 7840 12096 7892 12102
rect 7840 12038 7892 12044
rect 7852 11354 7880 12038
rect 7840 11348 7892 11354
rect 7840 11290 7892 11296
rect 7472 11144 7524 11150
rect 7472 11086 7524 11092
rect 7196 10668 7248 10674
rect 7196 10610 7248 10616
rect 7208 8974 7236 10610
rect 7484 10198 7512 11086
rect 7840 11076 7892 11082
rect 7840 11018 7892 11024
rect 7564 11008 7616 11014
rect 7564 10950 7616 10956
rect 7576 10266 7604 10950
rect 7564 10260 7616 10266
rect 7564 10202 7616 10208
rect 7472 10192 7524 10198
rect 7472 10134 7524 10140
rect 7852 9586 7880 11018
rect 7932 10464 7984 10470
rect 7932 10406 7984 10412
rect 7944 10062 7972 10406
rect 8036 10062 8064 12174
rect 8220 11898 8248 15098
rect 8392 15020 8444 15026
rect 8392 14962 8444 14968
rect 8404 13938 8432 14962
rect 8392 13932 8444 13938
rect 8392 13874 8444 13880
rect 8404 12434 8432 13874
rect 8312 12406 8432 12434
rect 8496 12434 8524 16662
rect 8576 16584 8628 16590
rect 8576 16526 8628 16532
rect 8588 15162 8616 16526
rect 8576 15156 8628 15162
rect 8576 15098 8628 15104
rect 8588 14006 8616 15098
rect 8680 14822 8708 20878
rect 8852 19712 8904 19718
rect 8852 19654 8904 19660
rect 8864 19446 8892 19654
rect 8852 19440 8904 19446
rect 8852 19382 8904 19388
rect 8760 19372 8812 19378
rect 8760 19314 8812 19320
rect 8772 15162 8800 19314
rect 8852 18692 8904 18698
rect 8852 18634 8904 18640
rect 8864 18068 8892 18634
rect 8956 18442 8984 22918
rect 9232 22094 9260 24262
rect 9312 23656 9364 23662
rect 9312 23598 9364 23604
rect 9324 23322 9352 23598
rect 9312 23316 9364 23322
rect 9312 23258 9364 23264
rect 9416 23118 9444 29990
rect 9600 29073 9628 30330
rect 9956 30320 10008 30326
rect 9956 30262 10008 30268
rect 9680 29572 9732 29578
rect 9680 29514 9732 29520
rect 9586 29064 9642 29073
rect 9586 28999 9642 29008
rect 9496 28688 9548 28694
rect 9496 28630 9548 28636
rect 9508 28150 9536 28630
rect 9496 28144 9548 28150
rect 9496 28086 9548 28092
rect 9496 27872 9548 27878
rect 9496 27814 9548 27820
rect 9508 27674 9536 27814
rect 9496 27668 9548 27674
rect 9496 27610 9548 27616
rect 9600 27606 9628 28999
rect 9692 28082 9720 29514
rect 9968 29510 9996 30262
rect 10048 30252 10100 30258
rect 10048 30194 10100 30200
rect 9956 29504 10008 29510
rect 9956 29446 10008 29452
rect 9968 28558 9996 29446
rect 9956 28552 10008 28558
rect 9956 28494 10008 28500
rect 9680 28076 9732 28082
rect 9680 28018 9732 28024
rect 9772 28076 9824 28082
rect 9772 28018 9824 28024
rect 9784 27878 9812 28018
rect 10060 27962 10088 30194
rect 10416 28484 10468 28490
rect 10416 28426 10468 28432
rect 10508 28484 10560 28490
rect 10508 28426 10560 28432
rect 10140 28008 10192 28014
rect 9968 27956 10140 27962
rect 9968 27950 10192 27956
rect 9968 27934 10180 27950
rect 9772 27872 9824 27878
rect 9772 27814 9824 27820
rect 9588 27600 9640 27606
rect 9588 27542 9640 27548
rect 9600 26518 9628 27542
rect 9588 26512 9640 26518
rect 9588 26454 9640 26460
rect 9680 25696 9732 25702
rect 9680 25638 9732 25644
rect 9692 25498 9720 25638
rect 9680 25492 9732 25498
rect 9680 25434 9732 25440
rect 9588 25152 9640 25158
rect 9588 25094 9640 25100
rect 9600 24954 9628 25094
rect 9588 24948 9640 24954
rect 9588 24890 9640 24896
rect 9680 24880 9732 24886
rect 9680 24822 9732 24828
rect 9692 23798 9720 24822
rect 9680 23792 9732 23798
rect 9680 23734 9732 23740
rect 9404 23112 9456 23118
rect 9404 23054 9456 23060
rect 9680 23044 9732 23050
rect 9680 22986 9732 22992
rect 9692 22234 9720 22986
rect 9680 22228 9732 22234
rect 9680 22170 9732 22176
rect 9232 22066 9628 22094
rect 9600 21690 9628 22066
rect 9784 21894 9812 27814
rect 9864 27328 9916 27334
rect 9864 27270 9916 27276
rect 9876 27130 9904 27270
rect 9864 27124 9916 27130
rect 9864 27066 9916 27072
rect 9876 25362 9904 27066
rect 9864 25356 9916 25362
rect 9864 25298 9916 25304
rect 9968 25242 9996 27934
rect 10048 27396 10100 27402
rect 10048 27338 10100 27344
rect 10060 27130 10088 27338
rect 10048 27124 10100 27130
rect 10048 27066 10100 27072
rect 10048 25900 10100 25906
rect 10048 25842 10100 25848
rect 9876 25214 9996 25242
rect 9876 24750 9904 25214
rect 10060 24886 10088 25842
rect 10140 25288 10192 25294
rect 10140 25230 10192 25236
rect 10152 24954 10180 25230
rect 10140 24948 10192 24954
rect 10140 24890 10192 24896
rect 10048 24880 10100 24886
rect 10048 24822 10100 24828
rect 10428 24818 10456 28426
rect 10520 28218 10548 28426
rect 10508 28212 10560 28218
rect 10508 28154 10560 28160
rect 10508 25220 10560 25226
rect 10508 25162 10560 25168
rect 10520 24954 10548 25162
rect 10508 24948 10560 24954
rect 10508 24890 10560 24896
rect 10416 24812 10468 24818
rect 10416 24754 10468 24760
rect 9864 24744 9916 24750
rect 9864 24686 9916 24692
rect 9876 24313 9904 24686
rect 9862 24304 9918 24313
rect 9862 24239 9918 24248
rect 10048 23520 10100 23526
rect 10048 23462 10100 23468
rect 10060 23118 10088 23462
rect 9864 23112 9916 23118
rect 9864 23054 9916 23060
rect 10048 23112 10100 23118
rect 10048 23054 10100 23060
rect 9876 22778 9904 23054
rect 9864 22772 9916 22778
rect 9864 22714 9916 22720
rect 10048 22500 10100 22506
rect 10048 22442 10100 22448
rect 10060 22098 10088 22442
rect 10140 22432 10192 22438
rect 10140 22374 10192 22380
rect 10048 22092 10100 22098
rect 10048 22034 10100 22040
rect 10152 22094 10180 22374
rect 10612 22094 10640 31726
rect 10876 31476 10928 31482
rect 10876 31418 10928 31424
rect 10784 31272 10836 31278
rect 10784 31214 10836 31220
rect 10692 29504 10744 29510
rect 10692 29446 10744 29452
rect 10704 29238 10732 29446
rect 10692 29232 10744 29238
rect 10692 29174 10744 29180
rect 10796 29102 10824 31214
rect 10888 30598 10916 31418
rect 10876 30592 10928 30598
rect 10876 30534 10928 30540
rect 10784 29096 10836 29102
rect 10784 29038 10836 29044
rect 10888 22094 10916 30534
rect 10980 29646 11008 32778
rect 10968 29640 11020 29646
rect 10968 29582 11020 29588
rect 11072 28490 11100 35498
rect 11152 35080 11204 35086
rect 11152 35022 11204 35028
rect 11060 28484 11112 28490
rect 11060 28426 11112 28432
rect 11072 27470 11100 28426
rect 11060 27464 11112 27470
rect 11060 27406 11112 27412
rect 11072 25226 11100 27406
rect 11164 26586 11192 35022
rect 11244 28144 11296 28150
rect 11242 28112 11244 28121
rect 11296 28112 11298 28121
rect 11242 28047 11298 28056
rect 11152 26580 11204 26586
rect 11152 26522 11204 26528
rect 11152 26308 11204 26314
rect 11152 26250 11204 26256
rect 11060 25220 11112 25226
rect 11060 25162 11112 25168
rect 11072 24562 11100 25162
rect 11164 24698 11192 26250
rect 11164 24670 11284 24698
rect 11072 24534 11192 24562
rect 11164 23050 11192 24534
rect 11060 23044 11112 23050
rect 11060 22986 11112 22992
rect 11152 23044 11204 23050
rect 11152 22986 11204 22992
rect 11072 22778 11100 22986
rect 11256 22930 11284 24670
rect 11164 22902 11284 22930
rect 11060 22772 11112 22778
rect 11060 22714 11112 22720
rect 10152 22066 10640 22094
rect 10796 22066 10916 22094
rect 9772 21888 9824 21894
rect 9772 21830 9824 21836
rect 9864 21888 9916 21894
rect 9864 21830 9916 21836
rect 9588 21684 9640 21690
rect 9588 21626 9640 21632
rect 9678 21584 9734 21593
rect 9404 21548 9456 21554
rect 9404 21490 9456 21496
rect 9588 21548 9640 21554
rect 9678 21519 9680 21528
rect 9588 21490 9640 21496
rect 9732 21519 9734 21528
rect 9680 21490 9732 21496
rect 9416 21026 9444 21490
rect 9600 21434 9628 21490
rect 9600 21406 9720 21434
rect 9140 20998 9444 21026
rect 9140 20097 9168 20998
rect 9588 20936 9640 20942
rect 9588 20878 9640 20884
rect 9220 20868 9272 20874
rect 9220 20810 9272 20816
rect 9496 20868 9548 20874
rect 9496 20810 9548 20816
rect 9126 20088 9182 20097
rect 9126 20023 9182 20032
rect 9034 19408 9090 19417
rect 9034 19343 9036 19352
rect 9088 19343 9090 19352
rect 9036 19314 9088 19320
rect 8956 18414 9076 18442
rect 9048 18222 9076 18414
rect 9036 18216 9088 18222
rect 9036 18158 9088 18164
rect 8944 18080 8996 18086
rect 8864 18040 8944 18068
rect 8760 15156 8812 15162
rect 8760 15098 8812 15104
rect 8864 15042 8892 18040
rect 8944 18022 8996 18028
rect 8942 17912 8998 17921
rect 8942 17847 8998 17856
rect 8956 16590 8984 17847
rect 9048 17746 9076 18158
rect 9036 17740 9088 17746
rect 9036 17682 9088 17688
rect 9036 17196 9088 17202
rect 9036 17138 9088 17144
rect 9048 16726 9076 17138
rect 9036 16720 9088 16726
rect 9036 16662 9088 16668
rect 8944 16584 8996 16590
rect 8944 16526 8996 16532
rect 8956 15178 8984 16526
rect 8956 15150 9076 15178
rect 8772 15014 8892 15042
rect 8944 15020 8996 15026
rect 8668 14816 8720 14822
rect 8668 14758 8720 14764
rect 8680 14618 8708 14758
rect 8668 14612 8720 14618
rect 8668 14554 8720 14560
rect 8772 14346 8800 15014
rect 8944 14962 8996 14968
rect 8956 14822 8984 14962
rect 9048 14890 9076 15150
rect 9036 14884 9088 14890
rect 9036 14826 9088 14832
rect 8944 14816 8996 14822
rect 8944 14758 8996 14764
rect 8852 14612 8904 14618
rect 8852 14554 8904 14560
rect 8760 14340 8812 14346
rect 8760 14282 8812 14288
rect 8668 14272 8720 14278
rect 8668 14214 8720 14220
rect 8680 14074 8708 14214
rect 8668 14068 8720 14074
rect 8668 14010 8720 14016
rect 8576 14000 8628 14006
rect 8576 13942 8628 13948
rect 8576 13184 8628 13190
rect 8576 13126 8628 13132
rect 8588 12918 8616 13126
rect 8576 12912 8628 12918
rect 8576 12854 8628 12860
rect 8496 12406 8616 12434
rect 8312 12238 8340 12406
rect 8300 12232 8352 12238
rect 8300 12174 8352 12180
rect 8208 11892 8260 11898
rect 8208 11834 8260 11840
rect 8220 11218 8248 11834
rect 8312 11558 8340 12174
rect 8300 11552 8352 11558
rect 8300 11494 8352 11500
rect 8208 11212 8260 11218
rect 8208 11154 8260 11160
rect 8116 11076 8168 11082
rect 8116 11018 8168 11024
rect 7932 10056 7984 10062
rect 7932 9998 7984 10004
rect 8024 10056 8076 10062
rect 8024 9998 8076 10004
rect 8128 9586 8156 11018
rect 8220 10470 8248 11154
rect 8312 10470 8340 11494
rect 8588 11150 8616 12406
rect 8576 11144 8628 11150
rect 8576 11086 8628 11092
rect 8208 10464 8260 10470
rect 8208 10406 8260 10412
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8392 10192 8444 10198
rect 8392 10134 8444 10140
rect 8208 10124 8260 10130
rect 8208 10066 8260 10072
rect 8220 9654 8248 10066
rect 8404 10010 8432 10134
rect 8680 10130 8708 14010
rect 8864 12442 8892 14554
rect 8852 12436 8904 12442
rect 8956 12434 8984 14758
rect 9140 14550 9168 20023
rect 9232 18834 9260 20810
rect 9508 20618 9536 20810
rect 9600 20777 9628 20878
rect 9692 20806 9720 21406
rect 9784 21146 9812 21830
rect 9772 21140 9824 21146
rect 9772 21082 9824 21088
rect 9680 20800 9732 20806
rect 9586 20768 9642 20777
rect 9680 20742 9732 20748
rect 9586 20703 9642 20712
rect 9770 20632 9826 20641
rect 9508 20590 9770 20618
rect 9770 20567 9826 20576
rect 9680 19984 9732 19990
rect 9494 19952 9550 19961
rect 9680 19926 9732 19932
rect 9494 19887 9550 19896
rect 9508 19854 9536 19887
rect 9312 19848 9364 19854
rect 9312 19790 9364 19796
rect 9496 19848 9548 19854
rect 9496 19790 9548 19796
rect 9588 19848 9640 19854
rect 9588 19790 9640 19796
rect 9324 19310 9352 19790
rect 9600 19514 9628 19790
rect 9588 19508 9640 19514
rect 9588 19450 9640 19456
rect 9496 19372 9548 19378
rect 9496 19314 9548 19320
rect 9312 19304 9364 19310
rect 9312 19246 9364 19252
rect 9220 18828 9272 18834
rect 9220 18770 9272 18776
rect 9220 17332 9272 17338
rect 9220 17274 9272 17280
rect 9232 15162 9260 17274
rect 9220 15156 9272 15162
rect 9220 15098 9272 15104
rect 9128 14544 9180 14550
rect 9128 14486 9180 14492
rect 9036 14408 9088 14414
rect 9036 14350 9088 14356
rect 9048 13530 9076 14350
rect 9036 13524 9088 13530
rect 9036 13466 9088 13472
rect 9220 13320 9272 13326
rect 9220 13262 9272 13268
rect 8956 12406 9076 12434
rect 8852 12378 8904 12384
rect 8760 12232 8812 12238
rect 8760 12174 8812 12180
rect 8772 11898 8800 12174
rect 8760 11892 8812 11898
rect 8760 11834 8812 11840
rect 8668 10124 8720 10130
rect 8668 10066 8720 10072
rect 8404 9994 8524 10010
rect 8404 9988 8536 9994
rect 8404 9982 8484 9988
rect 8484 9930 8536 9936
rect 8208 9648 8260 9654
rect 8208 9590 8260 9596
rect 8496 9586 8524 9930
rect 7840 9580 7892 9586
rect 7840 9522 7892 9528
rect 8116 9580 8168 9586
rect 8116 9522 8168 9528
rect 8484 9580 8536 9586
rect 8484 9522 8536 9528
rect 7472 9444 7524 9450
rect 7472 9386 7524 9392
rect 8208 9444 8260 9450
rect 8208 9386 8260 9392
rect 7196 8968 7248 8974
rect 7196 8910 7248 8916
rect 7104 8628 7156 8634
rect 7104 8570 7156 8576
rect 6000 8560 6052 8566
rect 6000 8502 6052 8508
rect 5828 8452 5948 8480
rect 5540 8424 5592 8430
rect 5540 8366 5592 8372
rect 5632 8424 5684 8430
rect 5632 8366 5684 8372
rect 5724 8424 5776 8430
rect 5724 8366 5776 8372
rect 5552 8090 5580 8366
rect 5540 8084 5592 8090
rect 5540 8026 5592 8032
rect 5448 7404 5500 7410
rect 5448 7346 5500 7352
rect 5644 7342 5672 8366
rect 5736 7886 5764 8366
rect 5828 8090 5856 8452
rect 5908 8356 5960 8362
rect 5908 8298 5960 8304
rect 5816 8084 5868 8090
rect 5816 8026 5868 8032
rect 5920 7886 5948 8298
rect 5724 7880 5776 7886
rect 5724 7822 5776 7828
rect 5908 7880 5960 7886
rect 5908 7822 5960 7828
rect 6012 7410 6040 8502
rect 6276 8492 6328 8498
rect 6276 8434 6328 8440
rect 6288 8294 6316 8434
rect 6460 8356 6512 8362
rect 6460 8298 6512 8304
rect 6276 8288 6328 8294
rect 6276 8230 6328 8236
rect 6368 8084 6420 8090
rect 6472 8072 6500 8298
rect 6828 8288 6880 8294
rect 6828 8230 6880 8236
rect 6420 8044 6500 8072
rect 6368 8026 6420 8032
rect 6092 7744 6144 7750
rect 6092 7686 6144 7692
rect 6552 7744 6604 7750
rect 6552 7686 6604 7692
rect 6104 7546 6132 7686
rect 6564 7546 6592 7686
rect 6092 7540 6144 7546
rect 6092 7482 6144 7488
rect 6552 7540 6604 7546
rect 6552 7482 6604 7488
rect 6000 7404 6052 7410
rect 6000 7346 6052 7352
rect 5632 7336 5684 7342
rect 5632 7278 5684 7284
rect 6012 7002 6040 7346
rect 6840 7342 6868 8230
rect 6920 7948 6972 7954
rect 6920 7890 6972 7896
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 6000 6996 6052 7002
rect 6000 6938 6052 6944
rect 6460 6724 6512 6730
rect 6460 6666 6512 6672
rect 6472 5710 6500 6666
rect 6932 5778 6960 7890
rect 7196 7812 7248 7818
rect 7196 7754 7248 7760
rect 7208 7546 7236 7754
rect 7196 7540 7248 7546
rect 7196 7482 7248 7488
rect 7484 6254 7512 9386
rect 8024 8832 8076 8838
rect 8024 8774 8076 8780
rect 8036 7546 8064 8774
rect 8024 7540 8076 7546
rect 8024 7482 8076 7488
rect 8220 6798 8248 9386
rect 8484 8832 8536 8838
rect 8484 8774 8536 8780
rect 8668 8832 8720 8838
rect 8668 8774 8720 8780
rect 8496 8362 8524 8774
rect 8680 8498 8708 8774
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 8484 8356 8536 8362
rect 8484 8298 8536 8304
rect 8680 8294 8708 8434
rect 8668 8288 8720 8294
rect 8668 8230 8720 8236
rect 8680 8090 8708 8230
rect 8668 8084 8720 8090
rect 8668 8026 8720 8032
rect 8300 7880 8352 7886
rect 8300 7822 8352 7828
rect 8208 6792 8260 6798
rect 8208 6734 8260 6740
rect 8220 6322 8248 6734
rect 8312 6662 8340 7822
rect 8300 6656 8352 6662
rect 8300 6598 8352 6604
rect 8208 6316 8260 6322
rect 8208 6258 8260 6264
rect 7472 6248 7524 6254
rect 7472 6190 7524 6196
rect 7380 6112 7432 6118
rect 7380 6054 7432 6060
rect 8208 6112 8260 6118
rect 8208 6054 8260 6060
rect 6920 5772 6972 5778
rect 6920 5714 6972 5720
rect 6460 5704 6512 5710
rect 6460 5646 6512 5652
rect 5632 5636 5684 5642
rect 5632 5578 5684 5584
rect 5644 5370 5672 5578
rect 5632 5364 5684 5370
rect 5632 5306 5684 5312
rect 6932 4146 6960 5714
rect 7392 5370 7420 6054
rect 8220 5914 8248 6054
rect 8208 5908 8260 5914
rect 8208 5850 8260 5856
rect 8312 5710 8340 6598
rect 8300 5704 8352 5710
rect 8300 5646 8352 5652
rect 8208 5568 8260 5574
rect 8208 5510 8260 5516
rect 7380 5364 7432 5370
rect 7380 5306 7432 5312
rect 8220 5234 8248 5510
rect 8208 5228 8260 5234
rect 8208 5170 8260 5176
rect 8312 4298 8340 5646
rect 8312 4270 8432 4298
rect 8404 4214 8432 4270
rect 8392 4208 8444 4214
rect 8392 4150 8444 4156
rect 6920 4140 6972 4146
rect 6920 4082 6972 4088
rect 8392 2848 8444 2854
rect 8392 2790 8444 2796
rect 4214 2748 4522 2757
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 5368 2746 5488 2774
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2683 4522 2692
rect 5460 2446 5488 2746
rect 8404 2446 8432 2790
rect 8772 2650 8800 11834
rect 9048 11354 9076 12406
rect 9036 11348 9088 11354
rect 9036 11290 9088 11296
rect 8852 11212 8904 11218
rect 8852 11154 8904 11160
rect 8864 10674 8892 11154
rect 9048 11150 9076 11290
rect 9036 11144 9088 11150
rect 8956 11104 9036 11132
rect 8956 10810 8984 11104
rect 9036 11086 9088 11092
rect 8944 10804 8996 10810
rect 8944 10746 8996 10752
rect 8852 10668 8904 10674
rect 8852 10610 8904 10616
rect 9232 10146 9260 13262
rect 9324 11898 9352 19246
rect 9508 17270 9536 19314
rect 9588 17536 9640 17542
rect 9588 17478 9640 17484
rect 9496 17264 9548 17270
rect 9496 17206 9548 17212
rect 9600 16998 9628 17478
rect 9692 17270 9720 19926
rect 9784 17882 9812 20567
rect 9876 18834 9904 21830
rect 10048 21548 10100 21554
rect 10048 21490 10100 21496
rect 9956 21412 10008 21418
rect 9956 21354 10008 21360
rect 9968 20942 9996 21354
rect 10060 21321 10088 21490
rect 10046 21312 10102 21321
rect 10046 21247 10102 21256
rect 10152 21146 10180 22066
rect 10416 22024 10468 22030
rect 10416 21966 10468 21972
rect 10322 21584 10378 21593
rect 10232 21548 10284 21554
rect 10322 21519 10324 21528
rect 10232 21490 10284 21496
rect 10376 21519 10378 21528
rect 10324 21490 10376 21496
rect 10140 21140 10192 21146
rect 10140 21082 10192 21088
rect 9956 20936 10008 20942
rect 9956 20878 10008 20884
rect 10140 20936 10192 20942
rect 10140 20878 10192 20884
rect 9968 19854 9996 20878
rect 10048 20868 10100 20874
rect 10048 20810 10100 20816
rect 10060 20330 10088 20810
rect 10152 20754 10180 20878
rect 10244 20874 10272 21490
rect 10232 20868 10284 20874
rect 10232 20810 10284 20816
rect 10152 20726 10272 20754
rect 10138 20360 10194 20369
rect 10048 20324 10100 20330
rect 10138 20295 10194 20304
rect 10048 20266 10100 20272
rect 10060 19854 10088 20266
rect 10152 19854 10180 20295
rect 9956 19848 10008 19854
rect 9956 19790 10008 19796
rect 10048 19848 10100 19854
rect 10048 19790 10100 19796
rect 10140 19848 10192 19854
rect 10140 19790 10192 19796
rect 10244 19378 10272 20726
rect 9956 19372 10008 19378
rect 9956 19314 10008 19320
rect 10232 19372 10284 19378
rect 10232 19314 10284 19320
rect 9864 18828 9916 18834
rect 9864 18770 9916 18776
rect 9772 17876 9824 17882
rect 9772 17818 9824 17824
rect 9680 17264 9732 17270
rect 9680 17206 9732 17212
rect 9588 16992 9640 16998
rect 9588 16934 9640 16940
rect 9404 16516 9456 16522
rect 9404 16458 9456 16464
rect 9416 16250 9444 16458
rect 9404 16244 9456 16250
rect 9404 16186 9456 16192
rect 9496 15700 9548 15706
rect 9496 15642 9548 15648
rect 9404 14952 9456 14958
rect 9404 14894 9456 14900
rect 9416 13190 9444 14894
rect 9404 13184 9456 13190
rect 9404 13126 9456 13132
rect 9416 12238 9444 13126
rect 9508 12434 9536 15642
rect 9600 15094 9628 16934
rect 9680 16516 9732 16522
rect 9680 16458 9732 16464
rect 9588 15088 9640 15094
rect 9588 15030 9640 15036
rect 9586 14376 9642 14385
rect 9586 14311 9588 14320
rect 9640 14311 9642 14320
rect 9588 14282 9640 14288
rect 9586 13696 9642 13705
rect 9586 13631 9642 13640
rect 9600 13394 9628 13631
rect 9588 13388 9640 13394
rect 9588 13330 9640 13336
rect 9588 13184 9640 13190
rect 9588 13126 9640 13132
rect 9600 12714 9628 13126
rect 9692 12850 9720 16458
rect 9772 14816 9824 14822
rect 9772 14758 9824 14764
rect 9680 12844 9732 12850
rect 9680 12786 9732 12792
rect 9588 12708 9640 12714
rect 9588 12650 9640 12656
rect 9508 12406 9628 12434
rect 9404 12232 9456 12238
rect 9404 12174 9456 12180
rect 9312 11892 9364 11898
rect 9312 11834 9364 11840
rect 9312 11756 9364 11762
rect 9312 11698 9364 11704
rect 9324 11286 9352 11698
rect 9496 11620 9548 11626
rect 9496 11562 9548 11568
rect 9508 11286 9536 11562
rect 9312 11280 9364 11286
rect 9312 11222 9364 11228
rect 9496 11280 9548 11286
rect 9496 11222 9548 11228
rect 9404 11144 9456 11150
rect 9404 11086 9456 11092
rect 9416 10810 9444 11086
rect 9404 10804 9456 10810
rect 9404 10746 9456 10752
rect 8956 10118 9260 10146
rect 8956 10062 8984 10118
rect 8944 10056 8996 10062
rect 8944 9998 8996 10004
rect 8956 9586 8984 9998
rect 9496 9920 9548 9926
rect 9496 9862 9548 9868
rect 9312 9648 9364 9654
rect 9312 9590 9364 9596
rect 8944 9580 8996 9586
rect 8944 9522 8996 9528
rect 8852 8084 8904 8090
rect 8852 8026 8904 8032
rect 8864 7886 8892 8026
rect 8852 7880 8904 7886
rect 8852 7822 8904 7828
rect 8852 6384 8904 6390
rect 8852 6326 8904 6332
rect 8864 6118 8892 6326
rect 8852 6112 8904 6118
rect 8852 6054 8904 6060
rect 8864 5370 8892 6054
rect 8852 5364 8904 5370
rect 8852 5306 8904 5312
rect 8760 2644 8812 2650
rect 8760 2586 8812 2592
rect 8956 2514 8984 9522
rect 9324 9489 9352 9590
rect 9310 9480 9366 9489
rect 9310 9415 9366 9424
rect 9220 8628 9272 8634
rect 9220 8570 9272 8576
rect 9404 8628 9456 8634
rect 9404 8570 9456 8576
rect 9232 7886 9260 8570
rect 9416 7954 9444 8570
rect 9404 7948 9456 7954
rect 9404 7890 9456 7896
rect 9220 7880 9272 7886
rect 9220 7822 9272 7828
rect 9416 7410 9444 7890
rect 9404 7404 9456 7410
rect 9404 7346 9456 7352
rect 9508 6798 9536 9862
rect 9600 8566 9628 12406
rect 9588 8560 9640 8566
rect 9588 8502 9640 8508
rect 9600 8378 9628 8502
rect 9692 8480 9720 12786
rect 9784 10130 9812 14758
rect 9864 14408 9916 14414
rect 9864 14350 9916 14356
rect 9876 12986 9904 14350
rect 9968 13938 9996 19314
rect 10336 18714 10364 21490
rect 10428 20602 10456 21966
rect 10416 20596 10468 20602
rect 10416 20538 10468 20544
rect 10796 20058 10824 22066
rect 11164 21690 11192 22902
rect 11348 22094 11376 35974
rect 11440 34678 11468 36042
rect 11428 34672 11480 34678
rect 11428 34614 11480 34620
rect 11716 34490 11744 36042
rect 11440 34462 11744 34490
rect 11440 32910 11468 34462
rect 11520 34400 11572 34406
rect 11520 34342 11572 34348
rect 11532 33998 11560 34342
rect 11808 34066 11836 36110
rect 12452 36106 12480 37606
rect 12440 36100 12492 36106
rect 12440 36042 12492 36048
rect 12440 35488 12492 35494
rect 12440 35430 12492 35436
rect 12452 35018 12480 35430
rect 12440 35012 12492 35018
rect 12440 34954 12492 34960
rect 12164 34740 12216 34746
rect 12164 34682 12216 34688
rect 11888 34672 11940 34678
rect 11888 34614 11940 34620
rect 11796 34060 11848 34066
rect 11796 34002 11848 34008
rect 11520 33992 11572 33998
rect 11520 33934 11572 33940
rect 11612 33312 11664 33318
rect 11612 33254 11664 33260
rect 11624 33114 11652 33254
rect 11612 33108 11664 33114
rect 11612 33050 11664 33056
rect 11704 33040 11756 33046
rect 11704 32982 11756 32988
rect 11428 32904 11480 32910
rect 11428 32846 11480 32852
rect 11440 30258 11468 32846
rect 11612 32768 11664 32774
rect 11612 32710 11664 32716
rect 11624 32570 11652 32710
rect 11612 32564 11664 32570
rect 11612 32506 11664 32512
rect 11612 32428 11664 32434
rect 11612 32370 11664 32376
rect 11624 32230 11652 32370
rect 11612 32224 11664 32230
rect 11612 32166 11664 32172
rect 11624 31890 11652 32166
rect 11612 31884 11664 31890
rect 11612 31826 11664 31832
rect 11520 31680 11572 31686
rect 11520 31622 11572 31628
rect 11532 31346 11560 31622
rect 11612 31476 11664 31482
rect 11612 31418 11664 31424
rect 11624 31346 11652 31418
rect 11520 31340 11572 31346
rect 11520 31282 11572 31288
rect 11612 31340 11664 31346
rect 11612 31282 11664 31288
rect 11428 30252 11480 30258
rect 11428 30194 11480 30200
rect 11440 26926 11468 30194
rect 11624 28966 11652 31282
rect 11716 31226 11744 32982
rect 11808 32570 11836 34002
rect 11900 32910 11928 34614
rect 12072 34196 12124 34202
rect 12072 34138 12124 34144
rect 11980 33856 12032 33862
rect 11980 33798 12032 33804
rect 11992 33522 12020 33798
rect 11980 33516 12032 33522
rect 11980 33458 12032 33464
rect 11888 32904 11940 32910
rect 12084 32858 12112 34138
rect 12176 33046 12204 34682
rect 12256 34604 12308 34610
rect 12256 34546 12308 34552
rect 12164 33040 12216 33046
rect 12164 32982 12216 32988
rect 12162 32872 12218 32881
rect 11940 32852 12020 32858
rect 11888 32846 12020 32852
rect 11900 32830 12020 32846
rect 12084 32842 12162 32858
rect 11796 32564 11848 32570
rect 11796 32506 11848 32512
rect 11808 32178 11836 32506
rect 11808 32150 11928 32178
rect 11796 31748 11848 31754
rect 11796 31690 11848 31696
rect 11808 31414 11836 31690
rect 11796 31408 11848 31414
rect 11796 31350 11848 31356
rect 11900 31346 11928 32150
rect 11992 31482 12020 32830
rect 12072 32836 12162 32842
rect 12124 32830 12162 32836
rect 12162 32807 12218 32816
rect 12072 32778 12124 32784
rect 12268 32774 12296 34546
rect 12452 34542 12480 34954
rect 12440 34536 12492 34542
rect 12440 34478 12492 34484
rect 12256 32768 12308 32774
rect 12256 32710 12308 32716
rect 12348 32768 12400 32774
rect 12348 32710 12400 32716
rect 11980 31476 12032 31482
rect 11980 31418 12032 31424
rect 11888 31340 11940 31346
rect 11888 31282 11940 31288
rect 11716 31198 11928 31226
rect 11704 30660 11756 30666
rect 11704 30602 11756 30608
rect 11716 30258 11744 30602
rect 11900 30258 11928 31198
rect 12268 30258 12296 32710
rect 12360 32570 12388 32710
rect 12348 32564 12400 32570
rect 12348 32506 12400 32512
rect 12348 31340 12400 31346
rect 12348 31282 12400 31288
rect 11704 30252 11756 30258
rect 11704 30194 11756 30200
rect 11888 30252 11940 30258
rect 12256 30252 12308 30258
rect 11888 30194 11940 30200
rect 12176 30212 12256 30240
rect 11520 28960 11572 28966
rect 11520 28902 11572 28908
rect 11612 28960 11664 28966
rect 11612 28902 11664 28908
rect 11532 28694 11560 28902
rect 11520 28688 11572 28694
rect 11520 28630 11572 28636
rect 11612 27328 11664 27334
rect 11612 27270 11664 27276
rect 11624 27130 11652 27270
rect 11612 27124 11664 27130
rect 11612 27066 11664 27072
rect 11428 26920 11480 26926
rect 11428 26862 11480 26868
rect 11900 26858 11928 30194
rect 12072 28688 12124 28694
rect 12072 28630 12124 28636
rect 11980 28416 12032 28422
rect 11980 28358 12032 28364
rect 11992 28150 12020 28358
rect 11980 28144 12032 28150
rect 11980 28086 12032 28092
rect 12084 28014 12112 28630
rect 11980 28008 12032 28014
rect 11980 27950 12032 27956
rect 12072 28008 12124 28014
rect 12072 27950 12124 27956
rect 11992 27878 12020 27950
rect 11980 27872 12032 27878
rect 11980 27814 12032 27820
rect 11992 27538 12020 27814
rect 11980 27532 12032 27538
rect 11980 27474 12032 27480
rect 11980 26920 12032 26926
rect 11980 26862 12032 26868
rect 11888 26852 11940 26858
rect 11888 26794 11940 26800
rect 11992 25838 12020 26862
rect 11980 25832 12032 25838
rect 11980 25774 12032 25780
rect 12084 25430 12112 27950
rect 12176 27112 12204 30212
rect 12256 30194 12308 30200
rect 12360 30054 12388 31282
rect 12256 30048 12308 30054
rect 12256 29990 12308 29996
rect 12348 30048 12400 30054
rect 12348 29990 12400 29996
rect 12268 29850 12296 29990
rect 12256 29844 12308 29850
rect 12256 29786 12308 29792
rect 12348 27396 12400 27402
rect 12348 27338 12400 27344
rect 12256 27124 12308 27130
rect 12176 27084 12256 27112
rect 12256 27066 12308 27072
rect 12072 25424 12124 25430
rect 12072 25366 12124 25372
rect 11796 25220 11848 25226
rect 11796 25162 11848 25168
rect 11520 23044 11572 23050
rect 11520 22986 11572 22992
rect 11428 22636 11480 22642
rect 11428 22578 11480 22584
rect 11440 22506 11468 22578
rect 11428 22500 11480 22506
rect 11428 22442 11480 22448
rect 11256 22066 11376 22094
rect 11152 21684 11204 21690
rect 11152 21626 11204 21632
rect 10968 21344 11020 21350
rect 10968 21286 11020 21292
rect 10980 20806 11008 21286
rect 10968 20800 11020 20806
rect 10968 20742 11020 20748
rect 10784 20052 10836 20058
rect 10784 19994 10836 20000
rect 10876 18828 10928 18834
rect 10876 18770 10928 18776
rect 10152 18686 10364 18714
rect 10048 18624 10100 18630
rect 10048 18566 10100 18572
rect 10060 17746 10088 18566
rect 10048 17740 10100 17746
rect 10048 17682 10100 17688
rect 10152 17338 10180 18686
rect 10324 18624 10376 18630
rect 10324 18566 10376 18572
rect 10232 18352 10284 18358
rect 10232 18294 10284 18300
rect 10140 17332 10192 17338
rect 10140 17274 10192 17280
rect 10244 15706 10272 18294
rect 10336 17678 10364 18566
rect 10506 18456 10562 18465
rect 10506 18391 10562 18400
rect 10520 18086 10548 18391
rect 10508 18080 10560 18086
rect 10888 18057 10916 18770
rect 10508 18022 10560 18028
rect 10874 18048 10930 18057
rect 10874 17983 10930 17992
rect 10874 17776 10930 17785
rect 10874 17711 10930 17720
rect 10324 17672 10376 17678
rect 10324 17614 10376 17620
rect 10508 17672 10560 17678
rect 10508 17614 10560 17620
rect 10336 17202 10364 17614
rect 10324 17196 10376 17202
rect 10324 17138 10376 17144
rect 10416 17196 10468 17202
rect 10416 17138 10468 17144
rect 10324 16040 10376 16046
rect 10324 15982 10376 15988
rect 10232 15700 10284 15706
rect 10232 15642 10284 15648
rect 10232 14816 10284 14822
rect 10232 14758 10284 14764
rect 10244 14482 10272 14758
rect 10232 14476 10284 14482
rect 10232 14418 10284 14424
rect 10140 14000 10192 14006
rect 10140 13942 10192 13948
rect 9956 13932 10008 13938
rect 9956 13874 10008 13880
rect 10152 13326 10180 13942
rect 10336 13530 10364 15982
rect 10428 13530 10456 17138
rect 10324 13524 10376 13530
rect 10324 13466 10376 13472
rect 10416 13524 10468 13530
rect 10416 13466 10468 13472
rect 10140 13320 10192 13326
rect 10060 13268 10140 13274
rect 10060 13262 10192 13268
rect 9956 13252 10008 13258
rect 9956 13194 10008 13200
rect 10060 13246 10180 13262
rect 9864 12980 9916 12986
rect 9864 12922 9916 12928
rect 9876 11218 9904 12922
rect 9864 11212 9916 11218
rect 9864 11154 9916 11160
rect 9772 10124 9824 10130
rect 9772 10066 9824 10072
rect 9876 9058 9904 11154
rect 9968 10266 9996 13194
rect 10060 12238 10088 13246
rect 10230 13016 10286 13025
rect 10230 12951 10286 12960
rect 10244 12850 10272 12951
rect 10232 12844 10284 12850
rect 10232 12786 10284 12792
rect 10140 12640 10192 12646
rect 10140 12582 10192 12588
rect 10048 12232 10100 12238
rect 10048 12174 10100 12180
rect 9956 10260 10008 10266
rect 9956 10202 10008 10208
rect 9956 9580 10008 9586
rect 9956 9522 10008 9528
rect 9968 9217 9996 9522
rect 10048 9376 10100 9382
rect 10048 9318 10100 9324
rect 9954 9208 10010 9217
rect 9954 9143 10010 9152
rect 9784 9042 9904 9058
rect 10060 9042 10088 9318
rect 9772 9036 9904 9042
rect 9824 9030 9904 9036
rect 9772 8978 9824 8984
rect 9876 8634 9904 9030
rect 10048 9036 10100 9042
rect 10048 8978 10100 8984
rect 10152 8634 10180 12582
rect 10232 12436 10284 12442
rect 10232 12378 10284 12384
rect 10244 12238 10272 12378
rect 10232 12232 10284 12238
rect 10232 12174 10284 12180
rect 10244 10606 10272 12174
rect 10336 11694 10364 13466
rect 10428 12986 10456 13466
rect 10416 12980 10468 12986
rect 10416 12922 10468 12928
rect 10520 12434 10548 17614
rect 10888 17610 10916 17711
rect 10876 17604 10928 17610
rect 10876 17546 10928 17552
rect 10888 17338 10916 17546
rect 10876 17332 10928 17338
rect 10876 17274 10928 17280
rect 10980 13802 11008 20742
rect 11150 19000 11206 19009
rect 11150 18935 11206 18944
rect 11164 18902 11192 18935
rect 11152 18896 11204 18902
rect 11152 18838 11204 18844
rect 11152 18148 11204 18154
rect 11152 18090 11204 18096
rect 11060 18080 11112 18086
rect 11060 18022 11112 18028
rect 11072 17678 11100 18022
rect 11164 17746 11192 18090
rect 11152 17740 11204 17746
rect 11152 17682 11204 17688
rect 11060 17672 11112 17678
rect 11060 17614 11112 17620
rect 11164 17134 11192 17682
rect 11256 17626 11284 22066
rect 11532 21026 11560 22986
rect 11612 22500 11664 22506
rect 11612 22442 11664 22448
rect 11624 21894 11652 22442
rect 11808 21894 11836 25162
rect 11980 25152 12032 25158
rect 11980 25094 12032 25100
rect 11992 24954 12020 25094
rect 11980 24948 12032 24954
rect 11980 24890 12032 24896
rect 12268 24886 12296 27066
rect 12360 26994 12388 27338
rect 12348 26988 12400 26994
rect 12348 26930 12400 26936
rect 12348 26852 12400 26858
rect 12348 26794 12400 26800
rect 12360 26382 12388 26794
rect 12348 26376 12400 26382
rect 12348 26318 12400 26324
rect 12348 25424 12400 25430
rect 12348 25366 12400 25372
rect 12360 25129 12388 25366
rect 12346 25120 12402 25129
rect 12346 25055 12402 25064
rect 12440 24948 12492 24954
rect 12440 24890 12492 24896
rect 12256 24880 12308 24886
rect 12256 24822 12308 24828
rect 12452 23186 12480 24890
rect 12440 23180 12492 23186
rect 12440 23122 12492 23128
rect 12452 22778 12480 23122
rect 12544 22778 12572 38898
rect 14004 38888 14056 38894
rect 14004 38830 14056 38836
rect 12808 38752 12860 38758
rect 12808 38694 12860 38700
rect 12716 38412 12768 38418
rect 12716 38354 12768 38360
rect 12624 36032 12676 36038
rect 12624 35974 12676 35980
rect 12636 34746 12664 35974
rect 12728 35834 12756 38354
rect 12820 38282 12848 38694
rect 13636 38480 13688 38486
rect 13636 38422 13688 38428
rect 13452 38344 13504 38350
rect 13452 38286 13504 38292
rect 12808 38276 12860 38282
rect 12808 38218 12860 38224
rect 13174 37904 13230 37913
rect 13174 37839 13176 37848
rect 13228 37839 13230 37848
rect 13176 37810 13228 37816
rect 13084 37800 13136 37806
rect 13084 37742 13136 37748
rect 12992 36576 13044 36582
rect 12992 36518 13044 36524
rect 13004 36106 13032 36518
rect 12808 36100 12860 36106
rect 12808 36042 12860 36048
rect 12992 36100 13044 36106
rect 12992 36042 13044 36048
rect 12716 35828 12768 35834
rect 12716 35770 12768 35776
rect 12820 35544 12848 36042
rect 12728 35516 12848 35544
rect 12624 34740 12676 34746
rect 12624 34682 12676 34688
rect 12728 34610 12756 35516
rect 13004 35442 13032 36042
rect 12820 35414 13032 35442
rect 12716 34604 12768 34610
rect 12716 34546 12768 34552
rect 12624 32292 12676 32298
rect 12624 32234 12676 32240
rect 12636 32201 12664 32234
rect 12622 32192 12678 32201
rect 12622 32127 12678 32136
rect 12716 29640 12768 29646
rect 12716 29582 12768 29588
rect 12728 29170 12756 29582
rect 12716 29164 12768 29170
rect 12716 29106 12768 29112
rect 12624 28960 12676 28966
rect 12624 28902 12676 28908
rect 12636 28082 12664 28902
rect 12624 28076 12676 28082
rect 12624 28018 12676 28024
rect 12636 27674 12664 28018
rect 12624 27668 12676 27674
rect 12624 27610 12676 27616
rect 12624 26376 12676 26382
rect 12624 26318 12676 26324
rect 12636 25294 12664 26318
rect 12624 25288 12676 25294
rect 12624 25230 12676 25236
rect 12728 24274 12756 29106
rect 12820 25242 12848 35414
rect 13096 31929 13124 37742
rect 13268 37732 13320 37738
rect 13268 37674 13320 37680
rect 13280 36174 13308 37674
rect 13268 36168 13320 36174
rect 13268 36110 13320 36116
rect 13176 35692 13228 35698
rect 13176 35634 13228 35640
rect 13360 35692 13412 35698
rect 13360 35634 13412 35640
rect 13188 33810 13216 35634
rect 13372 33862 13400 35634
rect 13268 33856 13320 33862
rect 13188 33804 13268 33810
rect 13188 33798 13320 33804
rect 13360 33856 13412 33862
rect 13360 33798 13412 33804
rect 13188 33782 13308 33798
rect 13188 33658 13216 33782
rect 13176 33652 13228 33658
rect 13176 33594 13228 33600
rect 13082 31920 13138 31929
rect 13082 31855 13138 31864
rect 12992 31680 13044 31686
rect 12992 31622 13044 31628
rect 13004 31482 13032 31622
rect 12992 31476 13044 31482
rect 12992 31418 13044 31424
rect 13004 30666 13032 31418
rect 12992 30660 13044 30666
rect 12992 30602 13044 30608
rect 12898 29064 12954 29073
rect 12898 28999 12900 29008
rect 12952 28999 12954 29008
rect 12900 28970 12952 28976
rect 12900 26784 12952 26790
rect 12900 26726 12952 26732
rect 12912 26586 12940 26726
rect 12900 26580 12952 26586
rect 12900 26522 12952 26528
rect 12992 25696 13044 25702
rect 12992 25638 13044 25644
rect 13004 25498 13032 25638
rect 12992 25492 13044 25498
rect 12992 25434 13044 25440
rect 12820 25214 12940 25242
rect 12808 25152 12860 25158
rect 12808 25094 12860 25100
rect 12820 24954 12848 25094
rect 12808 24948 12860 24954
rect 12808 24890 12860 24896
rect 12716 24268 12768 24274
rect 12716 24210 12768 24216
rect 12624 24064 12676 24070
rect 12624 24006 12676 24012
rect 12636 23497 12664 24006
rect 12728 23730 12756 24210
rect 12912 23866 12940 25214
rect 12990 24712 13046 24721
rect 12990 24647 13046 24656
rect 13004 24274 13032 24647
rect 12992 24268 13044 24274
rect 12992 24210 13044 24216
rect 12900 23860 12952 23866
rect 12900 23802 12952 23808
rect 13096 23730 13124 31855
rect 13188 31754 13216 33594
rect 13372 33590 13400 33798
rect 13360 33584 13412 33590
rect 13360 33526 13412 33532
rect 13176 31748 13228 31754
rect 13176 31690 13228 31696
rect 13188 30666 13216 31690
rect 13372 31482 13400 33526
rect 13464 31482 13492 38286
rect 13648 38010 13676 38422
rect 13636 38004 13688 38010
rect 13636 37946 13688 37952
rect 13820 37868 13872 37874
rect 13820 37810 13872 37816
rect 13728 36576 13780 36582
rect 13728 36518 13780 36524
rect 13740 36156 13768 36518
rect 13832 36378 13860 37810
rect 13820 36372 13872 36378
rect 13820 36314 13872 36320
rect 13820 36168 13872 36174
rect 13740 36128 13820 36156
rect 13820 36110 13872 36116
rect 13820 36032 13872 36038
rect 13820 35974 13872 35980
rect 13832 35698 13860 35974
rect 13728 35692 13780 35698
rect 13728 35634 13780 35640
rect 13820 35692 13872 35698
rect 13820 35634 13872 35640
rect 13636 34468 13688 34474
rect 13636 34410 13688 34416
rect 13648 34066 13676 34410
rect 13636 34060 13688 34066
rect 13636 34002 13688 34008
rect 13740 33862 13768 35634
rect 13728 33856 13780 33862
rect 13728 33798 13780 33804
rect 13636 31816 13688 31822
rect 13636 31758 13688 31764
rect 13360 31476 13412 31482
rect 13360 31418 13412 31424
rect 13452 31476 13504 31482
rect 13452 31418 13504 31424
rect 13360 31272 13412 31278
rect 13360 31214 13412 31220
rect 13372 30938 13400 31214
rect 13360 30932 13412 30938
rect 13360 30874 13412 30880
rect 13176 30660 13228 30666
rect 13176 30602 13228 30608
rect 13360 30592 13412 30598
rect 13360 30534 13412 30540
rect 13176 29504 13228 29510
rect 13176 29446 13228 29452
rect 13268 29504 13320 29510
rect 13268 29446 13320 29452
rect 13188 29034 13216 29446
rect 13176 29028 13228 29034
rect 13176 28970 13228 28976
rect 13176 27668 13228 27674
rect 13176 27610 13228 27616
rect 13188 25294 13216 27610
rect 13176 25288 13228 25294
rect 13176 25230 13228 25236
rect 13176 24608 13228 24614
rect 13176 24550 13228 24556
rect 12716 23724 12768 23730
rect 12716 23666 12768 23672
rect 12900 23724 12952 23730
rect 12900 23666 12952 23672
rect 13084 23724 13136 23730
rect 13084 23666 13136 23672
rect 12808 23520 12860 23526
rect 12622 23488 12678 23497
rect 12808 23462 12860 23468
rect 12622 23423 12678 23432
rect 12440 22772 12492 22778
rect 12440 22714 12492 22720
rect 12532 22772 12584 22778
rect 12532 22714 12584 22720
rect 12624 22636 12676 22642
rect 12624 22578 12676 22584
rect 11980 22568 12032 22574
rect 11980 22510 12032 22516
rect 12072 22568 12124 22574
rect 12072 22510 12124 22516
rect 11992 22234 12020 22510
rect 11980 22228 12032 22234
rect 11980 22170 12032 22176
rect 12084 22098 12112 22510
rect 12072 22092 12124 22098
rect 12636 22094 12664 22578
rect 12636 22066 12756 22094
rect 12072 22034 12124 22040
rect 12440 21956 12492 21962
rect 12440 21898 12492 21904
rect 11612 21888 11664 21894
rect 11612 21830 11664 21836
rect 11704 21888 11756 21894
rect 11704 21830 11756 21836
rect 11796 21888 11848 21894
rect 11796 21830 11848 21836
rect 12164 21888 12216 21894
rect 12164 21830 12216 21836
rect 11624 21350 11652 21830
rect 11612 21344 11664 21350
rect 11612 21286 11664 21292
rect 11440 20998 11560 21026
rect 11440 20262 11468 20998
rect 11520 20936 11572 20942
rect 11520 20878 11572 20884
rect 11428 20256 11480 20262
rect 11428 20198 11480 20204
rect 11440 19854 11468 20198
rect 11428 19848 11480 19854
rect 11428 19790 11480 19796
rect 11428 19712 11480 19718
rect 11428 19654 11480 19660
rect 11336 19168 11388 19174
rect 11336 19110 11388 19116
rect 11348 18834 11376 19110
rect 11336 18828 11388 18834
rect 11336 18770 11388 18776
rect 11348 18290 11376 18770
rect 11440 18766 11468 19654
rect 11532 19378 11560 20878
rect 11612 20392 11664 20398
rect 11612 20334 11664 20340
rect 11624 20058 11652 20334
rect 11612 20052 11664 20058
rect 11612 19994 11664 20000
rect 11520 19372 11572 19378
rect 11520 19314 11572 19320
rect 11428 18760 11480 18766
rect 11428 18702 11480 18708
rect 11336 18284 11388 18290
rect 11336 18226 11388 18232
rect 11428 18216 11480 18222
rect 11428 18158 11480 18164
rect 11440 17882 11468 18158
rect 11532 18086 11560 19314
rect 11520 18080 11572 18086
rect 11520 18022 11572 18028
rect 11428 17876 11480 17882
rect 11428 17818 11480 17824
rect 11624 17678 11652 19994
rect 11716 18442 11744 21830
rect 11808 19990 11836 21830
rect 11886 21584 11942 21593
rect 11886 21519 11888 21528
rect 11940 21519 11942 21528
rect 11888 21490 11940 21496
rect 12176 21486 12204 21830
rect 11980 21480 12032 21486
rect 11980 21422 12032 21428
rect 12164 21480 12216 21486
rect 12164 21422 12216 21428
rect 11992 20466 12020 21422
rect 12176 20806 12204 21422
rect 12164 20800 12216 20806
rect 12164 20742 12216 20748
rect 12452 20641 12480 21898
rect 12624 21888 12676 21894
rect 12624 21830 12676 21836
rect 12438 20632 12494 20641
rect 12438 20567 12494 20576
rect 11980 20460 12032 20466
rect 11980 20402 12032 20408
rect 11888 20256 11940 20262
rect 11888 20198 11940 20204
rect 12164 20256 12216 20262
rect 12164 20198 12216 20204
rect 11796 19984 11848 19990
rect 11796 19926 11848 19932
rect 11796 19712 11848 19718
rect 11796 19654 11848 19660
rect 11808 19514 11836 19654
rect 11796 19508 11848 19514
rect 11796 19450 11848 19456
rect 11796 19372 11848 19378
rect 11796 19314 11848 19320
rect 11808 18766 11836 19314
rect 11900 19310 11928 20198
rect 12176 20058 12204 20198
rect 12164 20052 12216 20058
rect 12164 19994 12216 20000
rect 11980 19848 12032 19854
rect 11980 19790 12032 19796
rect 11888 19304 11940 19310
rect 11888 19246 11940 19252
rect 11888 19168 11940 19174
rect 11888 19110 11940 19116
rect 11900 18766 11928 19110
rect 11796 18760 11848 18766
rect 11796 18702 11848 18708
rect 11888 18760 11940 18766
rect 11888 18702 11940 18708
rect 11716 18414 11836 18442
rect 11702 17912 11758 17921
rect 11702 17847 11758 17856
rect 11716 17746 11744 17847
rect 11704 17740 11756 17746
rect 11704 17682 11756 17688
rect 11612 17672 11664 17678
rect 11256 17598 11468 17626
rect 11612 17614 11664 17620
rect 11702 17640 11758 17649
rect 11152 17128 11204 17134
rect 11152 17070 11204 17076
rect 11244 16516 11296 16522
rect 11244 16458 11296 16464
rect 11060 16448 11112 16454
rect 11060 16390 11112 16396
rect 11072 16182 11100 16390
rect 11256 16250 11284 16458
rect 11244 16244 11296 16250
rect 11244 16186 11296 16192
rect 11060 16176 11112 16182
rect 11060 16118 11112 16124
rect 11244 15564 11296 15570
rect 11244 15506 11296 15512
rect 11152 15496 11204 15502
rect 11152 15438 11204 15444
rect 11060 15088 11112 15094
rect 11060 15030 11112 15036
rect 10968 13796 11020 13802
rect 10968 13738 11020 13744
rect 10428 12406 10548 12434
rect 10324 11688 10376 11694
rect 10324 11630 10376 11636
rect 10324 11552 10376 11558
rect 10324 11494 10376 11500
rect 10336 11354 10364 11494
rect 10324 11348 10376 11354
rect 10324 11290 10376 11296
rect 10232 10600 10284 10606
rect 10232 10542 10284 10548
rect 9864 8628 9916 8634
rect 9864 8570 9916 8576
rect 10140 8628 10192 8634
rect 10140 8570 10192 8576
rect 10244 8514 10272 10542
rect 10152 8486 10272 8514
rect 9692 8452 9904 8480
rect 9600 8350 9720 8378
rect 9692 7750 9720 8350
rect 9876 8090 9904 8452
rect 9864 8084 9916 8090
rect 9864 8026 9916 8032
rect 9680 7744 9732 7750
rect 9680 7686 9732 7692
rect 9772 7744 9824 7750
rect 9772 7686 9824 7692
rect 9784 7546 9812 7686
rect 9876 7546 9904 8026
rect 9772 7540 9824 7546
rect 9772 7482 9824 7488
rect 9864 7540 9916 7546
rect 9864 7482 9916 7488
rect 9496 6792 9548 6798
rect 9496 6734 9548 6740
rect 9036 6656 9088 6662
rect 9036 6598 9088 6604
rect 9048 5234 9076 6598
rect 9508 6458 9536 6734
rect 9496 6452 9548 6458
rect 9496 6394 9548 6400
rect 9404 6384 9456 6390
rect 9404 6326 9456 6332
rect 9312 6248 9364 6254
rect 9312 6190 9364 6196
rect 9324 5914 9352 6190
rect 9312 5908 9364 5914
rect 9312 5850 9364 5856
rect 9416 5710 9444 6326
rect 9772 6248 9824 6254
rect 9772 6190 9824 6196
rect 9496 6112 9548 6118
rect 9496 6054 9548 6060
rect 9508 5710 9536 6054
rect 9680 5840 9732 5846
rect 9680 5782 9732 5788
rect 9404 5704 9456 5710
rect 9404 5646 9456 5652
rect 9496 5704 9548 5710
rect 9496 5646 9548 5652
rect 9036 5228 9088 5234
rect 9036 5170 9088 5176
rect 9692 5166 9720 5782
rect 9784 5710 9812 6190
rect 9772 5704 9824 5710
rect 9772 5646 9824 5652
rect 9680 5160 9732 5166
rect 9680 5102 9732 5108
rect 9128 5024 9180 5030
rect 9128 4966 9180 4972
rect 9140 4282 9168 4966
rect 9692 4282 9720 5102
rect 9784 4622 9812 5646
rect 9864 5568 9916 5574
rect 9864 5510 9916 5516
rect 10048 5568 10100 5574
rect 10048 5510 10100 5516
rect 9876 5370 9904 5510
rect 9864 5364 9916 5370
rect 9864 5306 9916 5312
rect 10060 5234 10088 5510
rect 9864 5228 9916 5234
rect 9864 5170 9916 5176
rect 10048 5228 10100 5234
rect 10048 5170 10100 5176
rect 9876 4826 9904 5170
rect 9864 4820 9916 4826
rect 9864 4762 9916 4768
rect 9772 4616 9824 4622
rect 9772 4558 9824 4564
rect 9128 4276 9180 4282
rect 9128 4218 9180 4224
rect 9680 4276 9732 4282
rect 9680 4218 9732 4224
rect 10152 2650 10180 8486
rect 10428 8430 10456 12406
rect 11072 11830 11100 15030
rect 11164 14414 11192 15438
rect 11152 14408 11204 14414
rect 11152 14350 11204 14356
rect 11256 13530 11284 15506
rect 11440 15502 11468 17598
rect 11624 17338 11652 17614
rect 11702 17575 11704 17584
rect 11756 17575 11758 17584
rect 11704 17546 11756 17552
rect 11612 17332 11664 17338
rect 11612 17274 11664 17280
rect 11808 17202 11836 18414
rect 11900 17921 11928 18702
rect 11886 17912 11942 17921
rect 11886 17847 11942 17856
rect 11992 17762 12020 19790
rect 12176 19786 12204 19994
rect 12440 19848 12492 19854
rect 12440 19790 12492 19796
rect 12164 19780 12216 19786
rect 12164 19722 12216 19728
rect 12452 19446 12480 19790
rect 12532 19780 12584 19786
rect 12532 19722 12584 19728
rect 12544 19553 12572 19722
rect 12530 19544 12586 19553
rect 12530 19479 12586 19488
rect 12440 19440 12492 19446
rect 12440 19382 12492 19388
rect 12452 19334 12480 19382
rect 12544 19378 12572 19479
rect 12072 19304 12124 19310
rect 12072 19246 12124 19252
rect 12360 19306 12480 19334
rect 12532 19372 12584 19378
rect 12532 19314 12584 19320
rect 12084 18766 12112 19246
rect 12360 19242 12388 19306
rect 12348 19236 12400 19242
rect 12348 19178 12400 19184
rect 12256 19168 12308 19174
rect 12256 19110 12308 19116
rect 12072 18760 12124 18766
rect 12072 18702 12124 18708
rect 12084 18222 12112 18702
rect 12162 18592 12218 18601
rect 12162 18527 12218 18536
rect 12072 18216 12124 18222
rect 12072 18158 12124 18164
rect 12072 18080 12124 18086
rect 12072 18022 12124 18028
rect 11900 17734 12020 17762
rect 11900 17218 11928 17734
rect 11980 17604 12032 17610
rect 11980 17546 12032 17552
rect 11992 17338 12020 17546
rect 11980 17332 12032 17338
rect 11980 17274 12032 17280
rect 11796 17196 11848 17202
rect 11900 17190 12020 17218
rect 11796 17138 11848 17144
rect 11808 16998 11836 17138
rect 11796 16992 11848 16998
rect 11796 16934 11848 16940
rect 11428 15496 11480 15502
rect 11426 15464 11428 15473
rect 11888 15496 11940 15502
rect 11480 15464 11482 15473
rect 11888 15438 11940 15444
rect 11426 15399 11482 15408
rect 11612 15428 11664 15434
rect 11612 15370 11664 15376
rect 11244 13524 11296 13530
rect 11244 13466 11296 13472
rect 11152 13252 11204 13258
rect 11152 13194 11204 13200
rect 11164 12442 11192 13194
rect 11152 12436 11204 12442
rect 11152 12378 11204 12384
rect 11060 11824 11112 11830
rect 11060 11766 11112 11772
rect 10784 11756 10836 11762
rect 10784 11698 10836 11704
rect 10796 11218 10824 11698
rect 10876 11688 10928 11694
rect 10876 11630 10928 11636
rect 10784 11212 10836 11218
rect 10784 11154 10836 11160
rect 10796 10674 10824 11154
rect 10784 10668 10836 10674
rect 10784 10610 10836 10616
rect 10508 10260 10560 10266
rect 10508 10202 10560 10208
rect 10520 9586 10548 10202
rect 10508 9580 10560 9586
rect 10508 9522 10560 9528
rect 10888 9518 10916 11630
rect 11256 10606 11284 13466
rect 11520 10668 11572 10674
rect 11520 10610 11572 10616
rect 11244 10600 11296 10606
rect 11244 10542 11296 10548
rect 11532 10062 11560 10610
rect 11428 10056 11480 10062
rect 11428 9998 11480 10004
rect 11520 10056 11572 10062
rect 11520 9998 11572 10004
rect 11440 9722 11468 9998
rect 11428 9716 11480 9722
rect 11428 9658 11480 9664
rect 11624 9586 11652 15370
rect 11704 14408 11756 14414
rect 11704 14350 11756 14356
rect 11716 13258 11744 14350
rect 11900 13394 11928 15438
rect 11888 13388 11940 13394
rect 11888 13330 11940 13336
rect 11704 13252 11756 13258
rect 11704 13194 11756 13200
rect 11716 11150 11744 13194
rect 11900 12918 11928 13330
rect 11888 12912 11940 12918
rect 11888 12854 11940 12860
rect 11900 11762 11928 12854
rect 11992 12434 12020 17190
rect 12084 17134 12112 18022
rect 12072 17128 12124 17134
rect 12072 17070 12124 17076
rect 12176 16046 12204 18527
rect 12268 18358 12296 19110
rect 12256 18352 12308 18358
rect 12256 18294 12308 18300
rect 12532 18284 12584 18290
rect 12532 18226 12584 18232
rect 12544 17882 12572 18226
rect 12440 17876 12492 17882
rect 12440 17818 12492 17824
rect 12532 17876 12584 17882
rect 12532 17818 12584 17824
rect 12254 17776 12310 17785
rect 12254 17711 12256 17720
rect 12308 17711 12310 17720
rect 12256 17682 12308 17688
rect 12348 17672 12400 17678
rect 12348 17614 12400 17620
rect 12360 17338 12388 17614
rect 12452 17338 12480 17818
rect 12544 17649 12572 17818
rect 12530 17640 12586 17649
rect 12530 17575 12586 17584
rect 12348 17332 12400 17338
rect 12348 17274 12400 17280
rect 12440 17332 12492 17338
rect 12440 17274 12492 17280
rect 12544 17202 12572 17575
rect 12532 17196 12584 17202
rect 12532 17138 12584 17144
rect 12256 16448 12308 16454
rect 12256 16390 12308 16396
rect 12268 16114 12296 16390
rect 12636 16182 12664 21830
rect 12728 18465 12756 22066
rect 12820 22030 12848 23462
rect 12808 22024 12860 22030
rect 12808 21966 12860 21972
rect 12808 21480 12860 21486
rect 12808 21422 12860 21428
rect 12714 18456 12770 18465
rect 12714 18391 12770 18400
rect 12716 18080 12768 18086
rect 12716 18022 12768 18028
rect 12728 17814 12756 18022
rect 12716 17808 12768 17814
rect 12716 17750 12768 17756
rect 12716 17672 12768 17678
rect 12716 17614 12768 17620
rect 12728 17338 12756 17614
rect 12716 17332 12768 17338
rect 12716 17274 12768 17280
rect 12624 16176 12676 16182
rect 12346 16144 12402 16153
rect 12256 16108 12308 16114
rect 12624 16118 12676 16124
rect 12346 16079 12348 16088
rect 12256 16050 12308 16056
rect 12400 16079 12402 16088
rect 12348 16050 12400 16056
rect 12164 16040 12216 16046
rect 12268 16017 12296 16050
rect 12532 16040 12584 16046
rect 12164 15982 12216 15988
rect 12254 16008 12310 16017
rect 12532 15982 12584 15988
rect 12254 15943 12310 15952
rect 12544 15881 12572 15982
rect 12530 15872 12586 15881
rect 12530 15807 12586 15816
rect 12544 15706 12572 15807
rect 12532 15700 12584 15706
rect 12532 15642 12584 15648
rect 12440 15428 12492 15434
rect 12440 15370 12492 15376
rect 12452 15162 12480 15370
rect 12440 15156 12492 15162
rect 12440 15098 12492 15104
rect 12072 15088 12124 15094
rect 12072 15030 12124 15036
rect 12084 14482 12112 15030
rect 12532 14952 12584 14958
rect 12532 14894 12584 14900
rect 12256 14884 12308 14890
rect 12256 14826 12308 14832
rect 12072 14476 12124 14482
rect 12072 14418 12124 14424
rect 12268 12782 12296 14826
rect 12544 14482 12572 14894
rect 12532 14476 12584 14482
rect 12532 14418 12584 14424
rect 12440 13932 12492 13938
rect 12440 13874 12492 13880
rect 12256 12776 12308 12782
rect 12256 12718 12308 12724
rect 11992 12406 12112 12434
rect 11888 11756 11940 11762
rect 11888 11698 11940 11704
rect 11980 11756 12032 11762
rect 11980 11698 12032 11704
rect 11992 11354 12020 11698
rect 11980 11348 12032 11354
rect 11980 11290 12032 11296
rect 11704 11144 11756 11150
rect 11704 11086 11756 11092
rect 11612 9580 11664 9586
rect 11612 9522 11664 9528
rect 10876 9512 10928 9518
rect 10876 9454 10928 9460
rect 10508 9376 10560 9382
rect 10508 9318 10560 9324
rect 10520 9042 10548 9318
rect 10508 9036 10560 9042
rect 10508 8978 10560 8984
rect 10416 8424 10468 8430
rect 10416 8366 10468 8372
rect 10600 8424 10652 8430
rect 10600 8366 10652 8372
rect 10612 7954 10640 8366
rect 10600 7948 10652 7954
rect 10600 7890 10652 7896
rect 10888 7886 10916 9454
rect 11624 9178 11652 9522
rect 11612 9172 11664 9178
rect 11612 9114 11664 9120
rect 11716 8974 11744 11086
rect 11704 8968 11756 8974
rect 11704 8910 11756 8916
rect 11060 8832 11112 8838
rect 11060 8774 11112 8780
rect 10876 7880 10928 7886
rect 10876 7822 10928 7828
rect 10692 6792 10744 6798
rect 10692 6734 10744 6740
rect 10232 6316 10284 6322
rect 10232 6258 10284 6264
rect 10244 4622 10272 6258
rect 10704 5846 10732 6734
rect 11072 6390 11100 8774
rect 11152 8492 11204 8498
rect 11152 8434 11204 8440
rect 11796 8492 11848 8498
rect 11796 8434 11848 8440
rect 11164 7206 11192 8434
rect 11808 7478 11836 8434
rect 12084 7478 12112 12406
rect 12268 12238 12296 12718
rect 12256 12232 12308 12238
rect 12256 12174 12308 12180
rect 12256 11688 12308 11694
rect 12256 11630 12308 11636
rect 12268 10674 12296 11630
rect 12452 11150 12480 13874
rect 12544 13394 12572 14418
rect 12532 13388 12584 13394
rect 12532 13330 12584 13336
rect 12544 12306 12572 13330
rect 12716 13184 12768 13190
rect 12716 13126 12768 13132
rect 12728 12850 12756 13126
rect 12716 12844 12768 12850
rect 12716 12786 12768 12792
rect 12532 12300 12584 12306
rect 12532 12242 12584 12248
rect 12544 11218 12572 12242
rect 12532 11212 12584 11218
rect 12532 11154 12584 11160
rect 12440 11144 12492 11150
rect 12440 11086 12492 11092
rect 12256 10668 12308 10674
rect 12256 10610 12308 10616
rect 12268 8430 12296 10610
rect 12544 9518 12572 11154
rect 12532 9512 12584 9518
rect 12532 9454 12584 9460
rect 12544 9194 12572 9454
rect 12544 9166 12664 9194
rect 12636 8566 12664 9166
rect 12716 8968 12768 8974
rect 12716 8910 12768 8916
rect 12728 8634 12756 8910
rect 12716 8628 12768 8634
rect 12716 8570 12768 8576
rect 12624 8560 12676 8566
rect 12624 8502 12676 8508
rect 12348 8492 12400 8498
rect 12532 8492 12584 8498
rect 12400 8452 12480 8480
rect 12348 8434 12400 8440
rect 12256 8424 12308 8430
rect 12256 8366 12308 8372
rect 12268 7954 12296 8366
rect 12256 7948 12308 7954
rect 12256 7890 12308 7896
rect 11796 7472 11848 7478
rect 11796 7414 11848 7420
rect 12072 7472 12124 7478
rect 12072 7414 12124 7420
rect 11888 7336 11940 7342
rect 11888 7278 11940 7284
rect 11152 7200 11204 7206
rect 11152 7142 11204 7148
rect 11164 6934 11192 7142
rect 11152 6928 11204 6934
rect 11152 6870 11204 6876
rect 11060 6384 11112 6390
rect 11060 6326 11112 6332
rect 10784 5908 10836 5914
rect 10784 5850 10836 5856
rect 10692 5840 10744 5846
rect 10692 5782 10744 5788
rect 10704 5710 10732 5782
rect 10692 5704 10744 5710
rect 10692 5646 10744 5652
rect 10416 5636 10468 5642
rect 10416 5578 10468 5584
rect 10428 5302 10456 5578
rect 10692 5568 10744 5574
rect 10796 5556 10824 5850
rect 10744 5528 10824 5556
rect 11704 5568 11756 5574
rect 10692 5510 10744 5516
rect 11704 5510 11756 5516
rect 11716 5302 11744 5510
rect 11900 5370 11928 7278
rect 12084 7018 12112 7414
rect 12268 7342 12296 7890
rect 12348 7812 12400 7818
rect 12452 7800 12480 8452
rect 12532 8434 12584 8440
rect 12544 8090 12572 8434
rect 12532 8084 12584 8090
rect 12532 8026 12584 8032
rect 12532 7812 12584 7818
rect 12452 7772 12532 7800
rect 12348 7754 12400 7760
rect 12532 7754 12584 7760
rect 12256 7336 12308 7342
rect 12256 7278 12308 7284
rect 12084 6990 12296 7018
rect 12360 7002 12388 7754
rect 12820 7410 12848 21422
rect 12912 19990 12940 23666
rect 13188 22094 13216 24550
rect 13004 22066 13216 22094
rect 12900 19984 12952 19990
rect 12900 19926 12952 19932
rect 12898 19544 12954 19553
rect 12898 19479 12954 19488
rect 12912 17814 12940 19479
rect 12900 17808 12952 17814
rect 12900 17750 12952 17756
rect 12912 15094 12940 17750
rect 13004 16794 13032 22066
rect 13176 20528 13228 20534
rect 13176 20470 13228 20476
rect 13188 19514 13216 20470
rect 13176 19508 13228 19514
rect 13096 19468 13176 19496
rect 12992 16788 13044 16794
rect 12992 16730 13044 16736
rect 13096 16522 13124 19468
rect 13176 19450 13228 19456
rect 13280 17218 13308 29446
rect 13372 28218 13400 30534
rect 13464 30394 13492 31418
rect 13544 31136 13596 31142
rect 13544 31078 13596 31084
rect 13452 30388 13504 30394
rect 13452 30330 13504 30336
rect 13556 29646 13584 31078
rect 13648 30938 13676 31758
rect 13636 30932 13688 30938
rect 13636 30874 13688 30880
rect 13740 30666 13768 33798
rect 13912 31680 13964 31686
rect 13912 31622 13964 31628
rect 13728 30660 13780 30666
rect 13728 30602 13780 30608
rect 13636 30592 13688 30598
rect 13636 30534 13688 30540
rect 13648 30394 13676 30534
rect 13636 30388 13688 30394
rect 13636 30330 13688 30336
rect 13728 30048 13780 30054
rect 13728 29990 13780 29996
rect 13544 29640 13596 29646
rect 13544 29582 13596 29588
rect 13740 29102 13768 29990
rect 13820 29640 13872 29646
rect 13820 29582 13872 29588
rect 13728 29096 13780 29102
rect 13728 29038 13780 29044
rect 13360 28212 13412 28218
rect 13360 28154 13412 28160
rect 13372 27334 13400 28154
rect 13452 28076 13504 28082
rect 13452 28018 13504 28024
rect 13464 27470 13492 28018
rect 13636 27872 13688 27878
rect 13636 27814 13688 27820
rect 13452 27464 13504 27470
rect 13452 27406 13504 27412
rect 13360 27328 13412 27334
rect 13360 27270 13412 27276
rect 13464 24818 13492 27406
rect 13542 26616 13598 26625
rect 13542 26551 13598 26560
rect 13556 25838 13584 26551
rect 13648 26382 13676 27814
rect 13740 27538 13768 29038
rect 13728 27532 13780 27538
rect 13728 27474 13780 27480
rect 13832 26382 13860 29582
rect 13924 28218 13952 31622
rect 13912 28212 13964 28218
rect 13912 28154 13964 28160
rect 13912 27600 13964 27606
rect 13912 27542 13964 27548
rect 13636 26376 13688 26382
rect 13636 26318 13688 26324
rect 13820 26376 13872 26382
rect 13820 26318 13872 26324
rect 13924 25945 13952 27542
rect 13910 25936 13966 25945
rect 13820 25900 13872 25906
rect 13910 25871 13966 25880
rect 13820 25842 13872 25848
rect 13544 25832 13596 25838
rect 13544 25774 13596 25780
rect 13556 25294 13584 25774
rect 13728 25356 13780 25362
rect 13728 25298 13780 25304
rect 13544 25288 13596 25294
rect 13544 25230 13596 25236
rect 13452 24812 13504 24818
rect 13452 24754 13504 24760
rect 13556 23798 13584 25230
rect 13740 24954 13768 25298
rect 13728 24948 13780 24954
rect 13728 24890 13780 24896
rect 13544 23792 13596 23798
rect 13544 23734 13596 23740
rect 13726 23624 13782 23633
rect 13726 23559 13782 23568
rect 13740 23526 13768 23559
rect 13728 23520 13780 23526
rect 13728 23462 13780 23468
rect 13544 22636 13596 22642
rect 13544 22578 13596 22584
rect 13556 22030 13584 22578
rect 13544 22024 13596 22030
rect 13544 21966 13596 21972
rect 13542 21448 13598 21457
rect 13542 21383 13598 21392
rect 13556 19854 13584 21383
rect 13636 20596 13688 20602
rect 13636 20538 13688 20544
rect 13648 20233 13676 20538
rect 13634 20224 13690 20233
rect 13634 20159 13690 20168
rect 13544 19848 13596 19854
rect 13544 19790 13596 19796
rect 13452 19780 13504 19786
rect 13452 19722 13504 19728
rect 13360 19712 13412 19718
rect 13360 19654 13412 19660
rect 13372 19378 13400 19654
rect 13360 19372 13412 19378
rect 13360 19314 13412 19320
rect 13358 17912 13414 17921
rect 13358 17847 13360 17856
rect 13412 17847 13414 17856
rect 13360 17818 13412 17824
rect 13188 17190 13308 17218
rect 13084 16516 13136 16522
rect 13084 16458 13136 16464
rect 12900 15088 12952 15094
rect 12900 15030 12952 15036
rect 12992 15020 13044 15026
rect 12992 14962 13044 14968
rect 13004 14006 13032 14962
rect 12992 14000 13044 14006
rect 12992 13942 13044 13948
rect 13096 13326 13124 16458
rect 13084 13320 13136 13326
rect 13084 13262 13136 13268
rect 12992 11824 13044 11830
rect 12992 11766 13044 11772
rect 12900 11688 12952 11694
rect 12900 11630 12952 11636
rect 12912 11082 12940 11630
rect 12900 11076 12952 11082
rect 12900 11018 12952 11024
rect 13004 9994 13032 11766
rect 13096 10266 13124 13262
rect 13084 10260 13136 10266
rect 13084 10202 13136 10208
rect 13188 10130 13216 17190
rect 13360 15020 13412 15026
rect 13360 14962 13412 14968
rect 13268 14000 13320 14006
rect 13268 13942 13320 13948
rect 13280 10130 13308 13942
rect 13372 13938 13400 14962
rect 13360 13932 13412 13938
rect 13360 13874 13412 13880
rect 13372 13190 13400 13874
rect 13360 13184 13412 13190
rect 13360 13126 13412 13132
rect 13360 11144 13412 11150
rect 13360 11086 13412 11092
rect 13176 10124 13228 10130
rect 13176 10066 13228 10072
rect 13268 10124 13320 10130
rect 13268 10066 13320 10072
rect 12992 9988 13044 9994
rect 12992 9930 13044 9936
rect 13188 9722 13216 10066
rect 13176 9716 13228 9722
rect 13176 9658 13228 9664
rect 13280 9586 13308 10066
rect 13268 9580 13320 9586
rect 13268 9522 13320 9528
rect 13084 9376 13136 9382
rect 13084 9318 13136 9324
rect 13096 9178 13124 9318
rect 13084 9172 13136 9178
rect 13084 9114 13136 9120
rect 13372 8974 13400 11086
rect 13464 10062 13492 19722
rect 13544 19712 13596 19718
rect 13544 19654 13596 19660
rect 13556 19553 13584 19654
rect 13542 19544 13598 19553
rect 13542 19479 13598 19488
rect 13648 19174 13676 20159
rect 13728 19848 13780 19854
rect 13728 19790 13780 19796
rect 13636 19168 13688 19174
rect 13636 19110 13688 19116
rect 13740 17542 13768 19790
rect 13832 18426 13860 25842
rect 13910 23488 13966 23497
rect 13910 23423 13966 23432
rect 13924 23186 13952 23423
rect 14016 23202 14044 38830
rect 15568 38820 15620 38826
rect 15568 38762 15620 38768
rect 15580 38729 15608 38762
rect 15566 38720 15622 38729
rect 15566 38655 15622 38664
rect 17972 38554 18000 38898
rect 17960 38548 18012 38554
rect 17960 38490 18012 38496
rect 18512 38344 18564 38350
rect 18512 38286 18564 38292
rect 18524 38010 18552 38286
rect 19444 38010 19472 38898
rect 19616 38752 19668 38758
rect 22388 38729 22416 38898
rect 27080 38729 27108 38898
rect 27620 38752 27672 38758
rect 19616 38694 19668 38700
rect 22374 38720 22430 38729
rect 19628 38418 19656 38694
rect 22374 38655 22430 38664
rect 27066 38720 27122 38729
rect 27620 38694 27672 38700
rect 27066 38655 27122 38664
rect 22468 38548 22520 38554
rect 22468 38490 22520 38496
rect 19616 38412 19668 38418
rect 19616 38354 19668 38360
rect 21180 38344 21232 38350
rect 21180 38286 21232 38292
rect 21272 38344 21324 38350
rect 21272 38286 21324 38292
rect 20996 38208 21048 38214
rect 20996 38150 21048 38156
rect 21008 38010 21036 38150
rect 18512 38004 18564 38010
rect 18512 37946 18564 37952
rect 19432 38004 19484 38010
rect 19432 37946 19484 37952
rect 20996 38004 21048 38010
rect 20996 37946 21048 37952
rect 16948 37936 17000 37942
rect 20536 37936 20588 37942
rect 16948 37878 17000 37884
rect 14096 37868 14148 37874
rect 14096 37810 14148 37816
rect 14372 37868 14424 37874
rect 15292 37868 15344 37874
rect 14424 37828 14780 37856
rect 14372 37810 14424 37816
rect 14108 36582 14136 37810
rect 14096 36576 14148 36582
rect 14096 36518 14148 36524
rect 14280 36168 14332 36174
rect 14280 36110 14332 36116
rect 14292 35834 14320 36110
rect 14464 36032 14516 36038
rect 14464 35974 14516 35980
rect 14280 35828 14332 35834
rect 14280 35770 14332 35776
rect 14476 33998 14504 35974
rect 14648 34196 14700 34202
rect 14648 34138 14700 34144
rect 14464 33992 14516 33998
rect 14464 33934 14516 33940
rect 14660 33658 14688 34138
rect 14648 33652 14700 33658
rect 14648 33594 14700 33600
rect 14752 33522 14780 37828
rect 15292 37810 15344 37816
rect 15936 37868 15988 37874
rect 15936 37810 15988 37816
rect 16120 37868 16172 37874
rect 16120 37810 16172 37816
rect 16212 37868 16264 37874
rect 16396 37868 16448 37874
rect 16212 37810 16264 37816
rect 16316 37828 16396 37856
rect 14832 36576 14884 36582
rect 14832 36518 14884 36524
rect 14844 36242 14872 36518
rect 14832 36236 14884 36242
rect 14832 36178 14884 36184
rect 14844 34202 14872 36178
rect 15200 36168 15252 36174
rect 15200 36110 15252 36116
rect 14832 34196 14884 34202
rect 14832 34138 14884 34144
rect 14372 33516 14424 33522
rect 14372 33458 14424 33464
rect 14740 33516 14792 33522
rect 14740 33458 14792 33464
rect 14384 31686 14412 33458
rect 14556 31748 14608 31754
rect 14556 31690 14608 31696
rect 14372 31680 14424 31686
rect 14372 31622 14424 31628
rect 14568 30938 14596 31690
rect 14648 31136 14700 31142
rect 14648 31078 14700 31084
rect 14556 30932 14608 30938
rect 14556 30874 14608 30880
rect 14660 30734 14688 31078
rect 14752 30734 14780 33458
rect 14464 30728 14516 30734
rect 14464 30670 14516 30676
rect 14648 30728 14700 30734
rect 14648 30670 14700 30676
rect 14740 30728 14792 30734
rect 14740 30670 14792 30676
rect 14476 30598 14504 30670
rect 14096 30592 14148 30598
rect 14096 30534 14148 30540
rect 14372 30592 14424 30598
rect 14372 30534 14424 30540
rect 14464 30592 14516 30598
rect 14464 30534 14516 30540
rect 14108 29646 14136 30534
rect 14280 30116 14332 30122
rect 14280 30058 14332 30064
rect 14096 29640 14148 29646
rect 14096 29582 14148 29588
rect 14096 28144 14148 28150
rect 14096 28086 14148 28092
rect 14108 27606 14136 28086
rect 14188 27872 14240 27878
rect 14188 27814 14240 27820
rect 14200 27674 14228 27814
rect 14188 27668 14240 27674
rect 14188 27610 14240 27616
rect 14096 27600 14148 27606
rect 14096 27542 14148 27548
rect 14292 27418 14320 30058
rect 14384 27470 14412 30534
rect 14476 27878 14504 30534
rect 14556 30388 14608 30394
rect 14556 30330 14608 30336
rect 14568 28082 14596 30330
rect 14752 30122 14780 30670
rect 14844 30598 14872 34138
rect 15016 34128 15068 34134
rect 15016 34070 15068 34076
rect 14924 33856 14976 33862
rect 14924 33798 14976 33804
rect 14936 31634 14964 33798
rect 15028 33697 15056 34070
rect 15014 33688 15070 33697
rect 15014 33623 15070 33632
rect 15212 33561 15240 36110
rect 15304 36038 15332 37810
rect 15384 37732 15436 37738
rect 15384 37674 15436 37680
rect 15292 36032 15344 36038
rect 15292 35974 15344 35980
rect 15198 33552 15254 33561
rect 15198 33487 15254 33496
rect 14936 31606 15056 31634
rect 14832 30592 14884 30598
rect 14832 30534 14884 30540
rect 14924 30388 14976 30394
rect 14924 30330 14976 30336
rect 14832 30184 14884 30190
rect 14832 30126 14884 30132
rect 14740 30116 14792 30122
rect 14740 30058 14792 30064
rect 14844 29714 14872 30126
rect 14832 29708 14884 29714
rect 14832 29650 14884 29656
rect 14936 29578 14964 30330
rect 15028 30054 15056 31606
rect 15016 30048 15068 30054
rect 15016 29990 15068 29996
rect 14832 29572 14884 29578
rect 14832 29514 14884 29520
rect 14924 29572 14976 29578
rect 14924 29514 14976 29520
rect 14844 29306 14872 29514
rect 14832 29300 14884 29306
rect 14832 29242 14884 29248
rect 14648 28960 14700 28966
rect 14648 28902 14700 28908
rect 14660 28762 14688 28902
rect 14648 28756 14700 28762
rect 14648 28698 14700 28704
rect 14556 28076 14608 28082
rect 14556 28018 14608 28024
rect 14648 28076 14700 28082
rect 14648 28018 14700 28024
rect 14464 27872 14516 27878
rect 14464 27814 14516 27820
rect 14464 27668 14516 27674
rect 14464 27610 14516 27616
rect 14200 27390 14320 27418
rect 14372 27464 14424 27470
rect 14372 27406 14424 27412
rect 14096 27328 14148 27334
rect 14096 27270 14148 27276
rect 14108 24274 14136 27270
rect 14200 26466 14228 27390
rect 14280 26784 14332 26790
rect 14280 26726 14332 26732
rect 14292 26586 14320 26726
rect 14280 26580 14332 26586
rect 14280 26522 14332 26528
rect 14200 26450 14320 26466
rect 14200 26444 14332 26450
rect 14200 26438 14280 26444
rect 14280 26386 14332 26392
rect 14188 24812 14240 24818
rect 14188 24754 14240 24760
rect 14200 24614 14228 24754
rect 14188 24608 14240 24614
rect 14188 24550 14240 24556
rect 14096 24268 14148 24274
rect 14096 24210 14148 24216
rect 14292 23798 14320 26386
rect 14384 24868 14412 27406
rect 14476 26994 14504 27610
rect 14568 27334 14596 28018
rect 14660 27674 14688 28018
rect 14648 27668 14700 27674
rect 14648 27610 14700 27616
rect 14832 27464 14884 27470
rect 14832 27406 14884 27412
rect 14556 27328 14608 27334
rect 14556 27270 14608 27276
rect 14464 26988 14516 26994
rect 14464 26930 14516 26936
rect 14568 26466 14596 27270
rect 14648 26920 14700 26926
rect 14740 26920 14792 26926
rect 14648 26862 14700 26868
rect 14738 26888 14740 26897
rect 14792 26888 14794 26897
rect 14660 26586 14688 26862
rect 14738 26823 14794 26832
rect 14648 26580 14700 26586
rect 14648 26522 14700 26528
rect 14568 26438 14780 26466
rect 14844 26450 14872 27406
rect 14936 26994 14964 29514
rect 15028 28082 15056 29990
rect 15212 29753 15240 33487
rect 15396 29782 15424 37674
rect 15568 36712 15620 36718
rect 15568 36654 15620 36660
rect 15580 36242 15608 36654
rect 15752 36576 15804 36582
rect 15752 36518 15804 36524
rect 15568 36236 15620 36242
rect 15568 36178 15620 36184
rect 15764 36174 15792 36518
rect 15948 36378 15976 37810
rect 15936 36372 15988 36378
rect 15936 36314 15988 36320
rect 15752 36168 15804 36174
rect 15566 36136 15622 36145
rect 15476 36100 15528 36106
rect 15528 36080 15566 36088
rect 15752 36110 15804 36116
rect 15528 36071 15622 36080
rect 15528 36060 15608 36071
rect 15476 36042 15528 36048
rect 15660 36032 15712 36038
rect 15660 35974 15712 35980
rect 15672 33969 15700 35974
rect 15936 34944 15988 34950
rect 15936 34886 15988 34892
rect 15752 33992 15804 33998
rect 15658 33960 15714 33969
rect 15476 33924 15528 33930
rect 15752 33934 15804 33940
rect 15658 33895 15714 33904
rect 15476 33866 15528 33872
rect 15488 33810 15516 33866
rect 15566 33824 15622 33833
rect 15488 33782 15566 33810
rect 15566 33759 15622 33768
rect 15476 32428 15528 32434
rect 15476 32370 15528 32376
rect 15488 31346 15516 32370
rect 15672 31754 15700 33895
rect 15764 32434 15792 33934
rect 15844 32904 15896 32910
rect 15844 32846 15896 32852
rect 15752 32428 15804 32434
rect 15752 32370 15804 32376
rect 15856 31754 15884 32846
rect 15580 31726 15700 31754
rect 15764 31726 15884 31754
rect 15476 31340 15528 31346
rect 15476 31282 15528 31288
rect 15384 29776 15436 29782
rect 15198 29744 15254 29753
rect 15384 29718 15436 29724
rect 15198 29679 15254 29688
rect 15212 29646 15240 29679
rect 15200 29640 15252 29646
rect 15200 29582 15252 29588
rect 15212 28370 15240 29582
rect 15212 28342 15332 28370
rect 15016 28076 15068 28082
rect 15016 28018 15068 28024
rect 15304 27606 15332 28342
rect 15016 27600 15068 27606
rect 15016 27542 15068 27548
rect 15292 27600 15344 27606
rect 15292 27542 15344 27548
rect 14924 26988 14976 26994
rect 14924 26930 14976 26936
rect 15028 26466 15056 27542
rect 15396 27418 15424 29718
rect 15580 29646 15608 31726
rect 15764 31346 15792 31726
rect 15752 31340 15804 31346
rect 15752 31282 15804 31288
rect 15658 30152 15714 30161
rect 15658 30087 15714 30096
rect 15672 29646 15700 30087
rect 15568 29640 15620 29646
rect 15568 29582 15620 29588
rect 15660 29640 15712 29646
rect 15660 29582 15712 29588
rect 15580 27946 15608 29582
rect 15764 29458 15792 31282
rect 15844 30048 15896 30054
rect 15844 29990 15896 29996
rect 15856 29646 15884 29990
rect 15844 29640 15896 29646
rect 15842 29608 15844 29617
rect 15896 29608 15898 29617
rect 15842 29543 15898 29552
rect 15764 29430 15884 29458
rect 15752 28212 15804 28218
rect 15752 28154 15804 28160
rect 15568 27940 15620 27946
rect 15568 27882 15620 27888
rect 15476 27872 15528 27878
rect 15476 27814 15528 27820
rect 15304 27390 15424 27418
rect 15108 26852 15160 26858
rect 15108 26794 15160 26800
rect 15120 26586 15148 26794
rect 15304 26586 15332 27390
rect 15384 27328 15436 27334
rect 15384 27270 15436 27276
rect 15396 26858 15424 27270
rect 15488 27062 15516 27814
rect 15476 27056 15528 27062
rect 15476 26998 15528 27004
rect 15384 26852 15436 26858
rect 15384 26794 15436 26800
rect 15108 26580 15160 26586
rect 15108 26522 15160 26528
rect 15292 26580 15344 26586
rect 15292 26522 15344 26528
rect 15028 26450 15148 26466
rect 14464 26308 14516 26314
rect 14464 26250 14516 26256
rect 14476 24993 14504 26250
rect 14648 26240 14700 26246
rect 14648 26182 14700 26188
rect 14660 25838 14688 26182
rect 14752 26042 14780 26438
rect 14832 26444 14884 26450
rect 15028 26444 15160 26450
rect 15028 26438 15108 26444
rect 14832 26386 14884 26392
rect 15108 26386 15160 26392
rect 15304 26330 15332 26522
rect 15396 26450 15424 26794
rect 15384 26444 15436 26450
rect 15384 26386 15436 26392
rect 15580 26382 15608 27882
rect 15660 26988 15712 26994
rect 15660 26930 15712 26936
rect 15568 26376 15620 26382
rect 15120 26302 15332 26330
rect 15488 26336 15568 26364
rect 15120 26246 15148 26302
rect 15108 26240 15160 26246
rect 15108 26182 15160 26188
rect 14740 26036 14792 26042
rect 14740 25978 14792 25984
rect 14648 25832 14700 25838
rect 14648 25774 14700 25780
rect 14462 24984 14518 24993
rect 14462 24919 14518 24928
rect 14384 24840 14504 24868
rect 14372 24744 14424 24750
rect 14372 24686 14424 24692
rect 14384 24206 14412 24686
rect 14372 24200 14424 24206
rect 14372 24142 14424 24148
rect 14280 23792 14332 23798
rect 14278 23760 14280 23769
rect 14332 23760 14334 23769
rect 14188 23724 14240 23730
rect 14384 23730 14412 24142
rect 14476 23798 14504 24840
rect 14556 24268 14608 24274
rect 14556 24210 14608 24216
rect 14464 23792 14516 23798
rect 14464 23734 14516 23740
rect 14278 23695 14334 23704
rect 14372 23724 14424 23730
rect 14188 23666 14240 23672
rect 14372 23666 14424 23672
rect 14200 23322 14228 23666
rect 14188 23316 14240 23322
rect 14188 23258 14240 23264
rect 13912 23180 13964 23186
rect 14016 23174 14228 23202
rect 13912 23122 13964 23128
rect 14096 22500 14148 22506
rect 14096 22442 14148 22448
rect 13910 21720 13966 21729
rect 13910 21655 13966 21664
rect 13924 21418 13952 21655
rect 14004 21480 14056 21486
rect 14004 21422 14056 21428
rect 13912 21412 13964 21418
rect 13912 21354 13964 21360
rect 14016 21078 14044 21422
rect 14004 21072 14056 21078
rect 14004 21014 14056 21020
rect 13912 20324 13964 20330
rect 13912 20266 13964 20272
rect 13924 20058 13952 20266
rect 13912 20052 13964 20058
rect 13912 19994 13964 20000
rect 14004 19916 14056 19922
rect 14004 19858 14056 19864
rect 14016 18902 14044 19858
rect 14004 18896 14056 18902
rect 14004 18838 14056 18844
rect 13912 18624 13964 18630
rect 13912 18566 13964 18572
rect 13924 18426 13952 18566
rect 13820 18420 13872 18426
rect 13820 18362 13872 18368
rect 13912 18420 13964 18426
rect 13912 18362 13964 18368
rect 13820 18284 13872 18290
rect 14016 18272 14044 18838
rect 13872 18244 14044 18272
rect 13820 18226 13872 18232
rect 13728 17536 13780 17542
rect 13728 17478 13780 17484
rect 13544 17196 13596 17202
rect 13544 17138 13596 17144
rect 13556 14822 13584 17138
rect 13544 14816 13596 14822
rect 13544 14758 13596 14764
rect 13544 13184 13596 13190
rect 13544 13126 13596 13132
rect 13636 13184 13688 13190
rect 13636 13126 13688 13132
rect 13556 12918 13584 13126
rect 13648 12986 13676 13126
rect 13636 12980 13688 12986
rect 13636 12922 13688 12928
rect 13544 12912 13596 12918
rect 13544 12854 13596 12860
rect 13556 11898 13584 12854
rect 13740 12434 13768 17478
rect 13832 17338 13860 18226
rect 14108 17746 14136 22442
rect 14200 20874 14228 23174
rect 14280 23044 14332 23050
rect 14280 22986 14332 22992
rect 14292 22710 14320 22986
rect 14280 22704 14332 22710
rect 14280 22646 14332 22652
rect 14278 21040 14334 21049
rect 14384 21010 14412 23666
rect 14464 23044 14516 23050
rect 14464 22986 14516 22992
rect 14476 22642 14504 22986
rect 14464 22636 14516 22642
rect 14464 22578 14516 22584
rect 14568 22166 14596 24210
rect 14660 22574 14688 25774
rect 14752 23186 14780 25978
rect 14832 25764 14884 25770
rect 14832 25706 14884 25712
rect 14844 25362 14872 25706
rect 15016 25696 15068 25702
rect 15016 25638 15068 25644
rect 14832 25356 14884 25362
rect 14832 25298 14884 25304
rect 15028 25294 15056 25638
rect 15016 25288 15068 25294
rect 15016 25230 15068 25236
rect 15016 24948 15068 24954
rect 15016 24890 15068 24896
rect 14924 24812 14976 24818
rect 14924 24754 14976 24760
rect 14936 24342 14964 24754
rect 14924 24336 14976 24342
rect 14924 24278 14976 24284
rect 14936 24206 14964 24278
rect 14924 24200 14976 24206
rect 14924 24142 14976 24148
rect 14936 23730 14964 24142
rect 15028 24138 15056 24890
rect 15384 24812 15436 24818
rect 15384 24754 15436 24760
rect 15200 24608 15252 24614
rect 15200 24550 15252 24556
rect 15212 24342 15240 24550
rect 15396 24410 15424 24754
rect 15384 24404 15436 24410
rect 15384 24346 15436 24352
rect 15200 24336 15252 24342
rect 15200 24278 15252 24284
rect 15488 24274 15516 26336
rect 15568 26318 15620 26324
rect 15568 26036 15620 26042
rect 15568 25978 15620 25984
rect 15476 24268 15528 24274
rect 15476 24210 15528 24216
rect 15384 24200 15436 24206
rect 15580 24154 15608 25978
rect 15672 25362 15700 26930
rect 15660 25356 15712 25362
rect 15660 25298 15712 25304
rect 15384 24142 15436 24148
rect 15016 24132 15068 24138
rect 15016 24074 15068 24080
rect 15028 23798 15056 24074
rect 15016 23792 15068 23798
rect 15016 23734 15068 23740
rect 14924 23724 14976 23730
rect 14924 23666 14976 23672
rect 14740 23180 14792 23186
rect 14740 23122 14792 23128
rect 14648 22568 14700 22574
rect 14648 22510 14700 22516
rect 14832 22432 14884 22438
rect 14832 22374 14884 22380
rect 14556 22160 14608 22166
rect 14556 22102 14608 22108
rect 14648 22160 14700 22166
rect 14648 22102 14700 22108
rect 14556 22024 14608 22030
rect 14556 21966 14608 21972
rect 14464 21072 14516 21078
rect 14464 21014 14516 21020
rect 14278 20975 14334 20984
rect 14372 21004 14424 21010
rect 14188 20868 14240 20874
rect 14188 20810 14240 20816
rect 14292 20602 14320 20975
rect 14372 20946 14424 20952
rect 14280 20596 14332 20602
rect 14280 20538 14332 20544
rect 14372 20460 14424 20466
rect 14372 20402 14424 20408
rect 14280 20256 14332 20262
rect 14280 20198 14332 20204
rect 14292 19922 14320 20198
rect 14280 19916 14332 19922
rect 14280 19858 14332 19864
rect 14384 19378 14412 20402
rect 14476 19854 14504 21014
rect 14568 20942 14596 21966
rect 14660 21486 14688 22102
rect 14844 22030 14872 22374
rect 14832 22024 14884 22030
rect 14832 21966 14884 21972
rect 14936 21690 14964 23666
rect 15028 22438 15056 23734
rect 15396 23594 15424 24142
rect 15488 24126 15608 24154
rect 15384 23588 15436 23594
rect 15384 23530 15436 23536
rect 15108 23520 15160 23526
rect 15108 23462 15160 23468
rect 15016 22432 15068 22438
rect 15016 22374 15068 22380
rect 15120 22094 15148 23462
rect 15384 23112 15436 23118
rect 15384 23054 15436 23060
rect 15292 23044 15344 23050
rect 15292 22986 15344 22992
rect 15304 22778 15332 22986
rect 15292 22772 15344 22778
rect 15292 22714 15344 22720
rect 15200 22636 15252 22642
rect 15200 22578 15252 22584
rect 15028 22066 15148 22094
rect 14924 21684 14976 21690
rect 14924 21626 14976 21632
rect 14648 21480 14700 21486
rect 14648 21422 14700 21428
rect 14556 20936 14608 20942
rect 14556 20878 14608 20884
rect 14740 20936 14792 20942
rect 14740 20878 14792 20884
rect 14924 20936 14976 20942
rect 14924 20878 14976 20884
rect 14568 20602 14596 20878
rect 14556 20596 14608 20602
rect 14556 20538 14608 20544
rect 14648 20528 14700 20534
rect 14648 20470 14700 20476
rect 14464 19848 14516 19854
rect 14464 19790 14516 19796
rect 14554 19544 14610 19553
rect 14464 19508 14516 19514
rect 14554 19479 14610 19488
rect 14464 19450 14516 19456
rect 14372 19372 14424 19378
rect 14372 19314 14424 19320
rect 14188 18624 14240 18630
rect 14188 18566 14240 18572
rect 14200 18426 14228 18566
rect 14188 18420 14240 18426
rect 14188 18362 14240 18368
rect 14280 18284 14332 18290
rect 14280 18226 14332 18232
rect 14188 18080 14240 18086
rect 14188 18022 14240 18028
rect 14200 17814 14228 18022
rect 14188 17808 14240 17814
rect 14188 17750 14240 17756
rect 14096 17740 14148 17746
rect 14096 17682 14148 17688
rect 14004 17536 14056 17542
rect 14004 17478 14056 17484
rect 14016 17338 14044 17478
rect 13820 17332 13872 17338
rect 13820 17274 13872 17280
rect 14004 17332 14056 17338
rect 14004 17274 14056 17280
rect 13832 15434 13860 17274
rect 14108 16250 14136 17682
rect 14188 17672 14240 17678
rect 14188 17614 14240 17620
rect 14200 17066 14228 17614
rect 14292 17542 14320 18226
rect 14384 17610 14412 19314
rect 14372 17604 14424 17610
rect 14372 17546 14424 17552
rect 14280 17536 14332 17542
rect 14280 17478 14332 17484
rect 14188 17060 14240 17066
rect 14188 17002 14240 17008
rect 14200 16590 14228 17002
rect 14384 16697 14412 17546
rect 14476 17134 14504 19450
rect 14568 19378 14596 19479
rect 14660 19446 14688 20470
rect 14752 19990 14780 20878
rect 14830 20496 14886 20505
rect 14830 20431 14886 20440
rect 14844 20398 14872 20431
rect 14832 20392 14884 20398
rect 14832 20334 14884 20340
rect 14740 19984 14792 19990
rect 14740 19926 14792 19932
rect 14752 19514 14780 19926
rect 14740 19508 14792 19514
rect 14740 19450 14792 19456
rect 14648 19440 14700 19446
rect 14648 19382 14700 19388
rect 14556 19372 14608 19378
rect 14556 19314 14608 19320
rect 14660 19242 14688 19382
rect 14648 19236 14700 19242
rect 14648 19178 14700 19184
rect 14844 17746 14872 20334
rect 14936 19310 14964 20878
rect 14924 19304 14976 19310
rect 14924 19246 14976 19252
rect 14832 17740 14884 17746
rect 14832 17682 14884 17688
rect 14464 17128 14516 17134
rect 14464 17070 14516 17076
rect 14370 16688 14426 16697
rect 14370 16623 14426 16632
rect 14188 16584 14240 16590
rect 14188 16526 14240 16532
rect 14096 16244 14148 16250
rect 14096 16186 14148 16192
rect 14200 15994 14228 16526
rect 14108 15966 14228 15994
rect 14108 15502 14136 15966
rect 14188 15904 14240 15910
rect 14188 15846 14240 15852
rect 14200 15706 14228 15846
rect 14188 15700 14240 15706
rect 14188 15642 14240 15648
rect 14096 15496 14148 15502
rect 14096 15438 14148 15444
rect 13820 15428 13872 15434
rect 13820 15370 13872 15376
rect 14096 15020 14148 15026
rect 14096 14962 14148 14968
rect 14108 14618 14136 14962
rect 14096 14612 14148 14618
rect 14096 14554 14148 14560
rect 14004 14272 14056 14278
rect 14004 14214 14056 14220
rect 13648 12406 13768 12434
rect 13544 11892 13596 11898
rect 13544 11834 13596 11840
rect 13452 10056 13504 10062
rect 13452 9998 13504 10004
rect 13452 9376 13504 9382
rect 13452 9318 13504 9324
rect 13360 8968 13412 8974
rect 13360 8910 13412 8916
rect 13464 8838 13492 9318
rect 13544 9036 13596 9042
rect 13544 8978 13596 8984
rect 12992 8832 13044 8838
rect 12992 8774 13044 8780
rect 13452 8832 13504 8838
rect 13452 8774 13504 8780
rect 13004 8634 13032 8774
rect 13464 8634 13492 8774
rect 12992 8628 13044 8634
rect 12992 8570 13044 8576
rect 13452 8628 13504 8634
rect 13452 8570 13504 8576
rect 12992 8492 13044 8498
rect 12992 8434 13044 8440
rect 13004 8090 13032 8434
rect 12992 8084 13044 8090
rect 12992 8026 13044 8032
rect 13556 7954 13584 8978
rect 13544 7948 13596 7954
rect 13544 7890 13596 7896
rect 12900 7880 12952 7886
rect 12900 7822 12952 7828
rect 12808 7404 12860 7410
rect 12808 7346 12860 7352
rect 12268 6882 12296 6990
rect 12348 6996 12400 7002
rect 12348 6938 12400 6944
rect 12268 6854 12664 6882
rect 12360 6186 12480 6202
rect 12348 6180 12480 6186
rect 12400 6174 12480 6180
rect 12348 6122 12400 6128
rect 12452 5778 12480 6174
rect 12532 6112 12584 6118
rect 12532 6054 12584 6060
rect 12440 5772 12492 5778
rect 12440 5714 12492 5720
rect 12544 5658 12572 6054
rect 12452 5642 12572 5658
rect 12440 5636 12572 5642
rect 12492 5630 12572 5636
rect 12440 5578 12492 5584
rect 11888 5364 11940 5370
rect 11888 5306 11940 5312
rect 12164 5364 12216 5370
rect 12164 5306 12216 5312
rect 10416 5296 10468 5302
rect 10416 5238 10468 5244
rect 11704 5296 11756 5302
rect 11704 5238 11756 5244
rect 11152 5024 11204 5030
rect 11152 4966 11204 4972
rect 11164 4826 11192 4966
rect 11152 4820 11204 4826
rect 11152 4762 11204 4768
rect 12176 4690 12204 5306
rect 12452 4826 12480 5578
rect 12636 5216 12664 6854
rect 12820 6798 12848 7346
rect 12912 7206 12940 7822
rect 13544 7812 13596 7818
rect 13544 7754 13596 7760
rect 12900 7200 12952 7206
rect 12900 7142 12952 7148
rect 12912 6798 12940 7142
rect 13556 7002 13584 7754
rect 13648 7546 13676 12406
rect 13820 10736 13872 10742
rect 13820 10678 13872 10684
rect 13832 10470 13860 10678
rect 13820 10464 13872 10470
rect 13820 10406 13872 10412
rect 13728 9444 13780 9450
rect 13728 9386 13780 9392
rect 13740 9042 13768 9386
rect 13912 9376 13964 9382
rect 13912 9318 13964 9324
rect 13818 9208 13874 9217
rect 13924 9178 13952 9318
rect 13818 9143 13820 9152
rect 13872 9143 13874 9152
rect 13912 9172 13964 9178
rect 13820 9114 13872 9120
rect 13912 9114 13964 9120
rect 13728 9036 13780 9042
rect 13728 8978 13780 8984
rect 13912 8968 13964 8974
rect 13912 8910 13964 8916
rect 13924 8838 13952 8910
rect 13912 8832 13964 8838
rect 13912 8774 13964 8780
rect 13728 8084 13780 8090
rect 13728 8026 13780 8032
rect 13636 7540 13688 7546
rect 13636 7482 13688 7488
rect 13544 6996 13596 7002
rect 13544 6938 13596 6944
rect 12808 6792 12860 6798
rect 12808 6734 12860 6740
rect 12900 6792 12952 6798
rect 12900 6734 12952 6740
rect 13556 6322 13584 6938
rect 13740 6866 13768 8026
rect 14016 7954 14044 14214
rect 14096 11008 14148 11014
rect 14096 10950 14148 10956
rect 14108 10742 14136 10950
rect 14096 10736 14148 10742
rect 14096 10678 14148 10684
rect 14200 9674 14228 15642
rect 14384 15026 14412 16623
rect 14476 16454 14504 17070
rect 14464 16448 14516 16454
rect 14464 16390 14516 16396
rect 14476 16114 14504 16390
rect 14844 16114 14872 17682
rect 14464 16108 14516 16114
rect 14464 16050 14516 16056
rect 14740 16108 14792 16114
rect 14740 16050 14792 16056
rect 14832 16108 14884 16114
rect 14832 16050 14884 16056
rect 14372 15020 14424 15026
rect 14372 14962 14424 14968
rect 14384 14482 14412 14962
rect 14476 14890 14504 16050
rect 14752 15910 14780 16050
rect 14740 15904 14792 15910
rect 14740 15846 14792 15852
rect 14648 15496 14700 15502
rect 14648 15438 14700 15444
rect 14660 14958 14688 15438
rect 14740 15428 14792 15434
rect 14740 15370 14792 15376
rect 14648 14952 14700 14958
rect 14648 14894 14700 14900
rect 14752 14890 14780 15370
rect 14844 15026 14872 16050
rect 14832 15020 14884 15026
rect 14832 14962 14884 14968
rect 14464 14884 14516 14890
rect 14464 14826 14516 14832
rect 14740 14884 14792 14890
rect 14740 14826 14792 14832
rect 14372 14476 14424 14482
rect 14372 14418 14424 14424
rect 14476 14414 14504 14826
rect 14464 14408 14516 14414
rect 14464 14350 14516 14356
rect 14648 12640 14700 12646
rect 14648 12582 14700 12588
rect 14464 11824 14516 11830
rect 14464 11766 14516 11772
rect 14476 11354 14504 11766
rect 14464 11348 14516 11354
rect 14464 11290 14516 11296
rect 14660 11218 14688 12582
rect 14752 11694 14780 14826
rect 14844 14618 14872 14962
rect 14832 14612 14884 14618
rect 14832 14554 14884 14560
rect 14832 14408 14884 14414
rect 14832 14350 14884 14356
rect 14844 12918 14872 14350
rect 14832 12912 14884 12918
rect 14832 12854 14884 12860
rect 15028 12730 15056 22066
rect 15212 22030 15240 22578
rect 15396 22094 15424 23054
rect 15488 22522 15516 24126
rect 15568 24064 15620 24070
rect 15568 24006 15620 24012
rect 15580 23730 15608 24006
rect 15672 23866 15700 25298
rect 15764 24410 15792 28154
rect 15856 27878 15884 29430
rect 15844 27872 15896 27878
rect 15844 27814 15896 27820
rect 15856 27470 15884 27814
rect 15844 27464 15896 27470
rect 15844 27406 15896 27412
rect 15948 26042 15976 34886
rect 16132 32298 16160 37810
rect 16224 36174 16252 37810
rect 16212 36168 16264 36174
rect 16212 36110 16264 36116
rect 16224 35630 16252 36110
rect 16212 35624 16264 35630
rect 16212 35566 16264 35572
rect 16316 33998 16344 37828
rect 16396 37810 16448 37816
rect 16856 37868 16908 37874
rect 16856 37810 16908 37816
rect 16868 37738 16896 37810
rect 16856 37732 16908 37738
rect 16856 37674 16908 37680
rect 16488 37664 16540 37670
rect 16488 37606 16540 37612
rect 16500 37466 16528 37606
rect 16488 37460 16540 37466
rect 16488 37402 16540 37408
rect 16868 36174 16896 37674
rect 16960 36786 16988 37878
rect 17880 37874 18000 37890
rect 20536 37878 20588 37884
rect 17316 37868 17368 37874
rect 17316 37810 17368 37816
rect 17776 37868 17828 37874
rect 17776 37810 17828 37816
rect 17868 37868 18000 37874
rect 17920 37862 18000 37868
rect 17868 37810 17920 37816
rect 17224 37120 17276 37126
rect 17224 37062 17276 37068
rect 16948 36780 17000 36786
rect 16948 36722 17000 36728
rect 17040 36644 17092 36650
rect 17040 36586 17092 36592
rect 16672 36168 16724 36174
rect 16856 36168 16908 36174
rect 16724 36128 16804 36156
rect 16672 36110 16724 36116
rect 16488 34672 16540 34678
rect 16488 34614 16540 34620
rect 16500 33998 16528 34614
rect 16580 34604 16632 34610
rect 16580 34546 16632 34552
rect 16212 33992 16264 33998
rect 16212 33934 16264 33940
rect 16304 33992 16356 33998
rect 16304 33934 16356 33940
rect 16488 33992 16540 33998
rect 16488 33934 16540 33940
rect 16224 33318 16252 33934
rect 16212 33312 16264 33318
rect 16212 33254 16264 33260
rect 16224 32910 16252 33254
rect 16212 32904 16264 32910
rect 16212 32846 16264 32852
rect 16120 32292 16172 32298
rect 16120 32234 16172 32240
rect 16132 31346 16160 32234
rect 16316 31521 16344 33934
rect 16500 33658 16528 33934
rect 16488 33652 16540 33658
rect 16488 33594 16540 33600
rect 16592 33590 16620 34546
rect 16672 33924 16724 33930
rect 16672 33866 16724 33872
rect 16580 33584 16632 33590
rect 16580 33526 16632 33532
rect 16684 32484 16712 33866
rect 16776 33046 16804 36128
rect 16856 36110 16908 36116
rect 17052 36106 17080 36586
rect 16948 36100 17000 36106
rect 16948 36042 17000 36048
rect 17040 36100 17092 36106
rect 17040 36042 17092 36048
rect 16960 34678 16988 36042
rect 16948 34672 17000 34678
rect 16948 34614 17000 34620
rect 16856 34400 16908 34406
rect 16856 34342 16908 34348
rect 16948 34400 17000 34406
rect 16948 34342 17000 34348
rect 17040 34400 17092 34406
rect 17040 34342 17092 34348
rect 16868 34202 16896 34342
rect 16960 34202 16988 34342
rect 17052 34202 17080 34342
rect 16856 34196 16908 34202
rect 16856 34138 16908 34144
rect 16948 34196 17000 34202
rect 16948 34138 17000 34144
rect 17040 34196 17092 34202
rect 17040 34138 17092 34144
rect 16960 33918 17172 33946
rect 16960 33862 16988 33918
rect 17144 33862 17172 33918
rect 16948 33856 17000 33862
rect 16948 33798 17000 33804
rect 17040 33856 17092 33862
rect 17040 33798 17092 33804
rect 17132 33856 17184 33862
rect 17132 33798 17184 33804
rect 16856 33652 16908 33658
rect 16856 33594 16908 33600
rect 16764 33040 16816 33046
rect 16764 32982 16816 32988
rect 16868 32842 16896 33594
rect 16856 32836 16908 32842
rect 16856 32778 16908 32784
rect 16764 32496 16816 32502
rect 16684 32456 16764 32484
rect 16816 32456 16896 32484
rect 16764 32438 16816 32444
rect 16672 32224 16724 32230
rect 16672 32166 16724 32172
rect 16488 31748 16540 31754
rect 16488 31690 16540 31696
rect 16302 31512 16358 31521
rect 16212 31476 16264 31482
rect 16302 31447 16358 31456
rect 16212 31418 16264 31424
rect 16224 31346 16252 31418
rect 16028 31340 16080 31346
rect 16028 31282 16080 31288
rect 16120 31340 16172 31346
rect 16120 31282 16172 31288
rect 16212 31340 16264 31346
rect 16212 31282 16264 31288
rect 16040 29646 16068 31282
rect 16132 30546 16160 31282
rect 16316 30598 16344 31447
rect 16500 31346 16528 31690
rect 16488 31340 16540 31346
rect 16408 31300 16488 31328
rect 16304 30592 16356 30598
rect 16132 30518 16252 30546
rect 16304 30534 16356 30540
rect 16120 30048 16172 30054
rect 16120 29990 16172 29996
rect 16028 29640 16080 29646
rect 16028 29582 16080 29588
rect 16132 29170 16160 29990
rect 16120 29164 16172 29170
rect 16120 29106 16172 29112
rect 16224 28558 16252 30518
rect 16316 28994 16344 30534
rect 16408 30138 16436 31300
rect 16488 31282 16540 31288
rect 16488 31136 16540 31142
rect 16488 31078 16540 31084
rect 16500 30258 16528 31078
rect 16580 30728 16632 30734
rect 16580 30670 16632 30676
rect 16684 30682 16712 32166
rect 16868 31260 16896 32456
rect 16960 32230 16988 33798
rect 17052 33658 17080 33798
rect 17040 33652 17092 33658
rect 17040 33594 17092 33600
rect 17040 33380 17092 33386
rect 17040 33322 17092 33328
rect 16948 32224 17000 32230
rect 16948 32166 17000 32172
rect 16960 31686 16988 32166
rect 16948 31680 17000 31686
rect 16948 31622 17000 31628
rect 16948 31408 17000 31414
rect 17052 31396 17080 33322
rect 17130 32328 17186 32337
rect 17130 32263 17132 32272
rect 17184 32263 17186 32272
rect 17132 32234 17184 32240
rect 17236 31754 17264 37062
rect 17328 36174 17356 37810
rect 17788 37754 17816 37810
rect 17788 37726 17908 37754
rect 17776 37664 17828 37670
rect 17776 37606 17828 37612
rect 17788 37330 17816 37606
rect 17776 37324 17828 37330
rect 17776 37266 17828 37272
rect 17776 37188 17828 37194
rect 17776 37130 17828 37136
rect 17788 36378 17816 37130
rect 17776 36372 17828 36378
rect 17776 36314 17828 36320
rect 17316 36168 17368 36174
rect 17316 36110 17368 36116
rect 17592 36168 17644 36174
rect 17592 36110 17644 36116
rect 17328 35170 17356 36110
rect 17408 36032 17460 36038
rect 17406 36000 17408 36009
rect 17460 36000 17462 36009
rect 17406 35935 17462 35944
rect 17328 35142 17448 35170
rect 17316 35080 17368 35086
rect 17316 35022 17368 35028
rect 17328 34746 17356 35022
rect 17316 34740 17368 34746
rect 17316 34682 17368 34688
rect 17316 34604 17368 34610
rect 17316 34546 17368 34552
rect 17000 31368 17080 31396
rect 17144 31726 17264 31754
rect 16948 31350 17000 31356
rect 16868 31232 17080 31260
rect 16764 31136 16816 31142
rect 16764 31078 16816 31084
rect 16776 30870 16804 31078
rect 16764 30864 16816 30870
rect 16764 30806 16816 30812
rect 16948 30796 17000 30802
rect 16948 30738 17000 30744
rect 16488 30252 16540 30258
rect 16488 30194 16540 30200
rect 16408 30110 16528 30138
rect 16316 28966 16436 28994
rect 16120 28552 16172 28558
rect 16120 28494 16172 28500
rect 16212 28552 16264 28558
rect 16212 28494 16264 28500
rect 16132 28218 16160 28494
rect 16120 28212 16172 28218
rect 16120 28154 16172 28160
rect 16028 28076 16080 28082
rect 16028 28018 16080 28024
rect 15936 26036 15988 26042
rect 15936 25978 15988 25984
rect 16040 25294 16068 28018
rect 16304 27532 16356 27538
rect 16304 27474 16356 27480
rect 16212 27464 16264 27470
rect 16212 27406 16264 27412
rect 15936 25288 15988 25294
rect 15936 25230 15988 25236
rect 16028 25288 16080 25294
rect 16028 25230 16080 25236
rect 15844 24948 15896 24954
rect 15844 24890 15896 24896
rect 15752 24404 15804 24410
rect 15752 24346 15804 24352
rect 15856 24206 15884 24890
rect 15844 24200 15896 24206
rect 15844 24142 15896 24148
rect 15660 23860 15712 23866
rect 15660 23802 15712 23808
rect 15568 23724 15620 23730
rect 15568 23666 15620 23672
rect 15948 23526 15976 25230
rect 16120 24812 16172 24818
rect 16120 24754 16172 24760
rect 16028 23792 16080 23798
rect 16028 23734 16080 23740
rect 15936 23520 15988 23526
rect 15936 23462 15988 23468
rect 15844 23112 15896 23118
rect 15844 23054 15896 23060
rect 15936 23112 15988 23118
rect 15936 23054 15988 23060
rect 15752 22772 15804 22778
rect 15752 22714 15804 22720
rect 15488 22494 15608 22522
rect 15476 22094 15528 22098
rect 15396 22092 15528 22094
rect 15396 22080 15476 22092
rect 15304 22052 15476 22080
rect 15200 22024 15252 22030
rect 15200 21966 15252 21972
rect 15108 21684 15160 21690
rect 15108 21626 15160 21632
rect 15120 21010 15148 21626
rect 15108 21004 15160 21010
rect 15108 20946 15160 20952
rect 15108 20868 15160 20874
rect 15108 20810 15160 20816
rect 15120 20058 15148 20810
rect 15212 20602 15240 21966
rect 15304 21554 15332 22052
rect 15476 22034 15528 22040
rect 15476 21888 15528 21894
rect 15476 21830 15528 21836
rect 15488 21554 15516 21830
rect 15580 21593 15608 22494
rect 15764 22030 15792 22714
rect 15856 22030 15884 23054
rect 15948 22574 15976 23054
rect 15936 22568 15988 22574
rect 15936 22510 15988 22516
rect 16040 22166 16068 23734
rect 16132 23662 16160 24754
rect 16224 24664 16252 27406
rect 16316 24732 16344 27474
rect 16408 26228 16436 28966
rect 16500 28558 16528 30110
rect 16592 29850 16620 30670
rect 16684 30654 16804 30682
rect 16672 30592 16724 30598
rect 16672 30534 16724 30540
rect 16684 30297 16712 30534
rect 16670 30288 16726 30297
rect 16670 30223 16726 30232
rect 16684 30190 16712 30223
rect 16672 30184 16724 30190
rect 16672 30126 16724 30132
rect 16580 29844 16632 29850
rect 16580 29786 16632 29792
rect 16776 29510 16804 30654
rect 16960 30054 16988 30738
rect 16948 30048 17000 30054
rect 16948 29990 17000 29996
rect 17052 29510 17080 31232
rect 17144 30734 17172 31726
rect 17328 31657 17356 34546
rect 17420 33114 17448 35142
rect 17500 33856 17552 33862
rect 17500 33798 17552 33804
rect 17512 33561 17540 33798
rect 17498 33552 17554 33561
rect 17604 33538 17632 36110
rect 17684 36100 17736 36106
rect 17684 36042 17736 36048
rect 17696 34610 17724 36042
rect 17684 34604 17736 34610
rect 17684 34546 17736 34552
rect 17776 34536 17828 34542
rect 17776 34478 17828 34484
rect 17788 33998 17816 34478
rect 17684 33992 17736 33998
rect 17684 33934 17736 33940
rect 17776 33992 17828 33998
rect 17776 33934 17828 33940
rect 17696 33658 17724 33934
rect 17684 33652 17736 33658
rect 17684 33594 17736 33600
rect 17604 33510 17816 33538
rect 17498 33487 17554 33496
rect 17408 33108 17460 33114
rect 17408 33050 17460 33056
rect 17420 32026 17448 33050
rect 17684 33040 17736 33046
rect 17684 32982 17736 32988
rect 17592 32836 17644 32842
rect 17592 32778 17644 32784
rect 17604 32502 17632 32778
rect 17592 32496 17644 32502
rect 17592 32438 17644 32444
rect 17408 32020 17460 32026
rect 17408 31962 17460 31968
rect 17314 31648 17370 31657
rect 17314 31583 17370 31592
rect 17328 30870 17356 31583
rect 17420 31346 17448 31962
rect 17604 31822 17632 32438
rect 17592 31816 17644 31822
rect 17592 31758 17644 31764
rect 17604 31498 17632 31758
rect 17512 31470 17632 31498
rect 17696 31482 17724 32982
rect 17788 32450 17816 33510
rect 17880 33153 17908 37726
rect 17972 37330 18000 37862
rect 20352 37868 20404 37874
rect 20352 37810 20404 37816
rect 19340 37800 19392 37806
rect 19340 37742 19392 37748
rect 19984 37800 20036 37806
rect 19984 37742 20036 37748
rect 17960 37324 18012 37330
rect 17960 37266 18012 37272
rect 18604 37256 18656 37262
rect 18604 37198 18656 37204
rect 17960 36712 18012 36718
rect 17960 36654 18012 36660
rect 17972 36106 18000 36654
rect 18616 36310 18644 37198
rect 18972 37120 19024 37126
rect 18972 37062 19024 37068
rect 18696 36780 18748 36786
rect 18696 36722 18748 36728
rect 18604 36304 18656 36310
rect 18604 36246 18656 36252
rect 18708 36174 18736 36722
rect 18052 36168 18104 36174
rect 18696 36168 18748 36174
rect 18052 36110 18104 36116
rect 18248 36128 18696 36156
rect 17960 36100 18012 36106
rect 17960 36042 18012 36048
rect 17960 34672 18012 34678
rect 17960 34614 18012 34620
rect 17972 33930 18000 34614
rect 18064 34406 18092 36110
rect 18052 34400 18104 34406
rect 18052 34342 18104 34348
rect 18064 33998 18092 34342
rect 18052 33992 18104 33998
rect 18052 33934 18104 33940
rect 18144 33992 18196 33998
rect 18144 33934 18196 33940
rect 17960 33924 18012 33930
rect 17960 33866 18012 33872
rect 17972 33386 18000 33866
rect 17960 33380 18012 33386
rect 17960 33322 18012 33328
rect 18156 33318 18184 33934
rect 18144 33312 18196 33318
rect 18144 33254 18196 33260
rect 17866 33144 17922 33153
rect 17866 33079 17922 33088
rect 17880 32570 17908 33079
rect 18156 33046 18184 33254
rect 18144 33040 18196 33046
rect 18144 32982 18196 32988
rect 17960 32904 18012 32910
rect 17960 32846 18012 32852
rect 17868 32564 17920 32570
rect 17868 32506 17920 32512
rect 17972 32502 18000 32846
rect 17960 32496 18012 32502
rect 17788 32422 17908 32450
rect 18248 32450 18276 36128
rect 18696 36110 18748 36116
rect 18788 36100 18840 36106
rect 18788 36042 18840 36048
rect 18604 36032 18656 36038
rect 18604 35974 18656 35980
rect 18616 35766 18644 35974
rect 18604 35760 18656 35766
rect 18604 35702 18656 35708
rect 18696 35488 18748 35494
rect 18696 35430 18748 35436
rect 18420 33992 18472 33998
rect 18420 33934 18472 33940
rect 18328 33856 18380 33862
rect 18328 33798 18380 33804
rect 18340 33114 18368 33798
rect 18432 33590 18460 33934
rect 18604 33924 18656 33930
rect 18604 33866 18656 33872
rect 18512 33856 18564 33862
rect 18512 33798 18564 33804
rect 18420 33584 18472 33590
rect 18420 33526 18472 33532
rect 18420 33448 18472 33454
rect 18524 33436 18552 33798
rect 18616 33522 18644 33866
rect 18604 33516 18656 33522
rect 18604 33458 18656 33464
rect 18472 33408 18552 33436
rect 18420 33390 18472 33396
rect 18328 33108 18380 33114
rect 18328 33050 18380 33056
rect 18432 32910 18460 33390
rect 18604 32972 18656 32978
rect 18604 32914 18656 32920
rect 18420 32904 18472 32910
rect 18420 32846 18472 32852
rect 17960 32438 18012 32444
rect 17684 31476 17736 31482
rect 17408 31340 17460 31346
rect 17408 31282 17460 31288
rect 17316 30864 17368 30870
rect 17316 30806 17368 30812
rect 17132 30728 17184 30734
rect 17132 30670 17184 30676
rect 16764 29504 16816 29510
rect 17040 29504 17092 29510
rect 16816 29464 16988 29492
rect 16764 29446 16816 29452
rect 16856 29164 16908 29170
rect 16856 29106 16908 29112
rect 16488 28552 16540 28558
rect 16488 28494 16540 28500
rect 16580 28484 16632 28490
rect 16580 28426 16632 28432
rect 16592 28150 16620 28426
rect 16580 28144 16632 28150
rect 16580 28086 16632 28092
rect 16592 27674 16620 28086
rect 16672 28076 16724 28082
rect 16672 28018 16724 28024
rect 16764 28076 16816 28082
rect 16764 28018 16816 28024
rect 16684 27674 16712 28018
rect 16580 27668 16632 27674
rect 16580 27610 16632 27616
rect 16672 27668 16724 27674
rect 16672 27610 16724 27616
rect 16580 27532 16632 27538
rect 16580 27474 16632 27480
rect 16592 27130 16620 27474
rect 16776 27470 16804 28018
rect 16672 27464 16724 27470
rect 16672 27406 16724 27412
rect 16764 27464 16816 27470
rect 16764 27406 16816 27412
rect 16684 27130 16712 27406
rect 16580 27124 16632 27130
rect 16580 27066 16632 27072
rect 16672 27124 16724 27130
rect 16672 27066 16724 27072
rect 16488 26240 16540 26246
rect 16408 26200 16488 26228
rect 16488 26182 16540 26188
rect 16592 24818 16620 27066
rect 16868 26382 16896 29106
rect 16960 27130 16988 29464
rect 17040 29446 17092 29452
rect 16948 27124 17000 27130
rect 16948 27066 17000 27072
rect 16960 26926 16988 27066
rect 17052 26994 17080 29446
rect 17144 27470 17172 30670
rect 17224 30592 17276 30598
rect 17224 30534 17276 30540
rect 17236 30190 17264 30534
rect 17224 30184 17276 30190
rect 17224 30126 17276 30132
rect 17224 28416 17276 28422
rect 17224 28358 17276 28364
rect 17132 27464 17184 27470
rect 17132 27406 17184 27412
rect 17236 27130 17264 28358
rect 17328 27470 17356 30806
rect 17420 29170 17448 31282
rect 17512 29646 17540 31470
rect 17684 31418 17736 31424
rect 17592 31340 17644 31346
rect 17592 31282 17644 31288
rect 17604 30938 17632 31282
rect 17592 30932 17644 30938
rect 17592 30874 17644 30880
rect 17500 29640 17552 29646
rect 17500 29582 17552 29588
rect 17408 29164 17460 29170
rect 17408 29106 17460 29112
rect 17696 28994 17724 31418
rect 17880 31346 17908 32422
rect 17868 31340 17920 31346
rect 17868 31282 17920 31288
rect 17972 30734 18000 32438
rect 18156 32422 18276 32450
rect 18420 32428 18472 32434
rect 18156 31754 18184 32422
rect 18420 32370 18472 32376
rect 18236 32360 18288 32366
rect 18236 32302 18288 32308
rect 18144 31748 18196 31754
rect 18144 31690 18196 31696
rect 18144 31204 18196 31210
rect 18144 31146 18196 31152
rect 18052 31136 18104 31142
rect 18052 31078 18104 31084
rect 17960 30728 18012 30734
rect 17960 30670 18012 30676
rect 17960 30592 18012 30598
rect 17960 30534 18012 30540
rect 17972 29238 18000 30534
rect 18064 30258 18092 31078
rect 18156 30666 18184 31146
rect 18144 30660 18196 30666
rect 18144 30602 18196 30608
rect 18142 30288 18198 30297
rect 18052 30252 18104 30258
rect 18142 30223 18144 30232
rect 18052 30194 18104 30200
rect 18196 30223 18198 30232
rect 18144 30194 18196 30200
rect 18052 30048 18104 30054
rect 18052 29990 18104 29996
rect 18064 29782 18092 29990
rect 18052 29776 18104 29782
rect 18248 29730 18276 32302
rect 18432 32065 18460 32370
rect 18418 32056 18474 32065
rect 18418 31991 18474 32000
rect 18420 31340 18472 31346
rect 18420 31282 18472 31288
rect 18328 31136 18380 31142
rect 18328 31078 18380 31084
rect 18340 30433 18368 31078
rect 18326 30424 18382 30433
rect 18326 30359 18382 30368
rect 18432 30161 18460 31282
rect 18616 31124 18644 32914
rect 18708 32570 18736 35430
rect 18800 33862 18828 36042
rect 18880 35692 18932 35698
rect 18880 35634 18932 35640
rect 18892 35290 18920 35634
rect 18880 35284 18932 35290
rect 18880 35226 18932 35232
rect 18788 33856 18840 33862
rect 18788 33798 18840 33804
rect 18880 32904 18932 32910
rect 18880 32846 18932 32852
rect 18788 32836 18840 32842
rect 18788 32778 18840 32784
rect 18696 32564 18748 32570
rect 18696 32506 18748 32512
rect 18800 32416 18828 32778
rect 18892 32570 18920 32846
rect 18880 32564 18932 32570
rect 18880 32506 18932 32512
rect 18880 32428 18932 32434
rect 18800 32388 18880 32416
rect 18880 32370 18932 32376
rect 18696 31952 18748 31958
rect 18696 31894 18748 31900
rect 18878 31920 18934 31929
rect 18708 31482 18736 31894
rect 18878 31855 18934 31864
rect 18892 31822 18920 31855
rect 18788 31816 18840 31822
rect 18788 31758 18840 31764
rect 18880 31816 18932 31822
rect 18880 31758 18932 31764
rect 18800 31482 18828 31758
rect 18696 31476 18748 31482
rect 18696 31418 18748 31424
rect 18788 31476 18840 31482
rect 18788 31418 18840 31424
rect 18788 31340 18840 31346
rect 18984 31328 19012 37062
rect 19352 34950 19380 37742
rect 19892 37188 19944 37194
rect 19892 37130 19944 37136
rect 19708 36644 19760 36650
rect 19708 36586 19760 36592
rect 19340 34944 19392 34950
rect 19340 34886 19392 34892
rect 19720 34105 19748 36586
rect 19904 36378 19932 37130
rect 19892 36372 19944 36378
rect 19892 36314 19944 36320
rect 19800 36236 19852 36242
rect 19800 36178 19852 36184
rect 19812 35562 19840 36178
rect 19904 36106 19932 36314
rect 19892 36100 19944 36106
rect 19892 36042 19944 36048
rect 19800 35556 19852 35562
rect 19800 35498 19852 35504
rect 19706 34096 19762 34105
rect 19706 34031 19762 34040
rect 19338 33688 19394 33697
rect 19338 33623 19340 33632
rect 19392 33623 19394 33632
rect 19720 33640 19748 34031
rect 19720 33612 19840 33640
rect 19340 33594 19392 33600
rect 19708 33516 19760 33522
rect 19708 33458 19760 33464
rect 19064 33448 19116 33454
rect 19064 33390 19116 33396
rect 19340 33448 19392 33454
rect 19340 33390 19392 33396
rect 19616 33448 19668 33454
rect 19616 33390 19668 33396
rect 19076 33289 19104 33390
rect 19062 33280 19118 33289
rect 19062 33215 19118 33224
rect 19352 32978 19380 33390
rect 19524 33380 19576 33386
rect 19524 33322 19576 33328
rect 19340 32972 19392 32978
rect 19340 32914 19392 32920
rect 19536 32842 19564 33322
rect 19628 32978 19656 33390
rect 19720 33046 19748 33458
rect 19708 33040 19760 33046
rect 19708 32982 19760 32988
rect 19616 32972 19668 32978
rect 19616 32914 19668 32920
rect 19340 32836 19392 32842
rect 19340 32778 19392 32784
rect 19524 32836 19576 32842
rect 19524 32778 19576 32784
rect 19062 32328 19118 32337
rect 19062 32263 19064 32272
rect 19116 32263 19118 32272
rect 19064 32234 19116 32240
rect 19064 32020 19116 32026
rect 19064 31962 19116 31968
rect 18840 31300 19012 31328
rect 18788 31282 18840 31288
rect 18788 31136 18840 31142
rect 18616 31096 18788 31124
rect 18788 31078 18840 31084
rect 18512 30932 18564 30938
rect 18512 30874 18564 30880
rect 18524 30258 18552 30874
rect 18604 30660 18656 30666
rect 18604 30602 18656 30608
rect 18616 30258 18644 30602
rect 18800 30258 18828 31078
rect 18880 30864 18932 30870
rect 18880 30806 18932 30812
rect 19076 30818 19104 31962
rect 19156 31748 19208 31754
rect 19156 31690 19208 31696
rect 19168 30938 19196 31690
rect 19248 31340 19300 31346
rect 19248 31282 19300 31288
rect 19156 30932 19208 30938
rect 19156 30874 19208 30880
rect 18892 30394 18920 30806
rect 19076 30790 19196 30818
rect 19062 30696 19118 30705
rect 19062 30631 19064 30640
rect 19116 30631 19118 30640
rect 19064 30602 19116 30608
rect 18880 30388 18932 30394
rect 18880 30330 18932 30336
rect 19168 30326 19196 30790
rect 19260 30734 19288 31282
rect 19352 31249 19380 32778
rect 19432 31476 19484 31482
rect 19432 31418 19484 31424
rect 19338 31240 19394 31249
rect 19338 31175 19394 31184
rect 19444 30977 19472 31418
rect 19430 30968 19486 30977
rect 19430 30903 19486 30912
rect 19248 30728 19300 30734
rect 19248 30670 19300 30676
rect 19156 30320 19208 30326
rect 19156 30262 19208 30268
rect 18512 30252 18564 30258
rect 18512 30194 18564 30200
rect 18604 30252 18656 30258
rect 18604 30194 18656 30200
rect 18788 30252 18840 30258
rect 18788 30194 18840 30200
rect 18696 30184 18748 30190
rect 18418 30152 18474 30161
rect 18696 30126 18748 30132
rect 18418 30087 18474 30096
rect 18604 30116 18656 30122
rect 18604 30058 18656 30064
rect 18328 30048 18380 30054
rect 18328 29990 18380 29996
rect 18052 29718 18104 29724
rect 18156 29702 18276 29730
rect 18156 29646 18184 29702
rect 18340 29646 18368 29990
rect 18144 29640 18196 29646
rect 18144 29582 18196 29588
rect 18328 29640 18380 29646
rect 18328 29582 18380 29588
rect 17960 29232 18012 29238
rect 17960 29174 18012 29180
rect 17696 28966 17908 28994
rect 17880 28558 17908 28966
rect 17868 28552 17920 28558
rect 17868 28494 17920 28500
rect 18052 28552 18104 28558
rect 18052 28494 18104 28500
rect 17500 28212 17552 28218
rect 17500 28154 17552 28160
rect 17592 28212 17644 28218
rect 17592 28154 17644 28160
rect 17408 28144 17460 28150
rect 17406 28112 17408 28121
rect 17460 28112 17462 28121
rect 17406 28047 17462 28056
rect 17512 27470 17540 28154
rect 17316 27464 17368 27470
rect 17316 27406 17368 27412
rect 17408 27464 17460 27470
rect 17408 27406 17460 27412
rect 17500 27464 17552 27470
rect 17500 27406 17552 27412
rect 17316 27328 17368 27334
rect 17316 27270 17368 27276
rect 17420 27316 17448 27406
rect 17604 27316 17632 28154
rect 17880 28082 17908 28494
rect 17868 28076 17920 28082
rect 17868 28018 17920 28024
rect 17960 27396 18012 27402
rect 17960 27338 18012 27344
rect 17420 27288 17632 27316
rect 17776 27328 17828 27334
rect 17328 27130 17356 27270
rect 17224 27124 17276 27130
rect 17224 27066 17276 27072
rect 17316 27124 17368 27130
rect 17316 27066 17368 27072
rect 17040 26988 17092 26994
rect 17040 26930 17092 26936
rect 17144 26948 17356 26976
rect 16948 26920 17000 26926
rect 16948 26862 17000 26868
rect 16856 26376 16908 26382
rect 16856 26318 16908 26324
rect 16764 26240 16816 26246
rect 16764 26182 16816 26188
rect 16672 25152 16724 25158
rect 16672 25094 16724 25100
rect 16580 24812 16632 24818
rect 16580 24754 16632 24760
rect 16684 24750 16712 25094
rect 16672 24744 16724 24750
rect 16316 24704 16436 24732
rect 16224 24636 16344 24664
rect 16120 23656 16172 23662
rect 16120 23598 16172 23604
rect 16212 23520 16264 23526
rect 16212 23462 16264 23468
rect 16120 22976 16172 22982
rect 16120 22918 16172 22924
rect 16132 22642 16160 22918
rect 16120 22636 16172 22642
rect 16120 22578 16172 22584
rect 16028 22160 16080 22166
rect 16028 22102 16080 22108
rect 15752 22024 15804 22030
rect 15752 21966 15804 21972
rect 15844 22024 15896 22030
rect 16040 22001 16068 22102
rect 15844 21966 15896 21972
rect 16026 21992 16082 22001
rect 15566 21584 15622 21593
rect 15292 21548 15344 21554
rect 15292 21490 15344 21496
rect 15476 21548 15528 21554
rect 15566 21519 15622 21528
rect 15660 21548 15712 21554
rect 15476 21490 15528 21496
rect 15488 21350 15516 21490
rect 15384 21344 15436 21350
rect 15384 21286 15436 21292
rect 15476 21344 15528 21350
rect 15476 21286 15528 21292
rect 15396 21026 15424 21286
rect 15580 21078 15608 21519
rect 15660 21490 15712 21496
rect 15672 21350 15700 21490
rect 15660 21344 15712 21350
rect 15660 21286 15712 21292
rect 15568 21072 15620 21078
rect 15396 20998 15516 21026
rect 15568 21014 15620 21020
rect 15290 20632 15346 20641
rect 15200 20596 15252 20602
rect 15290 20567 15346 20576
rect 15200 20538 15252 20544
rect 15108 20052 15160 20058
rect 15108 19994 15160 20000
rect 15200 20052 15252 20058
rect 15200 19994 15252 20000
rect 15212 19854 15240 19994
rect 15200 19848 15252 19854
rect 15200 19790 15252 19796
rect 15106 18456 15162 18465
rect 15106 18391 15162 18400
rect 15120 18358 15148 18391
rect 15108 18352 15160 18358
rect 15108 18294 15160 18300
rect 15304 17882 15332 20567
rect 15396 18426 15424 20998
rect 15488 20924 15516 20998
rect 15568 20936 15620 20942
rect 15488 20896 15568 20924
rect 15568 20878 15620 20884
rect 15566 20632 15622 20641
rect 15566 20567 15622 20576
rect 15476 20392 15528 20398
rect 15476 20334 15528 20340
rect 15488 19990 15516 20334
rect 15580 20058 15608 20567
rect 15568 20052 15620 20058
rect 15568 19994 15620 20000
rect 15476 19984 15528 19990
rect 15476 19926 15528 19932
rect 15476 19508 15528 19514
rect 15476 19450 15528 19456
rect 15384 18420 15436 18426
rect 15384 18362 15436 18368
rect 15384 18216 15436 18222
rect 15384 18158 15436 18164
rect 15292 17876 15344 17882
rect 15292 17818 15344 17824
rect 15396 15026 15424 18158
rect 15488 15706 15516 19450
rect 15672 19334 15700 21286
rect 15764 21078 15792 21966
rect 15856 21434 15884 21966
rect 16026 21927 16082 21936
rect 16028 21888 16080 21894
rect 16132 21876 16160 22578
rect 16224 21962 16252 23462
rect 16316 23186 16344 24636
rect 16408 24342 16436 24704
rect 16672 24686 16724 24692
rect 16396 24336 16448 24342
rect 16396 24278 16448 24284
rect 16684 24206 16712 24686
rect 16672 24200 16724 24206
rect 16670 24168 16672 24177
rect 16724 24168 16726 24177
rect 16670 24103 16726 24112
rect 16672 23656 16724 23662
rect 16672 23598 16724 23604
rect 16304 23180 16356 23186
rect 16304 23122 16356 23128
rect 16684 22642 16712 23598
rect 16672 22636 16724 22642
rect 16672 22578 16724 22584
rect 16396 22568 16448 22574
rect 16448 22528 16528 22556
rect 16396 22510 16448 22516
rect 16304 22160 16356 22166
rect 16304 22102 16356 22108
rect 16212 21956 16264 21962
rect 16212 21898 16264 21904
rect 16080 21848 16160 21876
rect 16028 21830 16080 21836
rect 15856 21406 15976 21434
rect 15752 21072 15804 21078
rect 15752 21014 15804 21020
rect 15948 20942 15976 21406
rect 16040 21350 16068 21830
rect 16316 21690 16344 22102
rect 16500 22030 16528 22528
rect 16396 22024 16448 22030
rect 16396 21966 16448 21972
rect 16488 22024 16540 22030
rect 16488 21966 16540 21972
rect 16304 21684 16356 21690
rect 16304 21626 16356 21632
rect 16028 21344 16080 21350
rect 16028 21286 16080 21292
rect 16120 21344 16172 21350
rect 16120 21286 16172 21292
rect 15936 20936 15988 20942
rect 15936 20878 15988 20884
rect 15752 20868 15804 20874
rect 15752 20810 15804 20816
rect 15764 19514 15792 20810
rect 16040 20788 16068 21286
rect 16132 20942 16160 21286
rect 16120 20936 16172 20942
rect 16120 20878 16172 20884
rect 15948 20760 16068 20788
rect 15844 19712 15896 19718
rect 15844 19654 15896 19660
rect 15856 19514 15884 19654
rect 15752 19508 15804 19514
rect 15752 19450 15804 19456
rect 15844 19508 15896 19514
rect 15844 19450 15896 19456
rect 15672 19306 15884 19334
rect 15660 18760 15712 18766
rect 15660 18702 15712 18708
rect 15672 16658 15700 18702
rect 15752 18216 15804 18222
rect 15856 18204 15884 19306
rect 15948 18834 15976 20760
rect 16040 20534 16068 20760
rect 16212 20800 16264 20806
rect 16212 20742 16264 20748
rect 16304 20800 16356 20806
rect 16304 20742 16356 20748
rect 16028 20528 16080 20534
rect 16028 20470 16080 20476
rect 16028 19848 16080 19854
rect 16028 19790 16080 19796
rect 16040 19553 16068 19790
rect 16120 19712 16172 19718
rect 16224 19700 16252 20742
rect 16316 20398 16344 20742
rect 16304 20392 16356 20398
rect 16304 20334 16356 20340
rect 16304 20256 16356 20262
rect 16304 20198 16356 20204
rect 16316 19854 16344 20198
rect 16304 19848 16356 19854
rect 16304 19790 16356 19796
rect 16172 19672 16252 19700
rect 16120 19654 16172 19660
rect 16026 19544 16082 19553
rect 16026 19479 16082 19488
rect 15936 18828 15988 18834
rect 15936 18770 15988 18776
rect 15936 18216 15988 18222
rect 15856 18176 15936 18204
rect 15752 18158 15804 18164
rect 15936 18158 15988 18164
rect 15764 17338 15792 18158
rect 15844 17672 15896 17678
rect 15844 17614 15896 17620
rect 15752 17332 15804 17338
rect 15752 17274 15804 17280
rect 15764 17202 15792 17274
rect 15752 17196 15804 17202
rect 15752 17138 15804 17144
rect 15856 17066 15884 17614
rect 15844 17060 15896 17066
rect 15844 17002 15896 17008
rect 15660 16652 15712 16658
rect 15580 16612 15660 16640
rect 15476 15700 15528 15706
rect 15476 15642 15528 15648
rect 15580 15162 15608 16612
rect 15660 16594 15712 16600
rect 15856 16538 15884 17002
rect 15764 16510 15884 16538
rect 15764 15502 15792 16510
rect 15948 16436 15976 18158
rect 16040 17678 16068 19479
rect 16132 19446 16160 19654
rect 16120 19440 16172 19446
rect 16120 19382 16172 19388
rect 16132 18290 16160 19382
rect 16316 19174 16344 19790
rect 16408 19310 16436 21966
rect 16500 21554 16528 21966
rect 16488 21548 16540 21554
rect 16488 21490 16540 21496
rect 16684 21078 16712 22578
rect 16776 22166 16804 26182
rect 16856 25152 16908 25158
rect 16856 25094 16908 25100
rect 16868 24818 16896 25094
rect 16856 24812 16908 24818
rect 16856 24754 16908 24760
rect 16948 23044 17000 23050
rect 16948 22986 17000 22992
rect 16856 22636 16908 22642
rect 16856 22578 16908 22584
rect 16764 22160 16816 22166
rect 16764 22102 16816 22108
rect 16764 22024 16816 22030
rect 16762 21992 16764 22001
rect 16816 21992 16818 22001
rect 16762 21927 16818 21936
rect 16764 21412 16816 21418
rect 16764 21354 16816 21360
rect 16776 21146 16804 21354
rect 16764 21140 16816 21146
rect 16764 21082 16816 21088
rect 16672 21072 16724 21078
rect 16672 21014 16724 21020
rect 16578 20632 16634 20641
rect 16578 20567 16634 20576
rect 16592 20466 16620 20567
rect 16684 20482 16712 21014
rect 16580 20460 16632 20466
rect 16684 20454 16804 20482
rect 16580 20402 16632 20408
rect 16580 19984 16632 19990
rect 16580 19926 16632 19932
rect 16488 19848 16540 19854
rect 16488 19790 16540 19796
rect 16396 19304 16448 19310
rect 16396 19246 16448 19252
rect 16304 19168 16356 19174
rect 16304 19110 16356 19116
rect 16212 18624 16264 18630
rect 16212 18566 16264 18572
rect 16120 18284 16172 18290
rect 16120 18226 16172 18232
rect 16224 17746 16252 18566
rect 16212 17740 16264 17746
rect 16212 17682 16264 17688
rect 16028 17672 16080 17678
rect 16080 17632 16160 17660
rect 16028 17614 16080 17620
rect 16028 16788 16080 16794
rect 16028 16730 16080 16736
rect 15856 16408 15976 16436
rect 15856 15502 15884 16408
rect 15752 15496 15804 15502
rect 15752 15438 15804 15444
rect 15844 15496 15896 15502
rect 15844 15438 15896 15444
rect 15936 15496 15988 15502
rect 15936 15438 15988 15444
rect 15660 15428 15712 15434
rect 15660 15370 15712 15376
rect 15568 15156 15620 15162
rect 15568 15098 15620 15104
rect 15384 15020 15436 15026
rect 15384 14962 15436 14968
rect 15580 14618 15608 15098
rect 15568 14612 15620 14618
rect 15568 14554 15620 14560
rect 15292 14408 15344 14414
rect 15292 14350 15344 14356
rect 15108 14000 15160 14006
rect 15108 13942 15160 13948
rect 15120 13326 15148 13942
rect 15200 13932 15252 13938
rect 15200 13874 15252 13880
rect 15108 13320 15160 13326
rect 15108 13262 15160 13268
rect 15212 13258 15240 13874
rect 15304 13530 15332 14350
rect 15568 14340 15620 14346
rect 15568 14282 15620 14288
rect 15580 13870 15608 14282
rect 15568 13864 15620 13870
rect 15568 13806 15620 13812
rect 15672 13734 15700 15370
rect 15948 14618 15976 15438
rect 15936 14612 15988 14618
rect 15936 14554 15988 14560
rect 15660 13728 15712 13734
rect 15660 13670 15712 13676
rect 15292 13524 15344 13530
rect 15292 13466 15344 13472
rect 16040 13326 16068 16730
rect 16132 15094 16160 17632
rect 16212 17604 16264 17610
rect 16212 17546 16264 17552
rect 16224 17513 16252 17546
rect 16210 17504 16266 17513
rect 16210 17439 16266 17448
rect 16212 17332 16264 17338
rect 16212 17274 16264 17280
rect 16120 15088 16172 15094
rect 16120 15030 16172 15036
rect 16132 14278 16160 15030
rect 16224 15026 16252 17274
rect 16316 16454 16344 19110
rect 16500 18290 16528 19790
rect 16592 19786 16620 19926
rect 16776 19904 16804 20454
rect 16868 20058 16896 22578
rect 16960 22574 16988 22986
rect 16948 22568 17000 22574
rect 16948 22510 17000 22516
rect 17052 22030 17080 26930
rect 17144 26858 17172 26948
rect 17132 26852 17184 26858
rect 17132 26794 17184 26800
rect 17224 26852 17276 26858
rect 17224 26794 17276 26800
rect 17130 26752 17186 26761
rect 17130 26687 17186 26696
rect 17144 26042 17172 26687
rect 17236 26518 17264 26794
rect 17224 26512 17276 26518
rect 17224 26454 17276 26460
rect 17224 26376 17276 26382
rect 17224 26318 17276 26324
rect 17132 26036 17184 26042
rect 17132 25978 17184 25984
rect 17132 25900 17184 25906
rect 17132 25842 17184 25848
rect 17144 24682 17172 25842
rect 17236 25498 17264 26318
rect 17224 25492 17276 25498
rect 17224 25434 17276 25440
rect 17328 25294 17356 26948
rect 17420 25838 17448 27288
rect 17776 27270 17828 27276
rect 17684 26784 17736 26790
rect 17684 26726 17736 26732
rect 17696 26586 17724 26726
rect 17788 26625 17816 27270
rect 17774 26616 17830 26625
rect 17684 26580 17736 26586
rect 17774 26551 17830 26560
rect 17684 26522 17736 26528
rect 17592 26512 17644 26518
rect 17592 26454 17644 26460
rect 17604 26081 17632 26454
rect 17972 26194 18000 27338
rect 18064 26586 18092 28494
rect 18156 27470 18184 29582
rect 18512 29572 18564 29578
rect 18512 29514 18564 29520
rect 18420 29504 18472 29510
rect 18418 29472 18420 29481
rect 18472 29472 18474 29481
rect 18418 29407 18474 29416
rect 18234 29200 18290 29209
rect 18234 29135 18290 29144
rect 18144 27464 18196 27470
rect 18144 27406 18196 27412
rect 18144 26784 18196 26790
rect 18144 26726 18196 26732
rect 18052 26580 18104 26586
rect 18052 26522 18104 26528
rect 17788 26166 18000 26194
rect 17590 26072 17646 26081
rect 17590 26007 17646 26016
rect 17408 25832 17460 25838
rect 17408 25774 17460 25780
rect 17316 25288 17368 25294
rect 17316 25230 17368 25236
rect 17316 24880 17368 24886
rect 17316 24822 17368 24828
rect 17132 24676 17184 24682
rect 17132 24618 17184 24624
rect 17224 24676 17276 24682
rect 17224 24618 17276 24624
rect 17236 24342 17264 24618
rect 17224 24336 17276 24342
rect 17224 24278 17276 24284
rect 17236 24206 17264 24278
rect 17328 24256 17356 24822
rect 17420 24410 17448 25774
rect 17500 25152 17552 25158
rect 17500 25094 17552 25100
rect 17512 24750 17540 25094
rect 17604 24818 17632 26007
rect 17684 25152 17736 25158
rect 17684 25094 17736 25100
rect 17696 24954 17724 25094
rect 17684 24948 17736 24954
rect 17684 24890 17736 24896
rect 17592 24812 17644 24818
rect 17592 24754 17644 24760
rect 17500 24744 17552 24750
rect 17500 24686 17552 24692
rect 17408 24404 17460 24410
rect 17408 24346 17460 24352
rect 17512 24290 17540 24686
rect 17696 24682 17724 24890
rect 17684 24676 17736 24682
rect 17684 24618 17736 24624
rect 17512 24274 17724 24290
rect 17408 24268 17460 24274
rect 17328 24228 17408 24256
rect 17408 24210 17460 24216
rect 17512 24268 17736 24274
rect 17512 24262 17684 24268
rect 17224 24200 17276 24206
rect 17224 24142 17276 24148
rect 17236 23662 17264 24142
rect 17224 23656 17276 23662
rect 17224 23598 17276 23604
rect 17132 23112 17184 23118
rect 17132 23054 17184 23060
rect 17144 22642 17172 23054
rect 17236 23050 17264 23598
rect 17512 23526 17540 24262
rect 17684 24210 17736 24216
rect 17592 24200 17644 24206
rect 17592 24142 17644 24148
rect 17316 23520 17368 23526
rect 17316 23462 17368 23468
rect 17500 23520 17552 23526
rect 17500 23462 17552 23468
rect 17328 23118 17356 23462
rect 17604 23118 17632 24142
rect 17684 23656 17736 23662
rect 17684 23598 17736 23604
rect 17696 23118 17724 23598
rect 17316 23112 17368 23118
rect 17316 23054 17368 23060
rect 17592 23112 17644 23118
rect 17592 23054 17644 23060
rect 17684 23112 17736 23118
rect 17684 23054 17736 23060
rect 17224 23044 17276 23050
rect 17224 22986 17276 22992
rect 17132 22636 17184 22642
rect 17132 22578 17184 22584
rect 16948 22024 17000 22030
rect 16948 21966 17000 21972
rect 17040 22024 17092 22030
rect 17040 21966 17092 21972
rect 16960 21486 16988 21966
rect 16948 21480 17000 21486
rect 16948 21422 17000 21428
rect 16960 20942 16988 21422
rect 17052 21146 17080 21966
rect 17328 21690 17356 23054
rect 17604 22642 17632 23054
rect 17592 22636 17644 22642
rect 17592 22578 17644 22584
rect 17316 21684 17368 21690
rect 17604 21672 17632 22578
rect 17316 21626 17368 21632
rect 17512 21644 17632 21672
rect 17132 21548 17184 21554
rect 17132 21490 17184 21496
rect 17040 21140 17092 21146
rect 17040 21082 17092 21088
rect 17144 20942 17172 21490
rect 16948 20936 17000 20942
rect 16948 20878 17000 20884
rect 17132 20936 17184 20942
rect 17132 20878 17184 20884
rect 16856 20052 16908 20058
rect 16856 19994 16908 20000
rect 16776 19876 16896 19904
rect 16580 19780 16632 19786
rect 16580 19722 16632 19728
rect 16488 18284 16540 18290
rect 16488 18226 16540 18232
rect 16764 18284 16816 18290
rect 16764 18226 16816 18232
rect 16396 17672 16448 17678
rect 16396 17614 16448 17620
rect 16488 17672 16540 17678
rect 16488 17614 16540 17620
rect 16580 17672 16632 17678
rect 16580 17614 16632 17620
rect 16408 17542 16436 17614
rect 16500 17542 16528 17614
rect 16396 17536 16448 17542
rect 16396 17478 16448 17484
rect 16488 17536 16540 17542
rect 16488 17478 16540 17484
rect 16592 17338 16620 17614
rect 16580 17332 16632 17338
rect 16580 17274 16632 17280
rect 16396 17060 16448 17066
rect 16396 17002 16448 17008
rect 16408 16658 16436 17002
rect 16672 16992 16724 16998
rect 16672 16934 16724 16940
rect 16684 16794 16712 16934
rect 16580 16788 16632 16794
rect 16580 16730 16632 16736
rect 16672 16788 16724 16794
rect 16672 16730 16724 16736
rect 16592 16697 16620 16730
rect 16578 16688 16634 16697
rect 16396 16652 16448 16658
rect 16578 16623 16634 16632
rect 16396 16594 16448 16600
rect 16684 16590 16712 16730
rect 16672 16584 16724 16590
rect 16672 16526 16724 16532
rect 16580 16516 16632 16522
rect 16580 16458 16632 16464
rect 16304 16448 16356 16454
rect 16592 16402 16620 16458
rect 16304 16390 16356 16396
rect 16212 15020 16264 15026
rect 16212 14962 16264 14968
rect 16316 14958 16344 16390
rect 16500 16374 16620 16402
rect 16396 16108 16448 16114
rect 16396 16050 16448 16056
rect 16408 15570 16436 16050
rect 16500 15570 16528 16374
rect 16684 16250 16712 16526
rect 16672 16244 16724 16250
rect 16672 16186 16724 16192
rect 16776 16182 16804 18226
rect 16868 17202 16896 19876
rect 16960 18290 16988 20878
rect 17040 20800 17092 20806
rect 17040 20742 17092 20748
rect 17052 20641 17080 20742
rect 17038 20632 17094 20641
rect 17038 20567 17094 20576
rect 17144 18766 17172 20878
rect 17408 20868 17460 20874
rect 17408 20810 17460 20816
rect 17316 20460 17368 20466
rect 17316 20402 17368 20408
rect 17224 19236 17276 19242
rect 17224 19178 17276 19184
rect 17236 18970 17264 19178
rect 17224 18964 17276 18970
rect 17224 18906 17276 18912
rect 17132 18760 17184 18766
rect 17132 18702 17184 18708
rect 17040 18692 17092 18698
rect 17040 18634 17092 18640
rect 16948 18284 17000 18290
rect 16948 18226 17000 18232
rect 16960 17513 16988 18226
rect 17052 17610 17080 18634
rect 17144 18578 17172 18702
rect 17144 18550 17264 18578
rect 17130 18456 17186 18465
rect 17130 18391 17186 18400
rect 17040 17604 17092 17610
rect 17040 17546 17092 17552
rect 16946 17504 17002 17513
rect 16946 17439 17002 17448
rect 16856 17196 16908 17202
rect 16856 17138 16908 17144
rect 16764 16176 16816 16182
rect 16764 16118 16816 16124
rect 16764 15972 16816 15978
rect 16764 15914 16816 15920
rect 16672 15904 16724 15910
rect 16672 15846 16724 15852
rect 16396 15564 16448 15570
rect 16396 15506 16448 15512
rect 16488 15564 16540 15570
rect 16488 15506 16540 15512
rect 16408 15162 16436 15506
rect 16396 15156 16448 15162
rect 16396 15098 16448 15104
rect 16488 15156 16540 15162
rect 16488 15098 16540 15104
rect 16304 14952 16356 14958
rect 16304 14894 16356 14900
rect 16396 14816 16448 14822
rect 16396 14758 16448 14764
rect 16408 14482 16436 14758
rect 16396 14476 16448 14482
rect 16396 14418 16448 14424
rect 16500 14414 16528 15098
rect 16580 14816 16632 14822
rect 16580 14758 16632 14764
rect 16592 14618 16620 14758
rect 16580 14612 16632 14618
rect 16580 14554 16632 14560
rect 16684 14414 16712 15846
rect 16488 14408 16540 14414
rect 16488 14350 16540 14356
rect 16672 14408 16724 14414
rect 16672 14350 16724 14356
rect 16120 14272 16172 14278
rect 16120 14214 16172 14220
rect 16028 13320 16080 13326
rect 16028 13262 16080 13268
rect 15200 13252 15252 13258
rect 15200 13194 15252 13200
rect 15212 12986 15240 13194
rect 15476 13184 15528 13190
rect 15476 13126 15528 13132
rect 15200 12980 15252 12986
rect 15200 12922 15252 12928
rect 15292 12844 15344 12850
rect 15292 12786 15344 12792
rect 15028 12702 15240 12730
rect 15108 12640 15160 12646
rect 15028 12588 15108 12594
rect 15028 12582 15160 12588
rect 15028 12566 15148 12582
rect 15028 12434 15056 12566
rect 15212 12458 15240 12702
rect 14844 12406 15056 12434
rect 15120 12430 15240 12458
rect 14844 12238 14872 12406
rect 15120 12322 15148 12430
rect 15028 12294 15148 12322
rect 14832 12232 14884 12238
rect 14832 12174 14884 12180
rect 14832 11756 14884 11762
rect 14832 11698 14884 11704
rect 14740 11688 14792 11694
rect 14740 11630 14792 11636
rect 14844 11218 14872 11698
rect 14648 11212 14700 11218
rect 14648 11154 14700 11160
rect 14832 11212 14884 11218
rect 14832 11154 14884 11160
rect 15028 10690 15056 12294
rect 15108 12232 15160 12238
rect 15108 12174 15160 12180
rect 15120 11014 15148 12174
rect 15304 12102 15332 12786
rect 15292 12096 15344 12102
rect 15292 12038 15344 12044
rect 15292 11892 15344 11898
rect 15292 11834 15344 11840
rect 15108 11008 15160 11014
rect 15108 10950 15160 10956
rect 15120 10810 15148 10950
rect 15108 10804 15160 10810
rect 15108 10746 15160 10752
rect 15028 10662 15148 10690
rect 15304 10674 15332 11834
rect 14464 10260 14516 10266
rect 14464 10202 14516 10208
rect 14108 9646 14228 9674
rect 14004 7948 14056 7954
rect 14004 7890 14056 7896
rect 13728 6860 13780 6866
rect 13728 6802 13780 6808
rect 13544 6316 13596 6322
rect 13544 6258 13596 6264
rect 14108 5914 14136 9646
rect 14476 9110 14504 10202
rect 14464 9104 14516 9110
rect 14464 9046 14516 9052
rect 15016 8968 15068 8974
rect 15016 8910 15068 8916
rect 14740 8832 14792 8838
rect 14740 8774 14792 8780
rect 14924 8832 14976 8838
rect 14924 8774 14976 8780
rect 14188 7404 14240 7410
rect 14188 7346 14240 7352
rect 14464 7404 14516 7410
rect 14464 7346 14516 7352
rect 14096 5908 14148 5914
rect 14096 5850 14148 5856
rect 12992 5704 13044 5710
rect 12992 5646 13044 5652
rect 12900 5228 12952 5234
rect 12636 5188 12900 5216
rect 12900 5170 12952 5176
rect 12440 4820 12492 4826
rect 12440 4762 12492 4768
rect 12164 4684 12216 4690
rect 12164 4626 12216 4632
rect 10232 4616 10284 4622
rect 10232 4558 10284 4564
rect 12912 4554 12940 5170
rect 13004 5166 13032 5646
rect 14200 5642 14228 7346
rect 14476 6458 14504 7346
rect 14556 6656 14608 6662
rect 14556 6598 14608 6604
rect 14464 6452 14516 6458
rect 14464 6394 14516 6400
rect 14568 5710 14596 6598
rect 14556 5704 14608 5710
rect 14556 5646 14608 5652
rect 14188 5636 14240 5642
rect 14188 5578 14240 5584
rect 13636 5568 13688 5574
rect 13636 5510 13688 5516
rect 14372 5568 14424 5574
rect 14372 5510 14424 5516
rect 13648 5302 13676 5510
rect 13636 5296 13688 5302
rect 13636 5238 13688 5244
rect 12992 5160 13044 5166
rect 12992 5102 13044 5108
rect 12900 4548 12952 4554
rect 12900 4490 12952 4496
rect 14384 4146 14412 5510
rect 14464 4548 14516 4554
rect 14464 4490 14516 4496
rect 14476 4282 14504 4490
rect 14464 4276 14516 4282
rect 14464 4218 14516 4224
rect 14372 4140 14424 4146
rect 14372 4082 14424 4088
rect 12530 4040 12586 4049
rect 12530 3975 12586 3984
rect 13174 4040 13230 4049
rect 13174 3975 13230 3984
rect 12544 3058 12572 3975
rect 13188 3058 13216 3975
rect 12532 3052 12584 3058
rect 12532 2994 12584 3000
rect 13176 3052 13228 3058
rect 13176 2994 13228 3000
rect 12992 2848 13044 2854
rect 12992 2790 13044 2796
rect 10140 2644 10192 2650
rect 10140 2586 10192 2592
rect 8944 2508 8996 2514
rect 8944 2450 8996 2456
rect 13004 2446 13032 2790
rect 14752 2774 14780 8774
rect 14936 8430 14964 8774
rect 15028 8566 15056 8910
rect 15016 8560 15068 8566
rect 15016 8502 15068 8508
rect 14924 8424 14976 8430
rect 14924 8366 14976 8372
rect 14924 7268 14976 7274
rect 14924 7210 14976 7216
rect 14936 5778 14964 7210
rect 14924 5772 14976 5778
rect 14924 5714 14976 5720
rect 15120 3058 15148 10662
rect 15292 10668 15344 10674
rect 15292 10610 15344 10616
rect 15292 9716 15344 9722
rect 15292 9658 15344 9664
rect 15304 8974 15332 9658
rect 15382 9480 15438 9489
rect 15382 9415 15438 9424
rect 15396 9042 15424 9415
rect 15384 9036 15436 9042
rect 15384 8978 15436 8984
rect 15292 8968 15344 8974
rect 15292 8910 15344 8916
rect 15384 7744 15436 7750
rect 15384 7686 15436 7692
rect 15396 7546 15424 7686
rect 15384 7540 15436 7546
rect 15384 7482 15436 7488
rect 15292 7472 15344 7478
rect 15344 7420 15424 7426
rect 15292 7414 15424 7420
rect 15304 7398 15424 7414
rect 15292 7336 15344 7342
rect 15292 7278 15344 7284
rect 15200 6792 15252 6798
rect 15200 6734 15252 6740
rect 15212 6322 15240 6734
rect 15304 6322 15332 7278
rect 15396 6474 15424 7398
rect 15488 7274 15516 13126
rect 15844 12844 15896 12850
rect 15844 12786 15896 12792
rect 15856 12322 15884 12786
rect 15672 12300 15884 12322
rect 15672 12294 15752 12300
rect 15568 11552 15620 11558
rect 15568 11494 15620 11500
rect 15580 11150 15608 11494
rect 15568 11144 15620 11150
rect 15568 11086 15620 11092
rect 15672 10962 15700 12294
rect 15804 12294 15884 12300
rect 15752 12242 15804 12248
rect 15844 11824 15896 11830
rect 15844 11766 15896 11772
rect 15580 10934 15700 10962
rect 15752 11008 15804 11014
rect 15752 10950 15804 10956
rect 15580 9586 15608 10934
rect 15568 9580 15620 9586
rect 15568 9522 15620 9528
rect 15764 8974 15792 10950
rect 15856 9450 15884 11766
rect 16132 11354 16160 14214
rect 16684 13258 16712 14350
rect 16776 14074 16804 15914
rect 16764 14068 16816 14074
rect 16764 14010 16816 14016
rect 16868 13530 16896 17138
rect 16960 16454 16988 17439
rect 16948 16448 17000 16454
rect 16948 16390 17000 16396
rect 16960 14346 16988 16390
rect 17040 15020 17092 15026
rect 17040 14962 17092 14968
rect 17052 14618 17080 14962
rect 17040 14612 17092 14618
rect 17040 14554 17092 14560
rect 16948 14340 17000 14346
rect 16948 14282 17000 14288
rect 16856 13524 16908 13530
rect 16856 13466 16908 13472
rect 16764 13456 16816 13462
rect 16764 13398 16816 13404
rect 16672 13252 16724 13258
rect 16672 13194 16724 13200
rect 16488 12232 16540 12238
rect 16488 12174 16540 12180
rect 16120 11348 16172 11354
rect 16120 11290 16172 11296
rect 16132 10742 16160 11290
rect 16500 11014 16528 12174
rect 16488 11008 16540 11014
rect 16488 10950 16540 10956
rect 16120 10736 16172 10742
rect 16120 10678 16172 10684
rect 16028 9716 16080 9722
rect 16500 9704 16528 10950
rect 16672 10056 16724 10062
rect 16672 9998 16724 10004
rect 16500 9676 16620 9704
rect 16028 9658 16080 9664
rect 15936 9580 15988 9586
rect 15936 9522 15988 9528
rect 15948 9450 15976 9522
rect 15844 9444 15896 9450
rect 15844 9386 15896 9392
rect 15936 9444 15988 9450
rect 15936 9386 15988 9392
rect 15752 8968 15804 8974
rect 15752 8910 15804 8916
rect 15856 8922 15884 9386
rect 15476 7268 15528 7274
rect 15476 7210 15528 7216
rect 15568 7200 15620 7206
rect 15568 7142 15620 7148
rect 15580 7002 15608 7142
rect 15568 6996 15620 7002
rect 15568 6938 15620 6944
rect 15764 6866 15792 8910
rect 15856 8894 15976 8922
rect 16040 8906 16068 9658
rect 15948 7954 15976 8894
rect 16028 8900 16080 8906
rect 16592 8888 16620 9676
rect 16684 9586 16712 9998
rect 16776 9674 16804 13398
rect 16868 13258 16896 13466
rect 16960 13394 16988 14282
rect 16948 13388 17000 13394
rect 16948 13330 17000 13336
rect 16856 13252 16908 13258
rect 16856 13194 16908 13200
rect 16856 12844 16908 12850
rect 16856 12786 16908 12792
rect 16868 12442 16896 12786
rect 16856 12436 16908 12442
rect 16856 12378 16908 12384
rect 17144 10674 17172 18391
rect 17236 17678 17264 18550
rect 17328 17678 17356 20402
rect 17420 19854 17448 20810
rect 17408 19848 17460 19854
rect 17408 19790 17460 19796
rect 17420 19378 17448 19790
rect 17408 19372 17460 19378
rect 17408 19314 17460 19320
rect 17224 17672 17276 17678
rect 17224 17614 17276 17620
rect 17316 17672 17368 17678
rect 17316 17614 17368 17620
rect 17328 17202 17356 17614
rect 17512 17542 17540 21644
rect 17592 21548 17644 21554
rect 17592 21490 17644 21496
rect 17500 17536 17552 17542
rect 17500 17478 17552 17484
rect 17316 17196 17368 17202
rect 17316 17138 17368 17144
rect 17512 17134 17540 17478
rect 17500 17128 17552 17134
rect 17500 17070 17552 17076
rect 17408 16516 17460 16522
rect 17408 16458 17460 16464
rect 17316 16176 17368 16182
rect 17316 16118 17368 16124
rect 17328 14414 17356 16118
rect 17420 14618 17448 16458
rect 17512 16046 17540 17070
rect 17604 16590 17632 21490
rect 17696 20058 17724 23054
rect 17684 20052 17736 20058
rect 17684 19994 17736 20000
rect 17684 18760 17736 18766
rect 17684 18702 17736 18708
rect 17696 17882 17724 18702
rect 17684 17876 17736 17882
rect 17684 17818 17736 17824
rect 17684 16992 17736 16998
rect 17684 16934 17736 16940
rect 17592 16584 17644 16590
rect 17592 16526 17644 16532
rect 17696 16454 17724 16934
rect 17684 16448 17736 16454
rect 17684 16390 17736 16396
rect 17500 16040 17552 16046
rect 17500 15982 17552 15988
rect 17408 14612 17460 14618
rect 17408 14554 17460 14560
rect 17316 14408 17368 14414
rect 17316 14350 17368 14356
rect 17328 13938 17356 14350
rect 17512 14006 17540 15982
rect 17592 15972 17644 15978
rect 17592 15914 17644 15920
rect 17604 15026 17632 15914
rect 17788 15706 17816 26166
rect 17868 25900 17920 25906
rect 17868 25842 17920 25848
rect 18052 25900 18104 25906
rect 18052 25842 18104 25848
rect 17880 25242 17908 25842
rect 17880 25214 18000 25242
rect 17972 25158 18000 25214
rect 17960 25152 18012 25158
rect 17960 25094 18012 25100
rect 18064 24886 18092 25842
rect 18156 24954 18184 26726
rect 18248 25770 18276 29135
rect 18328 28960 18380 28966
rect 18328 28902 18380 28908
rect 18340 28626 18368 28902
rect 18328 28620 18380 28626
rect 18328 28562 18380 28568
rect 18328 28076 18380 28082
rect 18328 28018 18380 28024
rect 18340 27606 18368 28018
rect 18524 27606 18552 29514
rect 18616 29170 18644 30058
rect 18708 29850 18736 30126
rect 18696 29844 18748 29850
rect 18696 29786 18748 29792
rect 18696 29640 18748 29646
rect 18696 29582 18748 29588
rect 18708 29306 18736 29582
rect 18696 29300 18748 29306
rect 18696 29242 18748 29248
rect 18604 29164 18656 29170
rect 18656 29124 18736 29152
rect 18604 29106 18656 29112
rect 18604 28960 18656 28966
rect 18604 28902 18656 28908
rect 18328 27600 18380 27606
rect 18328 27542 18380 27548
rect 18512 27600 18564 27606
rect 18512 27542 18564 27548
rect 18512 27396 18564 27402
rect 18512 27338 18564 27344
rect 18524 27130 18552 27338
rect 18512 27124 18564 27130
rect 18512 27066 18564 27072
rect 18512 26920 18564 26926
rect 18512 26862 18564 26868
rect 18328 26512 18380 26518
rect 18328 26454 18380 26460
rect 18340 25974 18368 26454
rect 18328 25968 18380 25974
rect 18328 25910 18380 25916
rect 18236 25764 18288 25770
rect 18236 25706 18288 25712
rect 18524 25294 18552 26862
rect 18616 26790 18644 28902
rect 18708 27538 18736 29124
rect 18800 28218 18828 30194
rect 18972 29776 19024 29782
rect 18972 29718 19024 29724
rect 18880 29640 18932 29646
rect 18878 29608 18880 29617
rect 18932 29608 18934 29617
rect 18878 29543 18934 29552
rect 18880 29504 18932 29510
rect 18880 29446 18932 29452
rect 18892 29073 18920 29446
rect 18984 29238 19012 29718
rect 19064 29504 19116 29510
rect 19064 29446 19116 29452
rect 18972 29232 19024 29238
rect 18972 29174 19024 29180
rect 18878 29064 18934 29073
rect 18878 28999 18934 29008
rect 18788 28212 18840 28218
rect 18788 28154 18840 28160
rect 18880 28076 18932 28082
rect 18880 28018 18932 28024
rect 18696 27532 18748 27538
rect 18696 27474 18748 27480
rect 18708 27130 18736 27474
rect 18788 27328 18840 27334
rect 18788 27270 18840 27276
rect 18696 27124 18748 27130
rect 18696 27066 18748 27072
rect 18604 26784 18656 26790
rect 18604 26726 18656 26732
rect 18696 26376 18748 26382
rect 18800 26353 18828 27270
rect 18696 26318 18748 26324
rect 18786 26344 18842 26353
rect 18708 25906 18736 26318
rect 18786 26279 18842 26288
rect 18696 25900 18748 25906
rect 18696 25842 18748 25848
rect 18604 25764 18656 25770
rect 18604 25706 18656 25712
rect 18420 25288 18472 25294
rect 18420 25230 18472 25236
rect 18512 25288 18564 25294
rect 18512 25230 18564 25236
rect 18144 24948 18196 24954
rect 18144 24890 18196 24896
rect 18052 24880 18104 24886
rect 18052 24822 18104 24828
rect 17868 24336 17920 24342
rect 17868 24278 17920 24284
rect 17880 24177 17908 24278
rect 17866 24168 17922 24177
rect 17866 24103 17922 24112
rect 17960 24132 18012 24138
rect 17960 24074 18012 24080
rect 17868 23792 17920 23798
rect 17868 23734 17920 23740
rect 17880 23526 17908 23734
rect 17868 23520 17920 23526
rect 17868 23462 17920 23468
rect 17880 23118 17908 23462
rect 17972 23186 18000 24074
rect 18156 24070 18184 24890
rect 18432 24614 18460 25230
rect 18524 24886 18552 25230
rect 18512 24880 18564 24886
rect 18512 24822 18564 24828
rect 18420 24608 18472 24614
rect 18420 24550 18472 24556
rect 18432 24206 18460 24550
rect 18420 24200 18472 24206
rect 18420 24142 18472 24148
rect 18144 24064 18196 24070
rect 18144 24006 18196 24012
rect 18052 23520 18104 23526
rect 18050 23488 18052 23497
rect 18104 23488 18106 23497
rect 18050 23423 18106 23432
rect 17960 23180 18012 23186
rect 17960 23122 18012 23128
rect 17868 23112 17920 23118
rect 17868 23054 17920 23060
rect 18144 22500 18196 22506
rect 18144 22442 18196 22448
rect 17868 22092 17920 22098
rect 17868 22034 17920 22040
rect 17880 21690 17908 22034
rect 18052 22024 18104 22030
rect 18052 21966 18104 21972
rect 17868 21684 17920 21690
rect 17868 21626 17920 21632
rect 17868 21072 17920 21078
rect 17868 21014 17920 21020
rect 17880 20806 17908 21014
rect 17960 20936 18012 20942
rect 17960 20878 18012 20884
rect 17868 20800 17920 20806
rect 17868 20742 17920 20748
rect 17868 19848 17920 19854
rect 17972 19836 18000 20878
rect 18064 20505 18092 21966
rect 18156 21622 18184 22442
rect 18144 21616 18196 21622
rect 18144 21558 18196 21564
rect 18144 21480 18196 21486
rect 18144 21422 18196 21428
rect 18050 20496 18106 20505
rect 18156 20466 18184 21422
rect 18432 21146 18460 24142
rect 18524 22778 18552 24822
rect 18616 23866 18644 25706
rect 18788 24812 18840 24818
rect 18892 24800 18920 28018
rect 18972 27464 19024 27470
rect 18972 27406 19024 27412
rect 18984 27130 19012 27406
rect 18972 27124 19024 27130
rect 18972 27066 19024 27072
rect 18972 26920 19024 26926
rect 18970 26888 18972 26897
rect 19024 26888 19026 26897
rect 18970 26823 19026 26832
rect 19076 26738 19104 29446
rect 19168 28966 19196 30262
rect 19156 28960 19208 28966
rect 19156 28902 19208 28908
rect 19260 28150 19288 30670
rect 19432 30048 19484 30054
rect 19432 29990 19484 29996
rect 19338 29336 19394 29345
rect 19338 29271 19394 29280
rect 19352 28694 19380 29271
rect 19340 28688 19392 28694
rect 19340 28630 19392 28636
rect 19444 28506 19472 29990
rect 19352 28478 19472 28506
rect 19248 28144 19300 28150
rect 19248 28086 19300 28092
rect 19246 27976 19302 27985
rect 19246 27911 19302 27920
rect 19260 27878 19288 27911
rect 19248 27872 19300 27878
rect 19248 27814 19300 27820
rect 18984 26710 19104 26738
rect 18984 26382 19012 26710
rect 19154 26616 19210 26625
rect 19076 26574 19154 26602
rect 18972 26376 19024 26382
rect 18972 26318 19024 26324
rect 18972 26240 19024 26246
rect 18972 26182 19024 26188
rect 18984 25974 19012 26182
rect 18972 25968 19024 25974
rect 18972 25910 19024 25916
rect 18972 25424 19024 25430
rect 18972 25366 19024 25372
rect 18840 24772 18920 24800
rect 18788 24754 18840 24760
rect 18696 24200 18748 24206
rect 18696 24142 18748 24148
rect 18708 23866 18736 24142
rect 18604 23860 18656 23866
rect 18604 23802 18656 23808
rect 18696 23860 18748 23866
rect 18696 23802 18748 23808
rect 18512 22772 18564 22778
rect 18512 22714 18564 22720
rect 18800 22094 18828 24754
rect 18880 24608 18932 24614
rect 18880 24550 18932 24556
rect 18892 24206 18920 24550
rect 18880 24200 18932 24206
rect 18880 24142 18932 24148
rect 18984 23866 19012 25366
rect 19076 25362 19104 26574
rect 19154 26551 19210 26560
rect 19352 26518 19380 28478
rect 19536 28472 19564 32778
rect 19616 31680 19668 31686
rect 19616 31622 19668 31628
rect 19628 31346 19656 31622
rect 19812 31482 19840 33612
rect 19892 33380 19944 33386
rect 19892 33322 19944 33328
rect 19904 31686 19932 33322
rect 19996 33153 20024 37742
rect 20364 37466 20392 37810
rect 20548 37738 20576 37878
rect 20536 37732 20588 37738
rect 20536 37674 20588 37680
rect 20352 37460 20404 37466
rect 20352 37402 20404 37408
rect 20168 37256 20220 37262
rect 20168 37198 20220 37204
rect 20180 36009 20208 37198
rect 20720 37188 20772 37194
rect 20720 37130 20772 37136
rect 20732 36922 20760 37130
rect 20720 36916 20772 36922
rect 20720 36858 20772 36864
rect 20536 36100 20588 36106
rect 20536 36042 20588 36048
rect 20166 36000 20222 36009
rect 20166 35935 20222 35944
rect 20444 35760 20496 35766
rect 20444 35702 20496 35708
rect 20076 35692 20128 35698
rect 20076 35634 20128 35640
rect 19982 33144 20038 33153
rect 19982 33079 20038 33088
rect 19984 32904 20036 32910
rect 19984 32846 20036 32852
rect 19996 32774 20024 32846
rect 19984 32768 20036 32774
rect 19984 32710 20036 32716
rect 19984 32564 20036 32570
rect 19984 32506 20036 32512
rect 19892 31680 19944 31686
rect 19892 31622 19944 31628
rect 19800 31476 19852 31482
rect 19800 31418 19852 31424
rect 19996 31414 20024 32506
rect 19984 31408 20036 31414
rect 19984 31350 20036 31356
rect 19616 31340 19668 31346
rect 19616 31282 19668 31288
rect 19996 31113 20024 31350
rect 19982 31104 20038 31113
rect 19982 31039 20038 31048
rect 20088 30734 20116 35634
rect 20168 34060 20220 34066
rect 20168 34002 20220 34008
rect 20180 33561 20208 34002
rect 20260 33992 20312 33998
rect 20258 33960 20260 33969
rect 20312 33960 20314 33969
rect 20258 33895 20314 33904
rect 20352 33856 20404 33862
rect 20352 33798 20404 33804
rect 20260 33652 20312 33658
rect 20260 33594 20312 33600
rect 20166 33552 20222 33561
rect 20166 33487 20222 33496
rect 20272 32994 20300 33594
rect 20364 33522 20392 33798
rect 20352 33516 20404 33522
rect 20352 33458 20404 33464
rect 20456 33318 20484 35702
rect 20548 34202 20576 36042
rect 21008 35834 21036 37946
rect 21192 37806 21220 38286
rect 21284 38010 21312 38286
rect 22480 38162 22508 38490
rect 25778 38448 25834 38457
rect 27632 38418 27660 38694
rect 27724 38554 27752 38898
rect 29736 38820 29788 38826
rect 29736 38762 29788 38768
rect 27712 38548 27764 38554
rect 27712 38490 27764 38496
rect 25778 38383 25834 38392
rect 26056 38412 26108 38418
rect 25596 38276 25648 38282
rect 25596 38218 25648 38224
rect 23480 38208 23532 38214
rect 22480 38134 22600 38162
rect 23480 38150 23532 38156
rect 21272 38004 21324 38010
rect 21272 37946 21324 37952
rect 22572 37806 22600 38134
rect 23492 37874 23520 38150
rect 25608 38010 25636 38218
rect 25596 38004 25648 38010
rect 25596 37946 25648 37952
rect 25792 37942 25820 38383
rect 26056 38354 26108 38360
rect 27620 38412 27672 38418
rect 27620 38354 27672 38360
rect 29644 38412 29696 38418
rect 29644 38354 29696 38360
rect 26068 38282 26096 38354
rect 29552 38344 29604 38350
rect 29552 38286 29604 38292
rect 26056 38276 26108 38282
rect 26056 38218 26108 38224
rect 27528 38276 27580 38282
rect 27528 38218 27580 38224
rect 29276 38276 29328 38282
rect 29276 38218 29328 38224
rect 29460 38276 29512 38282
rect 29460 38218 29512 38224
rect 26516 38208 26568 38214
rect 26516 38150 26568 38156
rect 25780 37936 25832 37942
rect 25318 37904 25374 37913
rect 23020 37868 23072 37874
rect 23020 37810 23072 37816
rect 23480 37868 23532 37874
rect 23480 37810 23532 37816
rect 23664 37868 23716 37874
rect 23664 37810 23716 37816
rect 23940 37868 23992 37874
rect 23940 37810 23992 37816
rect 24124 37868 24176 37874
rect 25780 37878 25832 37884
rect 25318 37839 25320 37848
rect 24124 37810 24176 37816
rect 25372 37839 25374 37848
rect 25872 37868 25924 37874
rect 25320 37810 25372 37816
rect 25872 37810 25924 37816
rect 26424 37868 26476 37874
rect 26424 37810 26476 37816
rect 21180 37800 21232 37806
rect 21180 37742 21232 37748
rect 22468 37800 22520 37806
rect 22468 37742 22520 37748
rect 22560 37800 22612 37806
rect 22560 37742 22612 37748
rect 21192 37194 21220 37742
rect 22480 37262 22508 37742
rect 22468 37256 22520 37262
rect 22468 37198 22520 37204
rect 21180 37188 21232 37194
rect 21180 37130 21232 37136
rect 22376 37120 22428 37126
rect 22376 37062 22428 37068
rect 22388 36922 22416 37062
rect 22376 36916 22428 36922
rect 22376 36858 22428 36864
rect 22468 36916 22520 36922
rect 22468 36858 22520 36864
rect 22284 36712 22336 36718
rect 22284 36654 22336 36660
rect 22100 36168 22152 36174
rect 22100 36110 22152 36116
rect 21364 36100 21416 36106
rect 21364 36042 21416 36048
rect 20996 35828 21048 35834
rect 20916 35788 20996 35816
rect 20720 34944 20772 34950
rect 20720 34886 20772 34892
rect 20628 34400 20680 34406
rect 20628 34342 20680 34348
rect 20536 34196 20588 34202
rect 20536 34138 20588 34144
rect 20548 33998 20576 34138
rect 20640 33998 20668 34342
rect 20536 33992 20588 33998
rect 20536 33934 20588 33940
rect 20628 33992 20680 33998
rect 20628 33934 20680 33940
rect 20640 33386 20668 33934
rect 20732 33522 20760 34886
rect 20916 34678 20944 35788
rect 20996 35770 21048 35776
rect 21088 35692 21140 35698
rect 21008 35652 21088 35680
rect 20904 34672 20956 34678
rect 20904 34614 20956 34620
rect 20904 33992 20956 33998
rect 20902 33960 20904 33969
rect 20956 33960 20958 33969
rect 20902 33895 20958 33904
rect 20812 33856 20864 33862
rect 20812 33798 20864 33804
rect 20720 33516 20772 33522
rect 20720 33458 20772 33464
rect 20628 33380 20680 33386
rect 20628 33322 20680 33328
rect 20352 33312 20404 33318
rect 20352 33254 20404 33260
rect 20444 33312 20496 33318
rect 20444 33254 20496 33260
rect 20364 33114 20392 33254
rect 20352 33108 20404 33114
rect 20352 33050 20404 33056
rect 20536 33040 20588 33046
rect 20272 32966 20392 32994
rect 20536 32982 20588 32988
rect 20720 33040 20772 33046
rect 20720 32982 20772 32988
rect 20168 32904 20220 32910
rect 20168 32846 20220 32852
rect 20180 32230 20208 32846
rect 20168 32224 20220 32230
rect 20168 32166 20220 32172
rect 20260 31952 20312 31958
rect 20260 31894 20312 31900
rect 20076 30728 20128 30734
rect 20076 30670 20128 30676
rect 19892 30660 19944 30666
rect 19892 30602 19944 30608
rect 19904 30326 19932 30602
rect 20168 30592 20220 30598
rect 20168 30534 20220 30540
rect 19892 30320 19944 30326
rect 19892 30262 19944 30268
rect 20076 30320 20128 30326
rect 20076 30262 20128 30268
rect 19982 30016 20038 30025
rect 19982 29951 20038 29960
rect 19996 29782 20024 29951
rect 19984 29776 20036 29782
rect 19984 29718 20036 29724
rect 19708 29708 19760 29714
rect 19708 29650 19760 29656
rect 19616 28960 19668 28966
rect 19616 28902 19668 28908
rect 19628 28626 19656 28902
rect 19616 28620 19668 28626
rect 19616 28562 19668 28568
rect 19614 28520 19670 28529
rect 19536 28464 19614 28472
rect 19536 28444 19616 28464
rect 19432 28416 19484 28422
rect 19432 28358 19484 28364
rect 19444 28257 19472 28358
rect 19430 28248 19486 28257
rect 19430 28183 19486 28192
rect 19536 28082 19564 28444
rect 19668 28455 19670 28464
rect 19616 28426 19668 28432
rect 19614 28112 19670 28121
rect 19524 28076 19576 28082
rect 19614 28047 19616 28056
rect 19524 28018 19576 28024
rect 19668 28047 19670 28056
rect 19616 28018 19668 28024
rect 19628 26790 19656 28018
rect 19616 26784 19668 26790
rect 19616 26726 19668 26732
rect 19340 26512 19392 26518
rect 19340 26454 19392 26460
rect 19720 26382 19748 29650
rect 19800 29164 19852 29170
rect 19800 29106 19852 29112
rect 19812 28558 19840 29106
rect 20088 29050 20116 30262
rect 19904 29022 20116 29050
rect 19800 28552 19852 28558
rect 19800 28494 19852 28500
rect 19798 28248 19854 28257
rect 19798 28183 19854 28192
rect 19812 28082 19840 28183
rect 19800 28076 19852 28082
rect 19800 28018 19852 28024
rect 19904 27996 19932 29022
rect 19984 28960 20036 28966
rect 19984 28902 20036 28908
rect 20076 28960 20128 28966
rect 20076 28902 20128 28908
rect 19996 28150 20024 28902
rect 20088 28694 20116 28902
rect 20076 28688 20128 28694
rect 20076 28630 20128 28636
rect 20180 28558 20208 30534
rect 20272 30258 20300 31894
rect 20364 31657 20392 32966
rect 20442 32872 20498 32881
rect 20442 32807 20498 32816
rect 20456 32434 20484 32807
rect 20444 32428 20496 32434
rect 20444 32370 20496 32376
rect 20456 31686 20484 32370
rect 20444 31680 20496 31686
rect 20350 31648 20406 31657
rect 20444 31622 20496 31628
rect 20350 31583 20406 31592
rect 20352 31476 20404 31482
rect 20404 31436 20484 31464
rect 20352 31418 20404 31424
rect 20352 31272 20404 31278
rect 20352 31214 20404 31220
rect 20364 30734 20392 31214
rect 20352 30728 20404 30734
rect 20352 30670 20404 30676
rect 20260 30252 20312 30258
rect 20260 30194 20312 30200
rect 20260 30116 20312 30122
rect 20260 30058 20312 30064
rect 20272 29782 20300 30058
rect 20364 30036 20392 30670
rect 20456 30580 20484 31436
rect 20548 30734 20576 32982
rect 20628 31952 20680 31958
rect 20628 31894 20680 31900
rect 20640 31346 20668 31894
rect 20732 31346 20760 32982
rect 20824 32026 20852 33798
rect 20904 33380 20956 33386
rect 20904 33322 20956 33328
rect 20916 33114 20944 33322
rect 20904 33108 20956 33114
rect 20904 33050 20956 33056
rect 20904 32224 20956 32230
rect 20904 32166 20956 32172
rect 20812 32020 20864 32026
rect 20812 31962 20864 31968
rect 20824 31482 20852 31962
rect 20812 31476 20864 31482
rect 20812 31418 20864 31424
rect 20628 31340 20680 31346
rect 20628 31282 20680 31288
rect 20720 31340 20772 31346
rect 20720 31282 20772 31288
rect 20718 31240 20774 31249
rect 20916 31210 20944 32166
rect 20718 31175 20774 31184
rect 20904 31204 20956 31210
rect 20626 30968 20682 30977
rect 20626 30903 20682 30912
rect 20536 30728 20588 30734
rect 20536 30670 20588 30676
rect 20640 30666 20668 30903
rect 20732 30870 20760 31175
rect 20904 31146 20956 31152
rect 20720 30864 20772 30870
rect 20720 30806 20772 30812
rect 20628 30660 20680 30666
rect 20628 30602 20680 30608
rect 20456 30552 20576 30580
rect 20444 30048 20496 30054
rect 20364 30008 20444 30036
rect 20444 29990 20496 29996
rect 20352 29844 20404 29850
rect 20352 29786 20404 29792
rect 20260 29776 20312 29782
rect 20260 29718 20312 29724
rect 20260 28756 20312 28762
rect 20260 28698 20312 28704
rect 20272 28665 20300 28698
rect 20258 28656 20314 28665
rect 20258 28591 20314 28600
rect 20168 28552 20220 28558
rect 20168 28494 20220 28500
rect 19984 28144 20036 28150
rect 19984 28086 20036 28092
rect 20260 28008 20312 28014
rect 19904 27968 20024 27996
rect 19248 26376 19300 26382
rect 19248 26318 19300 26324
rect 19340 26376 19392 26382
rect 19340 26318 19392 26324
rect 19708 26376 19760 26382
rect 19708 26318 19760 26324
rect 19154 26072 19210 26081
rect 19154 26007 19210 26016
rect 19168 25974 19196 26007
rect 19156 25968 19208 25974
rect 19156 25910 19208 25916
rect 19156 25696 19208 25702
rect 19156 25638 19208 25644
rect 19064 25356 19116 25362
rect 19064 25298 19116 25304
rect 19076 24206 19104 25298
rect 19168 24410 19196 25638
rect 19260 24818 19288 26318
rect 19352 25906 19380 26318
rect 19432 26036 19484 26042
rect 19484 25996 19840 26024
rect 19432 25978 19484 25984
rect 19812 25906 19840 25996
rect 19340 25900 19392 25906
rect 19340 25842 19392 25848
rect 19432 25900 19484 25906
rect 19432 25842 19484 25848
rect 19800 25900 19852 25906
rect 19800 25842 19852 25848
rect 19892 25900 19944 25906
rect 19892 25842 19944 25848
rect 19338 25800 19394 25809
rect 19338 25735 19340 25744
rect 19392 25735 19394 25744
rect 19340 25706 19392 25712
rect 19444 25702 19472 25842
rect 19432 25696 19484 25702
rect 19432 25638 19484 25644
rect 19340 25288 19392 25294
rect 19340 25230 19392 25236
rect 19352 24993 19380 25230
rect 19444 25158 19472 25638
rect 19904 25430 19932 25842
rect 19892 25424 19944 25430
rect 19892 25366 19944 25372
rect 19524 25220 19576 25226
rect 19524 25162 19576 25168
rect 19432 25152 19484 25158
rect 19432 25094 19484 25100
rect 19338 24984 19394 24993
rect 19338 24919 19394 24928
rect 19248 24812 19300 24818
rect 19248 24754 19300 24760
rect 19156 24404 19208 24410
rect 19156 24346 19208 24352
rect 19064 24200 19116 24206
rect 19064 24142 19116 24148
rect 19156 24132 19208 24138
rect 19156 24074 19208 24080
rect 19064 24064 19116 24070
rect 19064 24006 19116 24012
rect 18972 23860 19024 23866
rect 18972 23802 19024 23808
rect 18800 22066 18920 22094
rect 18892 21622 18920 22066
rect 18880 21616 18932 21622
rect 18880 21558 18932 21564
rect 18972 21480 19024 21486
rect 18972 21422 19024 21428
rect 18328 21140 18380 21146
rect 18328 21082 18380 21088
rect 18420 21140 18472 21146
rect 18420 21082 18472 21088
rect 18234 21040 18290 21049
rect 18340 21026 18368 21082
rect 18340 21010 18736 21026
rect 18340 21004 18748 21010
rect 18340 20998 18696 21004
rect 18234 20975 18290 20984
rect 18050 20431 18106 20440
rect 18144 20460 18196 20466
rect 18144 20402 18196 20408
rect 18052 20256 18104 20262
rect 18052 20198 18104 20204
rect 17920 19808 18000 19836
rect 17868 19790 17920 19796
rect 17972 18086 18000 19808
rect 18064 18970 18092 20198
rect 18248 19990 18276 20975
rect 18696 20946 18748 20952
rect 18788 20936 18840 20942
rect 18788 20878 18840 20884
rect 18512 20800 18564 20806
rect 18512 20742 18564 20748
rect 18326 20632 18382 20641
rect 18326 20567 18382 20576
rect 18340 20534 18368 20567
rect 18328 20528 18380 20534
rect 18328 20470 18380 20476
rect 18524 20466 18552 20742
rect 18512 20460 18564 20466
rect 18512 20402 18564 20408
rect 18800 20398 18828 20878
rect 18604 20392 18656 20398
rect 18604 20334 18656 20340
rect 18788 20392 18840 20398
rect 18788 20334 18840 20340
rect 18420 20324 18472 20330
rect 18420 20266 18472 20272
rect 18236 19984 18288 19990
rect 18236 19926 18288 19932
rect 18144 19712 18196 19718
rect 18144 19654 18196 19660
rect 18052 18964 18104 18970
rect 18052 18906 18104 18912
rect 18052 18624 18104 18630
rect 18052 18566 18104 18572
rect 17960 18080 18012 18086
rect 17960 18022 18012 18028
rect 18064 17678 18092 18566
rect 18156 17678 18184 19654
rect 18328 19304 18380 19310
rect 18328 19246 18380 19252
rect 18340 19174 18368 19246
rect 18328 19168 18380 19174
rect 18328 19110 18380 19116
rect 18236 18964 18288 18970
rect 18236 18906 18288 18912
rect 18248 18290 18276 18906
rect 18340 18680 18368 19110
rect 18432 18970 18460 20266
rect 18510 19000 18566 19009
rect 18420 18964 18472 18970
rect 18510 18935 18566 18944
rect 18420 18906 18472 18912
rect 18524 18902 18552 18935
rect 18512 18896 18564 18902
rect 18512 18838 18564 18844
rect 18512 18760 18564 18766
rect 18512 18702 18564 18708
rect 18340 18652 18460 18680
rect 18236 18284 18288 18290
rect 18236 18226 18288 18232
rect 18248 18034 18276 18226
rect 18248 18006 18368 18034
rect 18234 17912 18290 17921
rect 18234 17847 18290 17856
rect 17960 17672 18012 17678
rect 17960 17614 18012 17620
rect 18052 17672 18104 17678
rect 18052 17614 18104 17620
rect 18144 17672 18196 17678
rect 18144 17614 18196 17620
rect 17972 17524 18000 17614
rect 17972 17496 18092 17524
rect 18064 17202 18092 17496
rect 18052 17196 18104 17202
rect 18052 17138 18104 17144
rect 17958 16688 18014 16697
rect 17958 16623 18014 16632
rect 17868 16176 17920 16182
rect 17868 16118 17920 16124
rect 17880 15978 17908 16118
rect 17868 15972 17920 15978
rect 17868 15914 17920 15920
rect 17776 15700 17828 15706
rect 17776 15642 17828 15648
rect 17868 15088 17920 15094
rect 17868 15030 17920 15036
rect 17592 15020 17644 15026
rect 17592 14962 17644 14968
rect 17684 15020 17736 15026
rect 17684 14962 17736 14968
rect 17500 14000 17552 14006
rect 17500 13942 17552 13948
rect 17316 13932 17368 13938
rect 17316 13874 17368 13880
rect 17408 13728 17460 13734
rect 17408 13670 17460 13676
rect 16948 10668 17000 10674
rect 16948 10610 17000 10616
rect 17132 10668 17184 10674
rect 17132 10610 17184 10616
rect 16960 10554 16988 10610
rect 16960 10526 17080 10554
rect 16776 9646 16896 9674
rect 16672 9580 16724 9586
rect 16672 9522 16724 9528
rect 16764 8900 16816 8906
rect 16592 8860 16764 8888
rect 16028 8842 16080 8848
rect 16764 8842 16816 8848
rect 16776 8498 16804 8842
rect 16764 8492 16816 8498
rect 16764 8434 16816 8440
rect 15936 7948 15988 7954
rect 15936 7890 15988 7896
rect 15752 6860 15804 6866
rect 15752 6802 15804 6808
rect 15396 6458 15516 6474
rect 15396 6452 15528 6458
rect 15396 6446 15476 6452
rect 15476 6394 15528 6400
rect 15384 6384 15436 6390
rect 15384 6326 15436 6332
rect 15200 6316 15252 6322
rect 15200 6258 15252 6264
rect 15292 6316 15344 6322
rect 15292 6258 15344 6264
rect 15212 5710 15240 6258
rect 15304 5914 15332 6258
rect 15292 5908 15344 5914
rect 15292 5850 15344 5856
rect 15200 5704 15252 5710
rect 15200 5646 15252 5652
rect 15212 5370 15240 5646
rect 15396 5574 15424 6326
rect 15764 5778 15792 6802
rect 16776 6730 16804 8434
rect 16868 7818 16896 9646
rect 16948 9580 17000 9586
rect 16948 9522 17000 9528
rect 16960 8362 16988 9522
rect 17052 9500 17080 10526
rect 17144 10266 17172 10610
rect 17132 10260 17184 10266
rect 17132 10202 17184 10208
rect 17132 9512 17184 9518
rect 17052 9472 17132 9500
rect 17132 9454 17184 9460
rect 17038 9208 17094 9217
rect 17144 9194 17172 9454
rect 17094 9166 17172 9194
rect 17038 9143 17094 9152
rect 17144 8498 17172 9166
rect 17420 8498 17448 13670
rect 17604 13462 17632 14962
rect 17696 14822 17724 14962
rect 17684 14816 17736 14822
rect 17684 14758 17736 14764
rect 17880 14074 17908 15030
rect 17972 14464 18000 16623
rect 18064 16538 18092 17138
rect 18248 16658 18276 17847
rect 18340 16998 18368 18006
rect 18432 17202 18460 18652
rect 18524 18426 18552 18702
rect 18512 18420 18564 18426
rect 18512 18362 18564 18368
rect 18616 18086 18644 20334
rect 18984 19854 19012 21422
rect 18972 19848 19024 19854
rect 18972 19790 19024 19796
rect 18984 18766 19012 19790
rect 18972 18760 19024 18766
rect 18970 18728 18972 18737
rect 19024 18728 19026 18737
rect 18696 18692 18748 18698
rect 18970 18663 19026 18672
rect 18696 18634 18748 18640
rect 18512 18080 18564 18086
rect 18512 18022 18564 18028
rect 18604 18080 18656 18086
rect 18604 18022 18656 18028
rect 18420 17196 18472 17202
rect 18420 17138 18472 17144
rect 18328 16992 18380 16998
rect 18328 16934 18380 16940
rect 18236 16652 18288 16658
rect 18236 16594 18288 16600
rect 18064 16510 18276 16538
rect 18052 16448 18104 16454
rect 18052 16390 18104 16396
rect 18144 16448 18196 16454
rect 18144 16390 18196 16396
rect 18064 16114 18092 16390
rect 18156 16114 18184 16390
rect 18248 16250 18276 16510
rect 18524 16454 18552 18022
rect 18602 17912 18658 17921
rect 18602 17847 18658 17856
rect 18616 17814 18644 17847
rect 18604 17808 18656 17814
rect 18604 17750 18656 17756
rect 18708 17746 18736 18634
rect 18788 18624 18840 18630
rect 18788 18566 18840 18572
rect 18696 17740 18748 17746
rect 18696 17682 18748 17688
rect 18800 17678 18828 18566
rect 18880 18284 18932 18290
rect 18880 18226 18932 18232
rect 18892 18193 18920 18226
rect 18878 18184 18934 18193
rect 18878 18119 18934 18128
rect 18788 17672 18840 17678
rect 18788 17614 18840 17620
rect 18604 17536 18656 17542
rect 18604 17478 18656 17484
rect 18880 17536 18932 17542
rect 18880 17478 18932 17484
rect 18972 17536 19024 17542
rect 18972 17478 19024 17484
rect 18616 16590 18644 17478
rect 18788 17128 18840 17134
rect 18788 17070 18840 17076
rect 18800 16590 18828 17070
rect 18604 16584 18656 16590
rect 18604 16526 18656 16532
rect 18788 16584 18840 16590
rect 18788 16526 18840 16532
rect 18696 16516 18748 16522
rect 18696 16458 18748 16464
rect 18512 16448 18564 16454
rect 18512 16390 18564 16396
rect 18236 16244 18288 16250
rect 18236 16186 18288 16192
rect 18052 16108 18104 16114
rect 18052 16050 18104 16056
rect 18144 16108 18196 16114
rect 18144 16050 18196 16056
rect 18604 15904 18656 15910
rect 18604 15846 18656 15852
rect 18616 15570 18644 15846
rect 18604 15564 18656 15570
rect 18604 15506 18656 15512
rect 18236 15496 18288 15502
rect 18236 15438 18288 15444
rect 18248 15026 18276 15438
rect 18616 15026 18644 15506
rect 18708 15434 18736 16458
rect 18892 16114 18920 17478
rect 18984 17270 19012 17478
rect 18972 17264 19024 17270
rect 18972 17206 19024 17212
rect 19076 16640 19104 24006
rect 19168 23730 19196 24074
rect 19248 24064 19300 24070
rect 19248 24006 19300 24012
rect 19260 23866 19288 24006
rect 19248 23860 19300 23866
rect 19248 23802 19300 23808
rect 19156 23724 19208 23730
rect 19156 23666 19208 23672
rect 19352 22166 19380 24919
rect 19536 24206 19564 25162
rect 19892 24676 19944 24682
rect 19892 24618 19944 24624
rect 19524 24200 19576 24206
rect 19524 24142 19576 24148
rect 19904 24070 19932 24618
rect 19996 24070 20024 27968
rect 20364 27996 20392 29786
rect 20456 28014 20484 29990
rect 20312 27968 20392 27996
rect 20444 28008 20496 28014
rect 20442 27976 20444 27985
rect 20496 27976 20498 27985
rect 20260 27950 20312 27956
rect 20168 27328 20220 27334
rect 20168 27270 20220 27276
rect 20076 26920 20128 26926
rect 20076 26862 20128 26868
rect 20088 26042 20116 26862
rect 20180 26314 20208 27270
rect 20168 26308 20220 26314
rect 20168 26250 20220 26256
rect 20076 26036 20128 26042
rect 20076 25978 20128 25984
rect 20168 25968 20220 25974
rect 20168 25910 20220 25916
rect 20076 25832 20128 25838
rect 20074 25800 20076 25809
rect 20128 25800 20130 25809
rect 20074 25735 20130 25744
rect 20180 25702 20208 25910
rect 20168 25696 20220 25702
rect 20168 25638 20220 25644
rect 20272 25294 20300 27950
rect 20442 27911 20498 27920
rect 20352 27872 20404 27878
rect 20352 27814 20404 27820
rect 20444 27872 20496 27878
rect 20444 27814 20496 27820
rect 20364 27538 20392 27814
rect 20352 27532 20404 27538
rect 20352 27474 20404 27480
rect 20350 26480 20406 26489
rect 20350 26415 20352 26424
rect 20404 26415 20406 26424
rect 20352 26386 20404 26392
rect 20352 26308 20404 26314
rect 20352 26250 20404 26256
rect 20364 25906 20392 26250
rect 20352 25900 20404 25906
rect 20352 25842 20404 25848
rect 20260 25288 20312 25294
rect 20260 25230 20312 25236
rect 20076 24812 20128 24818
rect 20076 24754 20128 24760
rect 20088 24274 20116 24754
rect 20260 24336 20312 24342
rect 20260 24278 20312 24284
rect 20352 24336 20404 24342
rect 20352 24278 20404 24284
rect 20076 24268 20128 24274
rect 20076 24210 20128 24216
rect 19892 24064 19944 24070
rect 19892 24006 19944 24012
rect 19984 24064 20036 24070
rect 19984 24006 20036 24012
rect 19904 23866 19932 24006
rect 19892 23860 19944 23866
rect 19892 23802 19944 23808
rect 19430 23760 19486 23769
rect 19996 23730 20024 24006
rect 19430 23695 19432 23704
rect 19484 23695 19486 23704
rect 19984 23724 20036 23730
rect 19432 23666 19484 23672
rect 19984 23666 20036 23672
rect 19708 23520 19760 23526
rect 19708 23462 19760 23468
rect 19720 23254 19748 23462
rect 19708 23248 19760 23254
rect 19708 23190 19760 23196
rect 19996 23186 20024 23666
rect 20088 23254 20116 24210
rect 20168 23860 20220 23866
rect 20168 23802 20220 23808
rect 20180 23322 20208 23802
rect 20272 23730 20300 24278
rect 20260 23724 20312 23730
rect 20260 23666 20312 23672
rect 20364 23594 20392 24278
rect 20352 23588 20404 23594
rect 20352 23530 20404 23536
rect 20168 23316 20220 23322
rect 20168 23258 20220 23264
rect 20076 23248 20128 23254
rect 20076 23190 20128 23196
rect 19984 23180 20036 23186
rect 19984 23122 20036 23128
rect 20364 23118 20392 23530
rect 20352 23112 20404 23118
rect 20352 23054 20404 23060
rect 19892 23044 19944 23050
rect 19892 22986 19944 22992
rect 19340 22160 19392 22166
rect 19246 22128 19302 22137
rect 19168 22086 19246 22114
rect 19168 21434 19196 22086
rect 19340 22102 19392 22108
rect 19246 22063 19302 22072
rect 19248 22024 19300 22030
rect 19248 21966 19300 21972
rect 19708 22024 19760 22030
rect 19708 21966 19760 21972
rect 19800 22024 19852 22030
rect 19800 21966 19852 21972
rect 19260 21554 19288 21966
rect 19340 21616 19392 21622
rect 19340 21558 19392 21564
rect 19248 21548 19300 21554
rect 19248 21490 19300 21496
rect 19168 21406 19288 21434
rect 19156 17808 19208 17814
rect 19156 17750 19208 17756
rect 19168 17270 19196 17750
rect 19260 17610 19288 21406
rect 19352 20466 19380 21558
rect 19720 21486 19748 21966
rect 19812 21622 19840 21966
rect 19800 21616 19852 21622
rect 19800 21558 19852 21564
rect 19708 21480 19760 21486
rect 19708 21422 19760 21428
rect 19798 21448 19854 21457
rect 19432 20936 19484 20942
rect 19432 20878 19484 20884
rect 19524 20936 19576 20942
rect 19524 20878 19576 20884
rect 19340 20460 19392 20466
rect 19340 20402 19392 20408
rect 19444 20262 19472 20878
rect 19536 20262 19564 20878
rect 19616 20324 19668 20330
rect 19616 20266 19668 20272
rect 19432 20256 19484 20262
rect 19432 20198 19484 20204
rect 19524 20256 19576 20262
rect 19524 20198 19576 20204
rect 19340 19712 19392 19718
rect 19340 19654 19392 19660
rect 19352 19310 19380 19654
rect 19444 19378 19472 20198
rect 19536 19718 19564 20198
rect 19628 19854 19656 20266
rect 19616 19848 19668 19854
rect 19616 19790 19668 19796
rect 19524 19712 19576 19718
rect 19524 19654 19576 19660
rect 19432 19372 19484 19378
rect 19432 19314 19484 19320
rect 19340 19304 19392 19310
rect 19340 19246 19392 19252
rect 19352 18952 19380 19246
rect 19352 18924 19472 18952
rect 19340 18828 19392 18834
rect 19340 18770 19392 18776
rect 19352 18170 19380 18770
rect 19444 18766 19472 18924
rect 19432 18760 19484 18766
rect 19432 18702 19484 18708
rect 19536 18204 19564 19654
rect 19616 19372 19668 19378
rect 19616 19314 19668 19320
rect 19628 18748 19656 19314
rect 19720 18970 19748 21422
rect 19798 21383 19854 21392
rect 19812 21350 19840 21383
rect 19800 21344 19852 21350
rect 19800 21286 19852 21292
rect 19800 19780 19852 19786
rect 19800 19722 19852 19728
rect 19812 19174 19840 19722
rect 19800 19168 19852 19174
rect 19800 19110 19852 19116
rect 19708 18964 19760 18970
rect 19708 18906 19760 18912
rect 19708 18760 19760 18766
rect 19628 18720 19708 18748
rect 19708 18702 19760 18708
rect 19798 18728 19854 18737
rect 19720 18426 19748 18702
rect 19798 18663 19854 18672
rect 19708 18420 19760 18426
rect 19708 18362 19760 18368
rect 19812 18290 19840 18663
rect 19800 18284 19852 18290
rect 19800 18226 19852 18232
rect 19536 18176 19657 18204
rect 19629 18170 19657 18176
rect 19352 18154 19472 18170
rect 19352 18148 19484 18154
rect 19352 18142 19432 18148
rect 19629 18142 19665 18170
rect 19484 18108 19564 18136
rect 19432 18090 19484 18096
rect 19536 17678 19564 18108
rect 19637 18034 19665 18142
rect 19628 18006 19665 18034
rect 19524 17672 19576 17678
rect 19524 17614 19576 17620
rect 19248 17604 19300 17610
rect 19248 17546 19300 17552
rect 19156 17264 19208 17270
rect 19156 17206 19208 17212
rect 18984 16612 19104 16640
rect 18880 16108 18932 16114
rect 18880 16050 18932 16056
rect 18880 15904 18932 15910
rect 18878 15872 18880 15881
rect 18932 15872 18934 15881
rect 18878 15807 18934 15816
rect 18696 15428 18748 15434
rect 18696 15370 18748 15376
rect 18788 15360 18840 15366
rect 18788 15302 18840 15308
rect 18236 15020 18288 15026
rect 18604 15020 18656 15026
rect 18288 14980 18368 15008
rect 18236 14962 18288 14968
rect 18052 14476 18104 14482
rect 17972 14436 18052 14464
rect 18052 14418 18104 14424
rect 17868 14068 17920 14074
rect 17868 14010 17920 14016
rect 17868 13728 17920 13734
rect 17868 13670 17920 13676
rect 17880 13530 17908 13670
rect 17868 13524 17920 13530
rect 17868 13466 17920 13472
rect 17592 13456 17644 13462
rect 17592 13398 17644 13404
rect 18236 13252 18288 13258
rect 18236 13194 18288 13200
rect 18248 12866 18276 13194
rect 18156 12838 18276 12866
rect 17684 12164 17736 12170
rect 17684 12106 17736 12112
rect 17592 12096 17644 12102
rect 17592 12038 17644 12044
rect 17604 11626 17632 12038
rect 17592 11620 17644 11626
rect 17592 11562 17644 11568
rect 17604 11354 17632 11562
rect 17592 11348 17644 11354
rect 17592 11290 17644 11296
rect 17498 10568 17554 10577
rect 17498 10503 17500 10512
rect 17552 10503 17554 10512
rect 17500 10474 17552 10480
rect 17696 9674 17724 12106
rect 18156 11558 18184 12838
rect 18340 12238 18368 14980
rect 18604 14962 18656 14968
rect 18696 14952 18748 14958
rect 18696 14894 18748 14900
rect 18420 13796 18472 13802
rect 18420 13738 18472 13744
rect 18432 13530 18460 13738
rect 18708 13682 18736 14894
rect 18800 14822 18828 15302
rect 18788 14816 18840 14822
rect 18788 14758 18840 14764
rect 18524 13654 18736 13682
rect 18420 13524 18472 13530
rect 18420 13466 18472 13472
rect 18420 13388 18472 13394
rect 18420 13330 18472 13336
rect 18432 13190 18460 13330
rect 18420 13184 18472 13190
rect 18420 13126 18472 13132
rect 18420 12844 18472 12850
rect 18420 12786 18472 12792
rect 18432 12306 18460 12786
rect 18420 12300 18472 12306
rect 18420 12242 18472 12248
rect 18328 12232 18380 12238
rect 18328 12174 18380 12180
rect 18144 11552 18196 11558
rect 18144 11494 18196 11500
rect 18052 10464 18104 10470
rect 18052 10406 18104 10412
rect 18064 10062 18092 10406
rect 18156 10130 18184 11494
rect 18340 11150 18368 12174
rect 18328 11144 18380 11150
rect 18328 11086 18380 11092
rect 18234 10976 18290 10985
rect 18234 10911 18290 10920
rect 18144 10124 18196 10130
rect 18144 10066 18196 10072
rect 18052 10056 18104 10062
rect 18052 9998 18104 10004
rect 17604 9646 17724 9674
rect 17604 9042 17632 9646
rect 18064 9586 18092 9998
rect 18052 9580 18104 9586
rect 18052 9522 18104 9528
rect 17592 9036 17644 9042
rect 17592 8978 17644 8984
rect 17132 8492 17184 8498
rect 17132 8434 17184 8440
rect 17408 8492 17460 8498
rect 17408 8434 17460 8440
rect 16948 8356 17000 8362
rect 16948 8298 17000 8304
rect 17224 8356 17276 8362
rect 17224 8298 17276 8304
rect 16856 7812 16908 7818
rect 16856 7754 16908 7760
rect 16764 6724 16816 6730
rect 16764 6666 16816 6672
rect 16488 6112 16540 6118
rect 16488 6054 16540 6060
rect 16304 5908 16356 5914
rect 16304 5850 16356 5856
rect 15752 5772 15804 5778
rect 15752 5714 15804 5720
rect 15936 5636 15988 5642
rect 15936 5578 15988 5584
rect 16120 5636 16172 5642
rect 16120 5578 16172 5584
rect 15384 5568 15436 5574
rect 15384 5510 15436 5516
rect 15200 5364 15252 5370
rect 15200 5306 15252 5312
rect 15396 5166 15424 5510
rect 15384 5160 15436 5166
rect 15384 5102 15436 5108
rect 15844 5160 15896 5166
rect 15844 5102 15896 5108
rect 15856 4826 15884 5102
rect 15844 4820 15896 4826
rect 15844 4762 15896 4768
rect 15948 4622 15976 5578
rect 16132 5302 16160 5578
rect 16120 5296 16172 5302
rect 16120 5238 16172 5244
rect 16316 4622 16344 5850
rect 16396 5024 16448 5030
rect 16396 4966 16448 4972
rect 16408 4826 16436 4966
rect 16396 4820 16448 4826
rect 16396 4762 16448 4768
rect 16500 4622 16528 6054
rect 16672 5160 16724 5166
rect 16672 5102 16724 5108
rect 16684 4826 16712 5102
rect 16672 4820 16724 4826
rect 16672 4762 16724 4768
rect 15936 4616 15988 4622
rect 15936 4558 15988 4564
rect 16304 4616 16356 4622
rect 16304 4558 16356 4564
rect 16488 4616 16540 4622
rect 16488 4558 16540 4564
rect 16776 4486 16804 6666
rect 17132 5704 17184 5710
rect 17132 5646 17184 5652
rect 17144 5370 17172 5646
rect 17132 5364 17184 5370
rect 17132 5306 17184 5312
rect 16764 4480 16816 4486
rect 16764 4422 16816 4428
rect 17236 3194 17264 8298
rect 17604 7886 17632 8978
rect 18156 8974 18184 10066
rect 18248 10062 18276 10911
rect 18340 10674 18368 11086
rect 18524 11082 18552 13654
rect 18696 13184 18748 13190
rect 18696 13126 18748 13132
rect 18708 13025 18736 13126
rect 18694 13016 18750 13025
rect 18694 12951 18750 12960
rect 18800 12238 18828 14758
rect 18892 13258 18920 15807
rect 18984 13802 19012 16612
rect 19064 16516 19116 16522
rect 19064 16458 19116 16464
rect 19076 16250 19104 16458
rect 19064 16244 19116 16250
rect 19064 16186 19116 16192
rect 19064 15632 19116 15638
rect 19064 15574 19116 15580
rect 19248 15632 19300 15638
rect 19248 15574 19300 15580
rect 19076 15162 19104 15574
rect 19156 15360 19208 15366
rect 19156 15302 19208 15308
rect 19064 15156 19116 15162
rect 19064 15098 19116 15104
rect 19076 15026 19104 15098
rect 19064 15020 19116 15026
rect 19064 14962 19116 14968
rect 18972 13796 19024 13802
rect 18972 13738 19024 13744
rect 18984 13258 19012 13738
rect 18880 13252 18932 13258
rect 18880 13194 18932 13200
rect 18972 13252 19024 13258
rect 18972 13194 19024 13200
rect 18892 12306 18920 13194
rect 18880 12300 18932 12306
rect 18880 12242 18932 12248
rect 18788 12232 18840 12238
rect 18788 12174 18840 12180
rect 19168 11830 19196 15302
rect 19260 14822 19288 15574
rect 19628 15434 19656 18006
rect 19800 17604 19852 17610
rect 19800 17546 19852 17552
rect 19812 17270 19840 17546
rect 19800 17264 19852 17270
rect 19800 17206 19852 17212
rect 19708 17196 19760 17202
rect 19708 17138 19760 17144
rect 19720 16114 19748 17138
rect 19708 16108 19760 16114
rect 19708 16050 19760 16056
rect 19616 15428 19668 15434
rect 19616 15370 19668 15376
rect 19628 15026 19656 15370
rect 19616 15020 19668 15026
rect 19616 14962 19668 14968
rect 19432 14952 19484 14958
rect 19432 14894 19484 14900
rect 19248 14816 19300 14822
rect 19248 14758 19300 14764
rect 19444 14278 19472 14894
rect 19524 14340 19576 14346
rect 19524 14282 19576 14288
rect 19432 14272 19484 14278
rect 19432 14214 19484 14220
rect 19248 13456 19300 13462
rect 19248 13398 19300 13404
rect 19340 13456 19392 13462
rect 19340 13398 19392 13404
rect 19260 13190 19288 13398
rect 19248 13184 19300 13190
rect 19248 13126 19300 13132
rect 19352 12238 19380 13398
rect 19444 12986 19472 14214
rect 19536 13326 19564 14282
rect 19708 13932 19760 13938
rect 19708 13874 19760 13880
rect 19616 13728 19668 13734
rect 19616 13670 19668 13676
rect 19524 13320 19576 13326
rect 19524 13262 19576 13268
rect 19432 12980 19484 12986
rect 19432 12922 19484 12928
rect 19536 12918 19564 13262
rect 19524 12912 19576 12918
rect 19524 12854 19576 12860
rect 19628 12646 19656 13670
rect 19720 13530 19748 13874
rect 19708 13524 19760 13530
rect 19708 13466 19760 13472
rect 19616 12640 19668 12646
rect 19616 12582 19668 12588
rect 19340 12232 19392 12238
rect 19340 12174 19392 12180
rect 19524 12096 19576 12102
rect 19524 12038 19576 12044
rect 19156 11824 19208 11830
rect 19156 11766 19208 11772
rect 18694 11656 18750 11665
rect 18694 11591 18696 11600
rect 18748 11591 18750 11600
rect 18696 11562 18748 11568
rect 18512 11076 18564 11082
rect 18512 11018 18564 11024
rect 18524 10674 18552 11018
rect 19168 10810 19196 11766
rect 19248 11552 19300 11558
rect 19248 11494 19300 11500
rect 19260 11286 19288 11494
rect 19248 11280 19300 11286
rect 19248 11222 19300 11228
rect 19536 11150 19564 12038
rect 19904 11286 19932 22986
rect 20364 22710 20392 23054
rect 20352 22704 20404 22710
rect 20352 22646 20404 22652
rect 20076 22024 20128 22030
rect 20076 21966 20128 21972
rect 20088 21622 20116 21966
rect 20076 21616 20128 21622
rect 20076 21558 20128 21564
rect 19984 21548 20036 21554
rect 19984 21490 20036 21496
rect 19996 21146 20024 21490
rect 20088 21350 20116 21558
rect 20352 21548 20404 21554
rect 20352 21490 20404 21496
rect 20260 21480 20312 21486
rect 20260 21422 20312 21428
rect 20076 21344 20128 21350
rect 20076 21286 20128 21292
rect 20166 21312 20222 21321
rect 20166 21247 20222 21256
rect 19984 21140 20036 21146
rect 19984 21082 20036 21088
rect 20076 20460 20128 20466
rect 20076 20402 20128 20408
rect 20088 19922 20116 20402
rect 20180 20262 20208 21247
rect 20168 20256 20220 20262
rect 20168 20198 20220 20204
rect 20076 19916 20128 19922
rect 20076 19858 20128 19864
rect 19984 19848 20036 19854
rect 19984 19790 20036 19796
rect 20272 19836 20300 21422
rect 20364 20942 20392 21490
rect 20352 20936 20404 20942
rect 20352 20878 20404 20884
rect 20352 20800 20404 20806
rect 20352 20742 20404 20748
rect 20364 20466 20392 20742
rect 20352 20460 20404 20466
rect 20352 20402 20404 20408
rect 20352 19848 20404 19854
rect 20272 19808 20352 19836
rect 19996 19514 20024 19790
rect 20076 19712 20128 19718
rect 20076 19654 20128 19660
rect 19984 19508 20036 19514
rect 19984 19450 20036 19456
rect 19984 18760 20036 18766
rect 19984 18702 20036 18708
rect 19996 18290 20024 18702
rect 20088 18698 20116 19654
rect 20076 18692 20128 18698
rect 20076 18634 20128 18640
rect 19984 18284 20036 18290
rect 19984 18226 20036 18232
rect 19996 18086 20024 18226
rect 20088 18193 20116 18634
rect 20166 18456 20222 18465
rect 20166 18391 20168 18400
rect 20220 18391 20222 18400
rect 20168 18362 20220 18368
rect 20074 18184 20130 18193
rect 20074 18119 20130 18128
rect 19984 18080 20036 18086
rect 19984 18022 20036 18028
rect 19996 17116 20024 18022
rect 20088 17678 20116 18119
rect 20272 18086 20300 19808
rect 20352 19790 20404 19796
rect 20352 18624 20404 18630
rect 20352 18566 20404 18572
rect 20364 18086 20392 18566
rect 20456 18086 20484 27814
rect 20548 26194 20576 30552
rect 20640 30326 20668 30602
rect 21008 30598 21036 35652
rect 21088 35634 21140 35640
rect 21180 35692 21232 35698
rect 21180 35634 21232 35640
rect 21088 32496 21140 32502
rect 21088 32438 21140 32444
rect 21100 31793 21128 32438
rect 21086 31784 21142 31793
rect 21086 31719 21142 31728
rect 21192 31634 21220 35634
rect 21272 34672 21324 34678
rect 21272 34614 21324 34620
rect 21284 33658 21312 34614
rect 21272 33652 21324 33658
rect 21272 33594 21324 33600
rect 21376 33590 21404 36042
rect 21548 35624 21600 35630
rect 21548 35566 21600 35572
rect 21456 35488 21508 35494
rect 21456 35430 21508 35436
rect 21468 33697 21496 35430
rect 21454 33688 21510 33697
rect 21454 33623 21510 33632
rect 21560 33590 21588 35566
rect 21824 35488 21876 35494
rect 21824 35430 21876 35436
rect 21836 35018 21864 35430
rect 21824 35012 21876 35018
rect 21824 34954 21876 34960
rect 21836 34678 21864 34954
rect 21824 34672 21876 34678
rect 21824 34614 21876 34620
rect 22112 34610 22140 36110
rect 22296 35698 22324 36654
rect 22480 35834 22508 36858
rect 22468 35828 22520 35834
rect 22468 35770 22520 35776
rect 22192 35692 22244 35698
rect 22192 35634 22244 35640
rect 22284 35692 22336 35698
rect 22284 35634 22336 35640
rect 22376 35692 22428 35698
rect 22376 35634 22428 35640
rect 22100 34604 22152 34610
rect 22100 34546 22152 34552
rect 22008 34400 22060 34406
rect 22008 34342 22060 34348
rect 21916 33992 21968 33998
rect 21916 33934 21968 33940
rect 21928 33658 21956 33934
rect 21916 33652 21968 33658
rect 21916 33594 21968 33600
rect 21364 33584 21416 33590
rect 21364 33526 21416 33532
rect 21548 33584 21600 33590
rect 21548 33526 21600 33532
rect 21456 33312 21508 33318
rect 21456 33254 21508 33260
rect 21468 32910 21496 33254
rect 21456 32904 21508 32910
rect 21456 32846 21508 32852
rect 21364 32428 21416 32434
rect 21100 31606 21220 31634
rect 21284 32388 21364 32416
rect 21100 30598 21128 31606
rect 21180 31340 21232 31346
rect 21284 31328 21312 32388
rect 21364 32370 21416 32376
rect 21364 31680 21416 31686
rect 21364 31622 21416 31628
rect 21232 31300 21312 31328
rect 21180 31282 21232 31288
rect 21192 30666 21220 31282
rect 21376 31278 21404 31622
rect 21468 31482 21496 32846
rect 21560 32842 21588 33526
rect 21824 33516 21876 33522
rect 21824 33458 21876 33464
rect 21548 32836 21600 32842
rect 21548 32778 21600 32784
rect 21560 31521 21588 32778
rect 21640 32496 21692 32502
rect 21638 32464 21640 32473
rect 21692 32464 21694 32473
rect 21638 32399 21694 32408
rect 21730 32056 21786 32065
rect 21730 31991 21786 32000
rect 21744 31822 21772 31991
rect 21732 31816 21784 31822
rect 21732 31758 21784 31764
rect 21836 31754 21864 33458
rect 21928 32910 21956 33594
rect 21916 32904 21968 32910
rect 21916 32846 21968 32852
rect 22020 32774 22048 34342
rect 22100 34196 22152 34202
rect 22100 34138 22152 34144
rect 22112 33658 22140 34138
rect 22100 33652 22152 33658
rect 22100 33594 22152 33600
rect 22204 32994 22232 35634
rect 22284 34672 22336 34678
rect 22284 34614 22336 34620
rect 22296 34377 22324 34614
rect 22282 34368 22338 34377
rect 22282 34303 22338 34312
rect 22284 33924 22336 33930
rect 22284 33866 22336 33872
rect 22112 32966 22232 32994
rect 22008 32768 22060 32774
rect 22008 32710 22060 32716
rect 22008 32020 22060 32026
rect 22008 31962 22060 31968
rect 22020 31822 22048 31962
rect 22112 31822 22140 32966
rect 22192 32904 22244 32910
rect 22192 32846 22244 32852
rect 22204 32230 22232 32846
rect 22296 32570 22324 33866
rect 22284 32564 22336 32570
rect 22284 32506 22336 32512
rect 22284 32360 22336 32366
rect 22284 32302 22336 32308
rect 22192 32224 22244 32230
rect 22192 32166 22244 32172
rect 21916 31816 21968 31822
rect 21916 31758 21968 31764
rect 22008 31816 22060 31822
rect 22008 31758 22060 31764
rect 22100 31816 22152 31822
rect 22100 31758 22152 31764
rect 21824 31748 21876 31754
rect 21824 31690 21876 31696
rect 21638 31648 21694 31657
rect 21638 31583 21694 31592
rect 21546 31512 21602 31521
rect 21456 31476 21508 31482
rect 21546 31447 21602 31456
rect 21652 31464 21680 31583
rect 21456 31418 21508 31424
rect 21560 31346 21588 31447
rect 21652 31436 21864 31464
rect 21730 31376 21786 31385
rect 21548 31340 21600 31346
rect 21730 31311 21786 31320
rect 21548 31282 21600 31288
rect 21744 31278 21772 31311
rect 21364 31272 21416 31278
rect 21364 31214 21416 31220
rect 21732 31272 21784 31278
rect 21732 31214 21784 31220
rect 21364 30728 21416 30734
rect 21364 30670 21416 30676
rect 21180 30660 21232 30666
rect 21180 30602 21232 30608
rect 20720 30592 20772 30598
rect 20720 30534 20772 30540
rect 20996 30592 21048 30598
rect 20996 30534 21048 30540
rect 21088 30592 21140 30598
rect 21088 30534 21140 30540
rect 20628 30320 20680 30326
rect 20628 30262 20680 30268
rect 20640 29850 20668 30262
rect 20628 29844 20680 29850
rect 20628 29786 20680 29792
rect 20732 29510 20760 30534
rect 20812 30320 20864 30326
rect 20812 30262 20864 30268
rect 20824 30054 20852 30262
rect 21008 30054 21036 30534
rect 20812 30048 20864 30054
rect 20812 29990 20864 29996
rect 20996 30048 21048 30054
rect 20996 29990 21048 29996
rect 21008 29646 21036 29990
rect 20812 29640 20864 29646
rect 20812 29582 20864 29588
rect 20996 29640 21048 29646
rect 20996 29582 21048 29588
rect 20720 29504 20772 29510
rect 20720 29446 20772 29452
rect 20824 29345 20852 29582
rect 21100 29510 21128 30534
rect 21088 29504 21140 29510
rect 21008 29464 21088 29492
rect 20810 29336 20866 29345
rect 20810 29271 20866 29280
rect 20824 29170 20852 29271
rect 20902 29200 20958 29209
rect 20812 29164 20864 29170
rect 20902 29135 20904 29144
rect 20812 29106 20864 29112
rect 20956 29135 20958 29144
rect 20904 29106 20956 29112
rect 21008 28994 21036 29464
rect 21088 29446 21140 29452
rect 21180 29504 21232 29510
rect 21180 29446 21232 29452
rect 21192 29170 21220 29446
rect 21180 29164 21232 29170
rect 21180 29106 21232 29112
rect 21086 29064 21142 29073
rect 21086 28999 21142 29008
rect 20916 28966 21036 28994
rect 20628 28076 20680 28082
rect 20628 28018 20680 28024
rect 20640 27402 20668 28018
rect 20628 27396 20680 27402
rect 20628 27338 20680 27344
rect 20720 26784 20772 26790
rect 20720 26726 20772 26732
rect 20626 26208 20682 26217
rect 20548 26166 20626 26194
rect 20626 26143 20682 26152
rect 20640 25974 20668 26143
rect 20628 25968 20680 25974
rect 20628 25910 20680 25916
rect 20732 25294 20760 26726
rect 20916 26518 20944 28966
rect 20996 28552 21048 28558
rect 20996 28494 21048 28500
rect 20904 26512 20956 26518
rect 20904 26454 20956 26460
rect 20812 26240 20864 26246
rect 20812 26182 20864 26188
rect 20824 26042 20852 26182
rect 20812 26036 20864 26042
rect 20812 25978 20864 25984
rect 20904 25968 20956 25974
rect 20824 25916 20904 25922
rect 20824 25910 20956 25916
rect 20824 25894 20944 25910
rect 21008 25906 21036 28494
rect 21100 28150 21128 28999
rect 21088 28144 21140 28150
rect 21088 28086 21140 28092
rect 21086 27976 21142 27985
rect 21086 27911 21142 27920
rect 20996 25900 21048 25906
rect 20720 25288 20772 25294
rect 20720 25230 20772 25236
rect 20628 25152 20680 25158
rect 20534 25120 20590 25129
rect 20628 25094 20680 25100
rect 20534 25055 20590 25064
rect 20548 24410 20576 25055
rect 20536 24404 20588 24410
rect 20536 24346 20588 24352
rect 20640 23118 20668 25094
rect 20824 24614 20852 25894
rect 20996 25842 21048 25848
rect 21100 25702 21128 27911
rect 21272 27464 21324 27470
rect 21272 27406 21324 27412
rect 21284 26450 21312 27406
rect 21272 26444 21324 26450
rect 21272 26386 21324 26392
rect 21180 25764 21232 25770
rect 21180 25706 21232 25712
rect 20996 25696 21048 25702
rect 20996 25638 21048 25644
rect 21088 25696 21140 25702
rect 21088 25638 21140 25644
rect 21008 25362 21036 25638
rect 20996 25356 21048 25362
rect 20996 25298 21048 25304
rect 20904 25220 20956 25226
rect 20904 25162 20956 25168
rect 20916 24886 20944 25162
rect 21192 24886 21220 25706
rect 21284 25294 21312 26386
rect 21272 25288 21324 25294
rect 21272 25230 21324 25236
rect 20904 24880 20956 24886
rect 20904 24822 20956 24828
rect 21180 24880 21232 24886
rect 21180 24822 21232 24828
rect 20812 24608 20864 24614
rect 20812 24550 20864 24556
rect 21376 24342 21404 30670
rect 21640 30592 21692 30598
rect 21640 30534 21692 30540
rect 21548 29572 21600 29578
rect 21548 29514 21600 29520
rect 21560 29102 21588 29514
rect 21652 29238 21680 30534
rect 21640 29232 21692 29238
rect 21640 29174 21692 29180
rect 21548 29096 21600 29102
rect 21548 29038 21600 29044
rect 21560 28762 21588 29038
rect 21548 28756 21600 28762
rect 21548 28698 21600 28704
rect 21548 28144 21600 28150
rect 21548 28086 21600 28092
rect 21456 28076 21508 28082
rect 21456 28018 21508 28024
rect 21468 27674 21496 28018
rect 21456 27668 21508 27674
rect 21456 27610 21508 27616
rect 21560 27538 21588 28086
rect 21548 27532 21600 27538
rect 21548 27474 21600 27480
rect 21744 27384 21772 31214
rect 21836 30818 21864 31436
rect 21928 30938 21956 31758
rect 22008 31680 22060 31686
rect 22008 31622 22060 31628
rect 22020 30938 22048 31622
rect 21916 30932 21968 30938
rect 21916 30874 21968 30880
rect 22008 30932 22060 30938
rect 22008 30874 22060 30880
rect 21836 30790 21956 30818
rect 21928 28098 21956 30790
rect 22112 29646 22140 31758
rect 22204 31482 22232 32166
rect 22296 31958 22324 32302
rect 22284 31952 22336 31958
rect 22284 31894 22336 31900
rect 22296 31822 22324 31894
rect 22388 31822 22416 35634
rect 22468 34196 22520 34202
rect 22468 34138 22520 34144
rect 22480 33998 22508 34138
rect 22468 33992 22520 33998
rect 22468 33934 22520 33940
rect 22572 33130 22600 37742
rect 22926 37360 22982 37369
rect 22836 37324 22888 37330
rect 22926 37295 22928 37304
rect 22836 37266 22888 37272
rect 22980 37295 22982 37304
rect 22928 37266 22980 37272
rect 22848 36174 22876 37266
rect 22836 36168 22888 36174
rect 22836 36110 22888 36116
rect 22652 36032 22704 36038
rect 22652 35974 22704 35980
rect 22664 35834 22692 35974
rect 22652 35828 22704 35834
rect 22652 35770 22704 35776
rect 22744 35692 22796 35698
rect 22744 35634 22796 35640
rect 22652 34400 22704 34406
rect 22652 34342 22704 34348
rect 22664 33998 22692 34342
rect 22652 33992 22704 33998
rect 22652 33934 22704 33940
rect 22480 33102 22600 33130
rect 22284 31816 22336 31822
rect 22284 31758 22336 31764
rect 22376 31816 22428 31822
rect 22376 31758 22428 31764
rect 22192 31476 22244 31482
rect 22192 31418 22244 31424
rect 22284 31408 22336 31414
rect 22284 31350 22336 31356
rect 22296 31113 22324 31350
rect 22282 31104 22338 31113
rect 22282 31039 22338 31048
rect 22282 29744 22338 29753
rect 22388 29730 22416 31758
rect 22338 29702 22416 29730
rect 22282 29679 22338 29688
rect 22100 29640 22152 29646
rect 22100 29582 22152 29588
rect 22112 29238 22140 29582
rect 22100 29232 22152 29238
rect 22100 29174 22152 29180
rect 22296 29170 22324 29679
rect 22480 29481 22508 33102
rect 22756 32434 22784 35634
rect 23032 35578 23060 37810
rect 23388 37256 23440 37262
rect 23388 37198 23440 37204
rect 23400 36922 23428 37198
rect 23388 36916 23440 36922
rect 23388 36858 23440 36864
rect 23492 36802 23520 37810
rect 23400 36774 23520 36802
rect 23296 36576 23348 36582
rect 23296 36518 23348 36524
rect 23204 36168 23256 36174
rect 23204 36110 23256 36116
rect 23216 35698 23244 36110
rect 23308 35698 23336 36518
rect 23112 35692 23164 35698
rect 23112 35634 23164 35640
rect 23204 35692 23256 35698
rect 23204 35634 23256 35640
rect 23296 35692 23348 35698
rect 23296 35634 23348 35640
rect 22836 35556 22888 35562
rect 22836 35498 22888 35504
rect 22940 35550 23060 35578
rect 22848 35222 22876 35498
rect 22836 35216 22888 35222
rect 22836 35158 22888 35164
rect 22836 34604 22888 34610
rect 22940 34592 22968 35550
rect 23020 35488 23072 35494
rect 23020 35430 23072 35436
rect 22888 34564 22968 34592
rect 22836 34546 22888 34552
rect 22848 33844 22876 34546
rect 22926 34096 22982 34105
rect 22926 34031 22982 34040
rect 22940 33998 22968 34031
rect 22928 33992 22980 33998
rect 22928 33934 22980 33940
rect 22928 33856 22980 33862
rect 22848 33816 22928 33844
rect 22928 33798 22980 33804
rect 22834 33552 22890 33561
rect 22834 33487 22890 33496
rect 22744 32428 22796 32434
rect 22664 32388 22744 32416
rect 22664 31822 22692 32388
rect 22744 32370 22796 32376
rect 22848 32314 22876 33487
rect 22940 33318 22968 33798
rect 22928 33312 22980 33318
rect 22928 33254 22980 33260
rect 23032 32434 23060 35430
rect 23124 34202 23152 35634
rect 23216 34678 23244 35634
rect 23204 34672 23256 34678
rect 23204 34614 23256 34620
rect 23112 34196 23164 34202
rect 23112 34138 23164 34144
rect 23124 32484 23152 34138
rect 23202 33824 23258 33833
rect 23202 33759 23258 33768
rect 23216 33590 23244 33759
rect 23204 33584 23256 33590
rect 23204 33526 23256 33532
rect 23204 32496 23256 32502
rect 23124 32456 23204 32484
rect 23204 32438 23256 32444
rect 22928 32428 22980 32434
rect 22928 32370 22980 32376
rect 23020 32428 23072 32434
rect 23020 32370 23072 32376
rect 22756 32286 22876 32314
rect 22756 31958 22784 32286
rect 22836 32224 22888 32230
rect 22836 32166 22888 32172
rect 22744 31952 22796 31958
rect 22744 31894 22796 31900
rect 22652 31816 22704 31822
rect 22652 31758 22704 31764
rect 22560 31680 22612 31686
rect 22560 31622 22612 31628
rect 22652 31680 22704 31686
rect 22652 31622 22704 31628
rect 22572 31278 22600 31622
rect 22664 31346 22692 31622
rect 22848 31346 22876 32166
rect 22652 31340 22704 31346
rect 22652 31282 22704 31288
rect 22836 31340 22888 31346
rect 22836 31282 22888 31288
rect 22560 31272 22612 31278
rect 22560 31214 22612 31220
rect 22652 31136 22704 31142
rect 22652 31078 22704 31084
rect 22560 30796 22612 30802
rect 22560 30738 22612 30744
rect 22466 29472 22522 29481
rect 22466 29407 22522 29416
rect 22572 29306 22600 30738
rect 22468 29300 22520 29306
rect 22468 29242 22520 29248
rect 22560 29300 22612 29306
rect 22560 29242 22612 29248
rect 22008 29164 22060 29170
rect 22008 29106 22060 29112
rect 22192 29164 22244 29170
rect 22192 29106 22244 29112
rect 22284 29164 22336 29170
rect 22284 29106 22336 29112
rect 22020 28694 22048 29106
rect 22008 28688 22060 28694
rect 22008 28630 22060 28636
rect 22204 28218 22232 29106
rect 22376 28416 22428 28422
rect 22376 28358 22428 28364
rect 22192 28212 22244 28218
rect 22192 28154 22244 28160
rect 21928 28070 22048 28098
rect 21916 28008 21968 28014
rect 21916 27950 21968 27956
rect 21928 27713 21956 27950
rect 21914 27704 21970 27713
rect 22020 27674 22048 28070
rect 21914 27639 21970 27648
rect 22008 27668 22060 27674
rect 22008 27610 22060 27616
rect 21824 27396 21876 27402
rect 21744 27356 21824 27384
rect 21824 27338 21876 27344
rect 21732 26988 21784 26994
rect 21732 26930 21784 26936
rect 21548 26240 21600 26246
rect 21548 26182 21600 26188
rect 21454 25800 21510 25809
rect 21454 25735 21510 25744
rect 21468 25294 21496 25735
rect 21560 25294 21588 26182
rect 21640 25696 21692 25702
rect 21640 25638 21692 25644
rect 21456 25288 21508 25294
rect 21456 25230 21508 25236
rect 21548 25288 21600 25294
rect 21548 25230 21600 25236
rect 21454 24984 21510 24993
rect 21454 24919 21456 24928
rect 21508 24919 21510 24928
rect 21456 24890 21508 24896
rect 21652 24886 21680 25638
rect 21744 25158 21772 26930
rect 21836 25294 21864 27338
rect 21916 26852 21968 26858
rect 21916 26794 21968 26800
rect 21928 26761 21956 26794
rect 21914 26752 21970 26761
rect 21914 26687 21970 26696
rect 22020 26382 22048 27610
rect 22204 27334 22232 28154
rect 22388 28082 22416 28358
rect 22480 28082 22508 29242
rect 22376 28076 22428 28082
rect 22376 28018 22428 28024
rect 22468 28076 22520 28082
rect 22468 28018 22520 28024
rect 22374 27840 22430 27849
rect 22374 27775 22430 27784
rect 22192 27328 22244 27334
rect 22192 27270 22244 27276
rect 22388 26994 22416 27775
rect 22376 26988 22428 26994
rect 22376 26930 22428 26936
rect 22664 26874 22692 31078
rect 22940 29782 22968 32370
rect 23032 32337 23060 32370
rect 23018 32328 23074 32337
rect 23018 32263 23074 32272
rect 23202 32328 23258 32337
rect 23202 32263 23204 32272
rect 23256 32263 23258 32272
rect 23204 32234 23256 32240
rect 23020 31952 23072 31958
rect 23308 31906 23336 35634
rect 23400 35562 23428 36774
rect 23572 36032 23624 36038
rect 23572 35974 23624 35980
rect 23584 35698 23612 35974
rect 23676 35766 23704 37810
rect 23848 37664 23900 37670
rect 23848 37606 23900 37612
rect 23860 37330 23888 37606
rect 23848 37324 23900 37330
rect 23848 37266 23900 37272
rect 23756 37188 23808 37194
rect 23756 37130 23808 37136
rect 23664 35760 23716 35766
rect 23664 35702 23716 35708
rect 23572 35692 23624 35698
rect 23572 35634 23624 35640
rect 23388 35556 23440 35562
rect 23388 35498 23440 35504
rect 23400 33998 23428 35498
rect 23480 35488 23532 35494
rect 23480 35430 23532 35436
rect 23492 35170 23520 35430
rect 23492 35154 23612 35170
rect 23492 35148 23624 35154
rect 23492 35142 23572 35148
rect 23572 35090 23624 35096
rect 23480 34944 23532 34950
rect 23480 34886 23532 34892
rect 23572 34944 23624 34950
rect 23572 34886 23624 34892
rect 23492 34649 23520 34886
rect 23478 34640 23534 34649
rect 23478 34575 23534 34584
rect 23480 34468 23532 34474
rect 23480 34410 23532 34416
rect 23388 33992 23440 33998
rect 23388 33934 23440 33940
rect 23492 33930 23520 34410
rect 23480 33924 23532 33930
rect 23480 33866 23532 33872
rect 23388 33856 23440 33862
rect 23388 33798 23440 33804
rect 23400 33425 23428 33798
rect 23492 33697 23520 33866
rect 23478 33688 23534 33697
rect 23478 33623 23534 33632
rect 23584 33454 23612 34886
rect 23768 34746 23796 37130
rect 23952 35816 23980 37810
rect 24032 37256 24084 37262
rect 24032 37198 24084 37204
rect 24044 36582 24072 37198
rect 24032 36576 24084 36582
rect 24032 36518 24084 36524
rect 24136 36106 24164 37810
rect 25228 37800 25280 37806
rect 25884 37754 25912 37810
rect 25228 37742 25280 37748
rect 24584 37664 24636 37670
rect 24584 37606 24636 37612
rect 24308 37256 24360 37262
rect 24308 37198 24360 37204
rect 24216 36644 24268 36650
rect 24216 36586 24268 36592
rect 24228 36310 24256 36586
rect 24216 36304 24268 36310
rect 24216 36246 24268 36252
rect 24124 36100 24176 36106
rect 24124 36042 24176 36048
rect 23952 35788 24072 35816
rect 23940 35692 23992 35698
rect 23940 35634 23992 35640
rect 23756 34740 23808 34746
rect 23756 34682 23808 34688
rect 23756 34400 23808 34406
rect 23756 34342 23808 34348
rect 23846 34368 23902 34377
rect 23664 34196 23716 34202
rect 23664 34138 23716 34144
rect 23676 33998 23704 34138
rect 23664 33992 23716 33998
rect 23664 33934 23716 33940
rect 23480 33448 23532 33454
rect 23386 33416 23442 33425
rect 23480 33390 23532 33396
rect 23572 33448 23624 33454
rect 23572 33390 23624 33396
rect 23676 33402 23704 33934
rect 23768 33522 23796 34342
rect 23846 34303 23902 34312
rect 23860 33998 23888 34303
rect 23848 33992 23900 33998
rect 23848 33934 23900 33940
rect 23848 33856 23900 33862
rect 23848 33798 23900 33804
rect 23860 33522 23888 33798
rect 23952 33561 23980 35634
rect 23938 33552 23994 33561
rect 23756 33516 23808 33522
rect 23756 33458 23808 33464
rect 23848 33516 23900 33522
rect 23938 33487 23994 33496
rect 23848 33458 23900 33464
rect 24044 33402 24072 35788
rect 24124 35488 24176 35494
rect 24124 35430 24176 35436
rect 24136 35222 24164 35430
rect 24124 35216 24176 35222
rect 24124 35158 24176 35164
rect 24124 34604 24176 34610
rect 24124 34546 24176 34552
rect 23386 33351 23442 33360
rect 23492 33114 23520 33390
rect 23676 33374 23888 33402
rect 23756 33312 23808 33318
rect 23756 33254 23808 33260
rect 23480 33108 23532 33114
rect 23480 33050 23532 33056
rect 23388 32904 23440 32910
rect 23388 32846 23440 32852
rect 23400 32570 23428 32846
rect 23388 32564 23440 32570
rect 23388 32506 23440 32512
rect 23020 31894 23072 31900
rect 22928 29776 22980 29782
rect 22928 29718 22980 29724
rect 22744 29504 22796 29510
rect 22744 29446 22796 29452
rect 22836 29504 22888 29510
rect 22836 29446 22888 29452
rect 22756 29306 22784 29446
rect 22744 29300 22796 29306
rect 22744 29242 22796 29248
rect 22742 28656 22798 28665
rect 22742 28591 22798 28600
rect 22756 28558 22784 28591
rect 22744 28552 22796 28558
rect 22744 28494 22796 28500
rect 22112 26846 22692 26874
rect 22008 26376 22060 26382
rect 22008 26318 22060 26324
rect 21824 25288 21876 25294
rect 21824 25230 21876 25236
rect 22008 25288 22060 25294
rect 22008 25230 22060 25236
rect 21732 25152 21784 25158
rect 21732 25094 21784 25100
rect 21836 24954 21864 25230
rect 21824 24948 21876 24954
rect 21824 24890 21876 24896
rect 21640 24880 21692 24886
rect 21640 24822 21692 24828
rect 21456 24404 21508 24410
rect 21456 24346 21508 24352
rect 21088 24336 21140 24342
rect 21088 24278 21140 24284
rect 21364 24336 21416 24342
rect 21364 24278 21416 24284
rect 20720 24200 20772 24206
rect 20720 24142 20772 24148
rect 20732 23730 20760 24142
rect 21100 23798 21128 24278
rect 21088 23792 21140 23798
rect 21088 23734 21140 23740
rect 20720 23724 20772 23730
rect 20720 23666 20772 23672
rect 20812 23724 20864 23730
rect 20812 23666 20864 23672
rect 20732 23322 20760 23666
rect 20824 23322 20852 23666
rect 21468 23662 21496 24346
rect 22020 23730 22048 25230
rect 22008 23724 22060 23730
rect 22008 23666 22060 23672
rect 21456 23656 21508 23662
rect 21456 23598 21508 23604
rect 20720 23316 20772 23322
rect 20720 23258 20772 23264
rect 20812 23316 20864 23322
rect 20812 23258 20864 23264
rect 20628 23112 20680 23118
rect 20628 23054 20680 23060
rect 22020 22982 22048 23666
rect 22008 22976 22060 22982
rect 22008 22918 22060 22924
rect 20720 22636 20772 22642
rect 20720 22578 20772 22584
rect 21916 22636 21968 22642
rect 21916 22578 21968 22584
rect 20536 21140 20588 21146
rect 20536 21082 20588 21088
rect 20548 20942 20576 21082
rect 20536 20936 20588 20942
rect 20536 20878 20588 20884
rect 20548 20448 20576 20878
rect 20628 20460 20680 20466
rect 20548 20420 20628 20448
rect 20628 20402 20680 20408
rect 20628 19848 20680 19854
rect 20628 19790 20680 19796
rect 20640 18834 20668 19790
rect 20732 18970 20760 22578
rect 20996 21548 21048 21554
rect 20996 21490 21048 21496
rect 21008 21026 21036 21490
rect 21928 21146 21956 22578
rect 22008 22024 22060 22030
rect 22008 21966 22060 21972
rect 22020 21146 22048 21966
rect 21088 21140 21140 21146
rect 21916 21140 21968 21146
rect 21140 21100 21404 21128
rect 21088 21082 21140 21088
rect 21008 21010 21220 21026
rect 20904 21004 20956 21010
rect 20904 20946 20956 20952
rect 21008 21004 21232 21010
rect 21008 20998 21180 21004
rect 20812 20868 20864 20874
rect 20812 20810 20864 20816
rect 20824 20058 20852 20810
rect 20916 20466 20944 20946
rect 21008 20466 21036 20998
rect 21180 20946 21232 20952
rect 21376 20942 21404 21100
rect 21916 21082 21968 21088
rect 22008 21140 22060 21146
rect 22008 21082 22060 21088
rect 21824 21072 21876 21078
rect 21824 21014 21876 21020
rect 21364 20936 21416 20942
rect 21364 20878 21416 20884
rect 21456 20936 21508 20942
rect 21456 20878 21508 20884
rect 21088 20868 21140 20874
rect 21088 20810 21140 20816
rect 21272 20868 21324 20874
rect 21272 20810 21324 20816
rect 21100 20602 21128 20810
rect 21088 20596 21140 20602
rect 21088 20538 21140 20544
rect 20904 20460 20956 20466
rect 20904 20402 20956 20408
rect 20996 20460 21048 20466
rect 20996 20402 21048 20408
rect 20812 20052 20864 20058
rect 21100 20040 21128 20538
rect 21284 20398 21312 20810
rect 21272 20392 21324 20398
rect 21272 20334 21324 20340
rect 21468 20330 21496 20878
rect 21456 20324 21508 20330
rect 21456 20266 21508 20272
rect 20812 19994 20864 20000
rect 20916 20012 21128 20040
rect 20916 19446 20944 20012
rect 21088 19916 21140 19922
rect 21088 19858 21140 19864
rect 20904 19440 20956 19446
rect 20904 19382 20956 19388
rect 20720 18964 20772 18970
rect 20720 18906 20772 18912
rect 20628 18828 20680 18834
rect 20628 18770 20680 18776
rect 20916 18714 20944 19382
rect 21100 18970 21128 19858
rect 21836 19854 21864 21014
rect 21928 20874 21956 21082
rect 21916 20868 21968 20874
rect 21916 20810 21968 20816
rect 22006 20360 22062 20369
rect 22006 20295 22062 20304
rect 21824 19848 21876 19854
rect 21824 19790 21876 19796
rect 22020 19514 22048 20295
rect 22008 19508 22060 19514
rect 22008 19450 22060 19456
rect 21732 19168 21784 19174
rect 21732 19110 21784 19116
rect 21088 18964 21140 18970
rect 21088 18906 21140 18912
rect 20548 18686 20944 18714
rect 20548 18290 20576 18686
rect 20628 18624 20680 18630
rect 20628 18566 20680 18572
rect 20536 18284 20588 18290
rect 20536 18226 20588 18232
rect 20260 18080 20312 18086
rect 20260 18022 20312 18028
rect 20352 18080 20404 18086
rect 20352 18022 20404 18028
rect 20444 18080 20496 18086
rect 20444 18022 20496 18028
rect 20364 17898 20392 18022
rect 20364 17870 20484 17898
rect 20260 17740 20312 17746
rect 20260 17682 20312 17688
rect 20076 17672 20128 17678
rect 20076 17614 20128 17620
rect 20168 17672 20220 17678
rect 20168 17614 20220 17620
rect 20180 17270 20208 17614
rect 20168 17264 20220 17270
rect 20168 17206 20220 17212
rect 20168 17128 20220 17134
rect 19996 17088 20168 17116
rect 19996 15892 20024 17088
rect 20168 17070 20220 17076
rect 20272 16776 20300 17682
rect 20456 17134 20484 17870
rect 20352 17128 20404 17134
rect 20352 17070 20404 17076
rect 20444 17128 20496 17134
rect 20444 17070 20496 17076
rect 20088 16748 20300 16776
rect 20088 16590 20116 16748
rect 20168 16652 20220 16658
rect 20168 16594 20220 16600
rect 20076 16584 20128 16590
rect 20076 16526 20128 16532
rect 20180 16164 20208 16594
rect 20364 16590 20392 17070
rect 20352 16584 20404 16590
rect 20352 16526 20404 16532
rect 20456 16538 20484 17070
rect 20548 16658 20576 18226
rect 20640 17746 20668 18566
rect 20812 17876 20864 17882
rect 20812 17818 20864 17824
rect 20628 17740 20680 17746
rect 20628 17682 20680 17688
rect 20824 17202 20852 17818
rect 21100 17338 21128 18906
rect 21744 18902 21772 19110
rect 22112 18970 22140 26846
rect 22192 26784 22244 26790
rect 22192 26726 22244 26732
rect 22204 25906 22232 26726
rect 22652 26512 22704 26518
rect 22652 26454 22704 26460
rect 22376 26376 22428 26382
rect 22376 26318 22428 26324
rect 22192 25900 22244 25906
rect 22192 25842 22244 25848
rect 22284 25696 22336 25702
rect 22284 25638 22336 25644
rect 22192 25288 22244 25294
rect 22192 25230 22244 25236
rect 22204 24614 22232 25230
rect 22192 24608 22244 24614
rect 22192 24550 22244 24556
rect 22192 24404 22244 24410
rect 22192 24346 22244 24352
rect 22204 24313 22232 24346
rect 22190 24304 22246 24313
rect 22190 24239 22246 24248
rect 22192 24064 22244 24070
rect 22192 24006 22244 24012
rect 22204 23594 22232 24006
rect 22192 23588 22244 23594
rect 22192 23530 22244 23536
rect 22296 23118 22324 25638
rect 22388 23186 22416 26318
rect 22664 25906 22692 26454
rect 22756 26353 22784 28494
rect 22742 26344 22798 26353
rect 22742 26279 22798 26288
rect 22848 26081 22876 29446
rect 22940 28098 22968 29718
rect 23032 29560 23060 31894
rect 23216 31878 23336 31906
rect 23216 31822 23244 31878
rect 23204 31816 23256 31822
rect 23124 31776 23204 31804
rect 23124 29850 23152 31776
rect 23388 31816 23440 31822
rect 23204 31758 23256 31764
rect 23308 31776 23388 31804
rect 23204 31680 23256 31686
rect 23204 31622 23256 31628
rect 23216 31346 23244 31622
rect 23308 31482 23336 31776
rect 23388 31758 23440 31764
rect 23296 31476 23348 31482
rect 23296 31418 23348 31424
rect 23386 31376 23442 31385
rect 23308 31346 23386 31362
rect 23204 31340 23256 31346
rect 23204 31282 23256 31288
rect 23296 31340 23386 31346
rect 23348 31334 23386 31340
rect 23386 31311 23442 31320
rect 23296 31282 23348 31288
rect 23308 30802 23336 31282
rect 23388 31272 23440 31278
rect 23388 31214 23440 31220
rect 23296 30796 23348 30802
rect 23296 30738 23348 30744
rect 23400 30734 23428 31214
rect 23388 30728 23440 30734
rect 23388 30670 23440 30676
rect 23386 30424 23442 30433
rect 23386 30359 23442 30368
rect 23112 29844 23164 29850
rect 23112 29786 23164 29792
rect 23204 29640 23256 29646
rect 23204 29582 23256 29588
rect 23294 29608 23350 29617
rect 23112 29572 23164 29578
rect 23032 29532 23112 29560
rect 23112 29514 23164 29520
rect 23110 29472 23166 29481
rect 23110 29407 23166 29416
rect 23020 29164 23072 29170
rect 23020 29106 23072 29112
rect 23032 28218 23060 29106
rect 23020 28212 23072 28218
rect 23020 28154 23072 28160
rect 22940 28070 23060 28098
rect 22928 28008 22980 28014
rect 22926 27976 22928 27985
rect 22980 27976 22982 27985
rect 22926 27911 22982 27920
rect 22834 26072 22890 26081
rect 22834 26007 22890 26016
rect 22652 25900 22704 25906
rect 22652 25842 22704 25848
rect 22560 25764 22612 25770
rect 22560 25706 22612 25712
rect 22652 25764 22704 25770
rect 22652 25706 22704 25712
rect 22572 25498 22600 25706
rect 22560 25492 22612 25498
rect 22560 25434 22612 25440
rect 22664 25430 22692 25706
rect 22940 25480 22968 27911
rect 23032 26625 23060 28070
rect 23018 26616 23074 26625
rect 23018 26551 23074 26560
rect 23020 26308 23072 26314
rect 23020 26250 23072 26256
rect 22848 25452 22968 25480
rect 22652 25424 22704 25430
rect 22652 25366 22704 25372
rect 22560 25220 22612 25226
rect 22560 25162 22612 25168
rect 22572 24886 22600 25162
rect 22560 24880 22612 24886
rect 22560 24822 22612 24828
rect 22572 24274 22600 24822
rect 22560 24268 22612 24274
rect 22560 24210 22612 24216
rect 22848 23769 22876 25452
rect 22928 25356 22980 25362
rect 22928 25298 22980 25304
rect 22940 24954 22968 25298
rect 22928 24948 22980 24954
rect 22928 24890 22980 24896
rect 22834 23760 22890 23769
rect 22834 23695 22890 23704
rect 22928 23724 22980 23730
rect 22928 23666 22980 23672
rect 22376 23180 22428 23186
rect 22376 23122 22428 23128
rect 22468 23180 22520 23186
rect 22468 23122 22520 23128
rect 22284 23112 22336 23118
rect 22284 23054 22336 23060
rect 22284 22976 22336 22982
rect 22284 22918 22336 22924
rect 22192 22636 22244 22642
rect 22192 22578 22244 22584
rect 22204 21690 22232 22578
rect 22192 21684 22244 21690
rect 22192 21626 22244 21632
rect 22192 21480 22244 21486
rect 22190 21448 22192 21457
rect 22244 21448 22246 21457
rect 22190 21383 22246 21392
rect 22192 20936 22244 20942
rect 22192 20878 22244 20884
rect 22100 18964 22152 18970
rect 22100 18906 22152 18912
rect 21732 18896 21784 18902
rect 22204 18850 22232 20878
rect 21732 18838 21784 18844
rect 22112 18822 22232 18850
rect 21640 18760 21692 18766
rect 21640 18702 21692 18708
rect 21180 18692 21232 18698
rect 21180 18634 21232 18640
rect 21192 17678 21220 18634
rect 21548 18080 21600 18086
rect 21548 18022 21600 18028
rect 21180 17672 21232 17678
rect 21180 17614 21232 17620
rect 21088 17332 21140 17338
rect 21088 17274 21140 17280
rect 20812 17196 20864 17202
rect 20812 17138 20864 17144
rect 20720 17060 20772 17066
rect 20720 17002 20772 17008
rect 20732 16726 20760 17002
rect 20720 16720 20772 16726
rect 20720 16662 20772 16668
rect 20536 16652 20588 16658
rect 20536 16594 20588 16600
rect 20628 16652 20680 16658
rect 20628 16594 20680 16600
rect 20456 16510 20576 16538
rect 20352 16176 20404 16182
rect 20180 16136 20352 16164
rect 20352 16118 20404 16124
rect 20444 16108 20496 16114
rect 20444 16050 20496 16056
rect 20352 15972 20404 15978
rect 20352 15914 20404 15920
rect 20168 15904 20220 15910
rect 19996 15864 20168 15892
rect 20168 15846 20220 15852
rect 20076 15428 20128 15434
rect 20076 15370 20128 15376
rect 20088 15026 20116 15370
rect 20180 15162 20208 15846
rect 20168 15156 20220 15162
rect 20168 15098 20220 15104
rect 20076 15020 20128 15026
rect 20076 14962 20128 14968
rect 19984 13320 20036 13326
rect 19984 13262 20036 13268
rect 20076 13320 20128 13326
rect 20076 13262 20128 13268
rect 19996 12646 20024 13262
rect 20088 12986 20116 13262
rect 20076 12980 20128 12986
rect 20076 12922 20128 12928
rect 20260 12708 20312 12714
rect 20260 12650 20312 12656
rect 19984 12640 20036 12646
rect 19984 12582 20036 12588
rect 20076 12164 20128 12170
rect 20076 12106 20128 12112
rect 19892 11280 19944 11286
rect 19892 11222 19944 11228
rect 20088 11150 20116 12106
rect 20272 11830 20300 12650
rect 20364 11898 20392 15914
rect 20456 14906 20484 16050
rect 20548 16046 20576 16510
rect 20536 16040 20588 16046
rect 20536 15982 20588 15988
rect 20548 15434 20576 15982
rect 20640 15570 20668 16594
rect 20732 16250 20760 16662
rect 20812 16584 20864 16590
rect 20812 16526 20864 16532
rect 20996 16584 21048 16590
rect 20996 16526 21048 16532
rect 20720 16244 20772 16250
rect 20720 16186 20772 16192
rect 20732 15910 20760 16186
rect 20824 15994 20852 16526
rect 20904 16448 20956 16454
rect 20904 16390 20956 16396
rect 20916 16114 20944 16390
rect 20904 16108 20956 16114
rect 20904 16050 20956 16056
rect 21008 16046 21036 16526
rect 20996 16040 21048 16046
rect 20824 15966 20944 15994
rect 20996 15982 21048 15988
rect 20720 15904 20772 15910
rect 20720 15846 20772 15852
rect 20628 15564 20680 15570
rect 20628 15506 20680 15512
rect 20536 15428 20588 15434
rect 20536 15370 20588 15376
rect 20456 14878 20668 14906
rect 20536 14816 20588 14822
rect 20536 14758 20588 14764
rect 20548 14550 20576 14758
rect 20640 14550 20668 14878
rect 20812 14816 20864 14822
rect 20812 14758 20864 14764
rect 20536 14544 20588 14550
rect 20536 14486 20588 14492
rect 20628 14544 20680 14550
rect 20628 14486 20680 14492
rect 20444 14340 20496 14346
rect 20444 14282 20496 14288
rect 20456 13938 20484 14282
rect 20548 14006 20576 14486
rect 20536 14000 20588 14006
rect 20536 13942 20588 13948
rect 20640 13954 20668 14486
rect 20444 13932 20496 13938
rect 20444 13874 20496 13880
rect 20456 13462 20484 13874
rect 20444 13456 20496 13462
rect 20444 13398 20496 13404
rect 20548 13326 20576 13942
rect 20640 13938 20760 13954
rect 20640 13932 20772 13938
rect 20640 13926 20720 13932
rect 20720 13874 20772 13880
rect 20628 13388 20680 13394
rect 20628 13330 20680 13336
rect 20536 13320 20588 13326
rect 20536 13262 20588 13268
rect 20352 11892 20404 11898
rect 20352 11834 20404 11840
rect 20260 11824 20312 11830
rect 20260 11766 20312 11772
rect 20536 11212 20588 11218
rect 20536 11154 20588 11160
rect 19524 11144 19576 11150
rect 19524 11086 19576 11092
rect 20076 11144 20128 11150
rect 20076 11086 20128 11092
rect 19156 10804 19208 10810
rect 19156 10746 19208 10752
rect 18328 10668 18380 10674
rect 18328 10610 18380 10616
rect 18512 10668 18564 10674
rect 18512 10610 18564 10616
rect 18524 10062 18552 10610
rect 18236 10056 18288 10062
rect 18236 9998 18288 10004
rect 18420 10056 18472 10062
rect 18420 9998 18472 10004
rect 18512 10056 18564 10062
rect 18512 9998 18564 10004
rect 18236 9512 18288 9518
rect 18236 9454 18288 9460
rect 18248 9178 18276 9454
rect 18236 9172 18288 9178
rect 18236 9114 18288 9120
rect 18144 8968 18196 8974
rect 18144 8910 18196 8916
rect 18432 8634 18460 9998
rect 18524 9586 18552 9998
rect 18696 9920 18748 9926
rect 18696 9862 18748 9868
rect 18708 9722 18736 9862
rect 18696 9716 18748 9722
rect 18696 9658 18748 9664
rect 18512 9580 18564 9586
rect 18512 9522 18564 9528
rect 18880 9512 18932 9518
rect 18878 9480 18880 9489
rect 18932 9480 18934 9489
rect 18878 9415 18934 9424
rect 18512 9376 18564 9382
rect 18512 9318 18564 9324
rect 18524 9110 18552 9318
rect 18512 9104 18564 9110
rect 18512 9046 18564 9052
rect 18420 8628 18472 8634
rect 18420 8570 18472 8576
rect 18970 8528 19026 8537
rect 19168 8498 19196 10746
rect 20088 9926 20116 11086
rect 20168 11008 20220 11014
rect 20220 10968 20300 10996
rect 20168 10950 20220 10956
rect 20168 10464 20220 10470
rect 20168 10406 20220 10412
rect 20180 10062 20208 10406
rect 20168 10056 20220 10062
rect 20168 9998 20220 10004
rect 20076 9920 20128 9926
rect 20076 9862 20128 9868
rect 19984 9648 20036 9654
rect 19984 9590 20036 9596
rect 19432 9512 19484 9518
rect 19432 9454 19484 9460
rect 18970 8463 18972 8472
rect 19024 8463 19026 8472
rect 19156 8492 19208 8498
rect 18972 8434 19024 8440
rect 19156 8434 19208 8440
rect 17592 7880 17644 7886
rect 17592 7822 17644 7828
rect 17776 7880 17828 7886
rect 17776 7822 17828 7828
rect 17316 7744 17368 7750
rect 17316 7686 17368 7692
rect 17328 6934 17356 7686
rect 17788 7410 17816 7822
rect 18512 7472 18564 7478
rect 18512 7414 18564 7420
rect 17776 7404 17828 7410
rect 17776 7346 17828 7352
rect 17788 7002 17816 7346
rect 17868 7200 17920 7206
rect 17868 7142 17920 7148
rect 18052 7200 18104 7206
rect 18052 7142 18104 7148
rect 17776 6996 17828 7002
rect 17776 6938 17828 6944
rect 17316 6928 17368 6934
rect 17316 6870 17368 6876
rect 17880 6866 17908 7142
rect 18064 7002 18092 7142
rect 18052 6996 18104 7002
rect 18052 6938 18104 6944
rect 18234 6896 18290 6905
rect 17868 6860 17920 6866
rect 18234 6831 18290 6840
rect 17868 6802 17920 6808
rect 17880 6458 17908 6802
rect 18248 6798 18276 6831
rect 18524 6798 18552 7414
rect 18696 7336 18748 7342
rect 18696 7278 18748 7284
rect 18236 6792 18288 6798
rect 18236 6734 18288 6740
rect 18512 6792 18564 6798
rect 18512 6734 18564 6740
rect 17868 6452 17920 6458
rect 17868 6394 17920 6400
rect 18248 6338 18276 6734
rect 18524 6390 18552 6734
rect 18708 6458 18736 7278
rect 18984 6798 19012 8434
rect 19168 7546 19196 8434
rect 19156 7540 19208 7546
rect 19156 7482 19208 7488
rect 18972 6792 19024 6798
rect 18972 6734 19024 6740
rect 18696 6452 18748 6458
rect 18696 6394 18748 6400
rect 18156 6322 18276 6338
rect 18512 6384 18564 6390
rect 18512 6326 18564 6332
rect 18984 6322 19012 6734
rect 18144 6316 18276 6322
rect 18196 6310 18276 6316
rect 18972 6316 19024 6322
rect 18144 6258 18196 6264
rect 18972 6258 19024 6264
rect 18144 6180 18196 6186
rect 18144 6122 18196 6128
rect 18156 5914 18184 6122
rect 18144 5908 18196 5914
rect 18144 5850 18196 5856
rect 19340 5772 19392 5778
rect 19340 5714 19392 5720
rect 19352 5302 19380 5714
rect 19340 5296 19392 5302
rect 19340 5238 19392 5244
rect 19444 4826 19472 9454
rect 19616 9376 19668 9382
rect 19616 9318 19668 9324
rect 19524 8968 19576 8974
rect 19524 8910 19576 8916
rect 19536 8566 19564 8910
rect 19524 8560 19576 8566
rect 19524 8502 19576 8508
rect 19524 8288 19576 8294
rect 19524 8230 19576 8236
rect 19536 7954 19564 8230
rect 19524 7948 19576 7954
rect 19524 7890 19576 7896
rect 19628 6458 19656 9318
rect 19996 8974 20024 9590
rect 20088 9450 20116 9862
rect 20180 9586 20208 9998
rect 20272 9586 20300 10968
rect 20548 10062 20576 11154
rect 20640 10062 20668 13330
rect 20824 12306 20852 14758
rect 20916 14414 20944 15966
rect 21008 15026 21036 15982
rect 21100 15706 21128 17274
rect 21560 16114 21588 18022
rect 21652 17882 21680 18702
rect 22112 17882 22140 18822
rect 22192 18624 22244 18630
rect 22192 18566 22244 18572
rect 21640 17876 21692 17882
rect 21640 17818 21692 17824
rect 22100 17876 22152 17882
rect 22100 17818 22152 17824
rect 21548 16108 21600 16114
rect 21548 16050 21600 16056
rect 22008 16108 22060 16114
rect 22008 16050 22060 16056
rect 21088 15700 21140 15706
rect 21088 15642 21140 15648
rect 22020 15502 22048 16050
rect 22008 15496 22060 15502
rect 22008 15438 22060 15444
rect 20996 15020 21048 15026
rect 20996 14962 21048 14968
rect 21916 15020 21968 15026
rect 21916 14962 21968 14968
rect 21824 14952 21876 14958
rect 21824 14894 21876 14900
rect 21272 14884 21324 14890
rect 21272 14826 21324 14832
rect 20904 14408 20956 14414
rect 20904 14350 20956 14356
rect 21088 14408 21140 14414
rect 21088 14350 21140 14356
rect 20916 13802 20944 14350
rect 21100 14074 21128 14350
rect 21088 14068 21140 14074
rect 21088 14010 21140 14016
rect 20904 13796 20956 13802
rect 20904 13738 20956 13744
rect 20916 13530 20944 13738
rect 20904 13524 20956 13530
rect 20904 13466 20956 13472
rect 21100 13326 21128 14010
rect 21088 13320 21140 13326
rect 21088 13262 21140 13268
rect 21088 13184 21140 13190
rect 21088 13126 21140 13132
rect 21180 13184 21232 13190
rect 21180 13126 21232 13132
rect 21100 12850 21128 13126
rect 21192 12986 21220 13126
rect 21180 12980 21232 12986
rect 21180 12922 21232 12928
rect 21088 12844 21140 12850
rect 21088 12786 21140 12792
rect 20812 12300 20864 12306
rect 20812 12242 20864 12248
rect 20904 12300 20956 12306
rect 20904 12242 20956 12248
rect 20810 10976 20866 10985
rect 20810 10911 20866 10920
rect 20824 10826 20852 10911
rect 20732 10810 20852 10826
rect 20720 10804 20852 10810
rect 20772 10798 20852 10804
rect 20720 10746 20772 10752
rect 20536 10056 20588 10062
rect 20628 10056 20680 10062
rect 20536 9998 20588 10004
rect 20626 10024 20628 10033
rect 20680 10024 20682 10033
rect 20548 9586 20576 9998
rect 20916 9994 20944 12242
rect 20996 11076 21048 11082
rect 20996 11018 21048 11024
rect 21008 10742 21036 11018
rect 20996 10736 21048 10742
rect 20996 10678 21048 10684
rect 21180 10600 21232 10606
rect 21180 10542 21232 10548
rect 21284 10554 21312 14826
rect 21836 14346 21864 14894
rect 21928 14482 21956 14962
rect 22204 14822 22232 18566
rect 22296 16726 22324 22918
rect 22388 22488 22416 23122
rect 22480 22642 22508 23122
rect 22940 23118 22968 23666
rect 22928 23112 22980 23118
rect 22928 23054 22980 23060
rect 22652 23044 22704 23050
rect 22652 22986 22704 22992
rect 22468 22636 22520 22642
rect 22468 22578 22520 22584
rect 22388 22460 22600 22488
rect 22376 22160 22428 22166
rect 22376 22102 22428 22108
rect 22388 22001 22416 22102
rect 22374 21992 22430 22001
rect 22374 21927 22430 21936
rect 22376 21888 22428 21894
rect 22376 21830 22428 21836
rect 22388 21078 22416 21830
rect 22376 21072 22428 21078
rect 22376 21014 22428 21020
rect 22376 20936 22428 20942
rect 22374 20904 22376 20913
rect 22428 20904 22430 20913
rect 22374 20839 22430 20848
rect 22466 19952 22522 19961
rect 22466 19887 22522 19896
rect 22480 19553 22508 19887
rect 22466 19544 22522 19553
rect 22466 19479 22522 19488
rect 22374 19408 22430 19417
rect 22480 19378 22508 19479
rect 22572 19378 22600 22460
rect 22664 22137 22692 22986
rect 22836 22976 22888 22982
rect 22836 22918 22888 22924
rect 22848 22642 22876 22918
rect 22940 22778 22968 23054
rect 22928 22772 22980 22778
rect 22928 22714 22980 22720
rect 22836 22636 22888 22642
rect 22836 22578 22888 22584
rect 22928 22636 22980 22642
rect 22928 22578 22980 22584
rect 22650 22128 22706 22137
rect 22650 22063 22706 22072
rect 22664 22030 22692 22063
rect 22652 22024 22704 22030
rect 22652 21966 22704 21972
rect 22744 22024 22796 22030
rect 22744 21966 22796 21972
rect 22756 21486 22784 21966
rect 22940 21554 22968 22578
rect 22928 21548 22980 21554
rect 22928 21490 22980 21496
rect 22744 21480 22796 21486
rect 22744 21422 22796 21428
rect 22834 21448 22890 21457
rect 22834 21383 22890 21392
rect 22848 21146 22876 21383
rect 22836 21140 22888 21146
rect 22836 21082 22888 21088
rect 22652 21004 22704 21010
rect 22652 20946 22704 20952
rect 22374 19343 22376 19352
rect 22428 19343 22430 19352
rect 22468 19372 22520 19378
rect 22376 19314 22428 19320
rect 22468 19314 22520 19320
rect 22560 19372 22612 19378
rect 22560 19314 22612 19320
rect 22374 19272 22430 19281
rect 22374 19207 22430 19216
rect 22388 18766 22416 19207
rect 22468 18964 22520 18970
rect 22468 18906 22520 18912
rect 22376 18760 22428 18766
rect 22376 18702 22428 18708
rect 22388 18290 22416 18702
rect 22480 18290 22508 18906
rect 22572 18290 22600 19314
rect 22664 18358 22692 20946
rect 22940 20602 22968 21490
rect 22928 20596 22980 20602
rect 22928 20538 22980 20544
rect 22834 20088 22890 20097
rect 22890 20032 22968 20040
rect 22834 20023 22836 20032
rect 22888 20012 22968 20032
rect 22836 19994 22888 20000
rect 22836 19780 22888 19786
rect 22836 19722 22888 19728
rect 22848 19514 22876 19722
rect 22940 19514 22968 20012
rect 22836 19508 22888 19514
rect 22836 19450 22888 19456
rect 22928 19508 22980 19514
rect 22928 19450 22980 19456
rect 22652 18352 22704 18358
rect 22652 18294 22704 18300
rect 22376 18284 22428 18290
rect 22376 18226 22428 18232
rect 22468 18284 22520 18290
rect 22468 18226 22520 18232
rect 22560 18284 22612 18290
rect 22560 18226 22612 18232
rect 22664 17882 22692 18294
rect 22742 17912 22798 17921
rect 22652 17876 22704 17882
rect 22742 17847 22798 17856
rect 22652 17818 22704 17824
rect 22468 17672 22520 17678
rect 22468 17614 22520 17620
rect 22480 16794 22508 17614
rect 22560 17196 22612 17202
rect 22560 17138 22612 17144
rect 22468 16788 22520 16794
rect 22468 16730 22520 16736
rect 22284 16720 22336 16726
rect 22284 16662 22336 16668
rect 22284 16584 22336 16590
rect 22284 16526 22336 16532
rect 22296 16250 22324 16526
rect 22468 16516 22520 16522
rect 22572 16504 22600 17138
rect 22520 16476 22600 16504
rect 22468 16458 22520 16464
rect 22284 16244 22336 16250
rect 22284 16186 22336 16192
rect 22192 14816 22244 14822
rect 22192 14758 22244 14764
rect 21916 14476 21968 14482
rect 21916 14418 21968 14424
rect 21824 14340 21876 14346
rect 21824 14282 21876 14288
rect 21364 13796 21416 13802
rect 21364 13738 21416 13744
rect 21376 13326 21404 13738
rect 21928 13326 21956 14418
rect 22100 13932 22152 13938
rect 22100 13874 22152 13880
rect 21364 13320 21416 13326
rect 21364 13262 21416 13268
rect 21732 13320 21784 13326
rect 21732 13262 21784 13268
rect 21916 13320 21968 13326
rect 21916 13262 21968 13268
rect 21376 12646 21404 13262
rect 21548 13184 21600 13190
rect 21548 13126 21600 13132
rect 21456 12844 21508 12850
rect 21456 12786 21508 12792
rect 21364 12640 21416 12646
rect 21364 12582 21416 12588
rect 21468 12238 21496 12786
rect 21560 12306 21588 13126
rect 21744 12986 21772 13262
rect 21732 12980 21784 12986
rect 21732 12922 21784 12928
rect 21928 12442 21956 13262
rect 22112 12850 22140 13874
rect 22480 13870 22508 16458
rect 22652 16448 22704 16454
rect 22652 16390 22704 16396
rect 22664 15570 22692 16390
rect 22756 15570 22784 17847
rect 23032 16182 23060 26250
rect 23124 26042 23152 29407
rect 23216 29306 23244 29582
rect 23294 29543 23350 29552
rect 23308 29510 23336 29543
rect 23296 29504 23348 29510
rect 23296 29446 23348 29452
rect 23204 29300 23256 29306
rect 23204 29242 23256 29248
rect 23204 28960 23256 28966
rect 23204 28902 23256 28908
rect 23216 28082 23244 28902
rect 23400 28200 23428 30359
rect 23492 29714 23520 33050
rect 23768 32774 23796 33254
rect 23572 32768 23624 32774
rect 23572 32710 23624 32716
rect 23756 32768 23808 32774
rect 23756 32710 23808 32716
rect 23584 32570 23612 32710
rect 23572 32564 23624 32570
rect 23572 32506 23624 32512
rect 23768 32434 23796 32710
rect 23756 32428 23808 32434
rect 23756 32370 23808 32376
rect 23572 31884 23624 31890
rect 23572 31826 23624 31832
rect 23584 30666 23612 31826
rect 23860 31754 23888 33374
rect 23952 33374 24072 33402
rect 23952 33153 23980 33374
rect 24032 33312 24084 33318
rect 24030 33280 24032 33289
rect 24084 33280 24086 33289
rect 24030 33215 24086 33224
rect 23938 33144 23994 33153
rect 24136 33130 24164 34546
rect 23938 33079 23994 33088
rect 24044 33102 24164 33130
rect 23952 31958 23980 33079
rect 23940 31952 23992 31958
rect 23940 31894 23992 31900
rect 23664 31748 23716 31754
rect 23664 31690 23716 31696
rect 23756 31748 23808 31754
rect 23860 31726 23980 31754
rect 23756 31690 23808 31696
rect 23572 30660 23624 30666
rect 23572 30602 23624 30608
rect 23480 29708 23532 29714
rect 23480 29650 23532 29656
rect 23572 29504 23624 29510
rect 23572 29446 23624 29452
rect 23584 29073 23612 29446
rect 23676 29238 23704 31690
rect 23768 31249 23796 31690
rect 23754 31240 23810 31249
rect 23754 31175 23810 31184
rect 23848 30388 23900 30394
rect 23848 30330 23900 30336
rect 23756 29640 23808 29646
rect 23756 29582 23808 29588
rect 23664 29232 23716 29238
rect 23664 29174 23716 29180
rect 23570 29064 23626 29073
rect 23570 28999 23626 29008
rect 23676 28948 23704 29174
rect 23308 28172 23428 28200
rect 23492 28920 23704 28948
rect 23204 28076 23256 28082
rect 23204 28018 23256 28024
rect 23308 26874 23336 28172
rect 23388 28076 23440 28082
rect 23388 28018 23440 28024
rect 23400 27878 23428 28018
rect 23388 27872 23440 27878
rect 23388 27814 23440 27820
rect 23400 27538 23428 27814
rect 23388 27532 23440 27538
rect 23388 27474 23440 27480
rect 23492 27062 23520 28920
rect 23572 28756 23624 28762
rect 23572 28698 23624 28704
rect 23584 28218 23612 28698
rect 23572 28212 23624 28218
rect 23572 28154 23624 28160
rect 23572 28008 23624 28014
rect 23572 27950 23624 27956
rect 23584 27674 23612 27950
rect 23768 27946 23796 29582
rect 23756 27940 23808 27946
rect 23756 27882 23808 27888
rect 23572 27668 23624 27674
rect 23572 27610 23624 27616
rect 23664 27600 23716 27606
rect 23664 27542 23716 27548
rect 23572 27464 23624 27470
rect 23572 27406 23624 27412
rect 23480 27056 23532 27062
rect 23480 26998 23532 27004
rect 23216 26846 23336 26874
rect 23112 26036 23164 26042
rect 23112 25978 23164 25984
rect 23110 25936 23166 25945
rect 23110 25871 23112 25880
rect 23164 25871 23166 25880
rect 23112 25842 23164 25848
rect 23112 24268 23164 24274
rect 23112 24210 23164 24216
rect 23124 23798 23152 24210
rect 23112 23792 23164 23798
rect 23112 23734 23164 23740
rect 23112 23112 23164 23118
rect 23112 23054 23164 23060
rect 23124 22166 23152 23054
rect 23112 22160 23164 22166
rect 23112 22102 23164 22108
rect 23112 21956 23164 21962
rect 23112 21898 23164 21904
rect 23124 21554 23152 21898
rect 23112 21548 23164 21554
rect 23112 21490 23164 21496
rect 23112 21344 23164 21350
rect 23112 21286 23164 21292
rect 23124 20806 23152 21286
rect 23112 20800 23164 20806
rect 23112 20742 23164 20748
rect 23110 20632 23166 20641
rect 23110 20567 23166 20576
rect 23124 20097 23152 20567
rect 23110 20088 23166 20097
rect 23110 20023 23166 20032
rect 23124 19854 23152 20023
rect 23112 19848 23164 19854
rect 23112 19790 23164 19796
rect 23124 17338 23152 19790
rect 23216 17882 23244 26846
rect 23388 25900 23440 25906
rect 23388 25842 23440 25848
rect 23400 24954 23428 25842
rect 23584 25158 23612 27406
rect 23676 25362 23704 27542
rect 23768 26382 23796 27882
rect 23756 26376 23808 26382
rect 23756 26318 23808 26324
rect 23756 26240 23808 26246
rect 23756 26182 23808 26188
rect 23768 26042 23796 26182
rect 23756 26036 23808 26042
rect 23756 25978 23808 25984
rect 23860 25702 23888 30330
rect 23952 28966 23980 31726
rect 24044 30598 24072 33102
rect 24124 32428 24176 32434
rect 24228 32416 24256 36246
rect 24176 32388 24256 32416
rect 24124 32370 24176 32376
rect 24032 30592 24084 30598
rect 24032 30534 24084 30540
rect 24030 30288 24086 30297
rect 24030 30223 24086 30232
rect 24044 29646 24072 30223
rect 24032 29640 24084 29646
rect 24032 29582 24084 29588
rect 24030 29336 24086 29345
rect 24030 29271 24086 29280
rect 24044 29238 24072 29271
rect 24032 29232 24084 29238
rect 24032 29174 24084 29180
rect 23940 28960 23992 28966
rect 23940 28902 23992 28908
rect 23952 28422 23980 28902
rect 23940 28416 23992 28422
rect 23940 28358 23992 28364
rect 24136 27470 24164 32370
rect 24320 32314 24348 37198
rect 24400 37120 24452 37126
rect 24400 37062 24452 37068
rect 24412 32450 24440 37062
rect 24596 36786 24624 37606
rect 24676 37460 24728 37466
rect 24676 37402 24728 37408
rect 24492 36780 24544 36786
rect 24492 36722 24544 36728
rect 24584 36780 24636 36786
rect 24584 36722 24636 36728
rect 24504 36378 24532 36722
rect 24688 36582 24716 37402
rect 25240 37369 25268 37742
rect 25792 37726 25912 37754
rect 26148 37800 26200 37806
rect 26148 37742 26200 37748
rect 25226 37360 25282 37369
rect 24860 37324 24912 37330
rect 25226 37295 25282 37304
rect 24860 37266 24912 37272
rect 24676 36576 24728 36582
rect 24676 36518 24728 36524
rect 24492 36372 24544 36378
rect 24492 36314 24544 36320
rect 24676 36168 24728 36174
rect 24676 36110 24728 36116
rect 24492 36100 24544 36106
rect 24492 36042 24544 36048
rect 24504 32910 24532 36042
rect 24584 33856 24636 33862
rect 24584 33798 24636 33804
rect 24596 32978 24624 33798
rect 24584 32972 24636 32978
rect 24584 32914 24636 32920
rect 24492 32904 24544 32910
rect 24492 32846 24544 32852
rect 24412 32422 24532 32450
rect 24228 32286 24348 32314
rect 24400 32360 24452 32366
rect 24504 32337 24532 32422
rect 24400 32302 24452 32308
rect 24490 32328 24546 32337
rect 24228 31822 24256 32286
rect 24308 32224 24360 32230
rect 24308 32166 24360 32172
rect 24320 32026 24348 32166
rect 24308 32020 24360 32026
rect 24308 31962 24360 31968
rect 24412 31958 24440 32302
rect 24490 32263 24546 32272
rect 24400 31952 24452 31958
rect 24400 31894 24452 31900
rect 24504 31822 24532 32263
rect 24216 31816 24268 31822
rect 24492 31816 24544 31822
rect 24216 31758 24268 31764
rect 24320 31776 24492 31804
rect 24228 30326 24256 31758
rect 24216 30320 24268 30326
rect 24216 30262 24268 30268
rect 24228 29170 24256 30262
rect 24216 29164 24268 29170
rect 24216 29106 24268 29112
rect 24216 29028 24268 29034
rect 24216 28970 24268 28976
rect 24228 28082 24256 28970
rect 24320 28762 24348 31776
rect 24492 31758 24544 31764
rect 24688 31770 24716 36110
rect 24872 35698 24900 37266
rect 25136 36848 25188 36854
rect 25136 36790 25188 36796
rect 24952 36576 25004 36582
rect 24952 36518 25004 36524
rect 24964 36009 24992 36518
rect 25044 36100 25096 36106
rect 25044 36042 25096 36048
rect 24950 36000 25006 36009
rect 24950 35935 25006 35944
rect 25056 35766 25084 36042
rect 25044 35760 25096 35766
rect 25044 35702 25096 35708
rect 24860 35692 24912 35698
rect 24860 35634 24912 35640
rect 25148 34921 25176 36790
rect 25596 36780 25648 36786
rect 25596 36722 25648 36728
rect 25228 36236 25280 36242
rect 25228 36178 25280 36184
rect 25240 35698 25268 36178
rect 25608 36174 25636 36722
rect 25688 36304 25740 36310
rect 25688 36246 25740 36252
rect 25596 36168 25648 36174
rect 25594 36136 25596 36145
rect 25648 36136 25650 36145
rect 25412 36100 25464 36106
rect 25594 36071 25650 36080
rect 25412 36042 25464 36048
rect 25228 35692 25280 35698
rect 25228 35634 25280 35640
rect 25320 35080 25372 35086
rect 25320 35022 25372 35028
rect 25134 34912 25190 34921
rect 25134 34847 25190 34856
rect 25228 34740 25280 34746
rect 25228 34682 25280 34688
rect 24768 34400 24820 34406
rect 24768 34342 24820 34348
rect 24780 34202 24808 34342
rect 24768 34196 24820 34202
rect 24768 34138 24820 34144
rect 25044 32768 25096 32774
rect 25044 32710 25096 32716
rect 24952 32224 25004 32230
rect 24952 32166 25004 32172
rect 24964 31822 24992 32166
rect 24768 31816 24820 31822
rect 24688 31764 24768 31770
rect 24688 31758 24820 31764
rect 24952 31816 25004 31822
rect 24952 31758 25004 31764
rect 24688 31742 24808 31758
rect 24584 31272 24636 31278
rect 24584 31214 24636 31220
rect 24492 30932 24544 30938
rect 24492 30874 24544 30880
rect 24400 30728 24452 30734
rect 24400 30670 24452 30676
rect 24412 29782 24440 30670
rect 24504 30394 24532 30874
rect 24596 30802 24624 31214
rect 24584 30796 24636 30802
rect 24584 30738 24636 30744
rect 24492 30388 24544 30394
rect 24492 30330 24544 30336
rect 24504 29850 24532 30330
rect 24492 29844 24544 29850
rect 24492 29786 24544 29792
rect 24400 29776 24452 29782
rect 24400 29718 24452 29724
rect 24308 28756 24360 28762
rect 24308 28698 24360 28704
rect 24412 28506 24440 29718
rect 24584 29640 24636 29646
rect 24582 29608 24584 29617
rect 24636 29608 24638 29617
rect 24582 29543 24638 29552
rect 24688 28994 24716 31742
rect 25056 30666 25084 32710
rect 25136 31816 25188 31822
rect 25136 31758 25188 31764
rect 25148 30938 25176 31758
rect 25136 30932 25188 30938
rect 25136 30874 25188 30880
rect 25044 30660 25096 30666
rect 25044 30602 25096 30608
rect 24858 30016 24914 30025
rect 24858 29951 24914 29960
rect 24768 29776 24820 29782
rect 24768 29718 24820 29724
rect 24780 29646 24808 29718
rect 24872 29646 24900 29951
rect 24768 29640 24820 29646
rect 24768 29582 24820 29588
rect 24860 29640 24912 29646
rect 24860 29582 24912 29588
rect 25056 29102 25084 30602
rect 25044 29096 25096 29102
rect 24858 29064 24914 29073
rect 25044 29038 25096 29044
rect 24858 28999 24860 29008
rect 24504 28966 24716 28994
rect 24912 28999 24914 29008
rect 24860 28970 24912 28976
rect 24504 28558 24532 28966
rect 24768 28756 24820 28762
rect 24768 28698 24820 28704
rect 24320 28478 24440 28506
rect 24492 28552 24544 28558
rect 24492 28494 24544 28500
rect 24676 28552 24728 28558
rect 24676 28494 24728 28500
rect 24216 28076 24268 28082
rect 24216 28018 24268 28024
rect 24216 27872 24268 27878
rect 24216 27814 24268 27820
rect 24228 27674 24256 27814
rect 24216 27668 24268 27674
rect 24216 27610 24268 27616
rect 24124 27464 24176 27470
rect 24124 27406 24176 27412
rect 24030 26072 24086 26081
rect 24030 26007 24086 26016
rect 24044 25838 24072 26007
rect 24320 25945 24348 28478
rect 24400 28416 24452 28422
rect 24400 28358 24452 28364
rect 24412 28082 24440 28358
rect 24400 28076 24452 28082
rect 24400 28018 24452 28024
rect 24504 27962 24532 28494
rect 24688 28218 24716 28494
rect 24780 28490 24808 28698
rect 24860 28552 24912 28558
rect 24858 28520 24860 28529
rect 24912 28520 24914 28529
rect 24768 28484 24820 28490
rect 24858 28455 24914 28464
rect 24768 28426 24820 28432
rect 24676 28212 24728 28218
rect 24676 28154 24728 28160
rect 24676 28076 24728 28082
rect 24676 28018 24728 28024
rect 24412 27934 24532 27962
rect 24306 25936 24362 25945
rect 24306 25871 24308 25880
rect 24360 25871 24362 25880
rect 24308 25842 24360 25848
rect 24032 25832 24084 25838
rect 24032 25774 24084 25780
rect 23848 25696 23900 25702
rect 23848 25638 23900 25644
rect 23664 25356 23716 25362
rect 23664 25298 23716 25304
rect 23572 25152 23624 25158
rect 23572 25094 23624 25100
rect 23388 24948 23440 24954
rect 23388 24890 23440 24896
rect 23676 24818 23704 25298
rect 23940 25220 23992 25226
rect 23940 25162 23992 25168
rect 23480 24812 23532 24818
rect 23480 24754 23532 24760
rect 23664 24812 23716 24818
rect 23664 24754 23716 24760
rect 23848 24812 23900 24818
rect 23848 24754 23900 24760
rect 23492 24206 23520 24754
rect 23664 24404 23716 24410
rect 23664 24346 23716 24352
rect 23480 24200 23532 24206
rect 23480 24142 23532 24148
rect 23388 23724 23440 23730
rect 23388 23666 23440 23672
rect 23296 23316 23348 23322
rect 23296 23258 23348 23264
rect 23308 22642 23336 23258
rect 23400 23118 23428 23666
rect 23492 23254 23520 24142
rect 23572 23656 23624 23662
rect 23572 23598 23624 23604
rect 23480 23248 23532 23254
rect 23480 23190 23532 23196
rect 23584 23118 23612 23598
rect 23388 23112 23440 23118
rect 23388 23054 23440 23060
rect 23572 23112 23624 23118
rect 23572 23054 23624 23060
rect 23296 22636 23348 22642
rect 23296 22578 23348 22584
rect 23296 21956 23348 21962
rect 23296 21898 23348 21904
rect 23308 21010 23336 21898
rect 23584 21622 23612 23054
rect 23676 22642 23704 24346
rect 23756 24200 23808 24206
rect 23756 24142 23808 24148
rect 23768 23730 23796 24142
rect 23756 23724 23808 23730
rect 23756 23666 23808 23672
rect 23768 22778 23796 23666
rect 23860 23186 23888 24754
rect 23952 24682 23980 25162
rect 24044 24721 24072 25774
rect 24308 25696 24360 25702
rect 24308 25638 24360 25644
rect 24320 24886 24348 25638
rect 24412 25294 24440 27934
rect 24492 27872 24544 27878
rect 24492 27814 24544 27820
rect 24504 26382 24532 27814
rect 24582 26480 24638 26489
rect 24582 26415 24638 26424
rect 24596 26382 24624 26415
rect 24492 26376 24544 26382
rect 24492 26318 24544 26324
rect 24584 26376 24636 26382
rect 24584 26318 24636 26324
rect 24688 26024 24716 28018
rect 24780 27849 24808 28426
rect 24766 27840 24822 27849
rect 24766 27775 24822 27784
rect 25056 27674 25084 29038
rect 25044 27668 25096 27674
rect 25044 27610 25096 27616
rect 25056 27470 25084 27610
rect 25044 27464 25096 27470
rect 25096 27424 25176 27452
rect 25044 27406 25096 27412
rect 24952 26988 25004 26994
rect 24952 26930 25004 26936
rect 24860 26920 24912 26926
rect 24860 26862 24912 26868
rect 24872 26772 24900 26862
rect 24780 26744 24900 26772
rect 24780 26058 24808 26744
rect 24964 26466 24992 26930
rect 25042 26480 25098 26489
rect 24964 26438 25042 26466
rect 24860 26308 24912 26314
rect 24860 26250 24912 26256
rect 24872 26217 24900 26250
rect 24858 26208 24914 26217
rect 24858 26143 24914 26152
rect 24780 26030 24900 26058
rect 24596 25996 24716 26024
rect 24492 25764 24544 25770
rect 24492 25706 24544 25712
rect 24400 25288 24452 25294
rect 24400 25230 24452 25236
rect 24504 24886 24532 25706
rect 24308 24880 24360 24886
rect 24308 24822 24360 24828
rect 24492 24880 24544 24886
rect 24492 24822 24544 24828
rect 24124 24744 24176 24750
rect 24030 24712 24086 24721
rect 23940 24676 23992 24682
rect 24124 24686 24176 24692
rect 24030 24647 24086 24656
rect 23940 24618 23992 24624
rect 24032 24608 24084 24614
rect 24032 24550 24084 24556
rect 24044 24342 24072 24550
rect 24032 24336 24084 24342
rect 24032 24278 24084 24284
rect 23940 24200 23992 24206
rect 23940 24142 23992 24148
rect 23848 23180 23900 23186
rect 23848 23122 23900 23128
rect 23756 22772 23808 22778
rect 23756 22714 23808 22720
rect 23664 22636 23716 22642
rect 23664 22578 23716 22584
rect 23676 22012 23704 22578
rect 23952 22506 23980 24142
rect 24136 23730 24164 24686
rect 24492 23792 24544 23798
rect 24492 23734 24544 23740
rect 24124 23724 24176 23730
rect 24124 23666 24176 23672
rect 24400 23656 24452 23662
rect 24306 23624 24362 23633
rect 24400 23598 24452 23604
rect 24306 23559 24308 23568
rect 24360 23559 24362 23568
rect 24308 23530 24360 23536
rect 24412 23118 24440 23598
rect 24504 23594 24532 23734
rect 24492 23588 24544 23594
rect 24492 23530 24544 23536
rect 24032 23112 24084 23118
rect 24032 23054 24084 23060
rect 24400 23112 24452 23118
rect 24400 23054 24452 23060
rect 24044 22642 24072 23054
rect 24124 22976 24176 22982
rect 24124 22918 24176 22924
rect 24032 22636 24084 22642
rect 24032 22578 24084 22584
rect 23940 22500 23992 22506
rect 23940 22442 23992 22448
rect 24044 22098 24072 22578
rect 24136 22574 24164 22918
rect 24124 22568 24176 22574
rect 24124 22510 24176 22516
rect 24032 22092 24084 22098
rect 24032 22034 24084 22040
rect 24596 22030 24624 25996
rect 24676 25900 24728 25906
rect 24676 25842 24728 25848
rect 24768 25900 24820 25906
rect 24768 25842 24820 25848
rect 24688 24342 24716 25842
rect 24780 25294 24808 25842
rect 24768 25288 24820 25294
rect 24768 25230 24820 25236
rect 24676 24336 24728 24342
rect 24676 24278 24728 24284
rect 24688 23746 24716 24278
rect 24872 24274 24900 26030
rect 24964 25498 24992 26438
rect 25042 26415 25098 26424
rect 25042 26072 25098 26081
rect 25042 26007 25098 26016
rect 24952 25492 25004 25498
rect 24952 25434 25004 25440
rect 24950 25392 25006 25401
rect 24950 25327 25006 25336
rect 24964 25294 24992 25327
rect 24952 25288 25004 25294
rect 24952 25230 25004 25236
rect 24860 24268 24912 24274
rect 24860 24210 24912 24216
rect 24688 23730 24808 23746
rect 24688 23724 24820 23730
rect 24688 23718 24768 23724
rect 24768 23666 24820 23672
rect 24766 22536 24822 22545
rect 24766 22471 24822 22480
rect 24780 22030 24808 22471
rect 24952 22432 25004 22438
rect 24952 22374 25004 22380
rect 23756 22024 23808 22030
rect 23676 21984 23756 22012
rect 23756 21966 23808 21972
rect 24584 22024 24636 22030
rect 24584 21966 24636 21972
rect 24768 22024 24820 22030
rect 24768 21966 24820 21972
rect 23572 21616 23624 21622
rect 23572 21558 23624 21564
rect 23296 21004 23348 21010
rect 23296 20946 23348 20952
rect 23768 20466 23796 21966
rect 24596 21078 24624 21966
rect 24676 21888 24728 21894
rect 24676 21830 24728 21836
rect 24584 21072 24636 21078
rect 24584 21014 24636 21020
rect 24688 21010 24716 21830
rect 24768 21616 24820 21622
rect 24768 21558 24820 21564
rect 24676 21004 24728 21010
rect 24676 20946 24728 20952
rect 24400 20936 24452 20942
rect 24400 20878 24452 20884
rect 24412 20602 24440 20878
rect 24400 20596 24452 20602
rect 24400 20538 24452 20544
rect 24412 20466 24440 20538
rect 24492 20528 24544 20534
rect 24492 20470 24544 20476
rect 23756 20460 23808 20466
rect 23676 20420 23756 20448
rect 23296 20256 23348 20262
rect 23296 20198 23348 20204
rect 23478 20224 23534 20233
rect 23308 19961 23336 20198
rect 23478 20159 23534 20168
rect 23492 20058 23520 20159
rect 23480 20052 23532 20058
rect 23480 19994 23532 20000
rect 23294 19952 23350 19961
rect 23294 19887 23296 19896
rect 23348 19887 23350 19896
rect 23296 19858 23348 19864
rect 23204 17876 23256 17882
rect 23204 17818 23256 17824
rect 23202 17640 23258 17649
rect 23202 17575 23258 17584
rect 23112 17332 23164 17338
rect 23112 17274 23164 17280
rect 23112 16720 23164 16726
rect 23112 16662 23164 16668
rect 23020 16176 23072 16182
rect 23020 16118 23072 16124
rect 22928 15904 22980 15910
rect 22928 15846 22980 15852
rect 22652 15564 22704 15570
rect 22652 15506 22704 15512
rect 22744 15564 22796 15570
rect 22744 15506 22796 15512
rect 22756 15314 22784 15506
rect 22940 15366 22968 15846
rect 23032 15502 23060 16118
rect 23020 15496 23072 15502
rect 23020 15438 23072 15444
rect 22664 15286 22784 15314
rect 22928 15360 22980 15366
rect 22928 15302 22980 15308
rect 22560 14000 22612 14006
rect 22560 13942 22612 13948
rect 22468 13864 22520 13870
rect 22468 13806 22520 13812
rect 22480 12850 22508 13806
rect 22100 12844 22152 12850
rect 22100 12786 22152 12792
rect 22468 12844 22520 12850
rect 22468 12786 22520 12792
rect 21916 12436 21968 12442
rect 21916 12378 21968 12384
rect 21548 12300 21600 12306
rect 21548 12242 21600 12248
rect 21456 12232 21508 12238
rect 21456 12174 21508 12180
rect 22112 12170 22140 12786
rect 22100 12164 22152 12170
rect 22100 12106 22152 12112
rect 22192 12096 22244 12102
rect 22192 12038 22244 12044
rect 22100 11348 22152 11354
rect 22100 11290 22152 11296
rect 22112 11082 22140 11290
rect 22204 11150 22232 12038
rect 22480 11286 22508 12786
rect 22284 11280 22336 11286
rect 22284 11222 22336 11228
rect 22468 11280 22520 11286
rect 22468 11222 22520 11228
rect 22192 11144 22244 11150
rect 22192 11086 22244 11092
rect 22100 11076 22152 11082
rect 22100 11018 22152 11024
rect 21824 11008 21876 11014
rect 21824 10950 21876 10956
rect 22098 10976 22154 10985
rect 21836 10826 21864 10950
rect 22098 10911 22154 10920
rect 21652 10798 21864 10826
rect 21652 10606 21680 10798
rect 22008 10736 22060 10742
rect 22006 10704 22008 10713
rect 22060 10704 22062 10713
rect 22006 10639 22062 10648
rect 21640 10600 21692 10606
rect 21088 10464 21140 10470
rect 21088 10406 21140 10412
rect 20626 9959 20682 9968
rect 20904 9988 20956 9994
rect 20904 9930 20956 9936
rect 20168 9580 20220 9586
rect 20168 9522 20220 9528
rect 20260 9580 20312 9586
rect 20260 9522 20312 9528
rect 20536 9580 20588 9586
rect 20536 9522 20588 9528
rect 20076 9444 20128 9450
rect 20076 9386 20128 9392
rect 20088 8974 20116 9386
rect 19984 8968 20036 8974
rect 19984 8910 20036 8916
rect 20076 8968 20128 8974
rect 20076 8910 20128 8916
rect 19892 8900 19944 8906
rect 19892 8842 19944 8848
rect 19708 8832 19760 8838
rect 19760 8792 19840 8820
rect 19708 8774 19760 8780
rect 19708 7880 19760 7886
rect 19708 7822 19760 7828
rect 19720 7410 19748 7822
rect 19708 7404 19760 7410
rect 19708 7346 19760 7352
rect 19812 6458 19840 8792
rect 19904 8566 19932 8842
rect 19996 8566 20024 8910
rect 20272 8906 20300 9522
rect 20812 9172 20864 9178
rect 20812 9114 20864 9120
rect 20260 8900 20312 8906
rect 20260 8842 20312 8848
rect 19892 8560 19944 8566
rect 19892 8502 19944 8508
rect 19984 8560 20036 8566
rect 19984 8502 20036 8508
rect 20824 8498 20852 9114
rect 20812 8492 20864 8498
rect 20812 8434 20864 8440
rect 20628 7948 20680 7954
rect 20628 7890 20680 7896
rect 20536 7744 20588 7750
rect 20536 7686 20588 7692
rect 20548 7206 20576 7686
rect 20640 7410 20668 7890
rect 20628 7404 20680 7410
rect 20628 7346 20680 7352
rect 20536 7200 20588 7206
rect 20536 7142 20588 7148
rect 19984 6860 20036 6866
rect 19984 6802 20036 6808
rect 19996 6458 20024 6802
rect 19616 6452 19668 6458
rect 19616 6394 19668 6400
rect 19800 6452 19852 6458
rect 19800 6394 19852 6400
rect 19984 6452 20036 6458
rect 19984 6394 20036 6400
rect 19524 6112 19576 6118
rect 19524 6054 19576 6060
rect 19536 5778 19564 6054
rect 19524 5772 19576 5778
rect 19524 5714 19576 5720
rect 19536 5302 19564 5714
rect 19628 5574 19656 6394
rect 19812 5778 19840 6394
rect 19800 5772 19852 5778
rect 19800 5714 19852 5720
rect 20548 5710 20576 7142
rect 20640 6798 20668 7346
rect 20628 6792 20680 6798
rect 20628 6734 20680 6740
rect 20076 5704 20128 5710
rect 20076 5646 20128 5652
rect 20444 5704 20496 5710
rect 20444 5646 20496 5652
rect 20536 5704 20588 5710
rect 20536 5646 20588 5652
rect 19616 5568 19668 5574
rect 19616 5510 19668 5516
rect 19524 5296 19576 5302
rect 19524 5238 19576 5244
rect 19892 5024 19944 5030
rect 19892 4966 19944 4972
rect 19432 4820 19484 4826
rect 19432 4762 19484 4768
rect 19904 4758 19932 4966
rect 19892 4752 19944 4758
rect 19892 4694 19944 4700
rect 20088 4554 20116 5646
rect 20456 5370 20484 5646
rect 20168 5364 20220 5370
rect 20168 5306 20220 5312
rect 20444 5364 20496 5370
rect 20444 5306 20496 5312
rect 20180 4826 20208 5306
rect 20168 4820 20220 4826
rect 20168 4762 20220 4768
rect 20548 4554 20576 5646
rect 20824 4622 20852 8434
rect 20916 8294 20944 9930
rect 21100 9654 21128 10406
rect 21192 10062 21220 10542
rect 21284 10526 21588 10554
rect 21640 10542 21692 10548
rect 21560 10470 21588 10526
rect 21456 10464 21508 10470
rect 21456 10406 21508 10412
rect 21548 10464 21600 10470
rect 21548 10406 21600 10412
rect 21468 10062 21496 10406
rect 21180 10056 21232 10062
rect 21180 9998 21232 10004
rect 21456 10056 21508 10062
rect 21456 9998 21508 10004
rect 21088 9648 21140 9654
rect 21088 9590 21140 9596
rect 21100 9178 21128 9590
rect 21088 9172 21140 9178
rect 21088 9114 21140 9120
rect 20904 8288 20956 8294
rect 20904 8230 20956 8236
rect 21100 7546 21128 9114
rect 21468 8566 21496 9998
rect 21456 8560 21508 8566
rect 21456 8502 21508 8508
rect 21468 7886 21496 8502
rect 21560 8430 21588 10406
rect 21652 10010 21680 10542
rect 22008 10464 22060 10470
rect 22008 10406 22060 10412
rect 22020 10266 22048 10406
rect 22008 10260 22060 10266
rect 22008 10202 22060 10208
rect 21916 10056 21968 10062
rect 21914 10024 21916 10033
rect 21968 10024 21970 10033
rect 21652 9982 21864 10010
rect 21652 9654 21680 9982
rect 21836 9926 21864 9982
rect 21914 9959 21970 9968
rect 22112 9926 22140 10911
rect 22192 10532 22244 10538
rect 22192 10474 22244 10480
rect 22204 10441 22232 10474
rect 22190 10432 22246 10441
rect 22190 10367 22246 10376
rect 22192 10192 22244 10198
rect 22192 10134 22244 10140
rect 21824 9920 21876 9926
rect 21824 9862 21876 9868
rect 22100 9920 22152 9926
rect 22100 9862 22152 9868
rect 21640 9648 21692 9654
rect 21640 9590 21692 9596
rect 22100 9172 22152 9178
rect 22100 9114 22152 9120
rect 21824 8492 21876 8498
rect 21824 8434 21876 8440
rect 22008 8492 22060 8498
rect 22008 8434 22060 8440
rect 21548 8424 21600 8430
rect 21836 8401 21864 8434
rect 21548 8366 21600 8372
rect 21822 8392 21878 8401
rect 21822 8327 21878 8336
rect 21836 7886 21864 8327
rect 21916 8288 21968 8294
rect 21916 8230 21968 8236
rect 21456 7880 21508 7886
rect 21456 7822 21508 7828
rect 21824 7880 21876 7886
rect 21824 7822 21876 7828
rect 21088 7540 21140 7546
rect 21088 7482 21140 7488
rect 21100 6882 21128 7482
rect 21272 7336 21324 7342
rect 21272 7278 21324 7284
rect 21284 7002 21312 7278
rect 21928 7206 21956 8230
rect 22020 7274 22048 8434
rect 22112 7750 22140 9114
rect 22204 9042 22232 10134
rect 22296 10062 22324 11222
rect 22376 10804 22428 10810
rect 22376 10746 22428 10752
rect 22388 10538 22416 10746
rect 22376 10532 22428 10538
rect 22376 10474 22428 10480
rect 22572 10266 22600 13942
rect 22664 10985 22692 15286
rect 22928 14612 22980 14618
rect 22928 14554 22980 14560
rect 22940 13870 22968 14554
rect 23124 13870 23152 16662
rect 23216 16658 23244 17575
rect 23308 17134 23336 19858
rect 23572 19712 23624 19718
rect 23572 19654 23624 19660
rect 23480 19372 23532 19378
rect 23480 19314 23532 19320
rect 23492 18834 23520 19314
rect 23584 18873 23612 19654
rect 23676 19378 23704 20420
rect 23756 20402 23808 20408
rect 24400 20460 24452 20466
rect 24400 20402 24452 20408
rect 23940 20256 23992 20262
rect 23940 20198 23992 20204
rect 24398 20224 24454 20233
rect 23952 20058 23980 20198
rect 24398 20159 24454 20168
rect 23940 20052 23992 20058
rect 23940 19994 23992 20000
rect 24412 19990 24440 20159
rect 24504 19990 24532 20470
rect 24676 20324 24728 20330
rect 24676 20266 24728 20272
rect 24400 19984 24452 19990
rect 24400 19926 24452 19932
rect 24492 19984 24544 19990
rect 24492 19926 24544 19932
rect 24688 19922 24716 20266
rect 23848 19916 23900 19922
rect 23848 19858 23900 19864
rect 24676 19916 24728 19922
rect 24676 19858 24728 19864
rect 23756 19440 23808 19446
rect 23756 19382 23808 19388
rect 23664 19372 23716 19378
rect 23664 19314 23716 19320
rect 23570 18864 23626 18873
rect 23480 18828 23532 18834
rect 23570 18799 23626 18808
rect 23480 18770 23532 18776
rect 23572 18284 23624 18290
rect 23572 18226 23624 18232
rect 23386 17912 23442 17921
rect 23386 17847 23442 17856
rect 23296 17128 23348 17134
rect 23296 17070 23348 17076
rect 23204 16652 23256 16658
rect 23204 16594 23256 16600
rect 23400 16590 23428 17847
rect 23480 17740 23532 17746
rect 23480 17682 23532 17688
rect 23492 17066 23520 17682
rect 23480 17060 23532 17066
rect 23480 17002 23532 17008
rect 23296 16584 23348 16590
rect 23296 16526 23348 16532
rect 23388 16584 23440 16590
rect 23388 16526 23440 16532
rect 23204 16516 23256 16522
rect 23204 16458 23256 16464
rect 23216 14346 23244 16458
rect 23308 16114 23336 16526
rect 23296 16108 23348 16114
rect 23296 16050 23348 16056
rect 23584 15434 23612 18226
rect 23664 18216 23716 18222
rect 23664 18158 23716 18164
rect 23676 17542 23704 18158
rect 23768 17678 23796 19382
rect 23860 19310 23888 19858
rect 24780 19854 24808 21558
rect 24860 21548 24912 21554
rect 24860 21490 24912 21496
rect 24872 21350 24900 21490
rect 24860 21344 24912 21350
rect 24860 21286 24912 21292
rect 24858 21176 24914 21185
rect 24964 21146 24992 22374
rect 25056 21298 25084 26007
rect 25148 25498 25176 27424
rect 25136 25492 25188 25498
rect 25136 25434 25188 25440
rect 25240 25344 25268 34682
rect 25332 33590 25360 35022
rect 25424 34202 25452 36042
rect 25596 35760 25648 35766
rect 25594 35728 25596 35737
rect 25648 35728 25650 35737
rect 25594 35663 25650 35672
rect 25504 35624 25556 35630
rect 25596 35624 25648 35630
rect 25504 35566 25556 35572
rect 25594 35592 25596 35601
rect 25648 35592 25650 35601
rect 25516 35086 25544 35566
rect 25594 35527 25650 35536
rect 25504 35080 25556 35086
rect 25504 35022 25556 35028
rect 25412 34196 25464 34202
rect 25412 34138 25464 34144
rect 25608 33998 25636 35527
rect 25700 34950 25728 36246
rect 25688 34944 25740 34950
rect 25688 34886 25740 34892
rect 25596 33992 25648 33998
rect 25596 33934 25648 33940
rect 25412 33856 25464 33862
rect 25412 33798 25464 33804
rect 25320 33584 25372 33590
rect 25320 33526 25372 33532
rect 25424 33402 25452 33798
rect 25504 33584 25556 33590
rect 25504 33526 25556 33532
rect 25332 33386 25452 33402
rect 25320 33380 25452 33386
rect 25372 33374 25452 33380
rect 25320 33322 25372 33328
rect 25412 33312 25464 33318
rect 25410 33280 25412 33289
rect 25464 33280 25466 33289
rect 25410 33215 25466 33224
rect 25410 32056 25466 32065
rect 25410 31991 25466 32000
rect 25424 31958 25452 31991
rect 25412 31952 25464 31958
rect 25412 31894 25464 31900
rect 25320 31816 25372 31822
rect 25320 31758 25372 31764
rect 25332 30122 25360 31758
rect 25516 31754 25544 33526
rect 25424 31726 25544 31754
rect 25424 31346 25452 31726
rect 25596 31680 25648 31686
rect 25596 31622 25648 31628
rect 25504 31408 25556 31414
rect 25504 31350 25556 31356
rect 25412 31340 25464 31346
rect 25412 31282 25464 31288
rect 25424 31142 25452 31282
rect 25412 31136 25464 31142
rect 25412 31078 25464 31084
rect 25320 30116 25372 30122
rect 25320 30058 25372 30064
rect 25332 28626 25360 30058
rect 25412 29504 25464 29510
rect 25412 29446 25464 29452
rect 25320 28620 25372 28626
rect 25320 28562 25372 28568
rect 25318 26208 25374 26217
rect 25318 26143 25374 26152
rect 25332 26042 25360 26143
rect 25320 26036 25372 26042
rect 25320 25978 25372 25984
rect 25320 25900 25372 25906
rect 25320 25842 25372 25848
rect 25332 25809 25360 25842
rect 25318 25800 25374 25809
rect 25318 25735 25374 25744
rect 25320 25696 25372 25702
rect 25320 25638 25372 25644
rect 25332 25498 25360 25638
rect 25320 25492 25372 25498
rect 25320 25434 25372 25440
rect 25240 25316 25360 25344
rect 25332 24800 25360 25316
rect 25240 24772 25360 24800
rect 25136 23724 25188 23730
rect 25136 23666 25188 23672
rect 25148 23186 25176 23666
rect 25136 23180 25188 23186
rect 25136 23122 25188 23128
rect 25134 21992 25190 22001
rect 25134 21927 25136 21936
rect 25188 21927 25190 21936
rect 25136 21898 25188 21904
rect 25056 21270 25176 21298
rect 24858 21111 24914 21120
rect 24952 21140 25004 21146
rect 24872 20942 24900 21111
rect 24952 21082 25004 21088
rect 25148 21026 25176 21270
rect 25056 20998 25176 21026
rect 25240 21026 25268 24772
rect 25320 24200 25372 24206
rect 25320 24142 25372 24148
rect 25332 23798 25360 24142
rect 25320 23792 25372 23798
rect 25320 23734 25372 23740
rect 25424 22642 25452 29446
rect 25516 27606 25544 31350
rect 25608 31346 25636 31622
rect 25596 31340 25648 31346
rect 25596 31282 25648 31288
rect 25596 30184 25648 30190
rect 25596 30126 25648 30132
rect 25608 30025 25636 30126
rect 25594 30016 25650 30025
rect 25594 29951 25650 29960
rect 25596 29164 25648 29170
rect 25596 29106 25648 29112
rect 25608 28762 25636 29106
rect 25596 28756 25648 28762
rect 25596 28698 25648 28704
rect 25596 28620 25648 28626
rect 25596 28562 25648 28568
rect 25504 27600 25556 27606
rect 25504 27542 25556 27548
rect 25504 26444 25556 26450
rect 25608 26432 25636 28562
rect 25700 27520 25728 34886
rect 25792 30376 25820 37726
rect 25964 37664 26016 37670
rect 25964 37606 26016 37612
rect 25872 36032 25924 36038
rect 25872 35974 25924 35980
rect 25884 35698 25912 35974
rect 25872 35692 25924 35698
rect 25872 35634 25924 35640
rect 25870 35184 25926 35193
rect 25870 35119 25926 35128
rect 25884 35086 25912 35119
rect 25872 35080 25924 35086
rect 25872 35022 25924 35028
rect 25976 34950 26004 37606
rect 26160 36310 26188 37742
rect 26436 37466 26464 37810
rect 26424 37460 26476 37466
rect 26424 37402 26476 37408
rect 26528 37330 26556 38150
rect 27540 38010 27568 38218
rect 28540 38208 28592 38214
rect 28540 38150 28592 38156
rect 27528 38004 27580 38010
rect 27528 37946 27580 37952
rect 26608 37868 26660 37874
rect 26608 37810 26660 37816
rect 26620 37466 26648 37810
rect 27068 37800 27120 37806
rect 27068 37742 27120 37748
rect 27988 37800 28040 37806
rect 27988 37742 28040 37748
rect 26608 37460 26660 37466
rect 26608 37402 26660 37408
rect 26516 37324 26568 37330
rect 26516 37266 26568 37272
rect 26148 36304 26200 36310
rect 26148 36246 26200 36252
rect 26528 36174 26556 37266
rect 26332 36168 26384 36174
rect 26332 36110 26384 36116
rect 26516 36168 26568 36174
rect 26516 36110 26568 36116
rect 26056 35692 26108 35698
rect 26240 35692 26292 35698
rect 26056 35634 26108 35640
rect 26160 35652 26240 35680
rect 25964 34944 26016 34950
rect 25964 34886 26016 34892
rect 25976 34746 26004 34886
rect 25964 34740 26016 34746
rect 25964 34682 26016 34688
rect 25964 33992 26016 33998
rect 26068 33980 26096 35634
rect 26160 35494 26188 35652
rect 26240 35634 26292 35640
rect 26344 35578 26372 36110
rect 26882 35728 26938 35737
rect 26516 35692 26568 35698
rect 26882 35663 26938 35672
rect 26516 35634 26568 35640
rect 26252 35550 26372 35578
rect 26422 35592 26478 35601
rect 26148 35488 26200 35494
rect 26148 35430 26200 35436
rect 26252 33998 26280 35550
rect 26528 35578 26556 35634
rect 26478 35550 26556 35578
rect 26422 35527 26478 35536
rect 26896 35494 26924 35663
rect 26608 35488 26660 35494
rect 26608 35430 26660 35436
rect 26884 35488 26936 35494
rect 26884 35430 26936 35436
rect 26620 35154 26648 35430
rect 26608 35148 26660 35154
rect 26608 35090 26660 35096
rect 26332 35080 26384 35086
rect 26332 35022 26384 35028
rect 26424 35080 26476 35086
rect 26424 35022 26476 35028
rect 26016 33952 26096 33980
rect 26240 33992 26292 33998
rect 25964 33934 26016 33940
rect 26240 33934 26292 33940
rect 25976 32774 26004 33934
rect 26148 33924 26200 33930
rect 26148 33866 26200 33872
rect 26160 33658 26188 33866
rect 26148 33652 26200 33658
rect 26148 33594 26200 33600
rect 26056 32972 26108 32978
rect 26056 32914 26108 32920
rect 25964 32768 26016 32774
rect 25964 32710 26016 32716
rect 25964 31136 26016 31142
rect 25964 31078 26016 31084
rect 25976 30648 26004 31078
rect 26068 30870 26096 32914
rect 26252 32314 26280 33934
rect 26344 32774 26372 35022
rect 26332 32768 26384 32774
rect 26332 32710 26384 32716
rect 26160 32286 26280 32314
rect 26160 31822 26188 32286
rect 26240 32224 26292 32230
rect 26240 32166 26292 32172
rect 26252 31822 26280 32166
rect 26148 31816 26200 31822
rect 26148 31758 26200 31764
rect 26240 31816 26292 31822
rect 26240 31758 26292 31764
rect 26148 31680 26200 31686
rect 26148 31622 26200 31628
rect 26240 31680 26292 31686
rect 26240 31622 26292 31628
rect 26056 30864 26108 30870
rect 26056 30806 26108 30812
rect 26160 30734 26188 31622
rect 26148 30728 26200 30734
rect 26148 30670 26200 30676
rect 25976 30620 26096 30648
rect 25792 30348 26004 30376
rect 25870 30152 25926 30161
rect 25870 30087 25872 30096
rect 25924 30087 25926 30096
rect 25872 30058 25924 30064
rect 25778 29880 25834 29889
rect 25778 29815 25834 29824
rect 25792 29646 25820 29815
rect 25780 29640 25832 29646
rect 25780 29582 25832 29588
rect 25870 29064 25926 29073
rect 25870 28999 25926 29008
rect 25700 27492 25820 27520
rect 25688 27396 25740 27402
rect 25688 27338 25740 27344
rect 25556 26404 25636 26432
rect 25504 26386 25556 26392
rect 25516 25906 25544 26386
rect 25700 26382 25728 27338
rect 25688 26376 25740 26382
rect 25688 26318 25740 26324
rect 25688 26240 25740 26246
rect 25688 26182 25740 26188
rect 25700 25906 25728 26182
rect 25504 25900 25556 25906
rect 25504 25842 25556 25848
rect 25688 25900 25740 25906
rect 25688 25842 25740 25848
rect 25504 25696 25556 25702
rect 25504 25638 25556 25644
rect 25412 22636 25464 22642
rect 25412 22578 25464 22584
rect 25412 22432 25464 22438
rect 25318 22400 25374 22409
rect 25412 22374 25464 22380
rect 25318 22335 25374 22344
rect 25332 22098 25360 22335
rect 25320 22092 25372 22098
rect 25320 22034 25372 22040
rect 25320 21616 25372 21622
rect 25320 21558 25372 21564
rect 25332 21146 25360 21558
rect 25320 21140 25372 21146
rect 25320 21082 25372 21088
rect 25240 20998 25360 21026
rect 24860 20936 24912 20942
rect 24860 20878 24912 20884
rect 24860 20800 24912 20806
rect 24860 20742 24912 20748
rect 24872 20466 24900 20742
rect 24860 20460 24912 20466
rect 24860 20402 24912 20408
rect 24860 20256 24912 20262
rect 24860 20198 24912 20204
rect 24950 20224 25006 20233
rect 24768 19848 24820 19854
rect 24768 19790 24820 19796
rect 24676 19780 24728 19786
rect 24676 19722 24728 19728
rect 24492 19712 24544 19718
rect 24492 19654 24544 19660
rect 24504 19446 24532 19654
rect 24492 19440 24544 19446
rect 24492 19382 24544 19388
rect 24688 19334 24716 19722
rect 23848 19304 23900 19310
rect 24688 19306 24808 19334
rect 23848 19246 23900 19252
rect 24216 19168 24268 19174
rect 24216 19110 24268 19116
rect 23848 18148 23900 18154
rect 23848 18090 23900 18096
rect 23756 17672 23808 17678
rect 23756 17614 23808 17620
rect 23664 17536 23716 17542
rect 23664 17478 23716 17484
rect 23768 16640 23796 17614
rect 23860 16658 23888 18090
rect 23676 16612 23796 16640
rect 23848 16652 23900 16658
rect 23572 15428 23624 15434
rect 23572 15370 23624 15376
rect 23296 14952 23348 14958
rect 23296 14894 23348 14900
rect 23308 14482 23336 14894
rect 23296 14476 23348 14482
rect 23296 14418 23348 14424
rect 23204 14340 23256 14346
rect 23204 14282 23256 14288
rect 23216 13870 23244 14282
rect 22928 13864 22980 13870
rect 22848 13824 22928 13852
rect 22744 13796 22796 13802
rect 22744 13738 22796 13744
rect 22756 13462 22784 13738
rect 22744 13456 22796 13462
rect 22744 13398 22796 13404
rect 22744 13184 22796 13190
rect 22744 13126 22796 13132
rect 22756 12986 22784 13126
rect 22744 12980 22796 12986
rect 22744 12922 22796 12928
rect 22848 12434 22876 13824
rect 23112 13864 23164 13870
rect 22928 13806 22980 13812
rect 23032 13824 23112 13852
rect 22928 13184 22980 13190
rect 22928 13126 22980 13132
rect 22756 12406 22876 12434
rect 22650 10976 22706 10985
rect 22650 10911 22706 10920
rect 22756 10674 22784 12406
rect 22836 12368 22888 12374
rect 22836 12310 22888 12316
rect 22848 10742 22876 12310
rect 22836 10736 22888 10742
rect 22836 10678 22888 10684
rect 22940 10674 22968 13126
rect 23032 12306 23060 13824
rect 23112 13806 23164 13812
rect 23204 13864 23256 13870
rect 23308 13852 23336 14418
rect 23388 13864 23440 13870
rect 23308 13824 23388 13852
rect 23204 13806 23256 13812
rect 23388 13806 23440 13812
rect 23112 13728 23164 13734
rect 23112 13670 23164 13676
rect 23124 13462 23152 13670
rect 23112 13456 23164 13462
rect 23112 13398 23164 13404
rect 23124 13190 23152 13398
rect 23204 13320 23256 13326
rect 23204 13262 23256 13268
rect 23112 13184 23164 13190
rect 23112 13126 23164 13132
rect 23112 12912 23164 12918
rect 23112 12854 23164 12860
rect 23020 12300 23072 12306
rect 23020 12242 23072 12248
rect 23032 10724 23060 12242
rect 23124 12186 23152 12854
rect 23216 12782 23244 13262
rect 23204 12776 23256 12782
rect 23204 12718 23256 12724
rect 23216 12306 23244 12718
rect 23204 12300 23256 12306
rect 23204 12242 23256 12248
rect 23124 12158 23244 12186
rect 23112 10736 23164 10742
rect 23032 10713 23112 10724
rect 23018 10704 23112 10713
rect 22652 10668 22704 10674
rect 22652 10610 22704 10616
rect 22744 10668 22796 10674
rect 22744 10610 22796 10616
rect 22928 10668 22980 10674
rect 23074 10696 23112 10704
rect 23112 10678 23164 10684
rect 23018 10639 23074 10648
rect 22928 10610 22980 10616
rect 22664 10266 22692 10610
rect 22744 10464 22796 10470
rect 22744 10406 22796 10412
rect 22756 10266 22784 10406
rect 22376 10260 22428 10266
rect 22376 10202 22428 10208
rect 22560 10260 22612 10266
rect 22560 10202 22612 10208
rect 22652 10260 22704 10266
rect 22652 10202 22704 10208
rect 22744 10260 22796 10266
rect 22744 10202 22796 10208
rect 22284 10056 22336 10062
rect 22284 9998 22336 10004
rect 22388 9722 22416 10202
rect 22376 9716 22428 9722
rect 22376 9658 22428 9664
rect 22282 9616 22338 9625
rect 22940 9586 22968 10610
rect 23112 10600 23164 10606
rect 23112 10542 23164 10548
rect 22282 9551 22338 9560
rect 22744 9580 22796 9586
rect 22296 9110 22324 9551
rect 22744 9522 22796 9528
rect 22928 9580 22980 9586
rect 22928 9522 22980 9528
rect 22756 9217 22784 9522
rect 22742 9208 22798 9217
rect 22572 9166 22742 9194
rect 22284 9104 22336 9110
rect 22284 9046 22336 9052
rect 22192 9036 22244 9042
rect 22192 8978 22244 8984
rect 22572 8974 22600 9166
rect 22742 9143 22798 9152
rect 22940 9110 22968 9522
rect 23124 9466 23152 10542
rect 23032 9450 23152 9466
rect 23020 9444 23152 9450
rect 23072 9438 23152 9444
rect 23020 9386 23072 9392
rect 22744 9104 22796 9110
rect 22650 9072 22706 9081
rect 22744 9046 22796 9052
rect 22928 9104 22980 9110
rect 22928 9046 22980 9052
rect 22650 9007 22706 9016
rect 22376 8968 22428 8974
rect 22376 8910 22428 8916
rect 22560 8968 22612 8974
rect 22560 8910 22612 8916
rect 22284 8900 22336 8906
rect 22284 8842 22336 8848
rect 22296 7954 22324 8842
rect 22388 8634 22416 8910
rect 22376 8628 22428 8634
rect 22376 8570 22428 8576
rect 22376 8288 22428 8294
rect 22664 8276 22692 9007
rect 22376 8230 22428 8236
rect 22572 8248 22692 8276
rect 22388 7954 22416 8230
rect 22284 7948 22336 7954
rect 22284 7890 22336 7896
rect 22376 7948 22428 7954
rect 22376 7890 22428 7896
rect 22376 7812 22428 7818
rect 22376 7754 22428 7760
rect 22100 7744 22152 7750
rect 22100 7686 22152 7692
rect 22284 7744 22336 7750
rect 22284 7686 22336 7692
rect 22296 7546 22324 7686
rect 22388 7546 22416 7754
rect 22468 7744 22520 7750
rect 22468 7686 22520 7692
rect 22284 7540 22336 7546
rect 22284 7482 22336 7488
rect 22376 7540 22428 7546
rect 22376 7482 22428 7488
rect 22480 7426 22508 7686
rect 22204 7410 22508 7426
rect 22100 7404 22152 7410
rect 22100 7346 22152 7352
rect 22192 7404 22508 7410
rect 22244 7398 22508 7404
rect 22192 7346 22244 7352
rect 22008 7268 22060 7274
rect 22008 7210 22060 7216
rect 21364 7200 21416 7206
rect 21364 7142 21416 7148
rect 21916 7200 21968 7206
rect 21916 7142 21968 7148
rect 21272 6996 21324 7002
rect 21272 6938 21324 6944
rect 21100 6854 21312 6882
rect 21284 6798 21312 6854
rect 21376 6798 21404 7142
rect 21272 6792 21324 6798
rect 21272 6734 21324 6740
rect 21364 6792 21416 6798
rect 21364 6734 21416 6740
rect 22112 6730 22140 7346
rect 22100 6724 22152 6730
rect 22100 6666 22152 6672
rect 22376 6656 22428 6662
rect 22376 6598 22428 6604
rect 20996 5568 21048 5574
rect 20996 5510 21048 5516
rect 21008 5302 21036 5510
rect 20996 5296 21048 5302
rect 20996 5238 21048 5244
rect 20904 5228 20956 5234
rect 20904 5170 20956 5176
rect 20916 4826 20944 5170
rect 20904 4820 20956 4826
rect 20904 4762 20956 4768
rect 20812 4616 20864 4622
rect 20812 4558 20864 4564
rect 20076 4548 20128 4554
rect 20076 4490 20128 4496
rect 20536 4548 20588 4554
rect 20536 4490 20588 4496
rect 21008 4282 21036 5238
rect 22388 5166 22416 6598
rect 22572 5914 22600 8248
rect 22756 8022 22784 9046
rect 23032 8974 23060 9386
rect 23112 9104 23164 9110
rect 23112 9046 23164 9052
rect 23020 8968 23072 8974
rect 23020 8910 23072 8916
rect 23124 8820 23152 9046
rect 22848 8792 23152 8820
rect 22652 8016 22704 8022
rect 22652 7958 22704 7964
rect 22744 8016 22796 8022
rect 22744 7958 22796 7964
rect 22664 7886 22692 7958
rect 22652 7880 22704 7886
rect 22652 7822 22704 7828
rect 22664 6322 22692 7822
rect 22744 7812 22796 7818
rect 22744 7754 22796 7760
rect 22756 6458 22784 7754
rect 22848 7460 22876 8792
rect 23020 8288 23072 8294
rect 23020 8230 23072 8236
rect 23032 7954 23060 8230
rect 23020 7948 23072 7954
rect 23020 7890 23072 7896
rect 23112 7812 23164 7818
rect 23112 7754 23164 7760
rect 23124 7546 23152 7754
rect 23216 7750 23244 12158
rect 23480 11756 23532 11762
rect 23480 11698 23532 11704
rect 23388 11552 23440 11558
rect 23388 11494 23440 11500
rect 23400 11354 23428 11494
rect 23492 11354 23520 11698
rect 23584 11694 23612 15370
rect 23676 14890 23704 16612
rect 23848 16594 23900 16600
rect 23756 16516 23808 16522
rect 23756 16458 23808 16464
rect 23768 16017 23796 16458
rect 23754 16008 23810 16017
rect 23754 15943 23810 15952
rect 24032 15904 24084 15910
rect 24032 15846 24084 15852
rect 23664 14884 23716 14890
rect 23664 14826 23716 14832
rect 23940 14544 23992 14550
rect 23940 14486 23992 14492
rect 23848 14272 23900 14278
rect 23848 14214 23900 14220
rect 23664 13864 23716 13870
rect 23664 13806 23716 13812
rect 23572 11688 23624 11694
rect 23572 11630 23624 11636
rect 23388 11348 23440 11354
rect 23388 11290 23440 11296
rect 23480 11348 23532 11354
rect 23480 11290 23532 11296
rect 23584 11286 23612 11630
rect 23572 11280 23624 11286
rect 23572 11222 23624 11228
rect 23388 11144 23440 11150
rect 23440 11104 23520 11132
rect 23388 11086 23440 11092
rect 23388 11008 23440 11014
rect 23388 10950 23440 10956
rect 23400 10742 23428 10950
rect 23388 10736 23440 10742
rect 23388 10678 23440 10684
rect 23400 9586 23428 10678
rect 23492 10470 23520 11104
rect 23676 10606 23704 13806
rect 23756 12640 23808 12646
rect 23756 12582 23808 12588
rect 23768 11762 23796 12582
rect 23756 11756 23808 11762
rect 23756 11698 23808 11704
rect 23664 10600 23716 10606
rect 23664 10542 23716 10548
rect 23572 10532 23624 10538
rect 23572 10474 23624 10480
rect 23480 10464 23532 10470
rect 23480 10406 23532 10412
rect 23388 9580 23440 9586
rect 23388 9522 23440 9528
rect 23296 9512 23348 9518
rect 23296 9454 23348 9460
rect 23308 8906 23336 9454
rect 23400 8974 23428 9522
rect 23584 9110 23612 10474
rect 23768 9994 23796 11698
rect 23860 10470 23888 14214
rect 23848 10464 23900 10470
rect 23848 10406 23900 10412
rect 23952 10146 23980 14486
rect 23860 10118 23980 10146
rect 23756 9988 23808 9994
rect 23756 9930 23808 9936
rect 23572 9104 23624 9110
rect 23572 9046 23624 9052
rect 23388 8968 23440 8974
rect 23388 8910 23440 8916
rect 23296 8900 23348 8906
rect 23296 8842 23348 8848
rect 23204 7744 23256 7750
rect 23204 7686 23256 7692
rect 23112 7540 23164 7546
rect 23112 7482 23164 7488
rect 22928 7472 22980 7478
rect 22848 7432 22928 7460
rect 22928 7414 22980 7420
rect 22744 6452 22796 6458
rect 22744 6394 22796 6400
rect 22940 6390 22968 7414
rect 23216 7002 23244 7686
rect 23308 7274 23336 8842
rect 23572 8832 23624 8838
rect 23572 8774 23624 8780
rect 23584 8634 23612 8774
rect 23572 8628 23624 8634
rect 23572 8570 23624 8576
rect 23572 8492 23624 8498
rect 23572 8434 23624 8440
rect 23478 8392 23534 8401
rect 23478 8327 23534 8336
rect 23296 7268 23348 7274
rect 23296 7210 23348 7216
rect 23204 6996 23256 7002
rect 23204 6938 23256 6944
rect 23492 6390 23520 8327
rect 23584 8090 23612 8434
rect 23572 8084 23624 8090
rect 23572 8026 23624 8032
rect 23584 7410 23612 8026
rect 23572 7404 23624 7410
rect 23572 7346 23624 7352
rect 23860 7002 23888 10118
rect 23940 10056 23992 10062
rect 23940 9998 23992 10004
rect 23952 9722 23980 9998
rect 24044 9722 24072 15846
rect 24228 15094 24256 19110
rect 24676 18692 24728 18698
rect 24676 18634 24728 18640
rect 24688 17746 24716 18634
rect 24676 17740 24728 17746
rect 24676 17682 24728 17688
rect 24688 17513 24716 17682
rect 24780 17678 24808 19306
rect 24872 18601 24900 20198
rect 24950 20159 25006 20168
rect 24964 19990 24992 20159
rect 24952 19984 25004 19990
rect 24952 19926 25004 19932
rect 24858 18592 24914 18601
rect 24858 18527 24914 18536
rect 25056 18290 25084 20998
rect 25226 20632 25282 20641
rect 25226 20567 25282 20576
rect 25240 20466 25268 20567
rect 25332 20466 25360 20998
rect 25228 20460 25280 20466
rect 25148 20420 25228 20448
rect 25148 19854 25176 20420
rect 25228 20402 25280 20408
rect 25320 20460 25372 20466
rect 25320 20402 25372 20408
rect 25320 20324 25372 20330
rect 25320 20266 25372 20272
rect 25332 19904 25360 20266
rect 25240 19876 25360 19904
rect 25136 19848 25188 19854
rect 25136 19790 25188 19796
rect 25240 19786 25268 19876
rect 25318 19816 25374 19825
rect 25228 19780 25280 19786
rect 25318 19751 25320 19760
rect 25228 19722 25280 19728
rect 25372 19751 25374 19760
rect 25320 19722 25372 19728
rect 25136 19508 25188 19514
rect 25136 19450 25188 19456
rect 25148 18630 25176 19450
rect 25136 18624 25188 18630
rect 25136 18566 25188 18572
rect 25240 18358 25268 19722
rect 25228 18352 25280 18358
rect 25228 18294 25280 18300
rect 24952 18284 25004 18290
rect 24952 18226 25004 18232
rect 25044 18284 25096 18290
rect 25044 18226 25096 18232
rect 24768 17672 24820 17678
rect 24768 17614 24820 17620
rect 24674 17504 24730 17513
rect 24674 17439 24730 17448
rect 24490 16552 24546 16561
rect 24490 16487 24546 16496
rect 24504 16153 24532 16487
rect 24490 16144 24546 16153
rect 24490 16079 24546 16088
rect 24676 16108 24728 16114
rect 24504 15706 24532 16079
rect 24676 16050 24728 16056
rect 24492 15700 24544 15706
rect 24492 15642 24544 15648
rect 24504 15502 24532 15642
rect 24688 15502 24716 16050
rect 24492 15496 24544 15502
rect 24492 15438 24544 15444
rect 24676 15496 24728 15502
rect 24676 15438 24728 15444
rect 24688 15366 24716 15438
rect 24676 15360 24728 15366
rect 24676 15302 24728 15308
rect 24216 15088 24268 15094
rect 24216 15030 24268 15036
rect 24124 14408 24176 14414
rect 24124 14350 24176 14356
rect 24492 14408 24544 14414
rect 24492 14350 24544 14356
rect 24136 13938 24164 14350
rect 24398 13968 24454 13977
rect 24124 13932 24176 13938
rect 24124 13874 24176 13880
rect 24320 13926 24398 13954
rect 24136 13326 24164 13874
rect 24320 13870 24348 13926
rect 24504 13938 24532 14350
rect 24398 13903 24454 13912
rect 24492 13932 24544 13938
rect 24492 13874 24544 13880
rect 24308 13864 24360 13870
rect 24308 13806 24360 13812
rect 24216 13796 24268 13802
rect 24216 13738 24268 13744
rect 24124 13320 24176 13326
rect 24124 13262 24176 13268
rect 24228 13138 24256 13738
rect 24136 13110 24256 13138
rect 24136 12073 24164 13110
rect 24320 12850 24348 13806
rect 24398 13424 24454 13433
rect 24398 13359 24454 13368
rect 24412 12918 24440 13359
rect 24492 13252 24544 13258
rect 24544 13212 24624 13240
rect 24492 13194 24544 13200
rect 24400 12912 24452 12918
rect 24400 12854 24452 12860
rect 24308 12844 24360 12850
rect 24308 12786 24360 12792
rect 24216 12436 24268 12442
rect 24216 12378 24268 12384
rect 24122 12064 24178 12073
rect 24122 11999 24178 12008
rect 23940 9716 23992 9722
rect 23940 9658 23992 9664
rect 24032 9716 24084 9722
rect 24032 9658 24084 9664
rect 24136 8480 24164 11999
rect 24228 11898 24256 12378
rect 24216 11892 24268 11898
rect 24216 11834 24268 11840
rect 24216 11756 24268 11762
rect 24320 11744 24348 12786
rect 24400 12776 24452 12782
rect 24400 12718 24452 12724
rect 24492 12776 24544 12782
rect 24492 12718 24544 12724
rect 24412 12442 24440 12718
rect 24400 12436 24452 12442
rect 24400 12378 24452 12384
rect 24268 11716 24348 11744
rect 24216 11698 24268 11704
rect 24320 11150 24348 11716
rect 24400 11756 24452 11762
rect 24504 11744 24532 12718
rect 24596 11762 24624 13212
rect 24688 12288 24716 15302
rect 24780 14890 24808 17614
rect 24860 16652 24912 16658
rect 24860 16594 24912 16600
rect 24872 16114 24900 16594
rect 24964 16454 24992 18226
rect 25228 16584 25280 16590
rect 25228 16526 25280 16532
rect 24952 16448 25004 16454
rect 24952 16390 25004 16396
rect 25136 16448 25188 16454
rect 25136 16390 25188 16396
rect 25148 16182 25176 16390
rect 25136 16176 25188 16182
rect 25136 16118 25188 16124
rect 24860 16108 24912 16114
rect 24860 16050 24912 16056
rect 25044 15904 25096 15910
rect 25044 15846 25096 15852
rect 24768 14884 24820 14890
rect 24768 14826 24820 14832
rect 25056 13938 25084 15846
rect 25148 15473 25176 16118
rect 25240 15978 25268 16526
rect 25228 15972 25280 15978
rect 25228 15914 25280 15920
rect 25240 15502 25268 15914
rect 25228 15496 25280 15502
rect 25134 15464 25190 15473
rect 25228 15438 25280 15444
rect 25134 15399 25190 15408
rect 25320 15428 25372 15434
rect 25320 15370 25372 15376
rect 24768 13932 24820 13938
rect 24768 13874 24820 13880
rect 25044 13932 25096 13938
rect 25044 13874 25096 13880
rect 24780 12714 24808 13874
rect 25044 13796 25096 13802
rect 25044 13738 25096 13744
rect 24860 13184 24912 13190
rect 24860 13126 24912 13132
rect 24872 12782 24900 13126
rect 24860 12776 24912 12782
rect 24860 12718 24912 12724
rect 24768 12708 24820 12714
rect 24768 12650 24820 12656
rect 24768 12300 24820 12306
rect 24688 12260 24768 12288
rect 24768 12242 24820 12248
rect 24780 11762 24808 12242
rect 25056 12238 25084 13738
rect 25228 12776 25280 12782
rect 25228 12718 25280 12724
rect 25136 12640 25188 12646
rect 25136 12582 25188 12588
rect 25148 12442 25176 12582
rect 25240 12442 25268 12718
rect 25136 12436 25188 12442
rect 25136 12378 25188 12384
rect 25228 12436 25280 12442
rect 25228 12378 25280 12384
rect 25044 12232 25096 12238
rect 25044 12174 25096 12180
rect 25056 11762 25084 12174
rect 25332 11830 25360 15370
rect 25424 12434 25452 22374
rect 25516 21690 25544 25638
rect 25688 24608 25740 24614
rect 25688 24550 25740 24556
rect 25700 24410 25728 24550
rect 25688 24404 25740 24410
rect 25688 24346 25740 24352
rect 25688 23112 25740 23118
rect 25792 23100 25820 27492
rect 25884 26042 25912 28999
rect 25872 26036 25924 26042
rect 25872 25978 25924 25984
rect 25976 24698 26004 30348
rect 26068 29646 26096 30620
rect 26148 30252 26200 30258
rect 26252 30240 26280 31622
rect 26332 31340 26384 31346
rect 26332 31282 26384 31288
rect 26344 31142 26372 31282
rect 26436 31260 26464 35022
rect 26792 34196 26844 34202
rect 26792 34138 26844 34144
rect 26516 33924 26568 33930
rect 26516 33866 26568 33872
rect 26528 33522 26556 33866
rect 26516 33516 26568 33522
rect 26516 33458 26568 33464
rect 26608 33516 26660 33522
rect 26608 33458 26660 33464
rect 26620 33114 26648 33458
rect 26608 33108 26660 33114
rect 26608 33050 26660 33056
rect 26700 32768 26752 32774
rect 26700 32710 26752 32716
rect 26516 32360 26568 32366
rect 26516 32302 26568 32308
rect 26528 31822 26556 32302
rect 26712 31929 26740 32710
rect 26698 31920 26754 31929
rect 26698 31855 26754 31864
rect 26516 31816 26568 31822
rect 26516 31758 26568 31764
rect 26804 31754 26832 34138
rect 26976 33992 27028 33998
rect 26976 33934 27028 33940
rect 26988 32026 27016 33934
rect 26976 32020 27028 32026
rect 26976 31962 27028 31968
rect 26988 31822 27016 31962
rect 26976 31816 27028 31822
rect 26976 31758 27028 31764
rect 26792 31748 26844 31754
rect 26792 31690 26844 31696
rect 26516 31272 26568 31278
rect 26436 31232 26516 31260
rect 26516 31214 26568 31220
rect 26332 31136 26384 31142
rect 26332 31078 26384 31084
rect 26424 30728 26476 30734
rect 26424 30670 26476 30676
rect 26200 30212 26280 30240
rect 26148 30194 26200 30200
rect 26056 29640 26108 29646
rect 26056 29582 26108 29588
rect 26160 28490 26188 30194
rect 26240 30048 26292 30054
rect 26240 29990 26292 29996
rect 26252 29730 26280 29990
rect 26252 29714 26372 29730
rect 26252 29708 26384 29714
rect 26252 29702 26332 29708
rect 26332 29650 26384 29656
rect 26436 29646 26464 30670
rect 26528 29782 26556 31214
rect 26700 31204 26752 31210
rect 26700 31146 26752 31152
rect 26608 31136 26660 31142
rect 26608 31078 26660 31084
rect 26620 30274 26648 31078
rect 26712 30433 26740 31146
rect 26792 31136 26844 31142
rect 26792 31078 26844 31084
rect 26804 30870 26832 31078
rect 26792 30864 26844 30870
rect 26792 30806 26844 30812
rect 26698 30424 26754 30433
rect 26698 30359 26754 30368
rect 26620 30246 26740 30274
rect 26608 30048 26660 30054
rect 26608 29990 26660 29996
rect 26620 29889 26648 29990
rect 26606 29880 26662 29889
rect 26606 29815 26662 29824
rect 26516 29776 26568 29782
rect 26516 29718 26568 29724
rect 26608 29776 26660 29782
rect 26608 29718 26660 29724
rect 26424 29640 26476 29646
rect 26424 29582 26476 29588
rect 26332 29572 26384 29578
rect 26252 29532 26332 29560
rect 26252 29170 26280 29532
rect 26332 29514 26384 29520
rect 26436 29306 26464 29582
rect 26528 29306 26556 29718
rect 26424 29300 26476 29306
rect 26424 29242 26476 29248
rect 26516 29300 26568 29306
rect 26516 29242 26568 29248
rect 26240 29164 26292 29170
rect 26240 29106 26292 29112
rect 26516 29164 26568 29170
rect 26516 29106 26568 29112
rect 26252 29073 26280 29106
rect 26238 29064 26294 29073
rect 26528 29034 26556 29106
rect 26238 28999 26294 29008
rect 26516 29028 26568 29034
rect 26516 28970 26568 28976
rect 26148 28484 26200 28490
rect 26148 28426 26200 28432
rect 26160 26314 26188 28426
rect 26620 27674 26648 29718
rect 26712 28121 26740 30246
rect 26882 30016 26938 30025
rect 26882 29951 26938 29960
rect 26896 29782 26924 29951
rect 26884 29776 26936 29782
rect 26884 29718 26936 29724
rect 27080 29034 27108 37742
rect 28000 37369 28028 37742
rect 27986 37360 28042 37369
rect 27986 37295 28042 37304
rect 27344 37256 27396 37262
rect 27344 37198 27396 37204
rect 27356 36174 27384 37198
rect 27896 37188 27948 37194
rect 27896 37130 27948 37136
rect 27528 37120 27580 37126
rect 27528 37062 27580 37068
rect 27436 36576 27488 36582
rect 27436 36518 27488 36524
rect 27160 36168 27212 36174
rect 27160 36110 27212 36116
rect 27252 36168 27304 36174
rect 27252 36110 27304 36116
rect 27344 36168 27396 36174
rect 27344 36110 27396 36116
rect 27172 34542 27200 36110
rect 27160 34536 27212 34542
rect 27160 34478 27212 34484
rect 27264 34406 27292 36110
rect 27356 35698 27384 36110
rect 27344 35692 27396 35698
rect 27344 35634 27396 35640
rect 27448 35630 27476 36518
rect 27436 35624 27488 35630
rect 27436 35566 27488 35572
rect 27540 35018 27568 37062
rect 27804 36916 27856 36922
rect 27804 36858 27856 36864
rect 27712 36780 27764 36786
rect 27712 36722 27764 36728
rect 27528 35012 27580 35018
rect 27528 34954 27580 34960
rect 27344 34944 27396 34950
rect 27344 34886 27396 34892
rect 27252 34400 27304 34406
rect 27252 34342 27304 34348
rect 27160 33856 27212 33862
rect 27160 33798 27212 33804
rect 27172 33590 27200 33798
rect 27160 33584 27212 33590
rect 27160 33526 27212 33532
rect 27252 32972 27304 32978
rect 27252 32914 27304 32920
rect 27160 31340 27212 31346
rect 27160 31282 27212 31288
rect 27172 30938 27200 31282
rect 27160 30932 27212 30938
rect 27160 30874 27212 30880
rect 27264 30734 27292 32914
rect 27356 32774 27384 34886
rect 27528 32904 27580 32910
rect 27528 32846 27580 32852
rect 27344 32768 27396 32774
rect 27344 32710 27396 32716
rect 27252 30728 27304 30734
rect 27252 30670 27304 30676
rect 27356 30580 27384 32710
rect 27540 32570 27568 32846
rect 27528 32564 27580 32570
rect 27528 32506 27580 32512
rect 27724 32502 27752 36722
rect 27816 35834 27844 36858
rect 27804 35828 27856 35834
rect 27804 35770 27856 35776
rect 27816 34950 27844 35770
rect 27804 34944 27856 34950
rect 27804 34886 27856 34892
rect 27804 33448 27856 33454
rect 27804 33390 27856 33396
rect 27816 32978 27844 33390
rect 27804 32972 27856 32978
rect 27804 32914 27856 32920
rect 27712 32496 27764 32502
rect 27712 32438 27764 32444
rect 27724 31754 27752 32438
rect 27908 32298 27936 37130
rect 28172 36780 28224 36786
rect 28172 36722 28224 36728
rect 28264 36780 28316 36786
rect 28264 36722 28316 36728
rect 28184 36258 28212 36722
rect 28276 36378 28304 36722
rect 28448 36576 28500 36582
rect 28448 36518 28500 36524
rect 28264 36372 28316 36378
rect 28264 36314 28316 36320
rect 28184 36230 28304 36258
rect 27988 36168 28040 36174
rect 27988 36110 28040 36116
rect 28000 35290 28028 36110
rect 28276 35630 28304 36230
rect 28460 36009 28488 36518
rect 28552 36174 28580 38150
rect 29000 37868 29052 37874
rect 29000 37810 29052 37816
rect 28632 37324 28684 37330
rect 28632 37266 28684 37272
rect 28908 37324 28960 37330
rect 28908 37266 28960 37272
rect 28644 36582 28672 37266
rect 28632 36576 28684 36582
rect 28632 36518 28684 36524
rect 28540 36168 28592 36174
rect 28540 36110 28592 36116
rect 28446 36000 28502 36009
rect 28446 35935 28502 35944
rect 28172 35624 28224 35630
rect 28172 35566 28224 35572
rect 28264 35624 28316 35630
rect 28264 35566 28316 35572
rect 27988 35284 28040 35290
rect 27988 35226 28040 35232
rect 28000 34474 28028 35226
rect 28184 35222 28212 35566
rect 28172 35216 28224 35222
rect 28172 35158 28224 35164
rect 28276 34610 28304 35566
rect 28356 35216 28408 35222
rect 28354 35184 28356 35193
rect 28408 35184 28410 35193
rect 28354 35119 28410 35128
rect 28552 34678 28580 36110
rect 28540 34672 28592 34678
rect 28540 34614 28592 34620
rect 28264 34604 28316 34610
rect 28264 34546 28316 34552
rect 27988 34468 28040 34474
rect 27988 34410 28040 34416
rect 28080 34400 28132 34406
rect 28080 34342 28132 34348
rect 28092 34202 28120 34342
rect 28080 34196 28132 34202
rect 28080 34138 28132 34144
rect 28552 33590 28580 34614
rect 28644 34066 28672 36518
rect 28724 36236 28776 36242
rect 28724 36178 28776 36184
rect 28736 35766 28764 36178
rect 28816 36168 28868 36174
rect 28814 36136 28816 36145
rect 28868 36136 28870 36145
rect 28814 36071 28870 36080
rect 28724 35760 28776 35766
rect 28724 35702 28776 35708
rect 28632 34060 28684 34066
rect 28632 34002 28684 34008
rect 28540 33584 28592 33590
rect 28540 33526 28592 33532
rect 28540 33312 28592 33318
rect 28540 33254 28592 33260
rect 28552 32842 28580 33254
rect 28080 32836 28132 32842
rect 28080 32778 28132 32784
rect 28540 32836 28592 32842
rect 28540 32778 28592 32784
rect 28092 32570 28120 32778
rect 28080 32564 28132 32570
rect 28080 32506 28132 32512
rect 28448 32360 28500 32366
rect 28448 32302 28500 32308
rect 27896 32292 27948 32298
rect 27896 32234 27948 32240
rect 27632 31726 27752 31754
rect 27632 31414 27660 31726
rect 27712 31680 27764 31686
rect 27712 31622 27764 31628
rect 27620 31408 27672 31414
rect 27620 31350 27672 31356
rect 27528 31340 27580 31346
rect 27528 31282 27580 31288
rect 27436 30728 27488 30734
rect 27436 30670 27488 30676
rect 27172 30552 27384 30580
rect 27068 29028 27120 29034
rect 27068 28970 27120 28976
rect 26976 28960 27028 28966
rect 26976 28902 27028 28908
rect 26698 28112 26754 28121
rect 26754 28070 26924 28098
rect 26698 28047 26754 28056
rect 26608 27668 26660 27674
rect 26608 27610 26660 27616
rect 26700 27668 26752 27674
rect 26700 27610 26752 27616
rect 26424 27532 26476 27538
rect 26424 27474 26476 27480
rect 26332 27396 26384 27402
rect 26332 27338 26384 27344
rect 26344 27130 26372 27338
rect 26332 27124 26384 27130
rect 26332 27066 26384 27072
rect 26436 27062 26464 27474
rect 26424 27056 26476 27062
rect 26424 26998 26476 27004
rect 26514 27024 26570 27033
rect 26238 26752 26294 26761
rect 26294 26710 26372 26738
rect 26238 26687 26294 26696
rect 26344 26382 26372 26710
rect 26332 26376 26384 26382
rect 26332 26318 26384 26324
rect 26148 26308 26200 26314
rect 26148 26250 26200 26256
rect 26240 26308 26292 26314
rect 26240 26250 26292 26256
rect 26056 26240 26108 26246
rect 26056 26182 26108 26188
rect 26068 25906 26096 26182
rect 26148 26036 26200 26042
rect 26148 25978 26200 25984
rect 26160 25945 26188 25978
rect 26146 25936 26202 25945
rect 26056 25900 26108 25906
rect 26146 25871 26202 25880
rect 26056 25842 26108 25848
rect 26054 25392 26110 25401
rect 26252 25378 26280 26250
rect 26436 25838 26464 26998
rect 26514 26959 26570 26968
rect 26528 25906 26556 26959
rect 26620 26382 26648 27610
rect 26712 26994 26740 27610
rect 26792 27396 26844 27402
rect 26792 27338 26844 27344
rect 26700 26988 26752 26994
rect 26700 26930 26752 26936
rect 26804 26518 26832 27338
rect 26792 26512 26844 26518
rect 26792 26454 26844 26460
rect 26608 26376 26660 26382
rect 26608 26318 26660 26324
rect 26698 26344 26754 26353
rect 26698 26279 26754 26288
rect 26516 25900 26568 25906
rect 26516 25842 26568 25848
rect 26424 25832 26476 25838
rect 26424 25774 26476 25780
rect 26332 25764 26384 25770
rect 26332 25706 26384 25712
rect 26110 25350 26280 25378
rect 26054 25327 26110 25336
rect 25740 23072 25820 23100
rect 25884 24670 26004 24698
rect 25688 23054 25740 23060
rect 25884 22778 25912 24670
rect 25964 24608 26016 24614
rect 25964 24550 26016 24556
rect 25976 24274 26004 24550
rect 26344 24410 26372 25706
rect 26436 25294 26464 25774
rect 26608 25696 26660 25702
rect 26608 25638 26660 25644
rect 26424 25288 26476 25294
rect 26424 25230 26476 25236
rect 26332 24404 26384 24410
rect 26332 24346 26384 24352
rect 25964 24268 26016 24274
rect 25964 24210 26016 24216
rect 26424 24268 26476 24274
rect 26424 24210 26476 24216
rect 26056 23724 26108 23730
rect 26056 23666 26108 23672
rect 26068 23322 26096 23666
rect 26056 23316 26108 23322
rect 26056 23258 26108 23264
rect 26332 23316 26384 23322
rect 26332 23258 26384 23264
rect 26148 23112 26200 23118
rect 25962 23080 26018 23089
rect 26148 23054 26200 23060
rect 25962 23015 25964 23024
rect 26016 23015 26018 23024
rect 25964 22986 26016 22992
rect 26056 22976 26108 22982
rect 26056 22918 26108 22924
rect 25872 22772 25924 22778
rect 25872 22714 25924 22720
rect 25594 22672 25650 22681
rect 25650 22630 25728 22658
rect 25594 22607 25650 22616
rect 25700 21690 25728 22630
rect 25780 22568 25832 22574
rect 25780 22510 25832 22516
rect 25792 22032 25820 22510
rect 25780 22026 25832 22032
rect 25780 21968 25832 21974
rect 26068 21894 26096 22918
rect 26160 22574 26188 23054
rect 26240 22976 26292 22982
rect 26240 22918 26292 22924
rect 26252 22778 26280 22918
rect 26240 22772 26292 22778
rect 26240 22714 26292 22720
rect 26148 22568 26200 22574
rect 26148 22510 26200 22516
rect 26240 22568 26292 22574
rect 26240 22510 26292 22516
rect 26160 22012 26188 22510
rect 26252 22234 26280 22510
rect 26240 22228 26292 22234
rect 26240 22170 26292 22176
rect 26240 22024 26292 22030
rect 26160 21984 26240 22012
rect 26240 21966 26292 21972
rect 26056 21888 26108 21894
rect 26056 21830 26108 21836
rect 25504 21684 25556 21690
rect 25504 21626 25556 21632
rect 25688 21684 25740 21690
rect 25688 21626 25740 21632
rect 25504 21548 25556 21554
rect 25504 21490 25556 21496
rect 25516 21434 25544 21490
rect 25516 21406 25636 21434
rect 25608 20074 25636 21406
rect 25700 21146 25728 21626
rect 25780 21616 25832 21622
rect 25778 21584 25780 21593
rect 25832 21584 25834 21593
rect 25778 21519 25834 21528
rect 25780 21344 25832 21350
rect 25780 21286 25832 21292
rect 25688 21140 25740 21146
rect 25688 21082 25740 21088
rect 25608 20046 25728 20074
rect 25596 19848 25648 19854
rect 25596 19790 25648 19796
rect 25608 18290 25636 19790
rect 25700 18698 25728 20046
rect 25792 19836 25820 21286
rect 25872 21140 25924 21146
rect 25872 21082 25924 21088
rect 25884 20534 25912 21082
rect 25872 20528 25924 20534
rect 25872 20470 25924 20476
rect 25964 20460 26016 20466
rect 26068 20448 26096 21830
rect 26016 20420 26096 20448
rect 26148 20460 26200 20466
rect 25964 20402 26016 20408
rect 26252 20448 26280 21966
rect 26200 20420 26280 20448
rect 26148 20402 26200 20408
rect 26056 20324 26108 20330
rect 26056 20266 26108 20272
rect 25964 20256 26016 20262
rect 25964 20198 26016 20204
rect 25976 19990 26004 20198
rect 25964 19984 26016 19990
rect 25964 19926 26016 19932
rect 25964 19848 26016 19854
rect 25792 19808 25964 19836
rect 25964 19790 26016 19796
rect 25778 19408 25834 19417
rect 25778 19343 25834 19352
rect 25792 19242 25820 19343
rect 25780 19236 25832 19242
rect 25780 19178 25832 19184
rect 25688 18692 25740 18698
rect 25688 18634 25740 18640
rect 25596 18284 25648 18290
rect 25596 18226 25648 18232
rect 25792 18222 25820 19178
rect 25976 18902 26004 19790
rect 26068 19689 26096 20266
rect 26160 19786 26188 20402
rect 26240 20324 26292 20330
rect 26240 20266 26292 20272
rect 26252 20058 26280 20266
rect 26344 20058 26372 23258
rect 26436 20058 26464 24210
rect 26620 22642 26648 25638
rect 26712 24750 26740 26279
rect 26700 24744 26752 24750
rect 26700 24686 26752 24692
rect 26804 24154 26832 26454
rect 26896 25106 26924 28070
rect 26988 25294 27016 28902
rect 26976 25288 27028 25294
rect 26976 25230 27028 25236
rect 26896 25078 27016 25106
rect 26884 24880 26936 24886
rect 26884 24822 26936 24828
rect 26896 24342 26924 24822
rect 26884 24336 26936 24342
rect 26884 24278 26936 24284
rect 26804 24138 26924 24154
rect 26804 24132 26936 24138
rect 26804 24126 26884 24132
rect 26884 24074 26936 24080
rect 26988 23798 27016 25078
rect 26976 23792 27028 23798
rect 26976 23734 27028 23740
rect 26700 23588 26752 23594
rect 26700 23530 26752 23536
rect 26516 22636 26568 22642
rect 26516 22578 26568 22584
rect 26608 22636 26660 22642
rect 26608 22578 26660 22584
rect 26528 21962 26556 22578
rect 26620 22098 26648 22578
rect 26608 22092 26660 22098
rect 26608 22034 26660 22040
rect 26516 21956 26568 21962
rect 26516 21898 26568 21904
rect 26528 21146 26556 21898
rect 26516 21140 26568 21146
rect 26516 21082 26568 21088
rect 26712 21010 26740 23530
rect 26988 23118 27016 23734
rect 27080 23730 27108 28970
rect 27172 27690 27200 30552
rect 27344 29504 27396 29510
rect 27344 29446 27396 29452
rect 27356 29306 27384 29446
rect 27344 29300 27396 29306
rect 27344 29242 27396 29248
rect 27172 27662 27292 27690
rect 27160 24812 27212 24818
rect 27160 24754 27212 24760
rect 27172 24274 27200 24754
rect 27160 24268 27212 24274
rect 27160 24210 27212 24216
rect 27068 23724 27120 23730
rect 27068 23666 27120 23672
rect 26976 23112 27028 23118
rect 26976 23054 27028 23060
rect 27160 23044 27212 23050
rect 27160 22986 27212 22992
rect 27172 22642 27200 22986
rect 27160 22636 27212 22642
rect 27160 22578 27212 22584
rect 27160 22228 27212 22234
rect 27160 22170 27212 22176
rect 27172 21350 27200 22170
rect 27264 22094 27292 27662
rect 27344 26784 27396 26790
rect 27344 26726 27396 26732
rect 27356 26246 27384 26726
rect 27344 26240 27396 26246
rect 27344 26182 27396 26188
rect 27344 25220 27396 25226
rect 27344 25162 27396 25168
rect 27356 24750 27384 25162
rect 27344 24744 27396 24750
rect 27344 24686 27396 24692
rect 27356 24410 27384 24686
rect 27344 24404 27396 24410
rect 27344 24346 27396 24352
rect 27448 24290 27476 30670
rect 27540 26518 27568 31282
rect 27724 31278 27752 31622
rect 27712 31272 27764 31278
rect 27712 31214 27764 31220
rect 27712 31136 27764 31142
rect 27710 31104 27712 31113
rect 27764 31104 27766 31113
rect 27710 31039 27766 31048
rect 27620 29708 27672 29714
rect 27620 29650 27672 29656
rect 27632 29510 27660 29650
rect 27620 29504 27672 29510
rect 27620 29446 27672 29452
rect 27528 26512 27580 26518
rect 27528 26454 27580 26460
rect 27632 26450 27660 29446
rect 27620 26444 27672 26450
rect 27620 26386 27672 26392
rect 27448 24262 27568 24290
rect 27436 23724 27488 23730
rect 27356 23684 27436 23712
rect 27356 22642 27384 23684
rect 27436 23666 27488 23672
rect 27540 23594 27568 24262
rect 27620 24132 27672 24138
rect 27620 24074 27672 24080
rect 27632 23594 27660 24074
rect 27724 23730 27752 31039
rect 27804 30796 27856 30802
rect 27804 30738 27856 30744
rect 27816 29510 27844 30738
rect 27804 29504 27856 29510
rect 27804 29446 27856 29452
rect 27908 27674 27936 32234
rect 28264 31816 28316 31822
rect 28264 31758 28316 31764
rect 27988 31680 28040 31686
rect 27988 31622 28040 31628
rect 28000 31414 28028 31622
rect 27988 31408 28040 31414
rect 27988 31350 28040 31356
rect 28276 30938 28304 31758
rect 28264 30932 28316 30938
rect 28264 30874 28316 30880
rect 28460 30598 28488 32302
rect 28552 30682 28580 32778
rect 28644 30802 28672 34002
rect 28736 33318 28764 35702
rect 28920 35086 28948 37266
rect 29012 36922 29040 37810
rect 29288 37262 29316 38218
rect 29472 38010 29500 38218
rect 29460 38004 29512 38010
rect 29460 37946 29512 37952
rect 29460 37800 29512 37806
rect 29460 37742 29512 37748
rect 29276 37256 29328 37262
rect 29276 37198 29328 37204
rect 29000 36916 29052 36922
rect 29000 36858 29052 36864
rect 29472 36802 29500 37742
rect 29564 37330 29592 38286
rect 29656 38010 29684 38354
rect 29644 38004 29696 38010
rect 29644 37946 29696 37952
rect 29552 37324 29604 37330
rect 29552 37266 29604 37272
rect 29368 36780 29420 36786
rect 29472 36774 29684 36802
rect 29368 36722 29420 36728
rect 28908 35080 28960 35086
rect 28908 35022 28960 35028
rect 28816 34944 28868 34950
rect 28816 34886 28868 34892
rect 28828 34746 28856 34886
rect 28816 34740 28868 34746
rect 28816 34682 28868 34688
rect 28816 34128 28868 34134
rect 28816 34070 28868 34076
rect 28828 33862 28856 34070
rect 28816 33856 28868 33862
rect 28816 33798 28868 33804
rect 28724 33312 28776 33318
rect 28724 33254 28776 33260
rect 28724 32768 28776 32774
rect 28724 32710 28776 32716
rect 28736 32434 28764 32710
rect 28724 32428 28776 32434
rect 28724 32370 28776 32376
rect 28736 31958 28764 32370
rect 28724 31952 28776 31958
rect 28724 31894 28776 31900
rect 28632 30796 28684 30802
rect 28632 30738 28684 30744
rect 28552 30654 28672 30682
rect 28448 30592 28500 30598
rect 28448 30534 28500 30540
rect 28460 29866 28488 30534
rect 28080 29844 28132 29850
rect 28460 29838 28580 29866
rect 28080 29786 28132 29792
rect 28092 29510 28120 29786
rect 28446 29608 28502 29617
rect 28446 29543 28448 29552
rect 28500 29543 28502 29552
rect 28448 29514 28500 29520
rect 28080 29504 28132 29510
rect 28080 29446 28132 29452
rect 28356 29504 28408 29510
rect 28356 29446 28408 29452
rect 27896 27668 27948 27674
rect 27896 27610 27948 27616
rect 27804 27328 27856 27334
rect 27804 27270 27856 27276
rect 27896 27328 27948 27334
rect 27896 27270 27948 27276
rect 27816 27130 27844 27270
rect 27804 27124 27856 27130
rect 27804 27066 27856 27072
rect 27908 26926 27936 27270
rect 27896 26920 27948 26926
rect 27896 26862 27948 26868
rect 27988 26444 28040 26450
rect 27988 26386 28040 26392
rect 27896 25900 27948 25906
rect 27896 25842 27948 25848
rect 27804 25696 27856 25702
rect 27804 25638 27856 25644
rect 27816 25430 27844 25638
rect 27804 25424 27856 25430
rect 27804 25366 27856 25372
rect 27908 25294 27936 25842
rect 27896 25288 27948 25294
rect 27896 25230 27948 25236
rect 27804 25220 27856 25226
rect 27804 25162 27856 25168
rect 27816 24721 27844 25162
rect 27802 24712 27858 24721
rect 27802 24647 27858 24656
rect 27896 24200 27948 24206
rect 27896 24142 27948 24148
rect 27712 23724 27764 23730
rect 27712 23666 27764 23672
rect 27908 23662 27936 24142
rect 27896 23656 27948 23662
rect 27896 23598 27948 23604
rect 27528 23588 27580 23594
rect 27528 23530 27580 23536
rect 27620 23588 27672 23594
rect 27620 23530 27672 23536
rect 27540 23338 27568 23530
rect 27540 23310 27660 23338
rect 27528 23248 27580 23254
rect 27528 23190 27580 23196
rect 27540 22778 27568 23190
rect 27632 23186 27660 23310
rect 27620 23180 27672 23186
rect 27620 23122 27672 23128
rect 28000 22778 28028 26386
rect 27528 22772 27580 22778
rect 27528 22714 27580 22720
rect 27988 22772 28040 22778
rect 27988 22714 28040 22720
rect 27344 22636 27396 22642
rect 27344 22578 27396 22584
rect 27436 22636 27488 22642
rect 27436 22578 27488 22584
rect 27264 22066 27384 22094
rect 27160 21344 27212 21350
rect 27160 21286 27212 21292
rect 27356 21146 27384 22066
rect 27448 21418 27476 22578
rect 27712 22228 27764 22234
rect 27712 22170 27764 22176
rect 27724 22030 27752 22170
rect 28092 22094 28120 29446
rect 28368 29306 28396 29446
rect 28356 29300 28408 29306
rect 28356 29242 28408 29248
rect 28448 27668 28500 27674
rect 28448 27610 28500 27616
rect 28172 27464 28224 27470
rect 28172 27406 28224 27412
rect 28184 26586 28212 27406
rect 28264 26784 28316 26790
rect 28264 26726 28316 26732
rect 28172 26580 28224 26586
rect 28172 26522 28224 26528
rect 28276 26489 28304 26726
rect 28262 26480 28318 26489
rect 28262 26415 28318 26424
rect 28276 26314 28304 26415
rect 28264 26308 28316 26314
rect 28264 26250 28316 26256
rect 28172 26240 28224 26246
rect 28172 26182 28224 26188
rect 28184 24818 28212 26182
rect 28276 25158 28304 26250
rect 28264 25152 28316 25158
rect 28264 25094 28316 25100
rect 28172 24812 28224 24818
rect 28172 24754 28224 24760
rect 28184 23866 28212 24754
rect 28356 24200 28408 24206
rect 28276 24160 28356 24188
rect 28172 23860 28224 23866
rect 28172 23802 28224 23808
rect 28172 22432 28224 22438
rect 28172 22374 28224 22380
rect 28000 22066 28120 22094
rect 27712 22024 27764 22030
rect 27712 21966 27764 21972
rect 27528 21888 27580 21894
rect 27528 21830 27580 21836
rect 27620 21888 27672 21894
rect 27896 21888 27948 21894
rect 27620 21830 27672 21836
rect 27816 21848 27896 21876
rect 27436 21412 27488 21418
rect 27436 21354 27488 21360
rect 27540 21146 27568 21830
rect 27632 21146 27660 21830
rect 27710 21584 27766 21593
rect 27710 21519 27712 21528
rect 27764 21519 27766 21528
rect 27712 21490 27764 21496
rect 27344 21140 27396 21146
rect 27344 21082 27396 21088
rect 27528 21140 27580 21146
rect 27528 21082 27580 21088
rect 27620 21140 27672 21146
rect 27620 21082 27672 21088
rect 27252 21072 27304 21078
rect 27252 21014 27304 21020
rect 26700 21004 26752 21010
rect 26700 20946 26752 20952
rect 26884 20936 26936 20942
rect 26884 20878 26936 20884
rect 27068 20936 27120 20942
rect 27068 20878 27120 20884
rect 26896 20097 26924 20878
rect 27080 20534 27108 20878
rect 27264 20806 27292 21014
rect 27344 20936 27396 20942
rect 27344 20878 27396 20884
rect 27528 20936 27580 20942
rect 27816 20924 27844 21848
rect 27896 21830 27948 21836
rect 27580 20896 27844 20924
rect 27528 20878 27580 20884
rect 27252 20800 27304 20806
rect 27252 20742 27304 20748
rect 27068 20528 27120 20534
rect 27068 20470 27120 20476
rect 26882 20088 26938 20097
rect 26240 20052 26292 20058
rect 26240 19994 26292 20000
rect 26332 20052 26384 20058
rect 26332 19994 26384 20000
rect 26424 20052 26476 20058
rect 26882 20023 26938 20032
rect 26424 19994 26476 20000
rect 26148 19780 26200 19786
rect 26148 19722 26200 19728
rect 26792 19780 26844 19786
rect 26792 19722 26844 19728
rect 26054 19680 26110 19689
rect 26054 19615 26110 19624
rect 26804 19174 26832 19722
rect 26792 19168 26844 19174
rect 26792 19110 26844 19116
rect 26804 18970 26832 19110
rect 26792 18964 26844 18970
rect 26792 18906 26844 18912
rect 25964 18896 26016 18902
rect 25964 18838 26016 18844
rect 25964 18624 26016 18630
rect 25964 18566 26016 18572
rect 25976 18290 26004 18566
rect 25964 18284 26016 18290
rect 25964 18226 26016 18232
rect 25780 18216 25832 18222
rect 25780 18158 25832 18164
rect 26240 18148 26292 18154
rect 26240 18090 26292 18096
rect 26252 17882 26280 18090
rect 26516 18080 26568 18086
rect 26516 18022 26568 18028
rect 26240 17876 26292 17882
rect 26240 17818 26292 17824
rect 26240 16652 26292 16658
rect 26240 16594 26292 16600
rect 26056 16584 26108 16590
rect 26056 16526 26108 16532
rect 25964 16516 26016 16522
rect 25964 16458 26016 16464
rect 25976 15502 26004 16458
rect 26068 15502 26096 16526
rect 26252 15502 26280 16594
rect 26424 16448 26476 16454
rect 26424 16390 26476 16396
rect 26436 16114 26464 16390
rect 26424 16108 26476 16114
rect 26424 16050 26476 16056
rect 25504 15496 25556 15502
rect 25504 15438 25556 15444
rect 25964 15496 26016 15502
rect 25964 15438 26016 15444
rect 26056 15496 26108 15502
rect 26056 15438 26108 15444
rect 26240 15496 26292 15502
rect 26240 15438 26292 15444
rect 25516 15366 25544 15438
rect 25504 15360 25556 15366
rect 25504 15302 25556 15308
rect 25688 15360 25740 15366
rect 25688 15302 25740 15308
rect 25700 15026 25728 15302
rect 26068 15162 26096 15438
rect 26056 15156 26108 15162
rect 26056 15098 26108 15104
rect 25688 15020 25740 15026
rect 25688 14962 25740 14968
rect 26424 15020 26476 15026
rect 26424 14962 26476 14968
rect 25596 14952 25648 14958
rect 25594 14920 25596 14929
rect 26148 14952 26200 14958
rect 25648 14920 25650 14929
rect 26148 14894 26200 14900
rect 25594 14855 25650 14864
rect 25596 14816 25648 14822
rect 25596 14758 25648 14764
rect 25608 13326 25636 14758
rect 26054 13968 26110 13977
rect 25780 13932 25832 13938
rect 26160 13938 26188 14894
rect 26332 14816 26384 14822
rect 26332 14758 26384 14764
rect 26240 14340 26292 14346
rect 26240 14282 26292 14288
rect 26054 13903 26056 13912
rect 25780 13874 25832 13880
rect 26108 13903 26110 13912
rect 26148 13932 26200 13938
rect 26056 13874 26108 13880
rect 26148 13874 26200 13880
rect 25792 13682 25820 13874
rect 26252 13818 26280 14282
rect 26344 14074 26372 14758
rect 26436 14278 26464 14962
rect 26424 14272 26476 14278
rect 26424 14214 26476 14220
rect 26332 14068 26384 14074
rect 26332 14010 26384 14016
rect 25976 13802 26280 13818
rect 25964 13796 26280 13802
rect 26016 13790 26280 13796
rect 25964 13738 26016 13744
rect 26056 13728 26108 13734
rect 25792 13654 26004 13682
rect 26240 13728 26292 13734
rect 26056 13670 26108 13676
rect 26160 13688 26240 13716
rect 25780 13388 25832 13394
rect 25780 13330 25832 13336
rect 25596 13320 25648 13326
rect 25596 13262 25648 13268
rect 25608 12850 25636 13262
rect 25596 12844 25648 12850
rect 25596 12786 25648 12792
rect 25424 12406 25636 12434
rect 25320 11824 25372 11830
rect 25320 11766 25372 11772
rect 24452 11716 24532 11744
rect 24584 11756 24636 11762
rect 24400 11698 24452 11704
rect 24768 11756 24820 11762
rect 24636 11716 24716 11744
rect 24584 11698 24636 11704
rect 24308 11144 24360 11150
rect 24308 11086 24360 11092
rect 24216 11076 24268 11082
rect 24216 11018 24268 11024
rect 24228 9586 24256 11018
rect 24216 9580 24268 9586
rect 24216 9522 24268 9528
rect 24320 9466 24348 11086
rect 24412 10674 24440 11698
rect 24584 11280 24636 11286
rect 24584 11222 24636 11228
rect 24400 10668 24452 10674
rect 24400 10610 24452 10616
rect 24492 10600 24544 10606
rect 24492 10542 24544 10548
rect 24400 10124 24452 10130
rect 24400 10066 24452 10072
rect 24412 9586 24440 10066
rect 24400 9580 24452 9586
rect 24400 9522 24452 9528
rect 24228 9450 24348 9466
rect 24216 9444 24348 9450
rect 24268 9438 24348 9444
rect 24216 9386 24268 9392
rect 24228 9042 24256 9386
rect 24308 9376 24360 9382
rect 24308 9318 24360 9324
rect 24216 9036 24268 9042
rect 24216 8978 24268 8984
rect 24320 8634 24348 9318
rect 24308 8628 24360 8634
rect 24308 8570 24360 8576
rect 24216 8492 24268 8498
rect 24136 8452 24216 8480
rect 24216 8434 24268 8440
rect 24032 7744 24084 7750
rect 24032 7686 24084 7692
rect 24044 7410 24072 7686
rect 24032 7404 24084 7410
rect 24032 7346 24084 7352
rect 23848 6996 23900 7002
rect 23848 6938 23900 6944
rect 23860 6662 23888 6938
rect 23572 6656 23624 6662
rect 23572 6598 23624 6604
rect 23848 6656 23900 6662
rect 23848 6598 23900 6604
rect 22928 6384 22980 6390
rect 22928 6326 22980 6332
rect 23480 6384 23532 6390
rect 23480 6326 23532 6332
rect 22652 6316 22704 6322
rect 22652 6258 22704 6264
rect 22560 5908 22612 5914
rect 22560 5850 22612 5856
rect 22664 5710 22692 6258
rect 22940 5710 22968 6326
rect 23112 6316 23164 6322
rect 23112 6258 23164 6264
rect 23020 6112 23072 6118
rect 23020 6054 23072 6060
rect 22652 5704 22704 5710
rect 22652 5646 22704 5652
rect 22928 5704 22980 5710
rect 22928 5646 22980 5652
rect 22928 5568 22980 5574
rect 22928 5510 22980 5516
rect 22652 5228 22704 5234
rect 22652 5170 22704 5176
rect 22376 5160 22428 5166
rect 22376 5102 22428 5108
rect 22664 4554 22692 5170
rect 22940 4690 22968 5510
rect 23032 5234 23060 6054
rect 23124 5710 23152 6258
rect 23296 6180 23348 6186
rect 23296 6122 23348 6128
rect 23204 5840 23256 5846
rect 23204 5782 23256 5788
rect 23112 5704 23164 5710
rect 23112 5646 23164 5652
rect 23124 5234 23152 5646
rect 23216 5234 23244 5782
rect 23308 5710 23336 6122
rect 23296 5704 23348 5710
rect 23296 5646 23348 5652
rect 23020 5228 23072 5234
rect 23020 5170 23072 5176
rect 23112 5228 23164 5234
rect 23112 5170 23164 5176
rect 23204 5228 23256 5234
rect 23204 5170 23256 5176
rect 23308 5098 23336 5646
rect 23296 5092 23348 5098
rect 23296 5034 23348 5040
rect 23388 5024 23440 5030
rect 23388 4966 23440 4972
rect 23400 4826 23428 4966
rect 23388 4820 23440 4826
rect 23492 4808 23520 6326
rect 23584 6322 23612 6598
rect 23572 6316 23624 6322
rect 23572 6258 23624 6264
rect 24228 5778 24256 8434
rect 24308 7744 24360 7750
rect 24308 7686 24360 7692
rect 24320 6322 24348 7686
rect 24504 7410 24532 10542
rect 24596 9382 24624 11222
rect 24584 9376 24636 9382
rect 24584 9318 24636 9324
rect 24688 9110 24716 11716
rect 24768 11698 24820 11704
rect 25044 11756 25096 11762
rect 25044 11698 25096 11704
rect 25056 11218 25084 11698
rect 25044 11212 25096 11218
rect 25044 11154 25096 11160
rect 25044 10124 25096 10130
rect 25044 10066 25096 10072
rect 24768 9444 24820 9450
rect 24820 9404 24900 9432
rect 24768 9386 24820 9392
rect 24676 9104 24728 9110
rect 24676 9046 24728 9052
rect 24872 8974 24900 9404
rect 25056 8974 25084 10066
rect 25318 9072 25374 9081
rect 25318 9007 25320 9016
rect 25372 9007 25374 9016
rect 25320 8978 25372 8984
rect 24860 8968 24912 8974
rect 24860 8910 24912 8916
rect 25044 8968 25096 8974
rect 25044 8910 25096 8916
rect 24584 8900 24636 8906
rect 24584 8842 24636 8848
rect 24596 7410 24624 8842
rect 25136 8832 25188 8838
rect 25136 8774 25188 8780
rect 24492 7404 24544 7410
rect 24492 7346 24544 7352
rect 24584 7404 24636 7410
rect 24584 7346 24636 7352
rect 25148 7206 25176 8774
rect 25332 8566 25360 8978
rect 25412 8900 25464 8906
rect 25412 8842 25464 8848
rect 25320 8560 25372 8566
rect 25320 8502 25372 8508
rect 25424 8498 25452 8842
rect 25412 8492 25464 8498
rect 25412 8434 25464 8440
rect 25424 8401 25452 8434
rect 25410 8392 25466 8401
rect 25410 8327 25466 8336
rect 25320 8288 25372 8294
rect 25320 8230 25372 8236
rect 25332 7478 25360 8230
rect 25320 7472 25372 7478
rect 25320 7414 25372 7420
rect 25228 7404 25280 7410
rect 25228 7346 25280 7352
rect 24768 7200 24820 7206
rect 24768 7142 24820 7148
rect 24860 7200 24912 7206
rect 24860 7142 24912 7148
rect 25044 7200 25096 7206
rect 25044 7142 25096 7148
rect 25136 7200 25188 7206
rect 25136 7142 25188 7148
rect 24780 6322 24808 7142
rect 24872 6866 24900 7142
rect 24860 6860 24912 6866
rect 24860 6802 24912 6808
rect 24952 6792 25004 6798
rect 24952 6734 25004 6740
rect 24964 6458 24992 6734
rect 24952 6452 25004 6458
rect 24952 6394 25004 6400
rect 24308 6316 24360 6322
rect 24308 6258 24360 6264
rect 24768 6316 24820 6322
rect 24768 6258 24820 6264
rect 24216 5772 24268 5778
rect 24216 5714 24268 5720
rect 23572 5704 23624 5710
rect 23572 5646 23624 5652
rect 23664 5704 23716 5710
rect 23664 5646 23716 5652
rect 24768 5704 24820 5710
rect 25056 5692 25084 7142
rect 25240 6458 25268 7346
rect 25412 7336 25464 7342
rect 25412 7278 25464 7284
rect 25424 7002 25452 7278
rect 25412 6996 25464 7002
rect 25412 6938 25464 6944
rect 25504 6724 25556 6730
rect 25504 6666 25556 6672
rect 25320 6656 25372 6662
rect 25320 6598 25372 6604
rect 25228 6452 25280 6458
rect 25228 6394 25280 6400
rect 25332 6390 25360 6598
rect 25320 6384 25372 6390
rect 25320 6326 25372 6332
rect 24820 5664 25084 5692
rect 24768 5646 24820 5652
rect 23584 5370 23612 5646
rect 23676 5370 23704 5646
rect 23756 5568 23808 5574
rect 23756 5510 23808 5516
rect 24400 5568 24452 5574
rect 24400 5510 24452 5516
rect 23572 5364 23624 5370
rect 23572 5306 23624 5312
rect 23664 5364 23716 5370
rect 23664 5306 23716 5312
rect 23572 4820 23624 4826
rect 23492 4780 23572 4808
rect 23388 4762 23440 4768
rect 23572 4762 23624 4768
rect 23768 4690 23796 5510
rect 24412 5166 24440 5510
rect 25516 5234 25544 6666
rect 24860 5228 24912 5234
rect 24860 5170 24912 5176
rect 25504 5228 25556 5234
rect 25504 5170 25556 5176
rect 24400 5160 24452 5166
rect 24400 5102 24452 5108
rect 24400 5024 24452 5030
rect 24400 4966 24452 4972
rect 24412 4826 24440 4966
rect 24400 4820 24452 4826
rect 24400 4762 24452 4768
rect 24596 4814 24808 4842
rect 24596 4690 24624 4814
rect 24676 4752 24728 4758
rect 24676 4694 24728 4700
rect 22928 4684 22980 4690
rect 22928 4626 22980 4632
rect 23756 4684 23808 4690
rect 23756 4626 23808 4632
rect 24584 4684 24636 4690
rect 24584 4626 24636 4632
rect 22652 4548 22704 4554
rect 22652 4490 22704 4496
rect 23480 4548 23532 4554
rect 23480 4490 23532 4496
rect 24584 4548 24636 4554
rect 24688 4536 24716 4694
rect 24780 4604 24808 4814
rect 24872 4758 24900 5170
rect 25504 4820 25556 4826
rect 25504 4762 25556 4768
rect 24860 4752 24912 4758
rect 24860 4694 24912 4700
rect 25412 4684 25464 4690
rect 25412 4626 25464 4632
rect 24952 4616 25004 4622
rect 24780 4576 24952 4604
rect 24952 4558 25004 4564
rect 24636 4508 24716 4536
rect 24584 4490 24636 4496
rect 20996 4276 21048 4282
rect 20996 4218 21048 4224
rect 22664 4214 22692 4490
rect 23204 4480 23256 4486
rect 23388 4480 23440 4486
rect 23256 4440 23388 4468
rect 23204 4422 23256 4428
rect 23388 4422 23440 4428
rect 23492 4214 23520 4490
rect 25044 4480 25096 4486
rect 25044 4422 25096 4428
rect 25056 4214 25084 4422
rect 22652 4208 22704 4214
rect 22652 4150 22704 4156
rect 23480 4208 23532 4214
rect 23480 4150 23532 4156
rect 25044 4208 25096 4214
rect 25044 4150 25096 4156
rect 25424 4010 25452 4626
rect 25516 4146 25544 4762
rect 25504 4140 25556 4146
rect 25504 4082 25556 4088
rect 25412 4004 25464 4010
rect 25412 3946 25464 3952
rect 25516 3942 25544 4082
rect 25504 3936 25556 3942
rect 25504 3878 25556 3884
rect 17224 3188 17276 3194
rect 17224 3130 17276 3136
rect 25608 3058 25636 12406
rect 25792 10282 25820 13330
rect 25872 13320 25924 13326
rect 25872 13262 25924 13268
rect 25884 12986 25912 13262
rect 25872 12980 25924 12986
rect 25872 12922 25924 12928
rect 25976 12288 26004 13654
rect 26068 13394 26096 13670
rect 26056 13388 26108 13394
rect 26056 13330 26108 13336
rect 26160 13326 26188 13688
rect 26240 13670 26292 13676
rect 26238 13424 26294 13433
rect 26238 13359 26240 13368
rect 26292 13359 26294 13368
rect 26240 13330 26292 13336
rect 26148 13320 26200 13326
rect 26148 13262 26200 13268
rect 26240 13184 26292 13190
rect 26240 13126 26292 13132
rect 26148 12912 26200 12918
rect 26146 12880 26148 12889
rect 26200 12880 26202 12889
rect 26146 12815 26202 12824
rect 26252 12714 26280 13126
rect 26344 12850 26372 14010
rect 26424 13864 26476 13870
rect 26424 13806 26476 13812
rect 26436 13433 26464 13806
rect 26422 13424 26478 13433
rect 26422 13359 26478 13368
rect 26528 13326 26556 18022
rect 26896 17882 26924 20023
rect 27080 19786 27108 20470
rect 27356 20466 27384 20878
rect 28000 20602 28028 22066
rect 28184 21962 28212 22374
rect 28276 22166 28304 24160
rect 28356 24142 28408 24148
rect 28264 22160 28316 22166
rect 28264 22102 28316 22108
rect 28276 21962 28304 22102
rect 28356 22024 28408 22030
rect 28356 21966 28408 21972
rect 28172 21956 28224 21962
rect 28172 21898 28224 21904
rect 28264 21956 28316 21962
rect 28264 21898 28316 21904
rect 28184 21690 28212 21898
rect 28172 21684 28224 21690
rect 28172 21626 28224 21632
rect 27988 20596 28040 20602
rect 27988 20538 28040 20544
rect 28276 20534 28304 21898
rect 28264 20528 28316 20534
rect 28264 20470 28316 20476
rect 27344 20460 27396 20466
rect 27344 20402 27396 20408
rect 27620 20460 27672 20466
rect 27620 20402 27672 20408
rect 27160 20256 27212 20262
rect 27160 20198 27212 20204
rect 27172 19922 27200 20198
rect 27160 19916 27212 19922
rect 27160 19858 27212 19864
rect 27356 19854 27384 20402
rect 27632 20262 27660 20402
rect 27436 20256 27488 20262
rect 27436 20198 27488 20204
rect 27620 20256 27672 20262
rect 27620 20198 27672 20204
rect 27344 19848 27396 19854
rect 27264 19808 27344 19836
rect 27068 19780 27120 19786
rect 27068 19722 27120 19728
rect 27264 19378 27292 19808
rect 27344 19790 27396 19796
rect 27448 19553 27476 20198
rect 27620 19780 27672 19786
rect 27620 19722 27672 19728
rect 27434 19544 27490 19553
rect 27434 19479 27490 19488
rect 27252 19372 27304 19378
rect 27252 19314 27304 19320
rect 27344 19372 27396 19378
rect 27344 19314 27396 19320
rect 27356 18766 27384 19314
rect 27344 18760 27396 18766
rect 27344 18702 27396 18708
rect 26884 17876 26936 17882
rect 26884 17818 26936 17824
rect 27448 17678 27476 19479
rect 27528 19372 27580 19378
rect 27632 19360 27660 19722
rect 28262 19408 28318 19417
rect 27580 19332 27660 19360
rect 27528 19314 27580 19320
rect 27632 18358 27660 19332
rect 27804 19372 27856 19378
rect 27804 19314 27856 19320
rect 28172 19372 28224 19378
rect 28262 19343 28264 19352
rect 28172 19314 28224 19320
rect 28316 19343 28318 19352
rect 28264 19314 28316 19320
rect 27620 18352 27672 18358
rect 27620 18294 27672 18300
rect 27710 17776 27766 17785
rect 27710 17711 27712 17720
rect 27764 17711 27766 17720
rect 27712 17682 27764 17688
rect 27436 17672 27488 17678
rect 27436 17614 27488 17620
rect 27160 16448 27212 16454
rect 27160 16390 27212 16396
rect 27172 15910 27200 16390
rect 27252 16176 27304 16182
rect 27252 16118 27304 16124
rect 27160 15904 27212 15910
rect 27160 15846 27212 15852
rect 27172 15502 27200 15846
rect 27160 15496 27212 15502
rect 27160 15438 27212 15444
rect 26700 15360 26752 15366
rect 26700 15302 26752 15308
rect 26712 13938 26740 15302
rect 27160 15020 27212 15026
rect 27160 14962 27212 14968
rect 27172 14346 27200 14962
rect 27160 14340 27212 14346
rect 27160 14282 27212 14288
rect 27264 14074 27292 16118
rect 27344 16108 27396 16114
rect 27344 16050 27396 16056
rect 27356 15978 27384 16050
rect 27344 15972 27396 15978
rect 27344 15914 27396 15920
rect 27356 15706 27384 15914
rect 27344 15700 27396 15706
rect 27344 15642 27396 15648
rect 27344 15360 27396 15366
rect 27344 15302 27396 15308
rect 27356 15162 27384 15302
rect 27344 15156 27396 15162
rect 27344 15098 27396 15104
rect 27252 14068 27304 14074
rect 27252 14010 27304 14016
rect 26700 13932 26752 13938
rect 26700 13874 26752 13880
rect 26976 13728 27028 13734
rect 26976 13670 27028 13676
rect 27344 13728 27396 13734
rect 27344 13670 27396 13676
rect 26516 13320 26568 13326
rect 26516 13262 26568 13268
rect 26792 13320 26844 13326
rect 26792 13262 26844 13268
rect 26332 12844 26384 12850
rect 26332 12786 26384 12792
rect 26240 12708 26292 12714
rect 26240 12650 26292 12656
rect 26528 12374 26556 13262
rect 26700 13184 26752 13190
rect 26700 13126 26752 13132
rect 26712 12986 26740 13126
rect 26700 12980 26752 12986
rect 26700 12922 26752 12928
rect 26606 12880 26662 12889
rect 26662 12838 26740 12866
rect 26606 12815 26662 12824
rect 26516 12368 26568 12374
rect 26516 12310 26568 12316
rect 26148 12300 26200 12306
rect 25976 12260 26148 12288
rect 26148 12242 26200 12248
rect 26056 12096 26108 12102
rect 26056 12038 26108 12044
rect 26068 11558 26096 12038
rect 26056 11552 26108 11558
rect 26056 11494 26108 11500
rect 26068 11014 26096 11494
rect 26160 11150 26188 12242
rect 26424 12232 26476 12238
rect 26424 12174 26476 12180
rect 26436 11694 26464 12174
rect 26424 11688 26476 11694
rect 26424 11630 26476 11636
rect 26436 11150 26464 11630
rect 26528 11354 26556 12310
rect 26608 12096 26660 12102
rect 26608 12038 26660 12044
rect 26620 11762 26648 12038
rect 26608 11756 26660 11762
rect 26608 11698 26660 11704
rect 26712 11558 26740 12838
rect 26804 12442 26832 13262
rect 26884 13252 26936 13258
rect 26884 13194 26936 13200
rect 26896 12646 26924 13194
rect 26988 12986 27016 13670
rect 27068 13456 27120 13462
rect 27068 13398 27120 13404
rect 26976 12980 27028 12986
rect 26976 12922 27028 12928
rect 26884 12640 26936 12646
rect 26884 12582 26936 12588
rect 26792 12436 26844 12442
rect 26792 12378 26844 12384
rect 26792 12232 26844 12238
rect 26792 12174 26844 12180
rect 26804 11898 26832 12174
rect 26792 11892 26844 11898
rect 26792 11834 26844 11840
rect 26976 11688 27028 11694
rect 26976 11630 27028 11636
rect 26700 11552 26752 11558
rect 26700 11494 26752 11500
rect 26516 11348 26568 11354
rect 26516 11290 26568 11296
rect 26148 11144 26200 11150
rect 26148 11086 26200 11092
rect 26424 11144 26476 11150
rect 26424 11086 26476 11092
rect 26516 11144 26568 11150
rect 26516 11086 26568 11092
rect 26056 11008 26108 11014
rect 26056 10950 26108 10956
rect 25792 10254 26004 10282
rect 25976 10198 26004 10254
rect 25964 10192 26016 10198
rect 25964 10134 26016 10140
rect 26068 9081 26096 10950
rect 26424 10532 26476 10538
rect 26424 10474 26476 10480
rect 26240 10056 26292 10062
rect 26240 9998 26292 10004
rect 26148 9920 26200 9926
rect 26148 9862 26200 9868
rect 26160 9586 26188 9862
rect 26148 9580 26200 9586
rect 26148 9522 26200 9528
rect 26054 9072 26110 9081
rect 26054 9007 26110 9016
rect 25964 8968 26016 8974
rect 25964 8910 26016 8916
rect 25976 7342 26004 8910
rect 26252 8090 26280 9998
rect 26332 9172 26384 9178
rect 26332 9114 26384 9120
rect 26344 8838 26372 9114
rect 26332 8832 26384 8838
rect 26332 8774 26384 8780
rect 26240 8084 26292 8090
rect 26240 8026 26292 8032
rect 26252 7478 26280 8026
rect 26344 7478 26372 8774
rect 26436 7546 26464 10474
rect 26528 9382 26556 11086
rect 26792 11008 26844 11014
rect 26792 10950 26844 10956
rect 26804 10674 26832 10950
rect 26792 10668 26844 10674
rect 26792 10610 26844 10616
rect 26608 10464 26660 10470
rect 26608 10406 26660 10412
rect 26620 9602 26648 10406
rect 26620 9574 26740 9602
rect 26988 9586 27016 11630
rect 27080 11150 27108 13398
rect 27356 13394 27384 13670
rect 27344 13388 27396 13394
rect 27344 13330 27396 13336
rect 27448 13326 27476 17614
rect 27816 17202 27844 19314
rect 27988 18284 28040 18290
rect 27988 18226 28040 18232
rect 27896 18080 27948 18086
rect 27896 18022 27948 18028
rect 27908 17678 27936 18022
rect 28000 17882 28028 18226
rect 27988 17876 28040 17882
rect 27988 17818 28040 17824
rect 28184 17678 28212 19314
rect 28368 18630 28396 21966
rect 28460 21622 28488 27610
rect 28552 21894 28580 29838
rect 28644 29170 28672 30654
rect 28632 29164 28684 29170
rect 28632 29106 28684 29112
rect 28644 27130 28672 29106
rect 28632 27124 28684 27130
rect 28632 27066 28684 27072
rect 28724 25696 28776 25702
rect 28724 25638 28776 25644
rect 28736 25294 28764 25638
rect 28724 25288 28776 25294
rect 28724 25230 28776 25236
rect 28632 24812 28684 24818
rect 28632 24754 28684 24760
rect 28644 23866 28672 24754
rect 28724 24336 28776 24342
rect 28724 24278 28776 24284
rect 28632 23860 28684 23866
rect 28632 23802 28684 23808
rect 28736 23798 28764 24278
rect 28724 23792 28776 23798
rect 28724 23734 28776 23740
rect 28828 22094 28856 33798
rect 28920 31890 28948 35022
rect 29000 33584 29052 33590
rect 29000 33526 29052 33532
rect 28908 31884 28960 31890
rect 28908 31826 28960 31832
rect 28920 29782 28948 31826
rect 29012 31482 29040 33526
rect 29380 31754 29408 36722
rect 29656 36718 29684 36774
rect 29644 36712 29696 36718
rect 29644 36654 29696 36660
rect 29656 35494 29684 36654
rect 29644 35488 29696 35494
rect 29644 35430 29696 35436
rect 29550 33144 29606 33153
rect 29550 33079 29606 33088
rect 29460 31816 29512 31822
rect 29460 31758 29512 31764
rect 29196 31726 29408 31754
rect 29092 31680 29144 31686
rect 29092 31622 29144 31628
rect 29000 31476 29052 31482
rect 29000 31418 29052 31424
rect 29104 29782 29132 31622
rect 28908 29776 28960 29782
rect 28908 29718 28960 29724
rect 29092 29776 29144 29782
rect 29092 29718 29144 29724
rect 28920 29646 28948 29718
rect 29000 29708 29052 29714
rect 29000 29650 29052 29656
rect 28908 29640 28960 29646
rect 28908 29582 28960 29588
rect 28920 29016 28948 29582
rect 29012 29306 29040 29650
rect 29000 29300 29052 29306
rect 29000 29242 29052 29248
rect 29104 29034 29132 29718
rect 29092 29028 29144 29034
rect 28920 28988 29040 29016
rect 29012 27606 29040 28988
rect 29092 28970 29144 28976
rect 29092 28756 29144 28762
rect 29092 28698 29144 28704
rect 29104 28665 29132 28698
rect 29090 28656 29146 28665
rect 29090 28591 29146 28600
rect 29000 27600 29052 27606
rect 29000 27542 29052 27548
rect 29012 25294 29040 27542
rect 29092 26240 29144 26246
rect 29092 26182 29144 26188
rect 29104 25770 29132 26182
rect 29092 25764 29144 25770
rect 29092 25706 29144 25712
rect 29000 25288 29052 25294
rect 29000 25230 29052 25236
rect 29092 25152 29144 25158
rect 29092 25094 29144 25100
rect 29104 24954 29132 25094
rect 29092 24948 29144 24954
rect 29092 24890 29144 24896
rect 29196 23322 29224 31726
rect 29472 31142 29500 31758
rect 29460 31136 29512 31142
rect 29460 31078 29512 31084
rect 29472 30666 29500 31078
rect 29460 30660 29512 30666
rect 29460 30602 29512 30608
rect 29276 29504 29328 29510
rect 29276 29446 29328 29452
rect 29368 29504 29420 29510
rect 29368 29446 29420 29452
rect 29288 29306 29316 29446
rect 29276 29300 29328 29306
rect 29276 29242 29328 29248
rect 29276 28960 29328 28966
rect 29276 28902 29328 28908
rect 29288 28694 29316 28902
rect 29276 28688 29328 28694
rect 29276 28630 29328 28636
rect 29276 24744 29328 24750
rect 29276 24686 29328 24692
rect 29184 23316 29236 23322
rect 29184 23258 29236 23264
rect 29288 22234 29316 24686
rect 29276 22228 29328 22234
rect 29276 22170 29328 22176
rect 29380 22094 29408 29446
rect 29460 26852 29512 26858
rect 29460 26794 29512 26800
rect 29472 24886 29500 26794
rect 29460 24880 29512 24886
rect 29460 24822 29512 24828
rect 29564 24206 29592 33079
rect 29644 31340 29696 31346
rect 29644 31282 29696 31288
rect 29656 30938 29684 31282
rect 29644 30932 29696 30938
rect 29644 30874 29696 30880
rect 29748 27674 29776 38762
rect 33060 38554 33088 38898
rect 34934 38652 35242 38661
rect 34934 38650 34940 38652
rect 34996 38650 35020 38652
rect 35076 38650 35100 38652
rect 35156 38650 35180 38652
rect 35236 38650 35242 38652
rect 34996 38598 34998 38650
rect 35178 38598 35180 38650
rect 34934 38596 34940 38598
rect 34996 38596 35020 38598
rect 35076 38596 35100 38598
rect 35156 38596 35180 38598
rect 35236 38596 35242 38598
rect 34934 38587 35242 38596
rect 35636 38554 35664 38898
rect 37646 38856 37702 38865
rect 37646 38791 37648 38800
rect 37700 38791 37702 38800
rect 37922 38856 37978 38865
rect 37922 38791 37978 38800
rect 37648 38762 37700 38768
rect 37936 38554 37964 38791
rect 33048 38548 33100 38554
rect 33048 38490 33100 38496
rect 35624 38548 35676 38554
rect 35624 38490 35676 38496
rect 37924 38548 37976 38554
rect 37924 38490 37976 38496
rect 31668 38276 31720 38282
rect 31668 38218 31720 38224
rect 30380 38208 30432 38214
rect 30380 38150 30432 38156
rect 31116 38208 31168 38214
rect 31116 38150 31168 38156
rect 30392 37942 30420 38150
rect 30380 37936 30432 37942
rect 30380 37878 30432 37884
rect 30392 37210 30420 37878
rect 30932 37664 30984 37670
rect 30932 37606 30984 37612
rect 30944 37330 30972 37606
rect 30932 37324 30984 37330
rect 30932 37266 30984 37272
rect 30392 37194 30512 37210
rect 30104 37188 30156 37194
rect 30392 37188 30524 37194
rect 30392 37182 30472 37188
rect 30104 37130 30156 37136
rect 30472 37130 30524 37136
rect 30012 37120 30064 37126
rect 30012 37062 30064 37068
rect 30024 36922 30052 37062
rect 30012 36916 30064 36922
rect 30012 36858 30064 36864
rect 29828 36304 29880 36310
rect 29828 36246 29880 36252
rect 29840 35698 29868 36246
rect 30024 36174 30052 36858
rect 30116 36718 30144 37130
rect 30104 36712 30156 36718
rect 30104 36654 30156 36660
rect 30116 36378 30144 36654
rect 30104 36372 30156 36378
rect 30104 36314 30156 36320
rect 30012 36168 30064 36174
rect 30012 36110 30064 36116
rect 30024 35698 30052 36110
rect 30748 36032 30800 36038
rect 30748 35974 30800 35980
rect 30760 35834 30788 35974
rect 30748 35828 30800 35834
rect 30748 35770 30800 35776
rect 30472 35760 30524 35766
rect 30472 35702 30524 35708
rect 29828 35692 29880 35698
rect 29828 35634 29880 35640
rect 30012 35692 30064 35698
rect 30012 35634 30064 35640
rect 30196 35692 30248 35698
rect 30196 35634 30248 35640
rect 29840 33930 29868 35634
rect 30104 35488 30156 35494
rect 30104 35430 30156 35436
rect 30012 34400 30064 34406
rect 30012 34342 30064 34348
rect 30024 33998 30052 34342
rect 30012 33992 30064 33998
rect 30012 33934 30064 33940
rect 29828 33924 29880 33930
rect 29828 33866 29880 33872
rect 29840 31822 29868 33866
rect 30012 33108 30064 33114
rect 30012 33050 30064 33056
rect 29828 31816 29880 31822
rect 29828 31758 29880 31764
rect 29840 30190 29868 31758
rect 30024 31686 30052 33050
rect 30012 31680 30064 31686
rect 30012 31622 30064 31628
rect 30116 30682 30144 35430
rect 30208 35290 30236 35634
rect 30196 35284 30248 35290
rect 30196 35226 30248 35232
rect 30380 35080 30432 35086
rect 30380 35022 30432 35028
rect 30196 34468 30248 34474
rect 30196 34410 30248 34416
rect 30208 33318 30236 34410
rect 30196 33312 30248 33318
rect 30196 33254 30248 33260
rect 30196 32768 30248 32774
rect 30196 32710 30248 32716
rect 30288 32768 30340 32774
rect 30288 32710 30340 32716
rect 30208 30705 30236 32710
rect 30300 32026 30328 32710
rect 30288 32020 30340 32026
rect 30288 31962 30340 31968
rect 30300 31890 30328 31962
rect 30288 31884 30340 31890
rect 30288 31826 30340 31832
rect 30024 30654 30144 30682
rect 30194 30696 30250 30705
rect 29828 30184 29880 30190
rect 29828 30126 29880 30132
rect 30024 29646 30052 30654
rect 30194 30631 30250 30640
rect 30300 30122 30328 31826
rect 30392 31754 30420 35022
rect 30484 33998 30512 35702
rect 31024 35488 31076 35494
rect 31024 35430 31076 35436
rect 30656 35284 30708 35290
rect 30656 35226 30708 35232
rect 30564 34400 30616 34406
rect 30564 34342 30616 34348
rect 30576 33998 30604 34342
rect 30668 34048 30696 35226
rect 31036 35154 31064 35430
rect 31024 35148 31076 35154
rect 31024 35090 31076 35096
rect 30932 34604 30984 34610
rect 30932 34546 30984 34552
rect 30944 34134 30972 34546
rect 30932 34128 30984 34134
rect 30932 34070 30984 34076
rect 30748 34060 30800 34066
rect 30668 34020 30748 34048
rect 30748 34002 30800 34008
rect 30472 33992 30524 33998
rect 30472 33934 30524 33940
rect 30564 33992 30616 33998
rect 30564 33934 30616 33940
rect 30484 33114 30512 33934
rect 30472 33108 30524 33114
rect 30472 33050 30524 33056
rect 30656 33040 30708 33046
rect 30656 32982 30708 32988
rect 30668 32366 30696 32982
rect 30656 32360 30708 32366
rect 30656 32302 30708 32308
rect 30392 31726 30512 31754
rect 30380 31680 30432 31686
rect 30380 31622 30432 31628
rect 30392 31142 30420 31622
rect 30380 31136 30432 31142
rect 30380 31078 30432 31084
rect 30380 30660 30432 30666
rect 30380 30602 30432 30608
rect 30392 30161 30420 30602
rect 30378 30152 30434 30161
rect 30288 30116 30340 30122
rect 30378 30087 30434 30096
rect 30288 30058 30340 30064
rect 29828 29640 29880 29646
rect 29826 29608 29828 29617
rect 30012 29640 30064 29646
rect 29880 29608 29882 29617
rect 30012 29582 30064 29588
rect 29826 29543 29882 29552
rect 30104 29572 30156 29578
rect 30104 29514 30156 29520
rect 29828 29300 29880 29306
rect 29828 29242 29880 29248
rect 29736 27668 29788 27674
rect 29736 27610 29788 27616
rect 29840 27418 29868 29242
rect 30012 29096 30064 29102
rect 30012 29038 30064 29044
rect 30024 28626 30052 29038
rect 30116 28966 30144 29514
rect 30288 29504 30340 29510
rect 30288 29446 30340 29452
rect 30380 29504 30432 29510
rect 30380 29446 30432 29452
rect 30300 29306 30328 29446
rect 30288 29300 30340 29306
rect 30288 29242 30340 29248
rect 30104 28960 30156 28966
rect 30104 28902 30156 28908
rect 30012 28620 30064 28626
rect 30012 28562 30064 28568
rect 30288 28620 30340 28626
rect 30288 28562 30340 28568
rect 30196 28416 30248 28422
rect 30196 28358 30248 28364
rect 30208 28014 30236 28358
rect 30196 28008 30248 28014
rect 29918 27976 29974 27985
rect 30196 27950 30248 27956
rect 29918 27911 29974 27920
rect 29748 27390 29868 27418
rect 29644 27328 29696 27334
rect 29644 27270 29696 27276
rect 29656 27130 29684 27270
rect 29644 27124 29696 27130
rect 29644 27066 29696 27072
rect 29748 25294 29776 27390
rect 29828 27328 29880 27334
rect 29828 27270 29880 27276
rect 29840 27130 29868 27270
rect 29828 27124 29880 27130
rect 29828 27066 29880 27072
rect 29736 25288 29788 25294
rect 29736 25230 29788 25236
rect 29748 24936 29776 25230
rect 29828 24948 29880 24954
rect 29748 24908 29828 24936
rect 29748 24206 29776 24908
rect 29828 24890 29880 24896
rect 29932 24206 29960 27911
rect 30012 27464 30064 27470
rect 30012 27406 30064 27412
rect 30024 26586 30052 27406
rect 30104 27328 30156 27334
rect 30104 27270 30156 27276
rect 30116 26790 30144 27270
rect 30104 26784 30156 26790
rect 30104 26726 30156 26732
rect 30012 26580 30064 26586
rect 30012 26522 30064 26528
rect 30116 26382 30144 26726
rect 30104 26376 30156 26382
rect 30104 26318 30156 26324
rect 30012 26240 30064 26246
rect 30012 26182 30064 26188
rect 30024 25974 30052 26182
rect 30012 25968 30064 25974
rect 30012 25910 30064 25916
rect 30208 24750 30236 27950
rect 30300 26450 30328 28562
rect 30392 28558 30420 29446
rect 30380 28552 30432 28558
rect 30380 28494 30432 28500
rect 30392 27470 30420 28494
rect 30380 27464 30432 27470
rect 30380 27406 30432 27412
rect 30484 26450 30512 31726
rect 30668 30938 30696 32302
rect 30760 31822 30788 34002
rect 30932 32904 30984 32910
rect 30932 32846 30984 32852
rect 30944 32434 30972 32846
rect 30840 32428 30892 32434
rect 30840 32370 30892 32376
rect 30932 32428 30984 32434
rect 30932 32370 30984 32376
rect 30748 31816 30800 31822
rect 30748 31758 30800 31764
rect 30656 30932 30708 30938
rect 30656 30874 30708 30880
rect 30656 30320 30708 30326
rect 30656 30262 30708 30268
rect 30564 30184 30616 30190
rect 30564 30126 30616 30132
rect 30576 29578 30604 30126
rect 30668 29646 30696 30262
rect 30656 29640 30708 29646
rect 30760 29628 30788 31758
rect 30852 31754 30880 32370
rect 31128 31754 31156 38150
rect 31208 37868 31260 37874
rect 31208 37810 31260 37816
rect 31220 36922 31248 37810
rect 31680 37806 31708 38218
rect 35594 38108 35902 38117
rect 35594 38106 35600 38108
rect 35656 38106 35680 38108
rect 35736 38106 35760 38108
rect 35816 38106 35840 38108
rect 35896 38106 35902 38108
rect 35656 38054 35658 38106
rect 35838 38054 35840 38106
rect 35594 38052 35600 38054
rect 35656 38052 35680 38054
rect 35736 38052 35760 38054
rect 35816 38052 35840 38054
rect 35896 38052 35902 38054
rect 35594 38043 35902 38052
rect 31668 37800 31720 37806
rect 31668 37742 31720 37748
rect 34934 37564 35242 37573
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37499 35242 37508
rect 32588 37256 32640 37262
rect 32588 37198 32640 37204
rect 31484 37188 31536 37194
rect 31484 37130 31536 37136
rect 31496 36922 31524 37130
rect 32496 37120 32548 37126
rect 32496 37062 32548 37068
rect 32508 36922 32536 37062
rect 31208 36916 31260 36922
rect 31208 36858 31260 36864
rect 31484 36916 31536 36922
rect 31484 36858 31536 36864
rect 32496 36916 32548 36922
rect 32496 36858 32548 36864
rect 32220 36712 32272 36718
rect 32220 36654 32272 36660
rect 32232 36378 32260 36654
rect 32220 36372 32272 36378
rect 32220 36314 32272 36320
rect 32404 36236 32456 36242
rect 32404 36178 32456 36184
rect 31852 36100 31904 36106
rect 31852 36042 31904 36048
rect 31392 35692 31444 35698
rect 31392 35634 31444 35640
rect 31404 34746 31432 35634
rect 31484 35624 31536 35630
rect 31484 35566 31536 35572
rect 31392 34740 31444 34746
rect 31392 34682 31444 34688
rect 31496 33998 31524 35566
rect 31864 35034 31892 36042
rect 32312 35216 32364 35222
rect 32312 35158 32364 35164
rect 31680 35006 31892 35034
rect 31680 34950 31708 35006
rect 31668 34944 31720 34950
rect 31668 34886 31720 34892
rect 31760 34944 31812 34950
rect 31760 34886 31812 34892
rect 31772 34678 31800 34886
rect 31760 34672 31812 34678
rect 31760 34614 31812 34620
rect 31484 33992 31536 33998
rect 31484 33934 31536 33940
rect 31208 32904 31260 32910
rect 31208 32846 31260 32852
rect 31220 32570 31248 32846
rect 31208 32564 31260 32570
rect 31208 32506 31260 32512
rect 31496 31822 31524 33934
rect 31576 33856 31628 33862
rect 31772 33844 31800 34614
rect 31864 34542 31892 35006
rect 31852 34536 31904 34542
rect 31852 34478 31904 34484
rect 31628 33816 31800 33844
rect 31576 33798 31628 33804
rect 31588 33658 31616 33798
rect 31576 33652 31628 33658
rect 31576 33594 31628 33600
rect 31864 33114 31892 34478
rect 32220 33856 32272 33862
rect 32220 33798 32272 33804
rect 31852 33108 31904 33114
rect 31852 33050 31904 33056
rect 31852 32768 31904 32774
rect 31852 32710 31904 32716
rect 31864 32298 31892 32710
rect 32048 32434 32168 32450
rect 32232 32434 32260 33798
rect 32324 33522 32352 35158
rect 32416 34542 32444 36178
rect 32600 35766 32628 37198
rect 37832 37120 37884 37126
rect 37832 37062 37884 37068
rect 35594 37020 35902 37029
rect 35594 37018 35600 37020
rect 35656 37018 35680 37020
rect 35736 37018 35760 37020
rect 35816 37018 35840 37020
rect 35896 37018 35902 37020
rect 35656 36966 35658 37018
rect 35838 36966 35840 37018
rect 35594 36964 35600 36966
rect 35656 36964 35680 36966
rect 35736 36964 35760 36966
rect 35816 36964 35840 36966
rect 35896 36964 35902 36966
rect 35594 36955 35902 36964
rect 37844 36825 37872 37062
rect 37830 36816 37886 36825
rect 33692 36780 33744 36786
rect 37830 36751 37886 36760
rect 33692 36722 33744 36728
rect 33140 36576 33192 36582
rect 33140 36518 33192 36524
rect 33152 36038 33180 36518
rect 33140 36032 33192 36038
rect 33140 35974 33192 35980
rect 33600 36032 33652 36038
rect 33600 35974 33652 35980
rect 32588 35760 32640 35766
rect 32588 35702 32640 35708
rect 32496 35012 32548 35018
rect 32496 34954 32548 34960
rect 32404 34536 32456 34542
rect 32404 34478 32456 34484
rect 32312 33516 32364 33522
rect 32312 33458 32364 33464
rect 32508 32910 32536 34954
rect 32496 32904 32548 32910
rect 32496 32846 32548 32852
rect 32600 32502 32628 35702
rect 33508 35692 33560 35698
rect 33508 35634 33560 35640
rect 32772 35488 32824 35494
rect 32772 35430 32824 35436
rect 33324 35488 33376 35494
rect 33324 35430 33376 35436
rect 32784 35290 32812 35430
rect 32772 35284 32824 35290
rect 32772 35226 32824 35232
rect 33336 35154 33364 35430
rect 33324 35148 33376 35154
rect 33324 35090 33376 35096
rect 33416 35148 33468 35154
rect 33416 35090 33468 35096
rect 33428 35018 33456 35090
rect 33416 35012 33468 35018
rect 33416 34954 33468 34960
rect 33324 34944 33376 34950
rect 33324 34886 33376 34892
rect 33336 34746 33364 34886
rect 33520 34746 33548 35634
rect 33324 34740 33376 34746
rect 33508 34740 33560 34746
rect 33376 34700 33456 34728
rect 33324 34682 33376 34688
rect 33324 34400 33376 34406
rect 33324 34342 33376 34348
rect 33232 33652 33284 33658
rect 33232 33594 33284 33600
rect 32956 32904 33008 32910
rect 32956 32846 33008 32852
rect 32588 32496 32640 32502
rect 32588 32438 32640 32444
rect 32048 32428 32180 32434
rect 32048 32422 32128 32428
rect 31852 32292 31904 32298
rect 31852 32234 31904 32240
rect 31864 32026 31892 32234
rect 31852 32020 31904 32026
rect 31852 31962 31904 31968
rect 31484 31816 31536 31822
rect 31484 31758 31536 31764
rect 31944 31816 31996 31822
rect 31944 31758 31996 31764
rect 30852 31726 31064 31754
rect 31128 31726 31248 31754
rect 30932 30660 30984 30666
rect 30932 30602 30984 30608
rect 30840 29640 30892 29646
rect 30760 29600 30840 29628
rect 30656 29582 30708 29588
rect 30840 29582 30892 29588
rect 30564 29572 30616 29578
rect 30564 29514 30616 29520
rect 30576 29209 30604 29514
rect 30562 29200 30618 29209
rect 30562 29135 30618 29144
rect 30576 28558 30604 29135
rect 30852 28558 30880 29582
rect 30564 28552 30616 28558
rect 30564 28494 30616 28500
rect 30748 28552 30800 28558
rect 30748 28494 30800 28500
rect 30840 28552 30892 28558
rect 30840 28494 30892 28500
rect 30576 27470 30604 28494
rect 30760 28218 30788 28494
rect 30748 28212 30800 28218
rect 30748 28154 30800 28160
rect 30852 27470 30880 28494
rect 30564 27464 30616 27470
rect 30564 27406 30616 27412
rect 30840 27464 30892 27470
rect 30840 27406 30892 27412
rect 30288 26444 30340 26450
rect 30288 26386 30340 26392
rect 30472 26444 30524 26450
rect 30472 26386 30524 26392
rect 30484 26353 30512 26386
rect 30470 26344 30526 26353
rect 30470 26279 30526 26288
rect 30288 26240 30340 26246
rect 30288 26182 30340 26188
rect 30300 25294 30328 26182
rect 30576 25430 30604 27406
rect 30748 27328 30800 27334
rect 30748 27270 30800 27276
rect 30760 26518 30788 27270
rect 30944 26897 30972 30602
rect 31036 30598 31064 31726
rect 31116 30728 31168 30734
rect 31116 30670 31168 30676
rect 31024 30592 31076 30598
rect 31024 30534 31076 30540
rect 31128 30326 31156 30670
rect 31116 30320 31168 30326
rect 31116 30262 31168 30268
rect 31116 30116 31168 30122
rect 31116 30058 31168 30064
rect 31128 29238 31156 30058
rect 31116 29232 31168 29238
rect 31116 29174 31168 29180
rect 31116 28416 31168 28422
rect 31116 28358 31168 28364
rect 31024 27464 31076 27470
rect 31024 27406 31076 27412
rect 30930 26888 30986 26897
rect 30930 26823 30986 26832
rect 30748 26512 30800 26518
rect 30748 26454 30800 26460
rect 31036 25498 31064 27406
rect 31024 25492 31076 25498
rect 31024 25434 31076 25440
rect 30564 25424 30616 25430
rect 30564 25366 30616 25372
rect 30288 25288 30340 25294
rect 30288 25230 30340 25236
rect 30380 25288 30432 25294
rect 30380 25230 30432 25236
rect 30196 24744 30248 24750
rect 30196 24686 30248 24692
rect 30300 24274 30328 25230
rect 30392 24868 30420 25230
rect 30656 25152 30708 25158
rect 30656 25094 30708 25100
rect 30472 24880 30524 24886
rect 30392 24840 30472 24868
rect 30392 24342 30420 24840
rect 30472 24822 30524 24828
rect 30380 24336 30432 24342
rect 30380 24278 30432 24284
rect 30288 24268 30340 24274
rect 30288 24210 30340 24216
rect 29552 24200 29604 24206
rect 29552 24142 29604 24148
rect 29736 24200 29788 24206
rect 29736 24142 29788 24148
rect 29828 24200 29880 24206
rect 29828 24142 29880 24148
rect 29920 24200 29972 24206
rect 29920 24142 29972 24148
rect 29840 24070 29868 24142
rect 29828 24064 29880 24070
rect 29828 24006 29880 24012
rect 30196 24064 30248 24070
rect 30196 24006 30248 24012
rect 29736 23112 29788 23118
rect 29736 23054 29788 23060
rect 29920 23112 29972 23118
rect 29920 23054 29972 23060
rect 29748 22438 29776 23054
rect 29932 22778 29960 23054
rect 30012 23044 30064 23050
rect 30012 22986 30064 22992
rect 29920 22772 29972 22778
rect 29920 22714 29972 22720
rect 29736 22432 29788 22438
rect 29736 22374 29788 22380
rect 28736 22066 28856 22094
rect 29012 22066 29408 22094
rect 28540 21888 28592 21894
rect 28540 21830 28592 21836
rect 28448 21616 28500 21622
rect 28448 21558 28500 21564
rect 28540 20460 28592 20466
rect 28540 20402 28592 20408
rect 28552 19922 28580 20402
rect 28540 19916 28592 19922
rect 28540 19858 28592 19864
rect 28736 19514 28764 22066
rect 28816 22024 28868 22030
rect 28816 21966 28868 21972
rect 28828 21418 28856 21966
rect 28816 21412 28868 21418
rect 28816 21354 28868 21360
rect 29012 20466 29040 22066
rect 29748 21622 29776 22374
rect 30024 22098 30052 22986
rect 30208 22642 30236 24006
rect 30472 23316 30524 23322
rect 30472 23258 30524 23264
rect 30196 22636 30248 22642
rect 30196 22578 30248 22584
rect 30012 22092 30064 22098
rect 30012 22034 30064 22040
rect 29828 22024 29880 22030
rect 30024 21978 30052 22034
rect 29880 21972 29960 21978
rect 29828 21966 29960 21972
rect 29840 21950 29960 21966
rect 30024 21950 30144 21978
rect 29828 21888 29880 21894
rect 29828 21830 29880 21836
rect 29736 21616 29788 21622
rect 29736 21558 29788 21564
rect 29644 21344 29696 21350
rect 29644 21286 29696 21292
rect 29368 20936 29420 20942
rect 29368 20878 29420 20884
rect 29000 20460 29052 20466
rect 29000 20402 29052 20408
rect 29012 19938 29040 20402
rect 28920 19922 29132 19938
rect 28920 19916 29144 19922
rect 28920 19910 29092 19916
rect 28920 19854 28948 19910
rect 29092 19858 29144 19864
rect 28908 19848 28960 19854
rect 28908 19790 28960 19796
rect 29276 19780 29328 19786
rect 29276 19722 29328 19728
rect 28724 19508 28776 19514
rect 28724 19450 28776 19456
rect 29288 19378 29316 19722
rect 29276 19372 29328 19378
rect 29276 19314 29328 19320
rect 28356 18624 28408 18630
rect 28356 18566 28408 18572
rect 29380 18290 29408 20878
rect 29656 20398 29684 21286
rect 29840 20874 29868 21830
rect 29828 20868 29880 20874
rect 29828 20810 29880 20816
rect 29644 20392 29696 20398
rect 29644 20334 29696 20340
rect 29552 20256 29604 20262
rect 29552 20198 29604 20204
rect 29564 19922 29592 20198
rect 29552 19916 29604 19922
rect 29552 19858 29604 19864
rect 29656 19854 29684 20334
rect 29932 19961 29960 21950
rect 30116 21622 30144 21950
rect 30104 21616 30156 21622
rect 30104 21558 30156 21564
rect 30484 21010 30512 23258
rect 30668 22692 30696 25094
rect 31128 24818 31156 28358
rect 31116 24812 31168 24818
rect 31116 24754 31168 24760
rect 31220 24698 31248 31726
rect 31300 30592 31352 30598
rect 31300 30534 31352 30540
rect 31312 30258 31340 30534
rect 31300 30252 31352 30258
rect 31300 30194 31352 30200
rect 31312 29646 31340 30194
rect 31300 29640 31352 29646
rect 31300 29582 31352 29588
rect 31300 29504 31352 29510
rect 31300 29446 31352 29452
rect 31312 29306 31340 29446
rect 31300 29300 31352 29306
rect 31300 29242 31352 29248
rect 31496 29238 31524 31758
rect 31668 31340 31720 31346
rect 31668 31282 31720 31288
rect 31680 30734 31708 31282
rect 31760 31136 31812 31142
rect 31760 31078 31812 31084
rect 31668 30728 31720 30734
rect 31668 30670 31720 30676
rect 31576 30660 31628 30666
rect 31576 30602 31628 30608
rect 31588 29238 31616 30602
rect 31484 29232 31536 29238
rect 31484 29174 31536 29180
rect 31576 29232 31628 29238
rect 31576 29174 31628 29180
rect 31496 28694 31524 29174
rect 31668 29028 31720 29034
rect 31668 28970 31720 28976
rect 31772 28994 31800 31078
rect 31956 30954 31984 31758
rect 32048 31142 32076 32422
rect 32128 32370 32180 32376
rect 32220 32428 32272 32434
rect 32220 32370 32272 32376
rect 32312 32360 32364 32366
rect 32312 32302 32364 32308
rect 32128 32292 32180 32298
rect 32128 32234 32180 32240
rect 32140 31754 32168 32234
rect 32140 31726 32260 31754
rect 32036 31136 32088 31142
rect 32036 31078 32088 31084
rect 31956 30926 32168 30954
rect 32140 30258 32168 30926
rect 32128 30252 32180 30258
rect 32128 30194 32180 30200
rect 31484 28688 31536 28694
rect 31390 28656 31446 28665
rect 31484 28630 31536 28636
rect 31390 28591 31446 28600
rect 31404 28558 31432 28591
rect 31392 28552 31444 28558
rect 31392 28494 31444 28500
rect 31576 27124 31628 27130
rect 31576 27066 31628 27072
rect 31392 26784 31444 26790
rect 31392 26726 31444 26732
rect 31404 26450 31432 26726
rect 31392 26444 31444 26450
rect 31392 26386 31444 26392
rect 31588 26314 31616 27066
rect 31576 26308 31628 26314
rect 31576 26250 31628 26256
rect 31680 26246 31708 28970
rect 31772 28966 31892 28994
rect 31760 28552 31812 28558
rect 31760 28494 31812 28500
rect 31772 28218 31800 28494
rect 31760 28212 31812 28218
rect 31760 28154 31812 28160
rect 31864 28082 31892 28966
rect 31852 28076 31904 28082
rect 31852 28018 31904 28024
rect 31944 28076 31996 28082
rect 31944 28018 31996 28024
rect 31852 27600 31904 27606
rect 31852 27542 31904 27548
rect 31760 27328 31812 27334
rect 31760 27270 31812 27276
rect 31668 26240 31720 26246
rect 31668 26182 31720 26188
rect 31772 25906 31800 27270
rect 31864 26450 31892 27542
rect 31956 27470 31984 28018
rect 31944 27464 31996 27470
rect 31944 27406 31996 27412
rect 32128 26988 32180 26994
rect 32128 26930 32180 26936
rect 31852 26444 31904 26450
rect 31852 26386 31904 26392
rect 31760 25900 31812 25906
rect 31760 25842 31812 25848
rect 31864 25838 31892 26386
rect 32140 26042 32168 26930
rect 32036 26036 32088 26042
rect 32036 25978 32088 25984
rect 32128 26036 32180 26042
rect 32128 25978 32180 25984
rect 31852 25832 31904 25838
rect 31852 25774 31904 25780
rect 32048 25702 32076 25978
rect 31300 25696 31352 25702
rect 31300 25638 31352 25644
rect 32036 25696 32088 25702
rect 32036 25638 32088 25644
rect 31312 24954 31340 25638
rect 31392 25152 31444 25158
rect 31392 25094 31444 25100
rect 31404 24954 31432 25094
rect 31300 24948 31352 24954
rect 31300 24890 31352 24896
rect 31392 24948 31444 24954
rect 31392 24890 31444 24896
rect 31576 24812 31628 24818
rect 31576 24754 31628 24760
rect 31128 24670 31248 24698
rect 30668 22664 30880 22692
rect 30656 22432 30708 22438
rect 30656 22374 30708 22380
rect 30564 22092 30616 22098
rect 30564 22034 30616 22040
rect 30576 21554 30604 22034
rect 30564 21548 30616 21554
rect 30564 21490 30616 21496
rect 30668 21010 30696 22374
rect 30472 21004 30524 21010
rect 30472 20946 30524 20952
rect 30656 21004 30708 21010
rect 30656 20946 30708 20952
rect 30380 20936 30432 20942
rect 30380 20878 30432 20884
rect 30104 20800 30156 20806
rect 30104 20742 30156 20748
rect 30288 20800 30340 20806
rect 30288 20742 30340 20748
rect 29918 19952 29974 19961
rect 29918 19887 29974 19896
rect 29644 19848 29696 19854
rect 29644 19790 29696 19796
rect 29828 19848 29880 19854
rect 29828 19790 29880 19796
rect 29552 19712 29604 19718
rect 29552 19654 29604 19660
rect 29736 19712 29788 19718
rect 29736 19654 29788 19660
rect 29564 19514 29592 19654
rect 29748 19514 29776 19654
rect 29840 19514 29868 19790
rect 29552 19508 29604 19514
rect 29552 19450 29604 19456
rect 29736 19508 29788 19514
rect 29736 19450 29788 19456
rect 29828 19508 29880 19514
rect 29828 19450 29880 19456
rect 29932 19394 29960 19887
rect 30116 19718 30144 20742
rect 30300 19854 30328 20742
rect 30392 20466 30420 20878
rect 30668 20466 30696 20946
rect 30380 20460 30432 20466
rect 30380 20402 30432 20408
rect 30656 20460 30708 20466
rect 30656 20402 30708 20408
rect 30288 19848 30340 19854
rect 30288 19790 30340 19796
rect 30104 19712 30156 19718
rect 30104 19654 30156 19660
rect 29460 19372 29512 19378
rect 29460 19314 29512 19320
rect 29840 19366 29960 19394
rect 28632 18284 28684 18290
rect 28632 18226 28684 18232
rect 29368 18284 29420 18290
rect 29368 18226 29420 18232
rect 28448 18148 28500 18154
rect 28448 18090 28500 18096
rect 27896 17672 27948 17678
rect 27896 17614 27948 17620
rect 28172 17672 28224 17678
rect 28172 17614 28224 17620
rect 28356 17672 28408 17678
rect 28356 17614 28408 17620
rect 28264 17604 28316 17610
rect 28264 17546 28316 17552
rect 28276 17338 28304 17546
rect 28368 17338 28396 17614
rect 28264 17332 28316 17338
rect 28264 17274 28316 17280
rect 28356 17332 28408 17338
rect 28356 17274 28408 17280
rect 27804 17196 27856 17202
rect 27804 17138 27856 17144
rect 27816 16794 27844 17138
rect 27804 16788 27856 16794
rect 27804 16730 27856 16736
rect 27620 15496 27672 15502
rect 27620 15438 27672 15444
rect 27632 13938 27660 15438
rect 28356 15360 28408 15366
rect 28356 15302 28408 15308
rect 27724 15162 28028 15178
rect 27712 15156 28028 15162
rect 27764 15150 28028 15156
rect 27712 15098 27764 15104
rect 28000 15094 28028 15150
rect 27988 15088 28040 15094
rect 27988 15030 28040 15036
rect 27896 15020 27948 15026
rect 27896 14962 27948 14968
rect 27804 14000 27856 14006
rect 27804 13942 27856 13948
rect 27620 13932 27672 13938
rect 27620 13874 27672 13880
rect 27816 13530 27844 13942
rect 27908 13530 27936 14962
rect 28368 14618 28396 15302
rect 28356 14612 28408 14618
rect 28356 14554 28408 14560
rect 28460 13530 28488 18090
rect 28644 17678 28672 18226
rect 29472 18086 29500 19314
rect 29644 19168 29696 19174
rect 29644 19110 29696 19116
rect 29550 18320 29606 18329
rect 29550 18255 29552 18264
rect 29604 18255 29606 18264
rect 29552 18226 29604 18232
rect 29460 18080 29512 18086
rect 29460 18022 29512 18028
rect 28632 17672 28684 17678
rect 28632 17614 28684 17620
rect 29184 17536 29236 17542
rect 29184 17478 29236 17484
rect 29196 17338 29224 17478
rect 29184 17332 29236 17338
rect 29184 17274 29236 17280
rect 28632 17264 28684 17270
rect 28632 17206 28684 17212
rect 28540 14884 28592 14890
rect 28540 14826 28592 14832
rect 28552 14074 28580 14826
rect 28540 14068 28592 14074
rect 28540 14010 28592 14016
rect 28540 13728 28592 13734
rect 28540 13670 28592 13676
rect 27804 13524 27856 13530
rect 27804 13466 27856 13472
rect 27896 13524 27948 13530
rect 27896 13466 27948 13472
rect 28172 13524 28224 13530
rect 28172 13466 28224 13472
rect 28448 13524 28500 13530
rect 28448 13466 28500 13472
rect 27618 13424 27674 13433
rect 27618 13359 27674 13368
rect 27436 13320 27488 13326
rect 27158 13288 27214 13297
rect 27214 13246 27292 13274
rect 27436 13262 27488 13268
rect 27158 13223 27214 13232
rect 27160 12640 27212 12646
rect 27160 12582 27212 12588
rect 27068 11144 27120 11150
rect 27068 11086 27120 11092
rect 27172 11082 27200 12582
rect 27160 11076 27212 11082
rect 27160 11018 27212 11024
rect 27172 9586 27200 11018
rect 27264 10674 27292 13246
rect 27632 11898 27660 13359
rect 27804 12368 27856 12374
rect 27804 12310 27856 12316
rect 27620 11892 27672 11898
rect 27620 11834 27672 11840
rect 27344 11756 27396 11762
rect 27344 11698 27396 11704
rect 27356 11354 27384 11698
rect 27528 11620 27580 11626
rect 27528 11562 27580 11568
rect 27344 11348 27396 11354
rect 27344 11290 27396 11296
rect 27540 10674 27568 11562
rect 27632 11354 27660 11834
rect 27816 11830 27844 12310
rect 28184 12102 28212 13466
rect 28264 13456 28316 13462
rect 28264 13398 28316 13404
rect 28172 12096 28224 12102
rect 28172 12038 28224 12044
rect 27804 11824 27856 11830
rect 27988 11824 28040 11830
rect 27856 11784 27936 11812
rect 27804 11766 27856 11772
rect 27710 11656 27766 11665
rect 27710 11591 27766 11600
rect 27724 11558 27752 11591
rect 27712 11552 27764 11558
rect 27712 11494 27764 11500
rect 27620 11348 27672 11354
rect 27620 11290 27672 11296
rect 27724 11286 27752 11494
rect 27712 11280 27764 11286
rect 27712 11222 27764 11228
rect 27724 11132 27752 11222
rect 27908 11150 27936 11784
rect 27988 11766 28040 11772
rect 27804 11144 27856 11150
rect 27724 11104 27804 11132
rect 27804 11086 27856 11092
rect 27896 11144 27948 11150
rect 27896 11086 27948 11092
rect 27620 11008 27672 11014
rect 27620 10950 27672 10956
rect 27632 10810 27660 10950
rect 27620 10804 27672 10810
rect 27620 10746 27672 10752
rect 27252 10668 27304 10674
rect 27252 10610 27304 10616
rect 27528 10668 27580 10674
rect 27528 10610 27580 10616
rect 27620 10464 27672 10470
rect 27620 10406 27672 10412
rect 27252 10260 27304 10266
rect 27252 10202 27304 10208
rect 26516 9376 26568 9382
rect 26516 9318 26568 9324
rect 26528 8974 26556 9318
rect 26516 8968 26568 8974
rect 26516 8910 26568 8916
rect 26516 8832 26568 8838
rect 26516 8774 26568 8780
rect 26528 8498 26556 8774
rect 26516 8492 26568 8498
rect 26516 8434 26568 8440
rect 26424 7540 26476 7546
rect 26424 7482 26476 7488
rect 26608 7540 26660 7546
rect 26608 7482 26660 7488
rect 26240 7472 26292 7478
rect 26240 7414 26292 7420
rect 26332 7472 26384 7478
rect 26332 7414 26384 7420
rect 25964 7336 26016 7342
rect 25964 7278 26016 7284
rect 26620 6866 26648 7482
rect 26608 6860 26660 6866
rect 26608 6802 26660 6808
rect 26056 6792 26108 6798
rect 26056 6734 26108 6740
rect 26240 6792 26292 6798
rect 26240 6734 26292 6740
rect 26068 6322 26096 6734
rect 26056 6316 26108 6322
rect 26056 6258 26108 6264
rect 26068 5098 26096 6258
rect 26252 5234 26280 6734
rect 26712 6662 26740 9574
rect 26976 9580 27028 9586
rect 26976 9522 27028 9528
rect 27160 9580 27212 9586
rect 27160 9522 27212 9528
rect 26896 9166 27108 9194
rect 26896 9042 26924 9166
rect 27080 9110 27108 9166
rect 26976 9104 27028 9110
rect 26976 9046 27028 9052
rect 27068 9104 27120 9110
rect 27068 9046 27120 9052
rect 26884 9036 26936 9042
rect 26884 8978 26936 8984
rect 26884 8900 26936 8906
rect 26884 8842 26936 8848
rect 26896 8566 26924 8842
rect 26988 8820 27016 9046
rect 27264 8974 27292 10202
rect 27632 10130 27660 10406
rect 27908 10266 27936 11086
rect 28000 10577 28028 11766
rect 28184 10674 28212 12038
rect 28276 10674 28304 13398
rect 28552 13326 28580 13670
rect 28356 13320 28408 13326
rect 28356 13262 28408 13268
rect 28540 13320 28592 13326
rect 28540 13262 28592 13268
rect 28172 10668 28224 10674
rect 28172 10610 28224 10616
rect 28264 10668 28316 10674
rect 28264 10610 28316 10616
rect 27986 10568 28042 10577
rect 27986 10503 28042 10512
rect 27896 10260 27948 10266
rect 27896 10202 27948 10208
rect 27620 10124 27672 10130
rect 27620 10066 27672 10072
rect 28276 10062 28304 10610
rect 28368 10441 28396 13262
rect 28448 12776 28500 12782
rect 28448 12718 28500 12724
rect 28460 12434 28488 12718
rect 28460 12406 28580 12434
rect 28552 10538 28580 12406
rect 28540 10532 28592 10538
rect 28540 10474 28592 10480
rect 28354 10432 28410 10441
rect 28354 10367 28410 10376
rect 28264 10056 28316 10062
rect 28264 9998 28316 10004
rect 27896 9920 27948 9926
rect 27896 9862 27948 9868
rect 27344 9580 27396 9586
rect 27344 9522 27396 9528
rect 27436 9580 27488 9586
rect 27436 9522 27488 9528
rect 27528 9580 27580 9586
rect 27528 9522 27580 9528
rect 27712 9580 27764 9586
rect 27712 9522 27764 9528
rect 27252 8968 27304 8974
rect 27252 8910 27304 8916
rect 27160 8832 27212 8838
rect 26988 8792 27160 8820
rect 27160 8774 27212 8780
rect 26884 8560 26936 8566
rect 26884 8502 26936 8508
rect 27356 8498 27384 9522
rect 27448 9450 27476 9522
rect 27436 9444 27488 9450
rect 27436 9386 27488 9392
rect 27540 9382 27568 9522
rect 27528 9376 27580 9382
rect 27528 9318 27580 9324
rect 27618 9072 27674 9081
rect 27618 9007 27674 9016
rect 27632 8974 27660 9007
rect 27620 8968 27672 8974
rect 27620 8910 27672 8916
rect 27724 8906 27752 9522
rect 27712 8900 27764 8906
rect 27712 8842 27764 8848
rect 27344 8492 27396 8498
rect 27344 8434 27396 8440
rect 27436 8492 27488 8498
rect 27620 8492 27672 8498
rect 27436 8434 27488 8440
rect 27540 8452 27620 8480
rect 27448 7546 27476 8434
rect 27436 7540 27488 7546
rect 27436 7482 27488 7488
rect 26976 6792 27028 6798
rect 26976 6734 27028 6740
rect 27436 6792 27488 6798
rect 27540 6780 27568 8452
rect 27620 8434 27672 8440
rect 27724 7546 27752 8842
rect 27804 8356 27856 8362
rect 27804 8298 27856 8304
rect 27620 7540 27672 7546
rect 27620 7482 27672 7488
rect 27712 7540 27764 7546
rect 27712 7482 27764 7488
rect 27488 6752 27568 6780
rect 27436 6734 27488 6740
rect 26700 6656 26752 6662
rect 26700 6598 26752 6604
rect 26240 5228 26292 5234
rect 26240 5170 26292 5176
rect 26988 5166 27016 6734
rect 27528 6248 27580 6254
rect 27528 6190 27580 6196
rect 27540 5846 27568 6190
rect 27632 6118 27660 7482
rect 27816 6866 27844 8298
rect 27804 6860 27856 6866
rect 27804 6802 27856 6808
rect 27804 6316 27856 6322
rect 27804 6258 27856 6264
rect 27712 6248 27764 6254
rect 27712 6190 27764 6196
rect 27620 6112 27672 6118
rect 27724 6100 27752 6190
rect 27672 6072 27752 6100
rect 27620 6054 27672 6060
rect 27528 5840 27580 5846
rect 27528 5782 27580 5788
rect 27632 5370 27660 6054
rect 27816 5914 27844 6258
rect 27804 5908 27856 5914
rect 27804 5850 27856 5856
rect 27620 5364 27672 5370
rect 27620 5306 27672 5312
rect 27620 5228 27672 5234
rect 27620 5170 27672 5176
rect 27712 5228 27764 5234
rect 27712 5170 27764 5176
rect 27804 5228 27856 5234
rect 27908 5216 27936 9862
rect 28080 9376 28132 9382
rect 28080 9318 28132 9324
rect 28092 9042 28120 9318
rect 28080 9036 28132 9042
rect 28080 8978 28132 8984
rect 28080 7268 28132 7274
rect 28080 7210 28132 7216
rect 27988 6792 28040 6798
rect 27988 6734 28040 6740
rect 28000 6458 28028 6734
rect 28092 6730 28120 7210
rect 28172 6792 28224 6798
rect 28172 6734 28224 6740
rect 28264 6792 28316 6798
rect 28264 6734 28316 6740
rect 28080 6724 28132 6730
rect 28080 6666 28132 6672
rect 27988 6452 28040 6458
rect 27988 6394 28040 6400
rect 27856 5188 27936 5216
rect 27804 5170 27856 5176
rect 26976 5160 27028 5166
rect 26976 5102 27028 5108
rect 26056 5092 26108 5098
rect 26056 5034 26108 5040
rect 26068 4826 26096 5034
rect 26056 4820 26108 4826
rect 26056 4762 26108 4768
rect 26988 4690 27016 5102
rect 27632 4826 27660 5170
rect 27620 4820 27672 4826
rect 27620 4762 27672 4768
rect 26976 4684 27028 4690
rect 26976 4626 27028 4632
rect 26332 4616 26384 4622
rect 26332 4558 26384 4564
rect 26344 4282 26372 4558
rect 27724 4486 27752 5170
rect 27816 4758 27844 5170
rect 27804 4752 27856 4758
rect 27804 4694 27856 4700
rect 28092 4690 28120 6666
rect 28184 6458 28212 6734
rect 28172 6452 28224 6458
rect 28172 6394 28224 6400
rect 28276 5166 28304 6734
rect 28368 6662 28396 10367
rect 28448 10260 28500 10266
rect 28448 10202 28500 10208
rect 28460 8974 28488 10202
rect 28448 8968 28500 8974
rect 28448 8910 28500 8916
rect 28460 6866 28488 8910
rect 28552 7954 28580 10474
rect 28540 7948 28592 7954
rect 28540 7890 28592 7896
rect 28540 7404 28592 7410
rect 28540 7346 28592 7352
rect 28552 6866 28580 7346
rect 28644 7342 28672 17206
rect 29184 17196 29236 17202
rect 29184 17138 29236 17144
rect 29196 16794 29224 17138
rect 29368 17060 29420 17066
rect 29368 17002 29420 17008
rect 29184 16788 29236 16794
rect 29184 16730 29236 16736
rect 29380 16522 29408 17002
rect 29368 16516 29420 16522
rect 29368 16458 29420 16464
rect 29184 16040 29236 16046
rect 29184 15982 29236 15988
rect 29196 15570 29224 15982
rect 29184 15564 29236 15570
rect 29184 15506 29236 15512
rect 28816 15020 28868 15026
rect 28816 14962 28868 14968
rect 28724 14952 28776 14958
rect 28722 14920 28724 14929
rect 28776 14920 28778 14929
rect 28828 14890 28856 14962
rect 29472 14958 29500 18022
rect 29656 17202 29684 19110
rect 29736 17672 29788 17678
rect 29736 17614 29788 17620
rect 29644 17196 29696 17202
rect 29644 17138 29696 17144
rect 29552 16108 29604 16114
rect 29552 16050 29604 16056
rect 29644 16108 29696 16114
rect 29644 16050 29696 16056
rect 29564 15570 29592 16050
rect 29552 15564 29604 15570
rect 29552 15506 29604 15512
rect 29656 15502 29684 16050
rect 29644 15496 29696 15502
rect 29644 15438 29696 15444
rect 29460 14952 29512 14958
rect 29460 14894 29512 14900
rect 28722 14855 28778 14864
rect 28816 14884 28868 14890
rect 28816 14826 28868 14832
rect 29184 14544 29236 14550
rect 29184 14486 29236 14492
rect 29196 13938 29224 14486
rect 29276 14068 29328 14074
rect 29276 14010 29328 14016
rect 28816 13932 28868 13938
rect 28816 13874 28868 13880
rect 29184 13932 29236 13938
rect 29184 13874 29236 13880
rect 28828 12288 28856 13874
rect 29000 13864 29052 13870
rect 29000 13806 29052 13812
rect 29012 13530 29040 13806
rect 29000 13524 29052 13530
rect 29000 13466 29052 13472
rect 29184 13524 29236 13530
rect 29184 13466 29236 13472
rect 29000 12708 29052 12714
rect 29000 12650 29052 12656
rect 29092 12708 29144 12714
rect 29092 12650 29144 12656
rect 28908 12300 28960 12306
rect 28828 12260 28908 12288
rect 28828 11762 28856 12260
rect 28908 12242 28960 12248
rect 28908 12096 28960 12102
rect 28906 12064 28908 12073
rect 28960 12064 28962 12073
rect 28906 11999 28962 12008
rect 29012 11762 29040 12650
rect 29104 11898 29132 12650
rect 29092 11892 29144 11898
rect 29092 11834 29144 11840
rect 28816 11756 28868 11762
rect 28816 11698 28868 11704
rect 29000 11756 29052 11762
rect 29000 11698 29052 11704
rect 29092 11552 29144 11558
rect 29092 11494 29144 11500
rect 29104 11150 29132 11494
rect 29196 11354 29224 13466
rect 29288 13326 29316 14010
rect 29368 13728 29420 13734
rect 29368 13670 29420 13676
rect 29380 13326 29408 13670
rect 29276 13320 29328 13326
rect 29276 13262 29328 13268
rect 29368 13320 29420 13326
rect 29368 13262 29420 13268
rect 29184 11348 29236 11354
rect 29184 11290 29236 11296
rect 29092 11144 29144 11150
rect 29092 11086 29144 11092
rect 28724 10804 28776 10810
rect 28724 10746 28776 10752
rect 28736 10538 28764 10746
rect 29092 10736 29144 10742
rect 29092 10678 29144 10684
rect 29000 10600 29052 10606
rect 29000 10542 29052 10548
rect 28724 10532 28776 10538
rect 28724 10474 28776 10480
rect 28724 10056 28776 10062
rect 28724 9998 28776 10004
rect 28816 10056 28868 10062
rect 28816 9998 28868 10004
rect 28736 9518 28764 9998
rect 28828 9722 28856 9998
rect 29012 9994 29040 10542
rect 29104 10198 29132 10678
rect 29092 10192 29144 10198
rect 29092 10134 29144 10140
rect 29000 9988 29052 9994
rect 29000 9930 29052 9936
rect 28816 9716 28868 9722
rect 28816 9658 28868 9664
rect 28724 9512 28776 9518
rect 28724 9454 28776 9460
rect 29104 8838 29132 10134
rect 29472 9692 29500 14894
rect 29644 13184 29696 13190
rect 29644 13126 29696 13132
rect 29656 12986 29684 13126
rect 29644 12980 29696 12986
rect 29644 12922 29696 12928
rect 29748 12442 29776 17614
rect 29736 12436 29788 12442
rect 29840 12434 29868 19366
rect 30300 19310 30328 19790
rect 30392 19514 30420 20402
rect 30656 20324 30708 20330
rect 30656 20266 30708 20272
rect 30668 20058 30696 20266
rect 30656 20052 30708 20058
rect 30656 19994 30708 20000
rect 30472 19780 30524 19786
rect 30472 19722 30524 19728
rect 30380 19508 30432 19514
rect 30380 19450 30432 19456
rect 30484 19310 30512 19722
rect 30288 19304 30340 19310
rect 30288 19246 30340 19252
rect 30472 19304 30524 19310
rect 30472 19246 30524 19252
rect 30378 18320 30434 18329
rect 30288 18284 30340 18290
rect 30378 18255 30380 18264
rect 30288 18226 30340 18232
rect 30432 18255 30434 18264
rect 30380 18226 30432 18232
rect 30012 17740 30064 17746
rect 30012 17682 30064 17688
rect 30024 15994 30052 17682
rect 30300 17678 30328 18226
rect 30484 18222 30512 19246
rect 30748 18692 30800 18698
rect 30748 18634 30800 18640
rect 30760 18426 30788 18634
rect 30748 18420 30800 18426
rect 30748 18362 30800 18368
rect 30852 18358 30880 22664
rect 31128 22409 31156 24670
rect 31208 24608 31260 24614
rect 31208 24550 31260 24556
rect 31220 24410 31248 24550
rect 31208 24404 31260 24410
rect 31208 24346 31260 24352
rect 31588 24342 31616 24754
rect 31576 24336 31628 24342
rect 31576 24278 31628 24284
rect 31484 24064 31536 24070
rect 31484 24006 31536 24012
rect 31496 23866 31524 24006
rect 31484 23860 31536 23866
rect 31484 23802 31536 23808
rect 31852 22976 31904 22982
rect 31852 22918 31904 22924
rect 31864 22574 31892 22918
rect 31944 22636 31996 22642
rect 31944 22578 31996 22584
rect 31852 22568 31904 22574
rect 31852 22510 31904 22516
rect 31114 22400 31170 22409
rect 31114 22335 31170 22344
rect 31206 22128 31262 22137
rect 31206 22063 31208 22072
rect 31260 22063 31262 22072
rect 31484 22092 31536 22098
rect 31208 22034 31260 22040
rect 31484 22034 31536 22040
rect 31116 22024 31168 22030
rect 31116 21966 31168 21972
rect 31128 21554 31156 21966
rect 31116 21548 31168 21554
rect 31116 21490 31168 21496
rect 30932 21344 30984 21350
rect 30932 21286 30984 21292
rect 30944 21146 30972 21286
rect 30932 21140 30984 21146
rect 30932 21082 30984 21088
rect 30944 20466 30972 21082
rect 30932 20460 30984 20466
rect 30932 20402 30984 20408
rect 31116 20460 31168 20466
rect 31116 20402 31168 20408
rect 31128 19417 31156 20402
rect 31208 20256 31260 20262
rect 31208 20198 31260 20204
rect 31220 19922 31248 20198
rect 31208 19916 31260 19922
rect 31208 19858 31260 19864
rect 31114 19408 31170 19417
rect 31114 19343 31170 19352
rect 30932 18624 30984 18630
rect 30932 18566 30984 18572
rect 30840 18352 30892 18358
rect 30840 18294 30892 18300
rect 30472 18216 30524 18222
rect 30472 18158 30524 18164
rect 30288 17672 30340 17678
rect 30288 17614 30340 17620
rect 30196 17536 30248 17542
rect 30196 17478 30248 17484
rect 30208 17338 30236 17478
rect 30196 17332 30248 17338
rect 30196 17274 30248 17280
rect 30300 16726 30328 17614
rect 30288 16720 30340 16726
rect 30288 16662 30340 16668
rect 30196 16584 30248 16590
rect 30196 16526 30248 16532
rect 30288 16584 30340 16590
rect 30288 16526 30340 16532
rect 30656 16584 30708 16590
rect 30656 16526 30708 16532
rect 30208 16250 30236 16526
rect 30196 16244 30248 16250
rect 30196 16186 30248 16192
rect 30300 16182 30328 16526
rect 30668 16454 30696 16526
rect 30656 16448 30708 16454
rect 30656 16390 30708 16396
rect 30748 16448 30800 16454
rect 30748 16390 30800 16396
rect 30760 16250 30788 16390
rect 30748 16244 30800 16250
rect 30748 16186 30800 16192
rect 30288 16176 30340 16182
rect 30288 16118 30340 16124
rect 29932 15966 30052 15994
rect 29932 12714 29960 15966
rect 30012 15904 30064 15910
rect 30196 15904 30248 15910
rect 30064 15864 30144 15892
rect 30012 15846 30064 15852
rect 29920 12708 29972 12714
rect 29920 12650 29972 12656
rect 30012 12640 30064 12646
rect 30012 12582 30064 12588
rect 29840 12406 29960 12434
rect 29736 12378 29788 12384
rect 29736 11756 29788 11762
rect 29736 11698 29788 11704
rect 29460 9686 29512 9692
rect 29748 9674 29776 11698
rect 29828 11688 29880 11694
rect 29828 11630 29880 11636
rect 29460 9628 29512 9634
rect 29564 9646 29776 9674
rect 29564 9586 29592 9646
rect 29460 9580 29512 9586
rect 29460 9522 29512 9528
rect 29552 9580 29604 9586
rect 29552 9522 29604 9528
rect 29184 9104 29236 9110
rect 29184 9046 29236 9052
rect 28816 8832 28868 8838
rect 28816 8774 28868 8780
rect 28908 8832 28960 8838
rect 28908 8774 28960 8780
rect 29000 8832 29052 8838
rect 29000 8774 29052 8780
rect 29092 8832 29144 8838
rect 29092 8774 29144 8780
rect 28724 7948 28776 7954
rect 28724 7890 28776 7896
rect 28632 7336 28684 7342
rect 28632 7278 28684 7284
rect 28448 6860 28500 6866
rect 28448 6802 28500 6808
rect 28540 6860 28592 6866
rect 28540 6802 28592 6808
rect 28632 6860 28684 6866
rect 28736 6848 28764 7890
rect 28684 6820 28764 6848
rect 28632 6802 28684 6808
rect 28448 6724 28500 6730
rect 28448 6666 28500 6672
rect 28356 6656 28408 6662
rect 28356 6598 28408 6604
rect 28460 5302 28488 6666
rect 28644 5914 28672 6802
rect 28828 6798 28856 8774
rect 28920 8634 28948 8774
rect 28908 8628 28960 8634
rect 28908 8570 28960 8576
rect 29012 8566 29040 8774
rect 29000 8560 29052 8566
rect 29000 8502 29052 8508
rect 29012 8294 29040 8502
rect 29000 8288 29052 8294
rect 29000 8230 29052 8236
rect 29196 7410 29224 9046
rect 29276 9036 29328 9042
rect 29328 8996 29408 9024
rect 29276 8978 29328 8984
rect 29276 8900 29328 8906
rect 29276 8842 29328 8848
rect 29288 8430 29316 8842
rect 29276 8424 29328 8430
rect 29276 8366 29328 8372
rect 29380 8090 29408 8996
rect 29472 8090 29500 9522
rect 29840 9466 29868 11630
rect 29932 9625 29960 12406
rect 30024 12238 30052 12582
rect 30012 12232 30064 12238
rect 30012 12174 30064 12180
rect 30116 11898 30144 15864
rect 30380 15904 30432 15910
rect 30196 15846 30248 15852
rect 30300 15864 30380 15892
rect 30208 14074 30236 15846
rect 30300 14385 30328 15864
rect 30380 15846 30432 15852
rect 30760 15706 30788 16186
rect 30748 15700 30800 15706
rect 30748 15642 30800 15648
rect 30748 15428 30800 15434
rect 30748 15370 30800 15376
rect 30472 15360 30524 15366
rect 30472 15302 30524 15308
rect 30484 15026 30512 15302
rect 30760 15026 30788 15370
rect 30472 15020 30524 15026
rect 30472 14962 30524 14968
rect 30748 15020 30800 15026
rect 30748 14962 30800 14968
rect 30840 15020 30892 15026
rect 30840 14962 30892 14968
rect 30380 14952 30432 14958
rect 30380 14894 30432 14900
rect 30286 14376 30342 14385
rect 30286 14311 30342 14320
rect 30392 14278 30420 14894
rect 30484 14346 30512 14962
rect 30760 14346 30788 14962
rect 30852 14482 30880 14962
rect 30840 14476 30892 14482
rect 30840 14418 30892 14424
rect 30472 14340 30524 14346
rect 30472 14282 30524 14288
rect 30748 14340 30800 14346
rect 30748 14282 30800 14288
rect 30288 14272 30340 14278
rect 30288 14214 30340 14220
rect 30380 14272 30432 14278
rect 30380 14214 30432 14220
rect 30196 14068 30248 14074
rect 30196 14010 30248 14016
rect 30300 13818 30328 14214
rect 30392 13938 30420 14214
rect 30380 13932 30432 13938
rect 30380 13874 30432 13880
rect 30472 13932 30524 13938
rect 30472 13874 30524 13880
rect 30300 13790 30420 13818
rect 30196 13728 30248 13734
rect 30196 13670 30248 13676
rect 30208 12220 30236 13670
rect 30288 13456 30340 13462
rect 30288 13398 30340 13404
rect 30300 12782 30328 13398
rect 30392 12850 30420 13790
rect 30484 13734 30512 13874
rect 30564 13864 30616 13870
rect 30564 13806 30616 13812
rect 30472 13728 30524 13734
rect 30472 13670 30524 13676
rect 30380 12844 30432 12850
rect 30380 12786 30432 12792
rect 30288 12776 30340 12782
rect 30288 12718 30340 12724
rect 30288 12232 30340 12238
rect 30208 12192 30288 12220
rect 30288 12174 30340 12180
rect 30104 11892 30156 11898
rect 30104 11834 30156 11840
rect 30104 11348 30156 11354
rect 30104 11290 30156 11296
rect 30012 11076 30064 11082
rect 30012 11018 30064 11024
rect 30024 10985 30052 11018
rect 30010 10976 30066 10985
rect 30010 10911 30066 10920
rect 30012 9648 30064 9654
rect 29918 9616 29974 9625
rect 30012 9590 30064 9596
rect 29918 9551 29974 9560
rect 29656 9438 29868 9466
rect 29656 9178 29684 9438
rect 29736 9376 29788 9382
rect 29736 9318 29788 9324
rect 29748 9178 29776 9318
rect 29644 9172 29696 9178
rect 29644 9114 29696 9120
rect 29736 9172 29788 9178
rect 29736 9114 29788 9120
rect 29826 9072 29882 9081
rect 29932 9058 29960 9551
rect 29882 9030 29960 9058
rect 29826 9007 29882 9016
rect 30024 8566 30052 9590
rect 30116 9450 30144 11290
rect 30300 11234 30328 12174
rect 30392 12102 30420 12786
rect 30380 12096 30432 12102
rect 30380 12038 30432 12044
rect 30472 12096 30524 12102
rect 30472 12038 30524 12044
rect 30392 11830 30420 12038
rect 30484 11898 30512 12038
rect 30472 11892 30524 11898
rect 30472 11834 30524 11840
rect 30380 11824 30432 11830
rect 30380 11766 30432 11772
rect 30380 11552 30432 11558
rect 30380 11494 30432 11500
rect 30392 11354 30420 11494
rect 30484 11354 30512 11834
rect 30380 11348 30432 11354
rect 30380 11290 30432 11296
rect 30472 11348 30524 11354
rect 30472 11290 30524 11296
rect 30300 11206 30420 11234
rect 30288 11144 30340 11150
rect 30288 11086 30340 11092
rect 30196 10668 30248 10674
rect 30300 10656 30328 11086
rect 30248 10628 30328 10656
rect 30196 10610 30248 10616
rect 30208 9674 30236 10610
rect 30288 10464 30340 10470
rect 30288 10406 30340 10412
rect 30300 10062 30328 10406
rect 30392 10198 30420 11206
rect 30576 10266 30604 13806
rect 30656 11688 30708 11694
rect 30656 11630 30708 11636
rect 30668 11354 30696 11630
rect 30656 11348 30708 11354
rect 30656 11290 30708 11296
rect 30656 11008 30708 11014
rect 30656 10950 30708 10956
rect 30564 10260 30616 10266
rect 30564 10202 30616 10208
rect 30386 10192 30438 10198
rect 30386 10134 30438 10140
rect 30668 10062 30696 10950
rect 30288 10056 30340 10062
rect 30656 10056 30708 10062
rect 30288 9998 30340 10004
rect 30392 10016 30656 10044
rect 30392 9722 30420 10016
rect 30656 9998 30708 10004
rect 30840 9920 30892 9926
rect 30840 9862 30892 9868
rect 30380 9716 30432 9722
rect 30208 9646 30328 9674
rect 30380 9658 30432 9664
rect 30104 9444 30156 9450
rect 30104 9386 30156 9392
rect 30116 8956 30144 9386
rect 30196 8968 30248 8974
rect 30116 8928 30196 8956
rect 30196 8910 30248 8916
rect 30208 8634 30236 8910
rect 30196 8628 30248 8634
rect 30196 8570 30248 8576
rect 30012 8560 30064 8566
rect 30012 8502 30064 8508
rect 29368 8084 29420 8090
rect 29368 8026 29420 8032
rect 29460 8084 29512 8090
rect 29460 8026 29512 8032
rect 29184 7404 29236 7410
rect 29184 7346 29236 7352
rect 28816 6792 28868 6798
rect 28816 6734 28868 6740
rect 28632 5908 28684 5914
rect 28632 5850 28684 5856
rect 29196 5778 29224 7346
rect 29380 5846 29408 8026
rect 29472 7410 29500 8026
rect 30012 7880 30064 7886
rect 30012 7822 30064 7828
rect 30024 7546 30052 7822
rect 30012 7540 30064 7546
rect 30012 7482 30064 7488
rect 29460 7404 29512 7410
rect 29460 7346 29512 7352
rect 30012 6792 30064 6798
rect 30012 6734 30064 6740
rect 29368 5840 29420 5846
rect 29368 5782 29420 5788
rect 29184 5772 29236 5778
rect 29184 5714 29236 5720
rect 28448 5296 28500 5302
rect 28448 5238 28500 5244
rect 28264 5160 28316 5166
rect 28264 5102 28316 5108
rect 29196 5098 29224 5714
rect 29380 5302 29408 5782
rect 30024 5710 30052 6734
rect 30012 5704 30064 5710
rect 30012 5646 30064 5652
rect 30300 5642 30328 9646
rect 30852 9586 30880 9862
rect 30748 9580 30800 9586
rect 30748 9522 30800 9528
rect 30840 9580 30892 9586
rect 30840 9522 30892 9528
rect 30760 9178 30788 9522
rect 30944 9450 30972 18566
rect 31128 18306 31156 19343
rect 31208 18760 31260 18766
rect 31392 18760 31444 18766
rect 31260 18720 31340 18748
rect 31208 18702 31260 18708
rect 31208 18624 31260 18630
rect 31208 18566 31260 18572
rect 31220 18426 31248 18566
rect 31208 18420 31260 18426
rect 31208 18362 31260 18368
rect 31036 18278 31156 18306
rect 31312 18290 31340 18720
rect 31392 18702 31444 18708
rect 31300 18284 31352 18290
rect 31036 15008 31064 18278
rect 31300 18226 31352 18232
rect 31116 18216 31168 18222
rect 31116 18158 31168 18164
rect 31128 16674 31156 18158
rect 31208 17876 31260 17882
rect 31208 17818 31260 17824
rect 31220 16794 31248 17818
rect 31312 17678 31340 18226
rect 31404 17882 31432 18702
rect 31496 18154 31524 22034
rect 31864 22030 31892 22510
rect 31956 22506 31984 22578
rect 31944 22500 31996 22506
rect 31944 22442 31996 22448
rect 31852 22024 31904 22030
rect 31852 21966 31904 21972
rect 31576 19848 31628 19854
rect 31576 19790 31628 19796
rect 31588 19310 31616 19790
rect 31576 19304 31628 19310
rect 31576 19246 31628 19252
rect 31956 18306 31984 22442
rect 32036 22432 32088 22438
rect 32036 22374 32088 22380
rect 32048 22030 32076 22374
rect 32232 22094 32260 31726
rect 32324 30258 32352 32302
rect 32968 31754 32996 32846
rect 33244 32434 33272 33594
rect 33140 32428 33192 32434
rect 33140 32370 33192 32376
rect 33232 32428 33284 32434
rect 33232 32370 33284 32376
rect 32876 31726 32996 31754
rect 32876 31346 32904 31726
rect 32864 31340 32916 31346
rect 32864 31282 32916 31288
rect 32496 31272 32548 31278
rect 32496 31214 32548 31220
rect 32508 30870 32536 31214
rect 32496 30864 32548 30870
rect 32496 30806 32548 30812
rect 32508 30258 32536 30806
rect 32876 30394 32904 31282
rect 33152 30954 33180 32370
rect 33060 30926 33180 30954
rect 32864 30388 32916 30394
rect 32864 30330 32916 30336
rect 33060 30326 33088 30926
rect 33336 30818 33364 34342
rect 33428 33998 33456 34700
rect 33508 34682 33560 34688
rect 33416 33992 33468 33998
rect 33416 33934 33468 33940
rect 33612 33658 33640 35974
rect 33704 35154 33732 36722
rect 34060 36576 34112 36582
rect 34060 36518 34112 36524
rect 34072 36378 34100 36518
rect 34934 36476 35242 36485
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36411 35242 36420
rect 34060 36372 34112 36378
rect 34060 36314 34112 36320
rect 35594 35932 35902 35941
rect 35594 35930 35600 35932
rect 35656 35930 35680 35932
rect 35736 35930 35760 35932
rect 35816 35930 35840 35932
rect 35896 35930 35902 35932
rect 35656 35878 35658 35930
rect 35838 35878 35840 35930
rect 35594 35876 35600 35878
rect 35656 35876 35680 35878
rect 35736 35876 35760 35878
rect 35816 35876 35840 35878
rect 35896 35876 35902 35878
rect 35594 35867 35902 35876
rect 34934 35388 35242 35397
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35323 35242 35332
rect 33692 35148 33744 35154
rect 33692 35090 33744 35096
rect 35594 34844 35902 34853
rect 35594 34842 35600 34844
rect 35656 34842 35680 34844
rect 35736 34842 35760 34844
rect 35816 34842 35840 34844
rect 35896 34842 35902 34844
rect 35656 34790 35658 34842
rect 35838 34790 35840 34842
rect 35594 34788 35600 34790
rect 35656 34788 35680 34790
rect 35736 34788 35760 34790
rect 35816 34788 35840 34790
rect 35896 34788 35902 34790
rect 35594 34779 35902 34788
rect 34152 34604 34204 34610
rect 34152 34546 34204 34552
rect 36912 34604 36964 34610
rect 36912 34546 36964 34552
rect 33876 33992 33928 33998
rect 33876 33934 33928 33940
rect 33888 33658 33916 33934
rect 34164 33658 34192 34546
rect 34934 34300 35242 34309
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34235 35242 34244
rect 35992 33924 36044 33930
rect 35992 33866 36044 33872
rect 36636 33924 36688 33930
rect 36636 33866 36688 33872
rect 34336 33856 34388 33862
rect 34336 33798 34388 33804
rect 33600 33652 33652 33658
rect 33600 33594 33652 33600
rect 33876 33652 33928 33658
rect 33876 33594 33928 33600
rect 34152 33652 34204 33658
rect 34152 33594 34204 33600
rect 34060 33448 34112 33454
rect 34060 33390 34112 33396
rect 33782 32464 33838 32473
rect 33782 32399 33838 32408
rect 33152 30802 33364 30818
rect 33140 30796 33364 30802
rect 33192 30790 33364 30796
rect 33508 30796 33560 30802
rect 33140 30738 33192 30744
rect 33508 30738 33560 30744
rect 33048 30320 33100 30326
rect 33048 30262 33100 30268
rect 32312 30252 32364 30258
rect 32312 30194 32364 30200
rect 32496 30252 32548 30258
rect 32496 30194 32548 30200
rect 32324 29306 32352 30194
rect 32496 30048 32548 30054
rect 32496 29990 32548 29996
rect 32956 30048 33008 30054
rect 32956 29990 33008 29996
rect 32508 29306 32536 29990
rect 32312 29300 32364 29306
rect 32312 29242 32364 29248
rect 32496 29300 32548 29306
rect 32496 29242 32548 29248
rect 32404 28960 32456 28966
rect 32404 28902 32456 28908
rect 32416 28626 32444 28902
rect 32404 28620 32456 28626
rect 32404 28562 32456 28568
rect 32680 28416 32732 28422
rect 32680 28358 32732 28364
rect 32692 28218 32720 28358
rect 32680 28212 32732 28218
rect 32680 28154 32732 28160
rect 32680 26036 32732 26042
rect 32680 25978 32732 25984
rect 32692 25838 32720 25978
rect 32680 25832 32732 25838
rect 32680 25774 32732 25780
rect 32692 24614 32720 25774
rect 32968 24970 32996 29990
rect 33048 29164 33100 29170
rect 33048 29106 33100 29112
rect 33060 28218 33088 29106
rect 33048 28212 33100 28218
rect 33048 28154 33100 28160
rect 33152 28014 33180 30738
rect 33324 30592 33376 30598
rect 33324 30534 33376 30540
rect 33232 30320 33284 30326
rect 33232 30262 33284 30268
rect 33244 29238 33272 30262
rect 33336 29510 33364 30534
rect 33520 29782 33548 30738
rect 33508 29776 33560 29782
rect 33508 29718 33560 29724
rect 33324 29504 33376 29510
rect 33324 29446 33376 29452
rect 33232 29232 33284 29238
rect 33232 29174 33284 29180
rect 33324 28620 33376 28626
rect 33324 28562 33376 28568
rect 33140 28008 33192 28014
rect 33140 27950 33192 27956
rect 33140 26988 33192 26994
rect 33140 26930 33192 26936
rect 33152 26586 33180 26930
rect 33140 26580 33192 26586
rect 33140 26522 33192 26528
rect 33232 26240 33284 26246
rect 33232 26182 33284 26188
rect 33244 25906 33272 26182
rect 33336 26042 33364 28562
rect 33692 27940 33744 27946
rect 33692 27882 33744 27888
rect 33704 27470 33732 27882
rect 33796 27606 33824 32399
rect 34072 31754 34100 33390
rect 34348 32910 34376 33798
rect 35594 33756 35902 33765
rect 35594 33754 35600 33756
rect 35656 33754 35680 33756
rect 35736 33754 35760 33756
rect 35816 33754 35840 33756
rect 35896 33754 35902 33756
rect 35656 33702 35658 33754
rect 35838 33702 35840 33754
rect 35594 33700 35600 33702
rect 35656 33700 35680 33702
rect 35736 33700 35760 33702
rect 35816 33700 35840 33702
rect 35896 33700 35902 33702
rect 35594 33691 35902 33700
rect 36004 33386 36032 33866
rect 36648 33522 36676 33866
rect 36924 33658 36952 34546
rect 37924 34536 37976 34542
rect 37924 34478 37976 34484
rect 37936 34105 37964 34478
rect 37922 34096 37978 34105
rect 37922 34031 37978 34040
rect 36912 33652 36964 33658
rect 36912 33594 36964 33600
rect 36636 33516 36688 33522
rect 36636 33458 36688 33464
rect 36728 33516 36780 33522
rect 36728 33458 36780 33464
rect 35992 33380 36044 33386
rect 35992 33322 36044 33328
rect 34796 33312 34848 33318
rect 34796 33254 34848 33260
rect 34808 33114 34836 33254
rect 34934 33212 35242 33221
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33147 35242 33156
rect 34796 33108 34848 33114
rect 34796 33050 34848 33056
rect 36004 32910 36032 33322
rect 34336 32904 34388 32910
rect 34336 32846 34388 32852
rect 35992 32904 36044 32910
rect 35992 32846 36044 32852
rect 36268 32768 36320 32774
rect 36268 32710 36320 32716
rect 35594 32668 35902 32677
rect 35594 32666 35600 32668
rect 35656 32666 35680 32668
rect 35736 32666 35760 32668
rect 35816 32666 35840 32668
rect 35896 32666 35902 32668
rect 35656 32614 35658 32666
rect 35838 32614 35840 32666
rect 35594 32612 35600 32614
rect 35656 32612 35680 32614
rect 35736 32612 35760 32614
rect 35816 32612 35840 32614
rect 35896 32612 35902 32614
rect 35594 32603 35902 32612
rect 36280 32502 36308 32710
rect 34612 32496 34664 32502
rect 34612 32438 34664 32444
rect 36268 32496 36320 32502
rect 36268 32438 36320 32444
rect 34624 31822 34652 32438
rect 34934 32124 35242 32133
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32059 35242 32068
rect 34612 31816 34664 31822
rect 34612 31758 34664 31764
rect 35440 31816 35492 31822
rect 35440 31758 35492 31764
rect 34072 31726 34284 31754
rect 34152 31272 34204 31278
rect 34152 31214 34204 31220
rect 34164 30938 34192 31214
rect 34152 30932 34204 30938
rect 34152 30874 34204 30880
rect 33968 30796 34020 30802
rect 33968 30738 34020 30744
rect 33980 28626 34008 30738
rect 34256 29782 34284 31726
rect 34520 31748 34572 31754
rect 34520 31690 34572 31696
rect 34532 31346 34560 31690
rect 34520 31340 34572 31346
rect 34520 31282 34572 31288
rect 34244 29776 34296 29782
rect 34244 29718 34296 29724
rect 34152 29640 34204 29646
rect 34152 29582 34204 29588
rect 34164 29306 34192 29582
rect 34152 29300 34204 29306
rect 34152 29242 34204 29248
rect 33968 28620 34020 28626
rect 33968 28562 34020 28568
rect 34060 28484 34112 28490
rect 34060 28426 34112 28432
rect 33876 28008 33928 28014
rect 33876 27950 33928 27956
rect 33784 27600 33836 27606
rect 33784 27542 33836 27548
rect 33692 27464 33744 27470
rect 33692 27406 33744 27412
rect 33600 27328 33652 27334
rect 33600 27270 33652 27276
rect 33612 27062 33640 27270
rect 33600 27056 33652 27062
rect 33600 26998 33652 27004
rect 33888 26450 33916 27950
rect 34072 27130 34100 28426
rect 34152 28416 34204 28422
rect 34152 28358 34204 28364
rect 34164 28082 34192 28358
rect 34152 28076 34204 28082
rect 34152 28018 34204 28024
rect 34256 27962 34284 29718
rect 34336 29572 34388 29578
rect 34336 29514 34388 29520
rect 34348 29238 34376 29514
rect 34520 29504 34572 29510
rect 34520 29446 34572 29452
rect 34336 29232 34388 29238
rect 34336 29174 34388 29180
rect 34164 27934 34284 27962
rect 34060 27124 34112 27130
rect 34060 27066 34112 27072
rect 33876 26444 33928 26450
rect 33876 26386 33928 26392
rect 33692 26240 33744 26246
rect 33692 26182 33744 26188
rect 33324 26036 33376 26042
rect 33324 25978 33376 25984
rect 33704 25974 33732 26182
rect 33692 25968 33744 25974
rect 33692 25910 33744 25916
rect 33232 25900 33284 25906
rect 33232 25842 33284 25848
rect 34164 25838 34192 27934
rect 34348 27606 34376 29174
rect 34532 29170 34560 29446
rect 34520 29164 34572 29170
rect 34520 29106 34572 29112
rect 34428 28484 34480 28490
rect 34428 28426 34480 28432
rect 34440 28218 34468 28426
rect 34520 28416 34572 28422
rect 34520 28358 34572 28364
rect 34428 28212 34480 28218
rect 34428 28154 34480 28160
rect 34532 28082 34560 28358
rect 34520 28076 34572 28082
rect 34520 28018 34572 28024
rect 34624 27946 34652 31758
rect 34796 31680 34848 31686
rect 34796 31622 34848 31628
rect 35256 31680 35308 31686
rect 35256 31622 35308 31628
rect 34808 31482 34836 31622
rect 34796 31476 34848 31482
rect 34796 31418 34848 31424
rect 35268 31278 35296 31622
rect 35256 31272 35308 31278
rect 35256 31214 35308 31220
rect 34934 31036 35242 31045
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30971 35242 30980
rect 35452 30938 35480 31758
rect 35594 31580 35902 31589
rect 35594 31578 35600 31580
rect 35656 31578 35680 31580
rect 35736 31578 35760 31580
rect 35816 31578 35840 31580
rect 35896 31578 35902 31580
rect 35656 31526 35658 31578
rect 35838 31526 35840 31578
rect 35594 31524 35600 31526
rect 35656 31524 35680 31526
rect 35736 31524 35760 31526
rect 35816 31524 35840 31526
rect 35896 31524 35902 31526
rect 35594 31515 35902 31524
rect 35992 31136 36044 31142
rect 35992 31078 36044 31084
rect 36544 31136 36596 31142
rect 36544 31078 36596 31084
rect 35440 30932 35492 30938
rect 35440 30874 35492 30880
rect 35594 30492 35902 30501
rect 35594 30490 35600 30492
rect 35656 30490 35680 30492
rect 35736 30490 35760 30492
rect 35816 30490 35840 30492
rect 35896 30490 35902 30492
rect 35656 30438 35658 30490
rect 35838 30438 35840 30490
rect 35594 30436 35600 30438
rect 35656 30436 35680 30438
rect 35736 30436 35760 30438
rect 35816 30436 35840 30438
rect 35896 30436 35902 30438
rect 35594 30427 35902 30436
rect 36004 30326 36032 31078
rect 36556 30666 36584 31078
rect 36544 30660 36596 30666
rect 36544 30602 36596 30608
rect 35992 30320 36044 30326
rect 35992 30262 36044 30268
rect 34934 29948 35242 29957
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29883 35242 29892
rect 34796 29640 34848 29646
rect 34796 29582 34848 29588
rect 34808 29306 34836 29582
rect 34980 29572 35032 29578
rect 34980 29514 35032 29520
rect 34796 29300 34848 29306
rect 34796 29242 34848 29248
rect 34992 29170 35020 29514
rect 36004 29510 36032 30262
rect 36648 29617 36676 33458
rect 36740 32570 36768 33458
rect 36728 32564 36780 32570
rect 36728 32506 36780 32512
rect 36634 29608 36690 29617
rect 36634 29543 36690 29552
rect 35992 29504 36044 29510
rect 35992 29446 36044 29452
rect 35594 29404 35902 29413
rect 35594 29402 35600 29404
rect 35656 29402 35680 29404
rect 35736 29402 35760 29404
rect 35816 29402 35840 29404
rect 35896 29402 35902 29404
rect 35656 29350 35658 29402
rect 35838 29350 35840 29402
rect 35594 29348 35600 29350
rect 35656 29348 35680 29350
rect 35736 29348 35760 29350
rect 35816 29348 35840 29350
rect 35896 29348 35902 29350
rect 35594 29339 35902 29348
rect 34980 29164 35032 29170
rect 34980 29106 35032 29112
rect 34704 29028 34756 29034
rect 34756 28976 34836 28994
rect 34704 28970 34836 28976
rect 34716 28966 34836 28970
rect 34704 28552 34756 28558
rect 34704 28494 34756 28500
rect 34716 28218 34744 28494
rect 34704 28212 34756 28218
rect 34704 28154 34756 28160
rect 34612 27940 34664 27946
rect 34612 27882 34664 27888
rect 34336 27600 34388 27606
rect 34336 27542 34388 27548
rect 34348 26042 34376 27542
rect 34704 26376 34756 26382
rect 34704 26318 34756 26324
rect 34716 26042 34744 26318
rect 34336 26036 34388 26042
rect 34336 25978 34388 25984
rect 34704 26036 34756 26042
rect 34704 25978 34756 25984
rect 34808 25888 34836 28966
rect 34934 28860 35242 28869
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28795 35242 28804
rect 36004 28490 36032 29446
rect 36648 29170 36676 29543
rect 36636 29164 36688 29170
rect 36636 29106 36688 29112
rect 36820 29164 36872 29170
rect 36820 29106 36872 29112
rect 35992 28484 36044 28490
rect 35992 28426 36044 28432
rect 35594 28316 35902 28325
rect 35594 28314 35600 28316
rect 35656 28314 35680 28316
rect 35736 28314 35760 28316
rect 35816 28314 35840 28316
rect 35896 28314 35902 28316
rect 35656 28262 35658 28314
rect 35838 28262 35840 28314
rect 35594 28260 35600 28262
rect 35656 28260 35680 28262
rect 35736 28260 35760 28262
rect 35816 28260 35840 28262
rect 35896 28260 35902 28262
rect 35594 28251 35902 28260
rect 34934 27772 35242 27781
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27707 35242 27716
rect 35594 27228 35902 27237
rect 35594 27226 35600 27228
rect 35656 27226 35680 27228
rect 35736 27226 35760 27228
rect 35816 27226 35840 27228
rect 35896 27226 35902 27228
rect 35656 27174 35658 27226
rect 35838 27174 35840 27226
rect 35594 27172 35600 27174
rect 35656 27172 35680 27174
rect 35736 27172 35760 27174
rect 35816 27172 35840 27174
rect 35896 27172 35902 27174
rect 35594 27163 35902 27172
rect 36004 26994 36032 28426
rect 35992 26988 36044 26994
rect 35992 26930 36044 26936
rect 35440 26920 35492 26926
rect 35440 26862 35492 26868
rect 34934 26684 35242 26693
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26619 35242 26628
rect 35452 26586 35480 26862
rect 35440 26580 35492 26586
rect 35440 26522 35492 26528
rect 34980 26376 35032 26382
rect 34980 26318 35032 26324
rect 34992 26042 35020 26318
rect 36004 26314 36032 26930
rect 35992 26308 36044 26314
rect 35992 26250 36044 26256
rect 36636 26308 36688 26314
rect 36636 26250 36688 26256
rect 35594 26140 35902 26149
rect 35594 26138 35600 26140
rect 35656 26138 35680 26140
rect 35736 26138 35760 26140
rect 35816 26138 35840 26140
rect 35896 26138 35902 26140
rect 35656 26086 35658 26138
rect 35838 26086 35840 26138
rect 35594 26084 35600 26086
rect 35656 26084 35680 26086
rect 35736 26084 35760 26086
rect 35816 26084 35840 26086
rect 35896 26084 35902 26086
rect 35594 26075 35902 26084
rect 34980 26036 35032 26042
rect 34980 25978 35032 25984
rect 34624 25860 34836 25888
rect 34152 25832 34204 25838
rect 34152 25774 34204 25780
rect 32968 24942 33180 24970
rect 33152 24818 33180 24942
rect 33048 24812 33100 24818
rect 33048 24754 33100 24760
rect 33140 24812 33192 24818
rect 33140 24754 33192 24760
rect 33784 24812 33836 24818
rect 33784 24754 33836 24760
rect 32680 24608 32732 24614
rect 32680 24550 32732 24556
rect 32956 24404 33008 24410
rect 32956 24346 33008 24352
rect 32864 24200 32916 24206
rect 32864 24142 32916 24148
rect 32404 24064 32456 24070
rect 32404 24006 32456 24012
rect 32588 24064 32640 24070
rect 32588 24006 32640 24012
rect 32416 23118 32444 24006
rect 32312 23112 32364 23118
rect 32312 23054 32364 23060
rect 32404 23112 32456 23118
rect 32404 23054 32456 23060
rect 32496 23112 32548 23118
rect 32496 23054 32548 23060
rect 32324 22250 32352 23054
rect 32416 22710 32444 23054
rect 32508 22778 32536 23054
rect 32496 22772 32548 22778
rect 32496 22714 32548 22720
rect 32404 22704 32456 22710
rect 32404 22646 32456 22652
rect 32496 22636 32548 22642
rect 32496 22578 32548 22584
rect 32508 22522 32536 22578
rect 32416 22494 32536 22522
rect 32416 22438 32444 22494
rect 32404 22432 32456 22438
rect 32404 22374 32456 22380
rect 32496 22432 32548 22438
rect 32496 22374 32548 22380
rect 32324 22222 32444 22250
rect 32416 22166 32444 22222
rect 32404 22160 32456 22166
rect 32404 22102 32456 22108
rect 32232 22066 32352 22094
rect 32036 22024 32088 22030
rect 32036 21966 32088 21972
rect 32220 21888 32272 21894
rect 32220 21830 32272 21836
rect 32232 21554 32260 21830
rect 32220 21548 32272 21554
rect 32220 21490 32272 21496
rect 32036 20528 32088 20534
rect 32036 20470 32088 20476
rect 32048 20058 32076 20470
rect 32324 20058 32352 22066
rect 32508 21842 32536 22374
rect 32600 22094 32628 24006
rect 32876 23866 32904 24142
rect 32864 23860 32916 23866
rect 32784 23820 32864 23848
rect 32784 23118 32812 23820
rect 32864 23802 32916 23808
rect 32772 23112 32824 23118
rect 32772 23054 32824 23060
rect 32968 22794 32996 24346
rect 33060 24342 33088 24754
rect 33232 24676 33284 24682
rect 33152 24636 33232 24664
rect 33048 24336 33100 24342
rect 33048 24278 33100 24284
rect 33060 23594 33088 24278
rect 33152 24206 33180 24636
rect 33232 24618 33284 24624
rect 33600 24676 33652 24682
rect 33600 24618 33652 24624
rect 33324 24608 33376 24614
rect 33324 24550 33376 24556
rect 33336 24206 33364 24550
rect 33508 24336 33560 24342
rect 33508 24278 33560 24284
rect 33140 24200 33192 24206
rect 33140 24142 33192 24148
rect 33324 24200 33376 24206
rect 33324 24142 33376 24148
rect 33140 24064 33192 24070
rect 33140 24006 33192 24012
rect 33152 23866 33180 24006
rect 33140 23860 33192 23866
rect 33140 23802 33192 23808
rect 33048 23588 33100 23594
rect 33048 23530 33100 23536
rect 33232 23520 33284 23526
rect 33232 23462 33284 23468
rect 32876 22766 32996 22794
rect 32876 22642 32904 22766
rect 33244 22642 33272 23462
rect 33324 23044 33376 23050
rect 33324 22986 33376 22992
rect 33336 22642 33364 22986
rect 32864 22636 32916 22642
rect 32864 22578 32916 22584
rect 33232 22636 33284 22642
rect 33232 22578 33284 22584
rect 33324 22636 33376 22642
rect 33324 22578 33376 22584
rect 32876 22234 32904 22578
rect 32956 22568 33008 22574
rect 32956 22510 33008 22516
rect 32864 22228 32916 22234
rect 32864 22170 32916 22176
rect 32862 22128 32918 22137
rect 32600 22066 32720 22094
rect 32692 22030 32720 22066
rect 32862 22063 32864 22072
rect 32916 22063 32918 22072
rect 32864 22034 32916 22040
rect 32680 22024 32732 22030
rect 32680 21966 32732 21972
rect 32508 21814 32720 21842
rect 32588 21684 32640 21690
rect 32588 21626 32640 21632
rect 32404 20868 32456 20874
rect 32404 20810 32456 20816
rect 32036 20052 32088 20058
rect 32036 19994 32088 20000
rect 32312 20052 32364 20058
rect 32312 19994 32364 20000
rect 32312 18624 32364 18630
rect 32312 18566 32364 18572
rect 31956 18278 32076 18306
rect 31944 18216 31996 18222
rect 31944 18158 31996 18164
rect 31484 18148 31536 18154
rect 31484 18090 31536 18096
rect 31392 17876 31444 17882
rect 31392 17818 31444 17824
rect 31300 17672 31352 17678
rect 31300 17614 31352 17620
rect 31956 17610 31984 18158
rect 32048 18086 32076 18278
rect 32036 18080 32088 18086
rect 32036 18022 32088 18028
rect 31944 17604 31996 17610
rect 31944 17546 31996 17552
rect 31956 17338 31984 17546
rect 31944 17332 31996 17338
rect 31944 17274 31996 17280
rect 31852 16992 31904 16998
rect 31852 16934 31904 16940
rect 31864 16794 31892 16934
rect 31208 16788 31260 16794
rect 31208 16730 31260 16736
rect 31852 16788 31904 16794
rect 31852 16730 31904 16736
rect 31128 16646 31248 16674
rect 31116 16584 31168 16590
rect 31116 16526 31168 16532
rect 31128 16182 31156 16526
rect 31116 16176 31168 16182
rect 31116 16118 31168 16124
rect 31220 15586 31248 16646
rect 31760 16652 31812 16658
rect 31760 16594 31812 16600
rect 31484 16584 31536 16590
rect 31484 16526 31536 16532
rect 31392 15904 31444 15910
rect 31392 15846 31444 15852
rect 31404 15706 31432 15846
rect 31392 15700 31444 15706
rect 31392 15642 31444 15648
rect 31220 15558 31432 15586
rect 31116 15020 31168 15026
rect 31036 14980 31116 15008
rect 31116 14962 31168 14968
rect 30932 9444 30984 9450
rect 30932 9386 30984 9392
rect 30748 9172 30800 9178
rect 30748 9114 30800 9120
rect 30654 9072 30710 9081
rect 30654 9007 30710 9016
rect 30380 8900 30432 8906
rect 30380 8842 30432 8848
rect 30392 7886 30420 8842
rect 30472 7948 30524 7954
rect 30472 7890 30524 7896
rect 30380 7880 30432 7886
rect 30380 7822 30432 7828
rect 30380 7336 30432 7342
rect 30380 7278 30432 7284
rect 30392 7002 30420 7278
rect 30380 6996 30432 7002
rect 30380 6938 30432 6944
rect 30484 6798 30512 7890
rect 30564 7880 30616 7886
rect 30564 7822 30616 7828
rect 30576 7206 30604 7822
rect 30668 7410 30696 9007
rect 30840 8832 30892 8838
rect 30840 8774 30892 8780
rect 30852 7886 30880 8774
rect 31024 8424 31076 8430
rect 31024 8366 31076 8372
rect 31036 7886 31064 8366
rect 30840 7880 30892 7886
rect 30840 7822 30892 7828
rect 31024 7880 31076 7886
rect 31024 7822 31076 7828
rect 30748 7812 30800 7818
rect 30748 7754 30800 7760
rect 30656 7404 30708 7410
rect 30656 7346 30708 7352
rect 30564 7200 30616 7206
rect 30564 7142 30616 7148
rect 30576 6866 30604 7142
rect 30564 6860 30616 6866
rect 30564 6802 30616 6808
rect 30760 6798 30788 7754
rect 30852 7002 30880 7822
rect 30840 6996 30892 7002
rect 30840 6938 30892 6944
rect 30472 6792 30524 6798
rect 30472 6734 30524 6740
rect 30748 6792 30800 6798
rect 30748 6734 30800 6740
rect 30484 5914 30512 6734
rect 31036 6458 31064 7822
rect 31128 7750 31156 14962
rect 31208 14816 31260 14822
rect 31208 14758 31260 14764
rect 31220 14414 31248 14758
rect 31300 14544 31352 14550
rect 31300 14486 31352 14492
rect 31208 14408 31260 14414
rect 31208 14350 31260 14356
rect 31208 13320 31260 13326
rect 31208 13262 31260 13268
rect 31220 12986 31248 13262
rect 31208 12980 31260 12986
rect 31208 12922 31260 12928
rect 31312 12850 31340 14486
rect 31404 14414 31432 15558
rect 31392 14408 31444 14414
rect 31392 14350 31444 14356
rect 31404 13954 31432 14350
rect 31496 14074 31524 16526
rect 31772 15910 31800 16594
rect 31760 15904 31812 15910
rect 31760 15846 31812 15852
rect 31668 14952 31720 14958
rect 31668 14894 31720 14900
rect 31680 14482 31708 14894
rect 31760 14612 31812 14618
rect 31760 14554 31812 14560
rect 31668 14476 31720 14482
rect 31668 14418 31720 14424
rect 31772 14414 31800 14554
rect 31760 14408 31812 14414
rect 31760 14350 31812 14356
rect 31484 14068 31536 14074
rect 31484 14010 31536 14016
rect 31404 13926 31524 13954
rect 31300 12844 31352 12850
rect 31300 12786 31352 12792
rect 31392 12844 31444 12850
rect 31392 12786 31444 12792
rect 31298 10976 31354 10985
rect 31298 10911 31354 10920
rect 31312 10742 31340 10911
rect 31300 10736 31352 10742
rect 31300 10678 31352 10684
rect 31404 9586 31432 12786
rect 31392 9580 31444 9586
rect 31392 9522 31444 9528
rect 31404 8634 31432 9522
rect 31392 8628 31444 8634
rect 31392 8570 31444 8576
rect 31496 8090 31524 13926
rect 31852 13728 31904 13734
rect 31852 13670 31904 13676
rect 31864 12986 31892 13670
rect 31852 12980 31904 12986
rect 31852 12922 31904 12928
rect 31760 12436 31812 12442
rect 31760 12378 31812 12384
rect 31772 11286 31800 12378
rect 32048 12238 32076 18022
rect 32324 17814 32352 18566
rect 32416 17814 32444 20810
rect 32600 20466 32628 21626
rect 32692 21554 32720 21814
rect 32680 21548 32732 21554
rect 32680 21490 32732 21496
rect 32588 20460 32640 20466
rect 32588 20402 32640 20408
rect 32864 18964 32916 18970
rect 32864 18906 32916 18912
rect 32680 18760 32732 18766
rect 32680 18702 32732 18708
rect 32772 18760 32824 18766
rect 32772 18702 32824 18708
rect 32692 18358 32720 18702
rect 32680 18352 32732 18358
rect 32680 18294 32732 18300
rect 32784 18290 32812 18702
rect 32772 18284 32824 18290
rect 32772 18226 32824 18232
rect 32496 18216 32548 18222
rect 32496 18158 32548 18164
rect 32588 18216 32640 18222
rect 32588 18158 32640 18164
rect 32508 17882 32536 18158
rect 32496 17876 32548 17882
rect 32496 17818 32548 17824
rect 32312 17808 32364 17814
rect 32312 17750 32364 17756
rect 32404 17808 32456 17814
rect 32404 17750 32456 17756
rect 32128 17196 32180 17202
rect 32128 17138 32180 17144
rect 32140 16794 32168 17138
rect 32324 17134 32352 17750
rect 32600 17746 32628 18158
rect 32588 17740 32640 17746
rect 32588 17682 32640 17688
rect 32496 17536 32548 17542
rect 32496 17478 32548 17484
rect 32404 17332 32456 17338
rect 32404 17274 32456 17280
rect 32416 17134 32444 17274
rect 32508 17270 32536 17478
rect 32496 17264 32548 17270
rect 32496 17206 32548 17212
rect 32508 17134 32536 17206
rect 32312 17128 32364 17134
rect 32312 17070 32364 17076
rect 32404 17128 32456 17134
rect 32404 17070 32456 17076
rect 32496 17128 32548 17134
rect 32496 17070 32548 17076
rect 32128 16788 32180 16794
rect 32128 16730 32180 16736
rect 32220 16040 32272 16046
rect 32220 15982 32272 15988
rect 32232 15706 32260 15982
rect 32220 15700 32272 15706
rect 32220 15642 32272 15648
rect 32232 15434 32260 15642
rect 32220 15428 32272 15434
rect 32220 15370 32272 15376
rect 32128 14272 32180 14278
rect 32128 14214 32180 14220
rect 32036 12232 32088 12238
rect 32036 12174 32088 12180
rect 32140 11354 32168 14214
rect 32324 12306 32352 17070
rect 32784 16522 32812 18226
rect 32876 17338 32904 18906
rect 32968 18748 32996 22510
rect 33140 22092 33192 22098
rect 33336 22080 33364 22578
rect 33192 22052 33364 22080
rect 33140 22034 33192 22040
rect 33336 21894 33364 22052
rect 33520 22030 33548 24278
rect 33612 23662 33640 24618
rect 33796 24206 33824 24754
rect 34164 24682 34192 25774
rect 34336 25288 34388 25294
rect 34336 25230 34388 25236
rect 34348 24954 34376 25230
rect 34336 24948 34388 24954
rect 34336 24890 34388 24896
rect 34152 24676 34204 24682
rect 34152 24618 34204 24624
rect 33784 24200 33836 24206
rect 33784 24142 33836 24148
rect 34624 23866 34652 25860
rect 34704 25764 34756 25770
rect 34704 25706 34756 25712
rect 34716 25430 34744 25706
rect 34796 25696 34848 25702
rect 34796 25638 34848 25644
rect 34704 25424 34756 25430
rect 34704 25366 34756 25372
rect 34612 23860 34664 23866
rect 34612 23802 34664 23808
rect 33600 23656 33652 23662
rect 33600 23598 33652 23604
rect 34624 23118 34652 23802
rect 34704 23656 34756 23662
rect 34704 23598 34756 23604
rect 34612 23112 34664 23118
rect 34612 23054 34664 23060
rect 34716 22778 34744 23598
rect 34808 23066 34836 25638
rect 34934 25596 35242 25605
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25531 35242 25540
rect 36004 25226 36032 26250
rect 36648 25906 36676 26250
rect 36636 25900 36688 25906
rect 36636 25842 36688 25848
rect 35992 25220 36044 25226
rect 35992 25162 36044 25168
rect 35594 25052 35902 25061
rect 35594 25050 35600 25052
rect 35656 25050 35680 25052
rect 35736 25050 35760 25052
rect 35816 25050 35840 25052
rect 35896 25050 35902 25052
rect 35656 24998 35658 25050
rect 35838 24998 35840 25050
rect 35594 24996 35600 24998
rect 35656 24996 35680 24998
rect 35736 24996 35760 24998
rect 35816 24996 35840 24998
rect 35896 24996 35902 24998
rect 35594 24987 35902 24996
rect 34934 24508 35242 24517
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24443 35242 24452
rect 35594 23964 35902 23973
rect 35594 23962 35600 23964
rect 35656 23962 35680 23964
rect 35736 23962 35760 23964
rect 35816 23962 35840 23964
rect 35896 23962 35902 23964
rect 35656 23910 35658 23962
rect 35838 23910 35840 23962
rect 35594 23908 35600 23910
rect 35656 23908 35680 23910
rect 35736 23908 35760 23910
rect 35816 23908 35840 23910
rect 35896 23908 35902 23910
rect 35594 23899 35902 23908
rect 35532 23724 35584 23730
rect 35532 23666 35584 23672
rect 35440 23588 35492 23594
rect 35440 23530 35492 23536
rect 34934 23420 35242 23429
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23355 35242 23364
rect 35452 23322 35480 23530
rect 35440 23316 35492 23322
rect 35440 23258 35492 23264
rect 35164 23248 35216 23254
rect 35162 23216 35164 23225
rect 35216 23216 35218 23225
rect 35162 23151 35218 23160
rect 35544 23118 35572 23666
rect 36084 23248 36136 23254
rect 36082 23216 36084 23225
rect 36136 23216 36138 23225
rect 35992 23180 36044 23186
rect 36082 23151 36138 23160
rect 35992 23122 36044 23128
rect 34980 23112 35032 23118
rect 34808 23038 34928 23066
rect 35532 23112 35584 23118
rect 34980 23054 35032 23060
rect 35268 23060 35532 23066
rect 35268 23054 35584 23060
rect 34900 22982 34928 23038
rect 34796 22976 34848 22982
rect 34796 22918 34848 22924
rect 34888 22976 34940 22982
rect 34888 22918 34940 22924
rect 34704 22772 34756 22778
rect 34704 22714 34756 22720
rect 34428 22636 34480 22642
rect 34428 22578 34480 22584
rect 33508 22024 33560 22030
rect 33508 21966 33560 21972
rect 34440 21962 34468 22578
rect 34808 22438 34836 22918
rect 34992 22642 35020 23054
rect 35268 23050 35572 23054
rect 35256 23044 35572 23050
rect 35308 23038 35572 23044
rect 35256 22986 35308 22992
rect 35440 22976 35492 22982
rect 35440 22918 35492 22924
rect 35452 22778 35480 22918
rect 35594 22876 35902 22885
rect 35594 22874 35600 22876
rect 35656 22874 35680 22876
rect 35736 22874 35760 22876
rect 35816 22874 35840 22876
rect 35896 22874 35902 22876
rect 35656 22822 35658 22874
rect 35838 22822 35840 22874
rect 35594 22820 35600 22822
rect 35656 22820 35680 22822
rect 35736 22820 35760 22822
rect 35816 22820 35840 22822
rect 35896 22820 35902 22822
rect 35594 22811 35902 22820
rect 35348 22772 35400 22778
rect 35348 22714 35400 22720
rect 35440 22772 35492 22778
rect 35440 22714 35492 22720
rect 34980 22636 35032 22642
rect 34980 22578 35032 22584
rect 34796 22432 34848 22438
rect 34796 22374 34848 22380
rect 34808 22030 34836 22374
rect 34934 22332 35242 22341
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22267 35242 22276
rect 35164 22092 35216 22098
rect 35164 22034 35216 22040
rect 35256 22092 35308 22098
rect 35256 22034 35308 22040
rect 34796 22024 34848 22030
rect 34796 21966 34848 21972
rect 34428 21956 34480 21962
rect 34428 21898 34480 21904
rect 33324 21888 33376 21894
rect 33324 21830 33376 21836
rect 34704 21888 34756 21894
rect 34704 21830 34756 21836
rect 33336 21554 33364 21830
rect 34716 21690 34744 21830
rect 35176 21690 35204 22034
rect 34704 21684 34756 21690
rect 34704 21626 34756 21632
rect 35164 21684 35216 21690
rect 35164 21626 35216 21632
rect 33324 21548 33376 21554
rect 33324 21490 33376 21496
rect 33508 21548 33560 21554
rect 33508 21490 33560 21496
rect 33600 21548 33652 21554
rect 33600 21490 33652 21496
rect 33520 21350 33548 21490
rect 33232 21344 33284 21350
rect 33232 21286 33284 21292
rect 33508 21344 33560 21350
rect 33508 21286 33560 21292
rect 33244 20398 33272 21286
rect 33612 21146 33640 21490
rect 35268 21486 35296 22034
rect 35360 21690 35388 22714
rect 36004 22710 36032 23122
rect 36084 22976 36136 22982
rect 36084 22918 36136 22924
rect 35992 22704 36044 22710
rect 35992 22646 36044 22652
rect 35440 22636 35492 22642
rect 35440 22578 35492 22584
rect 35348 21684 35400 21690
rect 35348 21626 35400 21632
rect 35452 21570 35480 22578
rect 36096 22522 36124 22918
rect 36096 22494 36216 22522
rect 36084 22432 36136 22438
rect 36084 22374 36136 22380
rect 36096 22250 36124 22374
rect 36004 22222 36124 22250
rect 35594 21788 35902 21797
rect 35594 21786 35600 21788
rect 35656 21786 35680 21788
rect 35736 21786 35760 21788
rect 35816 21786 35840 21788
rect 35896 21786 35902 21788
rect 35656 21734 35658 21786
rect 35838 21734 35840 21786
rect 35594 21732 35600 21734
rect 35656 21732 35680 21734
rect 35736 21732 35760 21734
rect 35816 21732 35840 21734
rect 35896 21732 35902 21734
rect 35594 21723 35902 21732
rect 35624 21616 35676 21622
rect 35452 21554 35572 21570
rect 35624 21558 35676 21564
rect 35452 21548 35584 21554
rect 35452 21542 35532 21548
rect 35532 21490 35584 21496
rect 35256 21480 35308 21486
rect 35256 21422 35308 21428
rect 34934 21244 35242 21253
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21179 35242 21188
rect 33600 21140 33652 21146
rect 33600 21082 33652 21088
rect 35256 21140 35308 21146
rect 35256 21082 35308 21088
rect 33232 20392 33284 20398
rect 33232 20334 33284 20340
rect 33140 20324 33192 20330
rect 33140 20266 33192 20272
rect 33152 19922 33180 20266
rect 33416 19984 33468 19990
rect 33416 19926 33468 19932
rect 33140 19916 33192 19922
rect 33140 19858 33192 19864
rect 33048 19848 33100 19854
rect 33048 19790 33100 19796
rect 33060 19446 33088 19790
rect 33048 19440 33100 19446
rect 33048 19382 33100 19388
rect 33152 19378 33180 19858
rect 33428 19718 33456 19926
rect 33416 19712 33468 19718
rect 33416 19654 33468 19660
rect 33140 19372 33192 19378
rect 33140 19314 33192 19320
rect 33140 19168 33192 19174
rect 33140 19110 33192 19116
rect 33152 18834 33180 19110
rect 33140 18828 33192 18834
rect 33140 18770 33192 18776
rect 33048 18760 33100 18766
rect 32968 18720 33048 18748
rect 33048 18702 33100 18708
rect 33060 18630 33088 18702
rect 33048 18624 33100 18630
rect 33048 18566 33100 18572
rect 33140 18624 33192 18630
rect 33140 18566 33192 18572
rect 33152 18358 33180 18566
rect 33140 18352 33192 18358
rect 33612 18329 33640 21082
rect 35070 21040 35126 21049
rect 35070 20975 35126 20984
rect 35084 20942 35112 20975
rect 35268 20942 35296 21082
rect 35072 20936 35124 20942
rect 35072 20878 35124 20884
rect 35256 20936 35308 20942
rect 35544 20890 35572 21490
rect 35636 21146 35664 21558
rect 35716 21344 35768 21350
rect 35716 21286 35768 21292
rect 35624 21140 35676 21146
rect 35624 21082 35676 21088
rect 35728 21078 35756 21286
rect 35716 21072 35768 21078
rect 35714 21040 35716 21049
rect 35768 21040 35770 21049
rect 35714 20975 35770 20984
rect 35256 20878 35308 20884
rect 34520 20868 34572 20874
rect 34520 20810 34572 20816
rect 35452 20862 35572 20890
rect 34532 20754 34560 20810
rect 34440 20726 34560 20754
rect 34440 20534 34468 20726
rect 35452 20602 35480 20862
rect 35594 20700 35902 20709
rect 35594 20698 35600 20700
rect 35656 20698 35680 20700
rect 35736 20698 35760 20700
rect 35816 20698 35840 20700
rect 35896 20698 35902 20700
rect 35656 20646 35658 20698
rect 35838 20646 35840 20698
rect 35594 20644 35600 20646
rect 35656 20644 35680 20646
rect 35736 20644 35760 20646
rect 35816 20644 35840 20646
rect 35896 20644 35902 20646
rect 35594 20635 35902 20644
rect 35440 20596 35492 20602
rect 35440 20538 35492 20544
rect 34428 20528 34480 20534
rect 34428 20470 34480 20476
rect 35900 20460 35952 20466
rect 36004 20448 36032 22222
rect 36084 22094 36136 22098
rect 36188 22094 36216 22494
rect 36452 22432 36504 22438
rect 36452 22374 36504 22380
rect 36268 22228 36320 22234
rect 36268 22170 36320 22176
rect 36084 22092 36216 22094
rect 36136 22066 36216 22092
rect 36084 22034 36136 22040
rect 36280 21554 36308 22170
rect 36464 22098 36492 22374
rect 36452 22092 36504 22098
rect 36648 22094 36676 25842
rect 36728 25220 36780 25226
rect 36728 25162 36780 25168
rect 36740 24954 36768 25162
rect 36728 24948 36780 24954
rect 36728 24890 36780 24896
rect 36648 22066 36768 22094
rect 36452 22034 36504 22040
rect 36360 21888 36412 21894
rect 36360 21830 36412 21836
rect 36372 21554 36400 21830
rect 36464 21554 36492 22034
rect 36268 21548 36320 21554
rect 36268 21490 36320 21496
rect 36360 21548 36412 21554
rect 36360 21490 36412 21496
rect 36452 21548 36504 21554
rect 36452 21490 36504 21496
rect 36176 21480 36228 21486
rect 36176 21422 36228 21428
rect 35952 20420 36032 20448
rect 35900 20402 35952 20408
rect 34428 20392 34480 20398
rect 34428 20334 34480 20340
rect 35808 20392 35860 20398
rect 35808 20334 35860 20340
rect 34152 19372 34204 19378
rect 34152 19314 34204 19320
rect 33968 18760 34020 18766
rect 33968 18702 34020 18708
rect 33140 18294 33192 18300
rect 33598 18320 33654 18329
rect 33598 18255 33654 18264
rect 32956 17672 33008 17678
rect 32956 17614 33008 17620
rect 32864 17332 32916 17338
rect 32864 17274 32916 17280
rect 32968 16998 32996 17614
rect 33612 17524 33640 18255
rect 33980 18086 34008 18702
rect 34164 18426 34192 19314
rect 34440 19242 34468 20334
rect 34520 20324 34572 20330
rect 34520 20266 34572 20272
rect 34428 19236 34480 19242
rect 34428 19178 34480 19184
rect 34440 18970 34468 19178
rect 34428 18964 34480 18970
rect 34428 18906 34480 18912
rect 34152 18420 34204 18426
rect 34152 18362 34204 18368
rect 33968 18080 34020 18086
rect 33968 18022 34020 18028
rect 33980 17678 34008 18022
rect 34060 17808 34112 17814
rect 34060 17750 34112 17756
rect 33968 17672 34020 17678
rect 33968 17614 34020 17620
rect 33784 17536 33836 17542
rect 33612 17496 33784 17524
rect 33784 17478 33836 17484
rect 33048 17332 33100 17338
rect 33048 17274 33100 17280
rect 32956 16992 33008 16998
rect 32956 16934 33008 16940
rect 32772 16516 32824 16522
rect 32772 16458 32824 16464
rect 32496 15904 32548 15910
rect 32496 15846 32548 15852
rect 32508 15706 32536 15846
rect 32496 15700 32548 15706
rect 32496 15642 32548 15648
rect 32404 13864 32456 13870
rect 32404 13806 32456 13812
rect 32416 13530 32444 13806
rect 32404 13524 32456 13530
rect 32404 13466 32456 13472
rect 32404 13252 32456 13258
rect 32404 13194 32456 13200
rect 32416 12850 32444 13194
rect 32404 12844 32456 12850
rect 32404 12786 32456 12792
rect 32508 12782 32536 15642
rect 32588 15360 32640 15366
rect 32588 15302 32640 15308
rect 32600 15162 32628 15302
rect 32588 15156 32640 15162
rect 32588 15098 32640 15104
rect 32588 13796 32640 13802
rect 32588 13738 32640 13744
rect 32600 13258 32628 13738
rect 32588 13252 32640 13258
rect 32588 13194 32640 13200
rect 32496 12776 32548 12782
rect 32496 12718 32548 12724
rect 32508 12434 32536 12718
rect 32416 12406 32536 12434
rect 32312 12300 32364 12306
rect 32312 12242 32364 12248
rect 32220 11688 32272 11694
rect 32220 11630 32272 11636
rect 32128 11348 32180 11354
rect 32128 11290 32180 11296
rect 31760 11280 31812 11286
rect 31760 11222 31812 11228
rect 31852 11144 31904 11150
rect 31852 11086 31904 11092
rect 31864 10674 31892 11086
rect 32128 10804 32180 10810
rect 32128 10746 32180 10752
rect 31852 10668 31904 10674
rect 31852 10610 31904 10616
rect 31576 9376 31628 9382
rect 31576 9318 31628 9324
rect 31668 9376 31720 9382
rect 31668 9318 31720 9324
rect 31588 9178 31616 9318
rect 31576 9172 31628 9178
rect 31576 9114 31628 9120
rect 31680 9058 31708 9318
rect 31588 9030 31708 9058
rect 31484 8084 31536 8090
rect 31484 8026 31536 8032
rect 31116 7744 31168 7750
rect 31116 7686 31168 7692
rect 31208 7744 31260 7750
rect 31208 7686 31260 7692
rect 31220 7546 31248 7686
rect 31208 7540 31260 7546
rect 31208 7482 31260 7488
rect 31588 7478 31616 9030
rect 31864 8974 31892 10610
rect 32140 10554 32168 10746
rect 32232 10674 32260 11630
rect 32312 11144 32364 11150
rect 32312 11086 32364 11092
rect 32324 10810 32352 11086
rect 32312 10804 32364 10810
rect 32312 10746 32364 10752
rect 32220 10668 32272 10674
rect 32220 10610 32272 10616
rect 32416 10554 32444 12406
rect 32600 12102 32628 13194
rect 32784 12442 32812 16458
rect 32864 15700 32916 15706
rect 32864 15642 32916 15648
rect 32876 15502 32904 15642
rect 32864 15496 32916 15502
rect 32864 15438 32916 15444
rect 32876 14074 32904 15438
rect 33060 15026 33088 17274
rect 33796 17270 33824 17478
rect 33980 17338 34008 17614
rect 33968 17332 34020 17338
rect 33968 17274 34020 17280
rect 33784 17264 33836 17270
rect 33784 17206 33836 17212
rect 33416 15496 33468 15502
rect 33416 15438 33468 15444
rect 33048 15020 33100 15026
rect 33048 14962 33100 14968
rect 32956 14952 33008 14958
rect 32956 14894 33008 14900
rect 32968 14618 32996 14894
rect 32956 14612 33008 14618
rect 32956 14554 33008 14560
rect 32864 14068 32916 14074
rect 32864 14010 32916 14016
rect 32956 13932 33008 13938
rect 32956 13874 33008 13880
rect 33232 13932 33284 13938
rect 33232 13874 33284 13880
rect 32864 13320 32916 13326
rect 32864 13262 32916 13268
rect 32968 13274 32996 13874
rect 33140 13728 33192 13734
rect 33140 13670 33192 13676
rect 33152 13326 33180 13670
rect 33244 13530 33272 13874
rect 33428 13530 33456 15438
rect 33796 14482 33824 17206
rect 34072 17134 34100 17750
rect 34532 17270 34560 20266
rect 34796 20256 34848 20262
rect 34796 20198 34848 20204
rect 34612 19780 34664 19786
rect 34612 19722 34664 19728
rect 34704 19780 34756 19786
rect 34704 19722 34756 19728
rect 34520 17264 34572 17270
rect 34520 17206 34572 17212
rect 34532 17134 34560 17206
rect 34060 17128 34112 17134
rect 34060 17070 34112 17076
rect 34520 17128 34572 17134
rect 34520 17070 34572 17076
rect 34520 16992 34572 16998
rect 34520 16934 34572 16940
rect 34532 15570 34560 16934
rect 34520 15564 34572 15570
rect 34520 15506 34572 15512
rect 34624 15502 34652 19722
rect 34716 16998 34744 19722
rect 34808 19718 34836 20198
rect 34934 20156 35242 20165
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20091 35242 20100
rect 35820 20058 35848 20334
rect 35808 20052 35860 20058
rect 35808 19994 35860 20000
rect 35164 19984 35216 19990
rect 35346 19952 35402 19961
rect 35164 19926 35216 19932
rect 35176 19854 35204 19926
rect 35268 19910 35346 19938
rect 35268 19854 35296 19910
rect 36188 19922 36216 21422
rect 35716 19916 35768 19922
rect 35346 19887 35402 19896
rect 35636 19876 35716 19904
rect 35164 19848 35216 19854
rect 35164 19790 35216 19796
rect 35256 19848 35308 19854
rect 35440 19848 35492 19854
rect 35256 19790 35308 19796
rect 35360 19808 35440 19836
rect 34796 19712 34848 19718
rect 34796 19654 34848 19660
rect 34808 19514 34836 19654
rect 34796 19508 34848 19514
rect 34796 19450 34848 19456
rect 34796 19304 34848 19310
rect 34796 19246 34848 19252
rect 34808 18850 34836 19246
rect 34934 19068 35242 19077
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 19003 35242 19012
rect 34808 18822 35020 18850
rect 35360 18834 35388 19808
rect 35440 19790 35492 19796
rect 35636 19700 35664 19876
rect 35716 19858 35768 19864
rect 36176 19916 36228 19922
rect 36176 19858 36228 19864
rect 35992 19848 36044 19854
rect 35992 19790 36044 19796
rect 35452 19672 35664 19700
rect 34992 18630 35020 18822
rect 35348 18828 35400 18834
rect 35348 18770 35400 18776
rect 34796 18624 34848 18630
rect 34796 18566 34848 18572
rect 34980 18624 35032 18630
rect 34980 18566 35032 18572
rect 35164 18624 35216 18630
rect 35164 18566 35216 18572
rect 34808 18426 34836 18566
rect 34796 18420 34848 18426
rect 34796 18362 34848 18368
rect 34992 18290 35020 18566
rect 35176 18290 35204 18566
rect 35452 18358 35480 19672
rect 35594 19612 35902 19621
rect 35594 19610 35600 19612
rect 35656 19610 35680 19612
rect 35736 19610 35760 19612
rect 35816 19610 35840 19612
rect 35896 19610 35902 19612
rect 35656 19558 35658 19610
rect 35838 19558 35840 19610
rect 35594 19556 35600 19558
rect 35656 19556 35680 19558
rect 35736 19556 35760 19558
rect 35816 19556 35840 19558
rect 35896 19556 35902 19558
rect 35594 19547 35902 19556
rect 36004 19394 36032 19790
rect 36084 19712 36136 19718
rect 36084 19654 36136 19660
rect 36096 19514 36124 19654
rect 36084 19508 36136 19514
rect 36084 19450 36136 19456
rect 36280 19394 36308 21490
rect 36372 19990 36400 21490
rect 36360 19984 36412 19990
rect 36360 19926 36412 19932
rect 36450 19952 36506 19961
rect 36450 19887 36452 19896
rect 36504 19887 36506 19896
rect 36452 19858 36504 19864
rect 36004 19366 36308 19394
rect 36004 19174 36032 19366
rect 35992 19168 36044 19174
rect 35992 19110 36044 19116
rect 36740 18834 36768 22066
rect 36832 21593 36860 29106
rect 37280 29028 37332 29034
rect 37280 28970 37332 28976
rect 37292 28218 37320 28970
rect 37280 28212 37332 28218
rect 37280 28154 37332 28160
rect 37556 27872 37608 27878
rect 37556 27814 37608 27820
rect 37568 22642 37596 27814
rect 37556 22636 37608 22642
rect 37556 22578 37608 22584
rect 37830 22536 37886 22545
rect 37830 22471 37832 22480
rect 37884 22471 37886 22480
rect 37832 22442 37884 22448
rect 37004 22432 37056 22438
rect 37004 22374 37056 22380
rect 37016 22094 37044 22374
rect 36924 22066 37044 22094
rect 36924 22030 36952 22066
rect 36912 22024 36964 22030
rect 36912 21966 36964 21972
rect 36818 21584 36874 21593
rect 36818 21519 36874 21528
rect 36728 18828 36780 18834
rect 36728 18770 36780 18776
rect 36832 18698 36860 21519
rect 37280 21480 37332 21486
rect 37280 21422 37332 21428
rect 36820 18692 36872 18698
rect 36820 18634 36872 18640
rect 35594 18524 35902 18533
rect 35594 18522 35600 18524
rect 35656 18522 35680 18524
rect 35736 18522 35760 18524
rect 35816 18522 35840 18524
rect 35896 18522 35902 18524
rect 35656 18470 35658 18522
rect 35838 18470 35840 18522
rect 35594 18468 35600 18470
rect 35656 18468 35680 18470
rect 35736 18468 35760 18470
rect 35816 18468 35840 18470
rect 35896 18468 35902 18470
rect 35594 18459 35902 18468
rect 35440 18352 35492 18358
rect 35440 18294 35492 18300
rect 34980 18284 35032 18290
rect 34980 18226 35032 18232
rect 35164 18284 35216 18290
rect 35164 18226 35216 18232
rect 34934 17980 35242 17989
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17915 35242 17924
rect 35594 17436 35902 17445
rect 35594 17434 35600 17436
rect 35656 17434 35680 17436
rect 35736 17434 35760 17436
rect 35816 17434 35840 17436
rect 35896 17434 35902 17436
rect 35656 17382 35658 17434
rect 35838 17382 35840 17434
rect 35594 17380 35600 17382
rect 35656 17380 35680 17382
rect 35736 17380 35760 17382
rect 35816 17380 35840 17382
rect 35896 17380 35902 17382
rect 35594 17371 35902 17380
rect 34704 16992 34756 16998
rect 34704 16934 34756 16940
rect 34796 16992 34848 16998
rect 34796 16934 34848 16940
rect 35348 16992 35400 16998
rect 35348 16934 35400 16940
rect 34704 16652 34756 16658
rect 34704 16594 34756 16600
rect 34716 15706 34744 16594
rect 34808 16522 34836 16934
rect 34934 16892 35242 16901
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16827 35242 16836
rect 35360 16810 35388 16934
rect 35268 16794 35388 16810
rect 35256 16788 35388 16794
rect 35308 16782 35388 16788
rect 35440 16788 35492 16794
rect 35256 16730 35308 16736
rect 35440 16730 35492 16736
rect 35072 16584 35124 16590
rect 35072 16526 35124 16532
rect 34796 16516 34848 16522
rect 34796 16458 34848 16464
rect 34808 16250 34836 16458
rect 35084 16250 35112 16526
rect 35164 16448 35216 16454
rect 35164 16390 35216 16396
rect 34796 16244 34848 16250
rect 34796 16186 34848 16192
rect 35072 16244 35124 16250
rect 35072 16186 35124 16192
rect 35084 15978 35112 16186
rect 35176 16114 35204 16390
rect 35164 16108 35216 16114
rect 35164 16050 35216 16056
rect 35268 16046 35296 16730
rect 35452 16250 35480 16730
rect 35594 16348 35902 16357
rect 35594 16346 35600 16348
rect 35656 16346 35680 16348
rect 35736 16346 35760 16348
rect 35816 16346 35840 16348
rect 35896 16346 35902 16348
rect 35656 16294 35658 16346
rect 35838 16294 35840 16346
rect 35594 16292 35600 16294
rect 35656 16292 35680 16294
rect 35736 16292 35760 16294
rect 35816 16292 35840 16294
rect 35896 16292 35902 16294
rect 35594 16283 35902 16292
rect 35440 16244 35492 16250
rect 35440 16186 35492 16192
rect 35256 16040 35308 16046
rect 35256 15982 35308 15988
rect 35072 15972 35124 15978
rect 35072 15914 35124 15920
rect 35348 15904 35400 15910
rect 35348 15846 35400 15852
rect 34934 15804 35242 15813
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15739 35242 15748
rect 35360 15706 35388 15846
rect 34704 15700 34756 15706
rect 34704 15642 34756 15648
rect 35348 15700 35400 15706
rect 35348 15642 35400 15648
rect 34796 15564 34848 15570
rect 34796 15506 34848 15512
rect 35348 15564 35400 15570
rect 35348 15506 35400 15512
rect 34612 15496 34664 15502
rect 34612 15438 34664 15444
rect 34808 15162 34836 15506
rect 34796 15156 34848 15162
rect 34796 15098 34848 15104
rect 34934 14716 35242 14725
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14651 35242 14660
rect 33784 14476 33836 14482
rect 33784 14418 33836 14424
rect 34060 14408 34112 14414
rect 34060 14350 34112 14356
rect 33508 13728 33560 13734
rect 33508 13670 33560 13676
rect 33232 13524 33284 13530
rect 33232 13466 33284 13472
rect 33416 13524 33468 13530
rect 33416 13466 33468 13472
rect 33520 13326 33548 13670
rect 33140 13320 33192 13326
rect 32876 12986 32904 13262
rect 32968 13258 33088 13274
rect 33140 13262 33192 13268
rect 33508 13320 33560 13326
rect 33508 13262 33560 13268
rect 33876 13320 33928 13326
rect 33876 13262 33928 13268
rect 32968 13252 33100 13258
rect 32968 13246 33048 13252
rect 33048 13194 33100 13200
rect 32864 12980 32916 12986
rect 32864 12922 32916 12928
rect 32772 12436 32824 12442
rect 32772 12378 32824 12384
rect 32680 12368 32732 12374
rect 32680 12310 32732 12316
rect 32588 12096 32640 12102
rect 32588 12038 32640 12044
rect 32692 11762 32720 12310
rect 32956 12232 33008 12238
rect 32956 12174 33008 12180
rect 32588 11756 32640 11762
rect 32588 11698 32640 11704
rect 32680 11756 32732 11762
rect 32680 11698 32732 11704
rect 32496 11144 32548 11150
rect 32496 11086 32548 11092
rect 32508 10606 32536 11086
rect 32600 10810 32628 11698
rect 32692 10810 32720 11698
rect 32772 11144 32824 11150
rect 32772 11086 32824 11092
rect 32588 10804 32640 10810
rect 32588 10746 32640 10752
rect 32680 10804 32732 10810
rect 32680 10746 32732 10752
rect 32784 10674 32812 11086
rect 32864 11008 32916 11014
rect 32864 10950 32916 10956
rect 32968 10962 32996 12174
rect 33060 11898 33088 13194
rect 33152 12986 33180 13262
rect 33140 12980 33192 12986
rect 33140 12922 33192 12928
rect 33888 12850 33916 13262
rect 33876 12844 33928 12850
rect 33876 12786 33928 12792
rect 33324 12776 33376 12782
rect 33324 12718 33376 12724
rect 33048 11892 33100 11898
rect 33048 11834 33100 11840
rect 33060 11150 33088 11834
rect 33048 11144 33100 11150
rect 33048 11086 33100 11092
rect 32772 10668 32824 10674
rect 32772 10610 32824 10616
rect 32140 10526 32444 10554
rect 32496 10600 32548 10606
rect 32496 10542 32548 10548
rect 32036 9444 32088 9450
rect 32036 9386 32088 9392
rect 32048 9042 32076 9386
rect 32036 9036 32088 9042
rect 32036 8978 32088 8984
rect 31760 8968 31812 8974
rect 31760 8910 31812 8916
rect 31852 8968 31904 8974
rect 31852 8910 31904 8916
rect 31668 8492 31720 8498
rect 31668 8434 31720 8440
rect 31680 7818 31708 8434
rect 31772 8090 31800 8910
rect 31944 8832 31996 8838
rect 31944 8774 31996 8780
rect 31956 8566 31984 8774
rect 32048 8634 32076 8978
rect 32036 8628 32088 8634
rect 32036 8570 32088 8576
rect 31944 8560 31996 8566
rect 31944 8502 31996 8508
rect 31760 8084 31812 8090
rect 31760 8026 31812 8032
rect 31668 7812 31720 7818
rect 31668 7754 31720 7760
rect 31576 7472 31628 7478
rect 31576 7414 31628 7420
rect 31772 7410 31800 8026
rect 31392 7404 31444 7410
rect 31392 7346 31444 7352
rect 31760 7404 31812 7410
rect 31760 7346 31812 7352
rect 31300 7336 31352 7342
rect 31300 7278 31352 7284
rect 31312 7002 31340 7278
rect 31404 7002 31432 7346
rect 31956 7002 31984 8502
rect 31300 6996 31352 7002
rect 31300 6938 31352 6944
rect 31392 6996 31444 7002
rect 31392 6938 31444 6944
rect 31944 6996 31996 7002
rect 31944 6938 31996 6944
rect 32140 6798 32168 10526
rect 32784 10266 32812 10610
rect 32772 10260 32824 10266
rect 32772 10202 32824 10208
rect 32784 9586 32812 10202
rect 32876 10062 32904 10950
rect 32968 10934 33088 10962
rect 32956 10464 33008 10470
rect 32956 10406 33008 10412
rect 32968 10130 32996 10406
rect 32956 10124 33008 10130
rect 32956 10066 33008 10072
rect 32864 10056 32916 10062
rect 32864 9998 32916 10004
rect 32876 9674 32904 9998
rect 32876 9646 32996 9674
rect 33060 9654 33088 10934
rect 33232 10736 33284 10742
rect 33232 10678 33284 10684
rect 33140 9716 33192 9722
rect 33140 9658 33192 9664
rect 32772 9580 32824 9586
rect 32772 9522 32824 9528
rect 32772 8968 32824 8974
rect 32772 8910 32824 8916
rect 32968 8956 32996 9646
rect 33048 9648 33100 9654
rect 33048 9590 33100 9596
rect 33152 9178 33180 9658
rect 33244 9382 33272 10678
rect 33232 9376 33284 9382
rect 33232 9318 33284 9324
rect 33140 9172 33192 9178
rect 33140 9114 33192 9120
rect 33244 9058 33272 9318
rect 33336 9178 33364 12718
rect 33600 12232 33652 12238
rect 33600 12174 33652 12180
rect 33612 10742 33640 12174
rect 33600 10736 33652 10742
rect 33600 10678 33652 10684
rect 33508 10668 33560 10674
rect 33508 10610 33560 10616
rect 33520 10266 33548 10610
rect 33508 10260 33560 10266
rect 33508 10202 33560 10208
rect 34072 10062 34100 14350
rect 34934 13628 35242 13637
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13563 35242 13572
rect 34934 12540 35242 12549
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12475 35242 12484
rect 34612 11620 34664 11626
rect 34612 11562 34664 11568
rect 34624 11354 34652 11562
rect 34934 11452 35242 11461
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11387 35242 11396
rect 34612 11348 34664 11354
rect 34612 11290 34664 11296
rect 35360 10810 35388 15506
rect 35594 15260 35902 15269
rect 35594 15258 35600 15260
rect 35656 15258 35680 15260
rect 35736 15258 35760 15260
rect 35816 15258 35840 15260
rect 35896 15258 35902 15260
rect 35656 15206 35658 15258
rect 35838 15206 35840 15258
rect 35594 15204 35600 15206
rect 35656 15204 35680 15206
rect 35736 15204 35760 15206
rect 35816 15204 35840 15206
rect 35896 15204 35902 15206
rect 35594 15195 35902 15204
rect 35594 14172 35902 14181
rect 35594 14170 35600 14172
rect 35656 14170 35680 14172
rect 35736 14170 35760 14172
rect 35816 14170 35840 14172
rect 35896 14170 35902 14172
rect 35656 14118 35658 14170
rect 35838 14118 35840 14170
rect 35594 14116 35600 14118
rect 35656 14116 35680 14118
rect 35736 14116 35760 14118
rect 35816 14116 35840 14118
rect 35896 14116 35902 14118
rect 35594 14107 35902 14116
rect 35594 13084 35902 13093
rect 35594 13082 35600 13084
rect 35656 13082 35680 13084
rect 35736 13082 35760 13084
rect 35816 13082 35840 13084
rect 35896 13082 35902 13084
rect 35656 13030 35658 13082
rect 35838 13030 35840 13082
rect 35594 13028 35600 13030
rect 35656 13028 35680 13030
rect 35736 13028 35760 13030
rect 35816 13028 35840 13030
rect 35896 13028 35902 13030
rect 35594 13019 35902 13028
rect 35594 11996 35902 12005
rect 35594 11994 35600 11996
rect 35656 11994 35680 11996
rect 35736 11994 35760 11996
rect 35816 11994 35840 11996
rect 35896 11994 35902 11996
rect 35656 11942 35658 11994
rect 35838 11942 35840 11994
rect 35594 11940 35600 11942
rect 35656 11940 35680 11942
rect 35736 11940 35760 11942
rect 35816 11940 35840 11942
rect 35896 11940 35902 11942
rect 35594 11931 35902 11940
rect 35594 10908 35902 10917
rect 35594 10906 35600 10908
rect 35656 10906 35680 10908
rect 35736 10906 35760 10908
rect 35816 10906 35840 10908
rect 35896 10906 35902 10908
rect 35656 10854 35658 10906
rect 35838 10854 35840 10906
rect 35594 10852 35600 10854
rect 35656 10852 35680 10854
rect 35736 10852 35760 10854
rect 35816 10852 35840 10854
rect 35896 10852 35902 10854
rect 35594 10843 35902 10852
rect 35348 10804 35400 10810
rect 35348 10746 35400 10752
rect 34428 10668 34480 10674
rect 34428 10610 34480 10616
rect 33968 10056 34020 10062
rect 33968 9998 34020 10004
rect 34060 10056 34112 10062
rect 34060 9998 34112 10004
rect 33980 9722 34008 9998
rect 33968 9716 34020 9722
rect 33968 9658 34020 9664
rect 33324 9172 33376 9178
rect 33324 9114 33376 9120
rect 33152 9030 33272 9058
rect 33152 8974 33180 9030
rect 33048 8968 33100 8974
rect 32968 8928 33048 8956
rect 32784 8634 32812 8910
rect 32864 8900 32916 8906
rect 32864 8842 32916 8848
rect 32772 8628 32824 8634
rect 32772 8570 32824 8576
rect 32588 8356 32640 8362
rect 32588 8298 32640 8304
rect 32496 6928 32548 6934
rect 32496 6870 32548 6876
rect 31760 6792 31812 6798
rect 31760 6734 31812 6740
rect 31852 6792 31904 6798
rect 31852 6734 31904 6740
rect 32128 6792 32180 6798
rect 32128 6734 32180 6740
rect 32220 6792 32272 6798
rect 32220 6734 32272 6740
rect 31024 6452 31076 6458
rect 31024 6394 31076 6400
rect 30472 5908 30524 5914
rect 30472 5850 30524 5856
rect 31772 5710 31800 6734
rect 31760 5704 31812 5710
rect 31760 5646 31812 5652
rect 31864 5658 31892 6734
rect 32232 6322 32260 6734
rect 32508 6458 32536 6870
rect 32600 6798 32628 8298
rect 32588 6792 32640 6798
rect 32588 6734 32640 6740
rect 32600 6458 32628 6734
rect 32680 6656 32732 6662
rect 32680 6598 32732 6604
rect 32496 6452 32548 6458
rect 32496 6394 32548 6400
rect 32588 6452 32640 6458
rect 32588 6394 32640 6400
rect 32692 6322 32720 6598
rect 32220 6316 32272 6322
rect 32220 6258 32272 6264
rect 32680 6316 32732 6322
rect 32680 6258 32732 6264
rect 32036 6112 32088 6118
rect 32036 6054 32088 6060
rect 32048 5914 32076 6054
rect 32232 5914 32260 6258
rect 32784 6186 32812 8570
rect 32876 6866 32904 8842
rect 32968 8480 32996 8928
rect 33048 8910 33100 8916
rect 33140 8968 33192 8974
rect 33140 8910 33192 8916
rect 33508 8968 33560 8974
rect 33508 8910 33560 8916
rect 33232 8832 33284 8838
rect 33232 8774 33284 8780
rect 33048 8492 33100 8498
rect 32968 8452 33048 8480
rect 33048 8434 33100 8440
rect 33244 8430 33272 8774
rect 33520 8634 33548 8910
rect 33508 8628 33560 8634
rect 33508 8570 33560 8576
rect 33232 8424 33284 8430
rect 33232 8366 33284 8372
rect 33048 8016 33100 8022
rect 33048 7958 33100 7964
rect 32864 6860 32916 6866
rect 32864 6802 32916 6808
rect 33060 6798 33088 7958
rect 34072 7274 34100 9998
rect 34060 7268 34112 7274
rect 34060 7210 34112 7216
rect 33048 6792 33100 6798
rect 33048 6734 33100 6740
rect 34440 6730 34468 10610
rect 34934 10364 35242 10373
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10299 35242 10308
rect 35594 9820 35902 9829
rect 35594 9818 35600 9820
rect 35656 9818 35680 9820
rect 35736 9818 35760 9820
rect 35816 9818 35840 9820
rect 35896 9818 35902 9820
rect 35656 9766 35658 9818
rect 35838 9766 35840 9818
rect 35594 9764 35600 9766
rect 35656 9764 35680 9766
rect 35736 9764 35760 9766
rect 35816 9764 35840 9766
rect 35896 9764 35902 9766
rect 35594 9755 35902 9764
rect 34934 9276 35242 9285
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9211 35242 9220
rect 36832 8906 36860 18634
rect 37096 18624 37148 18630
rect 37096 18566 37148 18572
rect 37108 18426 37136 18566
rect 37096 18420 37148 18426
rect 37096 18362 37148 18368
rect 37292 18358 37320 21422
rect 38384 20732 38436 20738
rect 38384 20674 38436 20680
rect 38396 20505 38424 20674
rect 38382 20496 38438 20505
rect 38382 20431 38438 20440
rect 37280 18352 37332 18358
rect 37280 18294 37332 18300
rect 37556 18080 37608 18086
rect 37556 18022 37608 18028
rect 35992 8900 36044 8906
rect 35992 8842 36044 8848
rect 36820 8900 36872 8906
rect 36820 8842 36872 8848
rect 35594 8732 35902 8741
rect 35594 8730 35600 8732
rect 35656 8730 35680 8732
rect 35736 8730 35760 8732
rect 35816 8730 35840 8732
rect 35896 8730 35902 8732
rect 35656 8678 35658 8730
rect 35838 8678 35840 8730
rect 35594 8676 35600 8678
rect 35656 8676 35680 8678
rect 35736 8676 35760 8678
rect 35816 8676 35840 8678
rect 35896 8676 35902 8678
rect 35594 8667 35902 8676
rect 36004 8566 36032 8842
rect 35992 8560 36044 8566
rect 35992 8502 36044 8508
rect 34934 8188 35242 8197
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8123 35242 8132
rect 35594 7644 35902 7653
rect 35594 7642 35600 7644
rect 35656 7642 35680 7644
rect 35736 7642 35760 7644
rect 35816 7642 35840 7644
rect 35896 7642 35902 7644
rect 35656 7590 35658 7642
rect 35838 7590 35840 7642
rect 35594 7588 35600 7590
rect 35656 7588 35680 7590
rect 35736 7588 35760 7590
rect 35816 7588 35840 7590
rect 35896 7588 35902 7590
rect 35594 7579 35902 7588
rect 34934 7100 35242 7109
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7035 35242 7044
rect 34428 6724 34480 6730
rect 34428 6666 34480 6672
rect 35594 6556 35902 6565
rect 35594 6554 35600 6556
rect 35656 6554 35680 6556
rect 35736 6554 35760 6556
rect 35816 6554 35840 6556
rect 35896 6554 35902 6556
rect 35656 6502 35658 6554
rect 35838 6502 35840 6554
rect 35594 6500 35600 6502
rect 35656 6500 35680 6502
rect 35736 6500 35760 6502
rect 35816 6500 35840 6502
rect 35896 6500 35902 6502
rect 35594 6491 35902 6500
rect 32772 6180 32824 6186
rect 32772 6122 32824 6128
rect 34934 6012 35242 6021
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5947 35242 5956
rect 32036 5908 32088 5914
rect 32036 5850 32088 5856
rect 32220 5908 32272 5914
rect 32220 5850 32272 5856
rect 32128 5704 32180 5710
rect 30196 5636 30248 5642
rect 30196 5578 30248 5584
rect 30288 5636 30340 5642
rect 30288 5578 30340 5584
rect 29460 5568 29512 5574
rect 29460 5510 29512 5516
rect 29368 5296 29420 5302
rect 29368 5238 29420 5244
rect 29184 5092 29236 5098
rect 29184 5034 29236 5040
rect 29196 4826 29224 5034
rect 29184 4820 29236 4826
rect 29184 4762 29236 4768
rect 29380 4758 29408 5238
rect 29472 5234 29500 5510
rect 29736 5364 29788 5370
rect 29788 5324 29868 5352
rect 29736 5306 29788 5312
rect 29840 5234 29868 5324
rect 29460 5228 29512 5234
rect 29460 5170 29512 5176
rect 29828 5228 29880 5234
rect 29828 5170 29880 5176
rect 30104 5228 30156 5234
rect 30104 5170 30156 5176
rect 29828 5092 29880 5098
rect 29828 5034 29880 5040
rect 29368 4752 29420 4758
rect 29368 4694 29420 4700
rect 27988 4684 28040 4690
rect 27988 4626 28040 4632
rect 28080 4684 28132 4690
rect 28080 4626 28132 4632
rect 27712 4480 27764 4486
rect 27712 4422 27764 4428
rect 28000 4282 28028 4626
rect 26332 4276 26384 4282
rect 26332 4218 26384 4224
rect 27988 4276 28040 4282
rect 27988 4218 28040 4224
rect 29840 4214 29868 5034
rect 30012 5024 30064 5030
rect 30012 4966 30064 4972
rect 30024 4826 30052 4966
rect 30012 4820 30064 4826
rect 30012 4762 30064 4768
rect 29828 4208 29880 4214
rect 29828 4150 29880 4156
rect 30116 4146 30144 5170
rect 30208 4622 30236 5578
rect 30300 5370 30328 5578
rect 30288 5364 30340 5370
rect 30288 5306 30340 5312
rect 30380 5296 30432 5302
rect 30380 5238 30432 5244
rect 30288 5024 30340 5030
rect 30288 4966 30340 4972
rect 30300 4826 30328 4966
rect 30288 4820 30340 4826
rect 30288 4762 30340 4768
rect 30392 4622 30420 5238
rect 31772 5234 31800 5646
rect 31864 5642 31984 5658
rect 32128 5646 32180 5652
rect 31864 5636 31996 5642
rect 31864 5630 31944 5636
rect 31944 5578 31996 5584
rect 31760 5228 31812 5234
rect 31760 5170 31812 5176
rect 30656 5092 30708 5098
rect 30656 5034 30708 5040
rect 30196 4616 30248 4622
rect 30196 4558 30248 4564
rect 30380 4616 30432 4622
rect 30380 4558 30432 4564
rect 30668 4214 30696 5034
rect 31956 4486 31984 5578
rect 32140 5370 32168 5646
rect 35594 5468 35902 5477
rect 35594 5466 35600 5468
rect 35656 5466 35680 5468
rect 35736 5466 35760 5468
rect 35816 5466 35840 5468
rect 35896 5466 35902 5468
rect 35656 5414 35658 5466
rect 35838 5414 35840 5466
rect 35594 5412 35600 5414
rect 35656 5412 35680 5414
rect 35736 5412 35760 5414
rect 35816 5412 35840 5414
rect 35896 5412 35902 5414
rect 35594 5403 35902 5412
rect 32128 5364 32180 5370
rect 32128 5306 32180 5312
rect 34934 4924 35242 4933
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4859 35242 4868
rect 31944 4480 31996 4486
rect 31944 4422 31996 4428
rect 35594 4380 35902 4389
rect 35594 4378 35600 4380
rect 35656 4378 35680 4380
rect 35736 4378 35760 4380
rect 35816 4378 35840 4380
rect 35896 4378 35902 4380
rect 35656 4326 35658 4378
rect 35838 4326 35840 4378
rect 35594 4324 35600 4326
rect 35656 4324 35680 4326
rect 35736 4324 35760 4326
rect 35816 4324 35840 4326
rect 35896 4324 35902 4326
rect 35594 4315 35902 4324
rect 30656 4208 30708 4214
rect 30656 4150 30708 4156
rect 30104 4140 30156 4146
rect 30104 4082 30156 4088
rect 34934 3836 35242 3845
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3771 35242 3780
rect 35594 3292 35902 3301
rect 35594 3290 35600 3292
rect 35656 3290 35680 3292
rect 35736 3290 35760 3292
rect 35816 3290 35840 3292
rect 35896 3290 35902 3292
rect 35656 3238 35658 3290
rect 35838 3238 35840 3290
rect 35594 3236 35600 3238
rect 35656 3236 35680 3238
rect 35736 3236 35760 3238
rect 35816 3236 35840 3238
rect 35896 3236 35902 3238
rect 35594 3227 35902 3236
rect 37568 3126 37596 18022
rect 38384 18012 38436 18018
rect 38384 17954 38436 17960
rect 38396 17785 38424 17954
rect 38382 17776 38438 17785
rect 38382 17711 38438 17720
rect 37832 15904 37884 15910
rect 37832 15846 37884 15852
rect 37844 15745 37872 15846
rect 37830 15736 37886 15745
rect 37830 15671 37886 15680
rect 37924 11076 37976 11082
rect 37924 11018 37976 11024
rect 37936 10985 37964 11018
rect 37922 10976 37978 10985
rect 37922 10911 37978 10920
rect 38292 8968 38344 8974
rect 38290 8936 38292 8945
rect 38344 8936 38346 8945
rect 38290 8871 38346 8880
rect 37556 3120 37608 3126
rect 37556 3062 37608 3068
rect 15108 3052 15160 3058
rect 15108 2994 15160 3000
rect 25596 3052 25648 3058
rect 25596 2994 25648 3000
rect 14924 2848 14976 2854
rect 14924 2790 14976 2796
rect 17408 2848 17460 2854
rect 17408 2790 17460 2796
rect 19800 2848 19852 2854
rect 19800 2790 19852 2796
rect 37188 2848 37240 2854
rect 37188 2790 37240 2796
rect 14660 2746 14780 2774
rect 1768 2440 1820 2446
rect 1768 2382 1820 2388
rect 2228 2440 2280 2446
rect 2228 2382 2280 2388
rect 5448 2440 5500 2446
rect 5448 2382 5500 2388
rect 8392 2440 8444 2446
rect 8392 2382 8444 2388
rect 8484 2440 8536 2446
rect 8484 2382 8536 2388
rect 12992 2440 13044 2446
rect 12992 2382 13044 2388
rect 20 2372 72 2378
rect 20 2314 72 2320
rect 2044 2372 2096 2378
rect 2044 2314 2096 2320
rect 3976 2372 4028 2378
rect 3976 2314 4028 2320
rect 6552 2372 6604 2378
rect 6552 2314 6604 2320
rect 32 800 60 2314
rect 2056 1170 2084 2314
rect 3988 1170 4016 2314
rect 4874 2204 5182 2213
rect 4874 2202 4880 2204
rect 4936 2202 4960 2204
rect 5016 2202 5040 2204
rect 5096 2202 5120 2204
rect 5176 2202 5182 2204
rect 4936 2150 4938 2202
rect 5118 2150 5120 2202
rect 4874 2148 4880 2150
rect 4936 2148 4960 2150
rect 5016 2148 5040 2150
rect 5096 2148 5120 2150
rect 5176 2148 5182 2150
rect 4874 2139 5182 2148
rect 6564 1170 6592 2314
rect 8496 1306 8524 2382
rect 14660 2378 14688 2746
rect 14936 2446 14964 2790
rect 17420 2446 17448 2790
rect 19812 2446 19840 2790
rect 34934 2748 35242 2757
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2683 35242 2692
rect 14924 2440 14976 2446
rect 14924 2382 14976 2388
rect 17408 2440 17460 2446
rect 17408 2382 17460 2388
rect 19800 2440 19852 2446
rect 19800 2382 19852 2388
rect 10968 2372 11020 2378
rect 10968 2314 11020 2320
rect 14648 2372 14700 2378
rect 14648 2314 14700 2320
rect 19432 2372 19484 2378
rect 19432 2314 19484 2320
rect 1964 1142 2084 1170
rect 3896 1142 4016 1170
rect 6472 1142 6592 1170
rect 8404 1278 8524 1306
rect 1964 800 1992 1142
rect 3896 800 3924 1142
rect 6472 800 6500 1142
rect 8404 800 8432 1278
rect 10980 800 11008 2314
rect 12900 2304 12952 2310
rect 12900 2246 12952 2252
rect 15016 2304 15068 2310
rect 15016 2246 15068 2252
rect 17408 2304 17460 2310
rect 17408 2246 17460 2252
rect 12912 800 12940 2246
rect 15028 1170 15056 2246
rect 14844 1142 15056 1170
rect 14844 800 14872 1142
rect 17420 800 17448 2246
rect 19444 1170 19472 2314
rect 26424 2304 26476 2310
rect 26424 2246 26476 2252
rect 19352 1142 19472 1170
rect 19352 800 19380 1142
rect 26436 800 26464 2246
rect 35594 2204 35902 2213
rect 35594 2202 35600 2204
rect 35656 2202 35680 2204
rect 35736 2202 35760 2204
rect 35816 2202 35840 2204
rect 35896 2202 35902 2204
rect 35656 2150 35658 2202
rect 35838 2150 35840 2202
rect 35594 2148 35600 2150
rect 35656 2148 35680 2150
rect 35736 2148 35760 2150
rect 35816 2148 35840 2150
rect 35896 2148 35902 2150
rect 35594 2139 35902 2148
rect 37200 1465 37228 2790
rect 37464 2440 37516 2446
rect 37464 2382 37516 2388
rect 37186 1456 37242 1465
rect 37186 1391 37242 1400
rect 37476 1306 37504 2382
rect 37384 1278 37504 1306
rect 37384 800 37412 1278
rect 18 0 74 800
rect 1950 0 2006 800
rect 3882 0 3938 800
rect 6458 0 6514 800
rect 8390 0 8446 800
rect 10966 0 11022 800
rect 12898 0 12954 800
rect 14830 0 14886 800
rect 17406 0 17462 800
rect 19338 0 19394 800
rect 21914 0 21970 800
rect 23846 0 23902 800
rect 26422 0 26478 800
rect 28354 0 28410 800
rect 30286 0 30342 800
rect 32862 0 32918 800
rect 34794 0 34850 800
rect 37370 0 37426 800
rect 39302 0 39358 800
<< via2 >>
rect 4880 39194 4936 39196
rect 4960 39194 5016 39196
rect 5040 39194 5096 39196
rect 5120 39194 5176 39196
rect 4880 39142 4926 39194
rect 4926 39142 4936 39194
rect 4960 39142 4990 39194
rect 4990 39142 5002 39194
rect 5002 39142 5016 39194
rect 5040 39142 5054 39194
rect 5054 39142 5066 39194
rect 5066 39142 5096 39194
rect 5120 39142 5130 39194
rect 5130 39142 5176 39194
rect 4880 39140 4936 39142
rect 4960 39140 5016 39142
rect 5040 39140 5096 39142
rect 5120 39140 5176 39142
rect 938 36760 994 36816
rect 4220 38650 4276 38652
rect 4300 38650 4356 38652
rect 4380 38650 4436 38652
rect 4460 38650 4516 38652
rect 4220 38598 4266 38650
rect 4266 38598 4276 38650
rect 4300 38598 4330 38650
rect 4330 38598 4342 38650
rect 4342 38598 4356 38650
rect 4380 38598 4394 38650
rect 4394 38598 4406 38650
rect 4406 38598 4436 38650
rect 4460 38598 4470 38650
rect 4470 38598 4516 38650
rect 4220 38596 4276 38598
rect 4300 38596 4356 38598
rect 4380 38596 4436 38598
rect 4460 38596 4516 38598
rect 5170 38392 5226 38448
rect 4880 38106 4936 38108
rect 4960 38106 5016 38108
rect 5040 38106 5096 38108
rect 5120 38106 5176 38108
rect 4880 38054 4926 38106
rect 4926 38054 4936 38106
rect 4960 38054 4990 38106
rect 4990 38054 5002 38106
rect 5002 38054 5016 38106
rect 5040 38054 5054 38106
rect 5054 38054 5066 38106
rect 5066 38054 5096 38106
rect 5120 38054 5130 38106
rect 5130 38054 5176 38106
rect 4880 38052 4936 38054
rect 4960 38052 5016 38054
rect 5040 38052 5096 38054
rect 5120 38052 5176 38054
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 4880 37018 4936 37020
rect 4960 37018 5016 37020
rect 5040 37018 5096 37020
rect 5120 37018 5176 37020
rect 4880 36966 4926 37018
rect 4926 36966 4936 37018
rect 4960 36966 4990 37018
rect 4990 36966 5002 37018
rect 5002 36966 5016 37018
rect 5040 36966 5054 37018
rect 5054 36966 5066 37018
rect 5066 36966 5096 37018
rect 5120 36966 5130 37018
rect 5130 36966 5176 37018
rect 4880 36964 4936 36966
rect 4960 36964 5016 36966
rect 5040 36964 5096 36966
rect 5120 36964 5176 36966
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 938 25200 994 25256
rect 1490 20576 1546 20632
rect 938 18400 994 18456
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4880 35930 4936 35932
rect 4960 35930 5016 35932
rect 5040 35930 5096 35932
rect 5120 35930 5176 35932
rect 4880 35878 4926 35930
rect 4926 35878 4936 35930
rect 4960 35878 4990 35930
rect 4990 35878 5002 35930
rect 5002 35878 5016 35930
rect 5040 35878 5054 35930
rect 5054 35878 5066 35930
rect 5066 35878 5096 35930
rect 5120 35878 5130 35930
rect 5130 35878 5176 35930
rect 4880 35876 4936 35878
rect 4960 35876 5016 35878
rect 5040 35876 5096 35878
rect 5120 35876 5176 35878
rect 4880 34842 4936 34844
rect 4960 34842 5016 34844
rect 5040 34842 5096 34844
rect 5120 34842 5176 34844
rect 4880 34790 4926 34842
rect 4926 34790 4936 34842
rect 4960 34790 4990 34842
rect 4990 34790 5002 34842
rect 5002 34790 5016 34842
rect 5040 34790 5054 34842
rect 5054 34790 5066 34842
rect 5066 34790 5096 34842
rect 5120 34790 5130 34842
rect 5130 34790 5176 34842
rect 4880 34788 4936 34790
rect 4960 34788 5016 34790
rect 5040 34788 5096 34790
rect 5120 34788 5176 34790
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4880 33754 4936 33756
rect 4960 33754 5016 33756
rect 5040 33754 5096 33756
rect 5120 33754 5176 33756
rect 4880 33702 4926 33754
rect 4926 33702 4936 33754
rect 4960 33702 4990 33754
rect 4990 33702 5002 33754
rect 5002 33702 5016 33754
rect 5040 33702 5054 33754
rect 5054 33702 5066 33754
rect 5066 33702 5096 33754
rect 5120 33702 5130 33754
rect 5130 33702 5176 33754
rect 4880 33700 4936 33702
rect 4960 33700 5016 33702
rect 5040 33700 5096 33702
rect 5120 33700 5176 33702
rect 4880 32666 4936 32668
rect 4960 32666 5016 32668
rect 5040 32666 5096 32668
rect 5120 32666 5176 32668
rect 4880 32614 4926 32666
rect 4926 32614 4936 32666
rect 4960 32614 4990 32666
rect 4990 32614 5002 32666
rect 5002 32614 5016 32666
rect 5040 32614 5054 32666
rect 5054 32614 5066 32666
rect 5066 32614 5096 32666
rect 5120 32614 5130 32666
rect 5130 32614 5176 32666
rect 4880 32612 4936 32614
rect 4960 32612 5016 32614
rect 5040 32612 5096 32614
rect 5120 32612 5176 32614
rect 4880 31578 4936 31580
rect 4960 31578 5016 31580
rect 5040 31578 5096 31580
rect 5120 31578 5176 31580
rect 4880 31526 4926 31578
rect 4926 31526 4936 31578
rect 4960 31526 4990 31578
rect 4990 31526 5002 31578
rect 5002 31526 5016 31578
rect 5040 31526 5054 31578
rect 5054 31526 5066 31578
rect 5066 31526 5096 31578
rect 5120 31526 5130 31578
rect 5130 31526 5176 31578
rect 4880 31524 4936 31526
rect 4960 31524 5016 31526
rect 5040 31524 5096 31526
rect 5120 31524 5176 31526
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4880 30490 4936 30492
rect 4960 30490 5016 30492
rect 5040 30490 5096 30492
rect 5120 30490 5176 30492
rect 4880 30438 4926 30490
rect 4926 30438 4936 30490
rect 4960 30438 4990 30490
rect 4990 30438 5002 30490
rect 5002 30438 5016 30490
rect 5040 30438 5054 30490
rect 5054 30438 5066 30490
rect 5066 30438 5096 30490
rect 5120 30438 5130 30490
rect 5130 30438 5176 30490
rect 4880 30436 4936 30438
rect 4960 30436 5016 30438
rect 5040 30436 5096 30438
rect 5120 30436 5176 30438
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4066 27240 4122 27296
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4880 29402 4936 29404
rect 4960 29402 5016 29404
rect 5040 29402 5096 29404
rect 5120 29402 5176 29404
rect 4880 29350 4926 29402
rect 4926 29350 4936 29402
rect 4960 29350 4990 29402
rect 4990 29350 5002 29402
rect 5002 29350 5016 29402
rect 5040 29350 5054 29402
rect 5054 29350 5066 29402
rect 5066 29350 5096 29402
rect 5120 29350 5130 29402
rect 5130 29350 5176 29402
rect 4880 29348 4936 29350
rect 4960 29348 5016 29350
rect 5040 29348 5096 29350
rect 5120 29348 5176 29350
rect 4880 28314 4936 28316
rect 4960 28314 5016 28316
rect 5040 28314 5096 28316
rect 5120 28314 5176 28316
rect 4880 28262 4926 28314
rect 4926 28262 4936 28314
rect 4960 28262 4990 28314
rect 4990 28262 5002 28314
rect 5002 28262 5016 28314
rect 5040 28262 5054 28314
rect 5054 28262 5066 28314
rect 5066 28262 5096 28314
rect 5120 28262 5130 28314
rect 5130 28262 5176 28314
rect 4880 28260 4936 28262
rect 4960 28260 5016 28262
rect 5040 28260 5096 28262
rect 5120 28260 5176 28262
rect 5630 29008 5686 29064
rect 4880 27226 4936 27228
rect 4960 27226 5016 27228
rect 5040 27226 5096 27228
rect 5120 27226 5176 27228
rect 4880 27174 4926 27226
rect 4926 27174 4936 27226
rect 4960 27174 4990 27226
rect 4990 27174 5002 27226
rect 5002 27174 5016 27226
rect 5040 27174 5054 27226
rect 5054 27174 5066 27226
rect 5066 27174 5096 27226
rect 5120 27174 5130 27226
rect 5130 27174 5176 27226
rect 4880 27172 4936 27174
rect 4960 27172 5016 27174
rect 5040 27172 5096 27174
rect 5120 27172 5176 27174
rect 4880 26138 4936 26140
rect 4960 26138 5016 26140
rect 5040 26138 5096 26140
rect 5120 26138 5176 26140
rect 4880 26086 4926 26138
rect 4926 26086 4936 26138
rect 4960 26086 4990 26138
rect 4990 26086 5002 26138
rect 5002 26086 5016 26138
rect 5040 26086 5054 26138
rect 5054 26086 5066 26138
rect 5066 26086 5096 26138
rect 5120 26086 5130 26138
rect 5130 26086 5176 26138
rect 4880 26084 4936 26086
rect 4960 26084 5016 26086
rect 5040 26084 5096 26086
rect 5120 26084 5176 26086
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4880 25050 4936 25052
rect 4960 25050 5016 25052
rect 5040 25050 5096 25052
rect 5120 25050 5176 25052
rect 4880 24998 4926 25050
rect 4926 24998 4936 25050
rect 4960 24998 4990 25050
rect 4990 24998 5002 25050
rect 5002 24998 5016 25050
rect 5040 24998 5054 25050
rect 5054 24998 5066 25050
rect 5066 24998 5096 25050
rect 5120 24998 5130 25050
rect 5130 24998 5176 25050
rect 4880 24996 4936 24998
rect 4960 24996 5016 24998
rect 5040 24996 5096 24998
rect 5120 24996 5176 24998
rect 2962 22636 3018 22672
rect 2962 22616 2964 22636
rect 2964 22616 3016 22636
rect 3016 22616 3018 22636
rect 938 15700 994 15736
rect 938 15680 940 15700
rect 940 15680 992 15700
rect 992 15680 994 15700
rect 1490 13640 1546 13696
rect 938 11600 994 11656
rect 938 8900 994 8936
rect 938 8880 940 8900
rect 940 8880 992 8900
rect 992 8880 994 8900
rect 1490 6840 1546 6896
rect 938 4120 994 4176
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 4880 23962 4936 23964
rect 4960 23962 5016 23964
rect 5040 23962 5096 23964
rect 5120 23962 5176 23964
rect 4880 23910 4926 23962
rect 4926 23910 4936 23962
rect 4960 23910 4990 23962
rect 4990 23910 5002 23962
rect 5002 23910 5016 23962
rect 5040 23910 5054 23962
rect 5054 23910 5066 23962
rect 5066 23910 5096 23962
rect 5120 23910 5130 23962
rect 5130 23910 5176 23962
rect 4880 23908 4936 23910
rect 4960 23908 5016 23910
rect 5040 23908 5096 23910
rect 5120 23908 5176 23910
rect 4894 23060 4896 23080
rect 4896 23060 4948 23080
rect 4948 23060 4950 23080
rect 4894 23024 4950 23060
rect 4880 22874 4936 22876
rect 4960 22874 5016 22876
rect 5040 22874 5096 22876
rect 5120 22874 5176 22876
rect 4880 22822 4926 22874
rect 4926 22822 4936 22874
rect 4960 22822 4990 22874
rect 4990 22822 5002 22874
rect 5002 22822 5016 22874
rect 5040 22822 5054 22874
rect 5054 22822 5066 22874
rect 5066 22822 5096 22874
rect 5120 22822 5130 22874
rect 5130 22822 5176 22874
rect 4880 22820 4936 22822
rect 4960 22820 5016 22822
rect 5040 22820 5096 22822
rect 5120 22820 5176 22822
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4880 21786 4936 21788
rect 4960 21786 5016 21788
rect 5040 21786 5096 21788
rect 5120 21786 5176 21788
rect 4880 21734 4926 21786
rect 4926 21734 4936 21786
rect 4960 21734 4990 21786
rect 4990 21734 5002 21786
rect 5002 21734 5016 21786
rect 5040 21734 5054 21786
rect 5054 21734 5066 21786
rect 5066 21734 5096 21786
rect 5120 21734 5130 21786
rect 5130 21734 5176 21786
rect 4880 21732 4936 21734
rect 4960 21732 5016 21734
rect 5040 21732 5096 21734
rect 5120 21732 5176 21734
rect 4880 20698 4936 20700
rect 4960 20698 5016 20700
rect 5040 20698 5096 20700
rect 5120 20698 5176 20700
rect 4880 20646 4926 20698
rect 4926 20646 4936 20698
rect 4960 20646 4990 20698
rect 4990 20646 5002 20698
rect 5002 20646 5016 20698
rect 5040 20646 5054 20698
rect 5054 20646 5066 20698
rect 5066 20646 5096 20698
rect 5120 20646 5130 20698
rect 5130 20646 5176 20698
rect 4880 20644 4936 20646
rect 4960 20644 5016 20646
rect 5040 20644 5096 20646
rect 5120 20644 5176 20646
rect 4986 19760 5042 19816
rect 5354 19760 5410 19816
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 3238 9580 3294 9616
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4434 16652 4490 16688
rect 4434 16632 4436 16652
rect 4436 16632 4488 16652
rect 4488 16632 4490 16652
rect 4880 19610 4936 19612
rect 4960 19610 5016 19612
rect 5040 19610 5096 19612
rect 5120 19610 5176 19612
rect 4880 19558 4926 19610
rect 4926 19558 4936 19610
rect 4960 19558 4990 19610
rect 4990 19558 5002 19610
rect 5002 19558 5016 19610
rect 5040 19558 5054 19610
rect 5054 19558 5066 19610
rect 5066 19558 5096 19610
rect 5120 19558 5130 19610
rect 5130 19558 5176 19610
rect 4880 19556 4936 19558
rect 4960 19556 5016 19558
rect 5040 19556 5096 19558
rect 5120 19556 5176 19558
rect 4880 18522 4936 18524
rect 4960 18522 5016 18524
rect 5040 18522 5096 18524
rect 5120 18522 5176 18524
rect 4880 18470 4926 18522
rect 4926 18470 4936 18522
rect 4960 18470 4990 18522
rect 4990 18470 5002 18522
rect 5002 18470 5016 18522
rect 5040 18470 5054 18522
rect 5054 18470 5066 18522
rect 5066 18470 5096 18522
rect 5120 18470 5130 18522
rect 5130 18470 5176 18522
rect 4880 18468 4936 18470
rect 4960 18468 5016 18470
rect 5040 18468 5096 18470
rect 5120 18468 5176 18470
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4880 17434 4936 17436
rect 4960 17434 5016 17436
rect 5040 17434 5096 17436
rect 5120 17434 5176 17436
rect 4880 17382 4926 17434
rect 4926 17382 4936 17434
rect 4960 17382 4990 17434
rect 4990 17382 5002 17434
rect 5002 17382 5016 17434
rect 5040 17382 5054 17434
rect 5054 17382 5066 17434
rect 5066 17382 5096 17434
rect 5120 17382 5130 17434
rect 5130 17382 5176 17434
rect 4880 17380 4936 17382
rect 4960 17380 5016 17382
rect 5040 17380 5096 17382
rect 5120 17380 5176 17382
rect 4880 16346 4936 16348
rect 4960 16346 5016 16348
rect 5040 16346 5096 16348
rect 5120 16346 5176 16348
rect 4880 16294 4926 16346
rect 4926 16294 4936 16346
rect 4960 16294 4990 16346
rect 4990 16294 5002 16346
rect 5002 16294 5016 16346
rect 5040 16294 5054 16346
rect 5054 16294 5066 16346
rect 5066 16294 5096 16346
rect 5120 16294 5130 16346
rect 5130 16294 5176 16346
rect 4880 16292 4936 16294
rect 4960 16292 5016 16294
rect 5040 16292 5096 16294
rect 5120 16292 5176 16294
rect 4880 15258 4936 15260
rect 4960 15258 5016 15260
rect 5040 15258 5096 15260
rect 5120 15258 5176 15260
rect 4880 15206 4926 15258
rect 4926 15206 4936 15258
rect 4960 15206 4990 15258
rect 4990 15206 5002 15258
rect 5002 15206 5016 15258
rect 5040 15206 5054 15258
rect 5054 15206 5066 15258
rect 5066 15206 5096 15258
rect 5120 15206 5130 15258
rect 5130 15206 5176 15258
rect 4880 15204 4936 15206
rect 4960 15204 5016 15206
rect 5040 15204 5096 15206
rect 5120 15204 5176 15206
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4880 14170 4936 14172
rect 4960 14170 5016 14172
rect 5040 14170 5096 14172
rect 5120 14170 5176 14172
rect 4880 14118 4926 14170
rect 4926 14118 4936 14170
rect 4960 14118 4990 14170
rect 4990 14118 5002 14170
rect 5002 14118 5016 14170
rect 5040 14118 5054 14170
rect 5054 14118 5066 14170
rect 5066 14118 5096 14170
rect 5120 14118 5130 14170
rect 5130 14118 5176 14170
rect 4880 14116 4936 14118
rect 4960 14116 5016 14118
rect 5040 14116 5096 14118
rect 5120 14116 5176 14118
rect 4880 13082 4936 13084
rect 4960 13082 5016 13084
rect 5040 13082 5096 13084
rect 5120 13082 5176 13084
rect 4880 13030 4926 13082
rect 4926 13030 4936 13082
rect 4960 13030 4990 13082
rect 4990 13030 5002 13082
rect 5002 13030 5016 13082
rect 5040 13030 5054 13082
rect 5054 13030 5066 13082
rect 5066 13030 5096 13082
rect 5120 13030 5130 13082
rect 5130 13030 5176 13082
rect 4880 13028 4936 13030
rect 4960 13028 5016 13030
rect 5040 13028 5096 13030
rect 5120 13028 5176 13030
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 5722 21120 5778 21176
rect 5630 20868 5686 20904
rect 5630 20848 5632 20868
rect 5632 20848 5684 20868
rect 5684 20848 5686 20868
rect 5998 18808 6054 18864
rect 4880 11994 4936 11996
rect 4960 11994 5016 11996
rect 5040 11994 5096 11996
rect 5120 11994 5176 11996
rect 4880 11942 4926 11994
rect 4926 11942 4936 11994
rect 4960 11942 4990 11994
rect 4990 11942 5002 11994
rect 5002 11942 5016 11994
rect 5040 11942 5054 11994
rect 5054 11942 5066 11994
rect 5066 11942 5096 11994
rect 5120 11942 5130 11994
rect 5130 11942 5176 11994
rect 4880 11940 4936 11942
rect 4960 11940 5016 11942
rect 5040 11940 5096 11942
rect 5120 11940 5176 11942
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4880 10906 4936 10908
rect 4960 10906 5016 10908
rect 5040 10906 5096 10908
rect 5120 10906 5176 10908
rect 4880 10854 4926 10906
rect 4926 10854 4936 10906
rect 4960 10854 4990 10906
rect 4990 10854 5002 10906
rect 5002 10854 5016 10906
rect 5040 10854 5054 10906
rect 5054 10854 5066 10906
rect 5066 10854 5096 10906
rect 5120 10854 5130 10906
rect 5130 10854 5176 10906
rect 4880 10852 4936 10854
rect 4960 10852 5016 10854
rect 5040 10852 5096 10854
rect 5120 10852 5176 10854
rect 3238 9560 3240 9580
rect 3240 9560 3292 9580
rect 3292 9560 3294 9580
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4880 9818 4936 9820
rect 4960 9818 5016 9820
rect 5040 9818 5096 9820
rect 5120 9818 5176 9820
rect 4880 9766 4926 9818
rect 4926 9766 4936 9818
rect 4960 9766 4990 9818
rect 4990 9766 5002 9818
rect 5002 9766 5016 9818
rect 5040 9766 5054 9818
rect 5054 9766 5066 9818
rect 5066 9766 5096 9818
rect 5120 9766 5130 9818
rect 5130 9766 5176 9818
rect 4880 9764 4936 9766
rect 4960 9764 5016 9766
rect 5040 9764 5096 9766
rect 5120 9764 5176 9766
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4158 9016 4214 9072
rect 4880 8730 4936 8732
rect 4960 8730 5016 8732
rect 5040 8730 5096 8732
rect 5120 8730 5176 8732
rect 4880 8678 4926 8730
rect 4926 8678 4936 8730
rect 4960 8678 4990 8730
rect 4990 8678 5002 8730
rect 5002 8678 5016 8730
rect 5040 8678 5054 8730
rect 5054 8678 5066 8730
rect 5066 8678 5096 8730
rect 5120 8678 5130 8730
rect 5130 8678 5176 8730
rect 4880 8676 4936 8678
rect 4960 8676 5016 8678
rect 5040 8676 5096 8678
rect 5120 8676 5176 8678
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4880 7642 4936 7644
rect 4960 7642 5016 7644
rect 5040 7642 5096 7644
rect 5120 7642 5176 7644
rect 4880 7590 4926 7642
rect 4926 7590 4936 7642
rect 4960 7590 4990 7642
rect 4990 7590 5002 7642
rect 5002 7590 5016 7642
rect 5040 7590 5054 7642
rect 5054 7590 5066 7642
rect 5066 7590 5096 7642
rect 5120 7590 5130 7642
rect 5130 7590 5176 7642
rect 4880 7588 4936 7590
rect 4960 7588 5016 7590
rect 5040 7588 5096 7590
rect 5120 7588 5176 7590
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4880 6554 4936 6556
rect 4960 6554 5016 6556
rect 5040 6554 5096 6556
rect 5120 6554 5176 6556
rect 4880 6502 4926 6554
rect 4926 6502 4936 6554
rect 4960 6502 4990 6554
rect 4990 6502 5002 6554
rect 5002 6502 5016 6554
rect 5040 6502 5054 6554
rect 5054 6502 5066 6554
rect 5066 6502 5096 6554
rect 5120 6502 5130 6554
rect 5130 6502 5176 6554
rect 4880 6500 4936 6502
rect 4960 6500 5016 6502
rect 5040 6500 5096 6502
rect 5120 6500 5176 6502
rect 4880 5466 4936 5468
rect 4960 5466 5016 5468
rect 5040 5466 5096 5468
rect 5120 5466 5176 5468
rect 4880 5414 4926 5466
rect 4926 5414 4936 5466
rect 4960 5414 4990 5466
rect 4990 5414 5002 5466
rect 5002 5414 5016 5466
rect 5040 5414 5054 5466
rect 5054 5414 5066 5466
rect 5066 5414 5096 5466
rect 5120 5414 5130 5466
rect 5130 5414 5176 5466
rect 4880 5412 4936 5414
rect 4960 5412 5016 5414
rect 5040 5412 5096 5414
rect 5120 5412 5176 5414
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4880 4378 4936 4380
rect 4960 4378 5016 4380
rect 5040 4378 5096 4380
rect 5120 4378 5176 4380
rect 4880 4326 4926 4378
rect 4926 4326 4936 4378
rect 4960 4326 4990 4378
rect 4990 4326 5002 4378
rect 5002 4326 5016 4378
rect 5040 4326 5054 4378
rect 5054 4326 5066 4378
rect 5066 4326 5096 4378
rect 5120 4326 5130 4378
rect 5130 4326 5176 4378
rect 4880 4324 4936 4326
rect 4960 4324 5016 4326
rect 5040 4324 5096 4326
rect 5120 4324 5176 4326
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4880 3290 4936 3292
rect 4960 3290 5016 3292
rect 5040 3290 5096 3292
rect 5120 3290 5176 3292
rect 4880 3238 4926 3290
rect 4926 3238 4936 3290
rect 4960 3238 4990 3290
rect 4990 3238 5002 3290
rect 5002 3238 5016 3290
rect 5040 3238 5054 3290
rect 5054 3238 5066 3290
rect 5066 3238 5096 3290
rect 5120 3238 5130 3290
rect 5130 3238 5176 3290
rect 4880 3236 4936 3238
rect 4960 3236 5016 3238
rect 5040 3236 5096 3238
rect 5120 3236 5176 3238
rect 35600 39194 35656 39196
rect 35680 39194 35736 39196
rect 35760 39194 35816 39196
rect 35840 39194 35896 39196
rect 35600 39142 35646 39194
rect 35646 39142 35656 39194
rect 35680 39142 35710 39194
rect 35710 39142 35722 39194
rect 35722 39142 35736 39194
rect 35760 39142 35774 39194
rect 35774 39142 35786 39194
rect 35786 39142 35816 39194
rect 35840 39142 35850 39194
rect 35850 39142 35896 39194
rect 35600 39140 35656 39142
rect 35680 39140 35736 39142
rect 35760 39140 35816 39142
rect 35840 39140 35896 39142
rect 8390 29280 8446 29336
rect 6550 19796 6552 19816
rect 6552 19796 6604 19816
rect 6604 19796 6606 19816
rect 6550 19760 6606 19796
rect 7930 23024 7986 23080
rect 7930 19760 7986 19816
rect 7930 16632 7986 16688
rect 8206 22500 8262 22536
rect 8206 22480 8208 22500
rect 8208 22480 8260 22500
rect 8260 22480 8262 22500
rect 11518 36116 11520 36136
rect 11520 36116 11572 36136
rect 11572 36116 11574 36136
rect 11518 36080 11574 36116
rect 8390 19660 8392 19680
rect 8392 19660 8444 19680
rect 8444 19660 8446 19680
rect 8390 19624 8446 19660
rect 6642 9424 6698 9480
rect 9586 29008 9642 29064
rect 9862 24248 9918 24304
rect 11242 28092 11244 28112
rect 11244 28092 11296 28112
rect 11296 28092 11298 28112
rect 11242 28056 11298 28092
rect 9678 21548 9734 21584
rect 9678 21528 9680 21548
rect 9680 21528 9732 21548
rect 9732 21528 9734 21548
rect 9126 20032 9182 20088
rect 9034 19372 9090 19408
rect 9034 19352 9036 19372
rect 9036 19352 9088 19372
rect 9088 19352 9090 19372
rect 8942 17856 8998 17912
rect 9586 20712 9642 20768
rect 9770 20576 9826 20632
rect 9494 19896 9550 19952
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 10046 21256 10102 21312
rect 10322 21548 10378 21584
rect 10322 21528 10324 21548
rect 10324 21528 10376 21548
rect 10376 21528 10378 21548
rect 10138 20304 10194 20360
rect 9586 14340 9642 14376
rect 9586 14320 9588 14340
rect 9588 14320 9640 14340
rect 9640 14320 9642 14340
rect 9586 13640 9642 13696
rect 9310 9424 9366 9480
rect 12162 32816 12218 32872
rect 10506 18400 10562 18456
rect 10874 17992 10930 18048
rect 10874 17720 10930 17776
rect 10230 12960 10286 13016
rect 9954 9152 10010 9208
rect 11150 18944 11206 19000
rect 12346 25064 12402 25120
rect 13174 37868 13230 37904
rect 13174 37848 13176 37868
rect 13176 37848 13228 37868
rect 13228 37848 13230 37868
rect 12622 32136 12678 32192
rect 13082 31864 13138 31920
rect 12898 29028 12954 29064
rect 12898 29008 12900 29028
rect 12900 29008 12952 29028
rect 12952 29008 12954 29028
rect 12990 24656 13046 24712
rect 12622 23432 12678 23488
rect 11886 21548 11942 21584
rect 11886 21528 11888 21548
rect 11888 21528 11940 21548
rect 11940 21528 11942 21548
rect 12438 20576 12494 20632
rect 11702 17856 11758 17912
rect 11702 17604 11758 17640
rect 11702 17584 11704 17604
rect 11704 17584 11756 17604
rect 11756 17584 11758 17604
rect 11886 17856 11942 17912
rect 12530 19488 12586 19544
rect 12162 18536 12218 18592
rect 11426 15444 11428 15464
rect 11428 15444 11480 15464
rect 11480 15444 11482 15464
rect 11426 15408 11482 15444
rect 12254 17740 12310 17776
rect 12254 17720 12256 17740
rect 12256 17720 12308 17740
rect 12308 17720 12310 17740
rect 12530 17584 12586 17640
rect 12714 18400 12770 18456
rect 12346 16108 12402 16144
rect 12346 16088 12348 16108
rect 12348 16088 12400 16108
rect 12400 16088 12402 16108
rect 12254 15952 12310 16008
rect 12530 15816 12586 15872
rect 12898 19488 12954 19544
rect 13542 26560 13598 26616
rect 13910 25880 13966 25936
rect 13726 23568 13782 23624
rect 13542 21392 13598 21448
rect 13634 20168 13690 20224
rect 13358 17876 13414 17912
rect 13358 17856 13360 17876
rect 13360 17856 13412 17876
rect 13412 17856 13414 17876
rect 13542 19488 13598 19544
rect 13910 23432 13966 23488
rect 15566 38664 15622 38720
rect 22374 38664 22430 38720
rect 27066 38664 27122 38720
rect 15014 33632 15070 33688
rect 15198 33496 15254 33552
rect 14738 26868 14740 26888
rect 14740 26868 14792 26888
rect 14792 26868 14794 26888
rect 14738 26832 14794 26868
rect 15566 36080 15622 36136
rect 15658 33904 15714 33960
rect 15566 33768 15622 33824
rect 15198 29688 15254 29744
rect 15658 30096 15714 30152
rect 15842 29588 15844 29608
rect 15844 29588 15896 29608
rect 15896 29588 15898 29608
rect 15842 29552 15898 29588
rect 14462 24928 14518 24984
rect 14278 23740 14280 23760
rect 14280 23740 14332 23760
rect 14332 23740 14334 23760
rect 14278 23704 14334 23740
rect 13910 21664 13966 21720
rect 14278 20984 14334 21040
rect 14554 19488 14610 19544
rect 14830 20440 14886 20496
rect 14370 16632 14426 16688
rect 13818 9172 13874 9208
rect 13818 9152 13820 9172
rect 13820 9152 13872 9172
rect 13872 9152 13874 9172
rect 16302 31456 16358 31512
rect 17130 32292 17186 32328
rect 17130 32272 17132 32292
rect 17132 32272 17184 32292
rect 17184 32272 17186 32292
rect 17406 35980 17408 36000
rect 17408 35980 17460 36000
rect 17460 35980 17462 36000
rect 17406 35944 17462 35980
rect 16670 30232 16726 30288
rect 17498 33496 17554 33552
rect 17314 31592 17370 31648
rect 17866 33088 17922 33144
rect 18142 30252 18198 30288
rect 18142 30232 18144 30252
rect 18144 30232 18196 30252
rect 18196 30232 18198 30252
rect 18418 32000 18474 32056
rect 18326 30368 18382 30424
rect 18878 31864 18934 31920
rect 19706 34040 19762 34096
rect 19338 33652 19394 33688
rect 19338 33632 19340 33652
rect 19340 33632 19392 33652
rect 19392 33632 19394 33652
rect 19062 33224 19118 33280
rect 19062 32292 19118 32328
rect 19062 32272 19064 32292
rect 19064 32272 19116 32292
rect 19116 32272 19118 32292
rect 19062 30660 19118 30696
rect 19062 30640 19064 30660
rect 19064 30640 19116 30660
rect 19116 30640 19118 30660
rect 19338 31184 19394 31240
rect 19430 30912 19486 30968
rect 18418 30096 18474 30152
rect 17406 28092 17408 28112
rect 17408 28092 17460 28112
rect 17460 28092 17462 28112
rect 17406 28056 17462 28092
rect 15566 21528 15622 21584
rect 15290 20576 15346 20632
rect 15106 18400 15162 18456
rect 15566 20576 15622 20632
rect 16026 21936 16082 21992
rect 16670 24148 16672 24168
rect 16672 24148 16724 24168
rect 16724 24148 16726 24168
rect 16670 24112 16726 24148
rect 16026 19488 16082 19544
rect 16762 21972 16764 21992
rect 16764 21972 16816 21992
rect 16816 21972 16818 21992
rect 16762 21936 16818 21972
rect 16578 20576 16634 20632
rect 16210 17448 16266 17504
rect 17130 26696 17186 26752
rect 17774 26560 17830 26616
rect 18418 29452 18420 29472
rect 18420 29452 18472 29472
rect 18472 29452 18474 29472
rect 18418 29416 18474 29452
rect 18234 29144 18290 29200
rect 17590 26016 17646 26072
rect 16578 16632 16634 16688
rect 17038 20576 17094 20632
rect 17130 18400 17186 18456
rect 16946 17448 17002 17504
rect 12530 3984 12586 4040
rect 13174 3984 13230 4040
rect 15382 9424 15438 9480
rect 18878 29588 18880 29608
rect 18880 29588 18932 29608
rect 18932 29588 18934 29608
rect 18878 29552 18934 29588
rect 18878 29008 18934 29064
rect 18786 26288 18842 26344
rect 17866 24112 17922 24168
rect 18050 23468 18052 23488
rect 18052 23468 18104 23488
rect 18104 23468 18106 23488
rect 18050 23432 18106 23468
rect 18050 20440 18106 20496
rect 18970 26868 18972 26888
rect 18972 26868 19024 26888
rect 19024 26868 19026 26888
rect 18970 26832 19026 26868
rect 19338 29280 19394 29336
rect 19246 27920 19302 27976
rect 19154 26560 19210 26616
rect 20166 35944 20222 36000
rect 19982 33088 20038 33144
rect 19982 31048 20038 31104
rect 20258 33940 20260 33960
rect 20260 33940 20312 33960
rect 20312 33940 20314 33960
rect 20258 33904 20314 33940
rect 20166 33496 20222 33552
rect 25778 38392 25834 38448
rect 25318 37868 25374 37904
rect 25318 37848 25320 37868
rect 25320 37848 25372 37868
rect 25372 37848 25374 37868
rect 20902 33940 20904 33960
rect 20904 33940 20956 33960
rect 20956 33940 20958 33960
rect 20902 33904 20958 33940
rect 19982 29960 20038 30016
rect 19614 28484 19670 28520
rect 19614 28464 19616 28484
rect 19616 28464 19668 28484
rect 19668 28464 19670 28484
rect 19430 28192 19486 28248
rect 19614 28076 19670 28112
rect 19614 28056 19616 28076
rect 19616 28056 19668 28076
rect 19668 28056 19670 28076
rect 19798 28192 19854 28248
rect 20442 32816 20498 32872
rect 20350 31592 20406 31648
rect 20718 31184 20774 31240
rect 20626 30912 20682 30968
rect 20258 28600 20314 28656
rect 19154 26016 19210 26072
rect 19338 25764 19394 25800
rect 19338 25744 19340 25764
rect 19340 25744 19392 25764
rect 19392 25744 19394 25764
rect 19338 24928 19394 24984
rect 18234 20984 18290 21040
rect 18326 20576 18382 20632
rect 18510 18944 18566 19000
rect 18234 17856 18290 17912
rect 17958 16632 18014 16688
rect 17038 9152 17094 9208
rect 18970 18708 18972 18728
rect 18972 18708 19024 18728
rect 19024 18708 19026 18728
rect 18970 18672 19026 18708
rect 18602 17856 18658 17912
rect 18878 18128 18934 18184
rect 20442 27956 20444 27976
rect 20444 27956 20496 27976
rect 20496 27956 20498 27976
rect 20074 25780 20076 25800
rect 20076 25780 20128 25800
rect 20128 25780 20130 25800
rect 20074 25744 20130 25780
rect 20442 27920 20498 27956
rect 20350 26444 20406 26480
rect 20350 26424 20352 26444
rect 20352 26424 20404 26444
rect 20404 26424 20406 26444
rect 19430 23724 19486 23760
rect 19430 23704 19432 23724
rect 19432 23704 19484 23724
rect 19484 23704 19486 23724
rect 19246 22072 19302 22128
rect 19798 21392 19854 21448
rect 19798 18672 19854 18728
rect 18878 15852 18880 15872
rect 18880 15852 18932 15872
rect 18932 15852 18934 15872
rect 18878 15816 18934 15852
rect 17498 10532 17554 10568
rect 17498 10512 17500 10532
rect 17500 10512 17552 10532
rect 17552 10512 17554 10532
rect 18234 10920 18290 10976
rect 18694 12960 18750 13016
rect 18694 11620 18750 11656
rect 18694 11600 18696 11620
rect 18696 11600 18748 11620
rect 18748 11600 18750 11620
rect 20166 21256 20222 21312
rect 20166 18420 20222 18456
rect 20166 18400 20168 18420
rect 20168 18400 20220 18420
rect 20220 18400 20222 18420
rect 20074 18128 20130 18184
rect 21086 31728 21142 31784
rect 21454 33632 21510 33688
rect 21638 32444 21640 32464
rect 21640 32444 21692 32464
rect 21692 32444 21694 32464
rect 21638 32408 21694 32444
rect 21730 32000 21786 32056
rect 22282 34312 22338 34368
rect 21638 31592 21694 31648
rect 21546 31456 21602 31512
rect 21730 31320 21786 31376
rect 20810 29280 20866 29336
rect 20902 29164 20958 29200
rect 20902 29144 20904 29164
rect 20904 29144 20956 29164
rect 20956 29144 20958 29164
rect 21086 29008 21142 29064
rect 20626 26152 20682 26208
rect 21086 27920 21142 27976
rect 20534 25064 20590 25120
rect 22926 37324 22982 37360
rect 22926 37304 22928 37324
rect 22928 37304 22980 37324
rect 22980 37304 22982 37324
rect 22282 31048 22338 31104
rect 22282 29688 22338 29744
rect 22926 34040 22982 34096
rect 22834 33496 22890 33552
rect 23202 33768 23258 33824
rect 22466 29416 22522 29472
rect 21914 27648 21970 27704
rect 21454 25744 21510 25800
rect 21454 24948 21510 24984
rect 21454 24928 21456 24948
rect 21456 24928 21508 24948
rect 21508 24928 21510 24948
rect 21914 26696 21970 26752
rect 22374 27784 22430 27840
rect 23018 32272 23074 32328
rect 23202 32292 23258 32328
rect 23202 32272 23204 32292
rect 23204 32272 23256 32292
rect 23256 32272 23258 32292
rect 23478 34584 23534 34640
rect 23478 33632 23534 33688
rect 23386 33360 23442 33416
rect 23846 34312 23902 34368
rect 23938 33496 23994 33552
rect 22742 28600 22798 28656
rect 22006 20304 22062 20360
rect 22190 24248 22246 24304
rect 22742 26288 22798 26344
rect 23386 31320 23442 31376
rect 23386 30368 23442 30424
rect 23110 29416 23166 29472
rect 22926 27956 22928 27976
rect 22928 27956 22980 27976
rect 22980 27956 22982 27976
rect 22926 27920 22982 27956
rect 22834 26016 22890 26072
rect 23018 26560 23074 26616
rect 22834 23704 22890 23760
rect 22190 21428 22192 21448
rect 22192 21428 22244 21448
rect 22244 21428 22246 21448
rect 22190 21392 22246 21428
rect 18878 9460 18880 9480
rect 18880 9460 18932 9480
rect 18932 9460 18934 9480
rect 18878 9424 18934 9460
rect 18970 8492 19026 8528
rect 18970 8472 18972 8492
rect 18972 8472 19024 8492
rect 19024 8472 19026 8492
rect 18234 6840 18290 6896
rect 20810 10920 20866 10976
rect 20626 10004 20628 10024
rect 20628 10004 20680 10024
rect 20680 10004 20682 10024
rect 20626 9968 20682 10004
rect 22374 21936 22430 21992
rect 22374 20884 22376 20904
rect 22376 20884 22428 20904
rect 22428 20884 22430 20904
rect 22374 20848 22430 20884
rect 22466 19896 22522 19952
rect 22466 19488 22522 19544
rect 22374 19372 22430 19408
rect 22650 22072 22706 22128
rect 22834 21392 22890 21448
rect 22374 19352 22376 19372
rect 22376 19352 22428 19372
rect 22428 19352 22430 19372
rect 22374 19216 22430 19272
rect 22834 20052 22890 20088
rect 22834 20032 22836 20052
rect 22836 20032 22888 20052
rect 22888 20032 22890 20052
rect 22742 17856 22798 17912
rect 23294 29552 23350 29608
rect 24030 33260 24032 33280
rect 24032 33260 24084 33280
rect 24084 33260 24086 33280
rect 24030 33224 24086 33260
rect 23938 33088 23994 33144
rect 23754 31184 23810 31240
rect 23570 29008 23626 29064
rect 23110 25900 23166 25936
rect 23110 25880 23112 25900
rect 23112 25880 23164 25900
rect 23164 25880 23166 25900
rect 23110 20576 23166 20632
rect 23110 20032 23166 20088
rect 24030 30232 24086 30288
rect 24030 29280 24086 29336
rect 25226 37304 25282 37360
rect 24490 32272 24546 32328
rect 24950 35944 25006 36000
rect 25594 36116 25596 36136
rect 25596 36116 25648 36136
rect 25648 36116 25650 36136
rect 25594 36080 25650 36116
rect 25134 34856 25190 34912
rect 24582 29588 24584 29608
rect 24584 29588 24636 29608
rect 24636 29588 24638 29608
rect 24582 29552 24638 29588
rect 24858 29960 24914 30016
rect 24858 29028 24914 29064
rect 24858 29008 24860 29028
rect 24860 29008 24912 29028
rect 24912 29008 24914 29028
rect 24030 26016 24086 26072
rect 24858 28500 24860 28520
rect 24860 28500 24912 28520
rect 24912 28500 24914 28520
rect 24858 28464 24914 28500
rect 24306 25900 24362 25936
rect 24306 25880 24308 25900
rect 24308 25880 24360 25900
rect 24360 25880 24362 25900
rect 24582 26424 24638 26480
rect 24766 27784 24822 27840
rect 24858 26152 24914 26208
rect 24030 24656 24086 24712
rect 24306 23588 24362 23624
rect 24306 23568 24308 23588
rect 24308 23568 24360 23588
rect 24360 23568 24362 23588
rect 25042 26424 25098 26480
rect 25042 26016 25098 26072
rect 24950 25336 25006 25392
rect 24766 22480 24822 22536
rect 23478 20168 23534 20224
rect 23294 19916 23350 19952
rect 23294 19896 23296 19916
rect 23296 19896 23348 19916
rect 23348 19896 23350 19916
rect 23202 17584 23258 17640
rect 22098 10920 22154 10976
rect 22006 10684 22008 10704
rect 22008 10684 22060 10704
rect 22060 10684 22062 10704
rect 22006 10648 22062 10684
rect 21914 10004 21916 10024
rect 21916 10004 21968 10024
rect 21968 10004 21970 10024
rect 21914 9968 21970 10004
rect 22190 10376 22246 10432
rect 21822 8336 21878 8392
rect 24398 20168 24454 20224
rect 23570 18808 23626 18864
rect 23386 17856 23442 17912
rect 24858 21120 24914 21176
rect 25594 35708 25596 35728
rect 25596 35708 25648 35728
rect 25648 35708 25650 35728
rect 25594 35672 25650 35708
rect 25594 35572 25596 35592
rect 25596 35572 25648 35592
rect 25648 35572 25650 35592
rect 25594 35536 25650 35572
rect 25410 33260 25412 33280
rect 25412 33260 25464 33280
rect 25464 33260 25466 33280
rect 25410 33224 25466 33260
rect 25410 32000 25466 32056
rect 25318 26152 25374 26208
rect 25318 25744 25374 25800
rect 25134 21956 25190 21992
rect 25134 21936 25136 21956
rect 25136 21936 25188 21956
rect 25188 21936 25190 21956
rect 25594 29960 25650 30016
rect 25870 35128 25926 35184
rect 26882 35672 26938 35728
rect 26422 35536 26478 35592
rect 25870 30116 25926 30152
rect 25870 30096 25872 30116
rect 25872 30096 25924 30116
rect 25924 30096 25926 30116
rect 25778 29824 25834 29880
rect 25870 29008 25926 29064
rect 25318 22344 25374 22400
rect 22650 10920 22706 10976
rect 23018 10648 23074 10704
rect 22282 9560 22338 9616
rect 22742 9152 22798 9208
rect 22650 9016 22706 9072
rect 23754 15952 23810 16008
rect 23478 8336 23534 8392
rect 24950 20168 25006 20224
rect 24858 18536 24914 18592
rect 25226 20576 25282 20632
rect 25318 19780 25374 19816
rect 25318 19760 25320 19780
rect 25320 19760 25372 19780
rect 25372 19760 25374 19780
rect 24674 17448 24730 17504
rect 24490 16496 24546 16552
rect 24490 16088 24546 16144
rect 24398 13912 24454 13968
rect 24398 13368 24454 13424
rect 24122 12008 24178 12064
rect 25134 15408 25190 15464
rect 26698 31864 26754 31920
rect 26698 30368 26754 30424
rect 26606 29824 26662 29880
rect 26238 29008 26294 29064
rect 26882 29960 26938 30016
rect 27986 37304 28042 37360
rect 28446 35944 28502 36000
rect 28354 35164 28356 35184
rect 28356 35164 28408 35184
rect 28408 35164 28410 35184
rect 28354 35128 28410 35164
rect 28814 36116 28816 36136
rect 28816 36116 28868 36136
rect 28868 36116 28870 36136
rect 28814 36080 28870 36116
rect 26698 28056 26754 28112
rect 26238 26696 26294 26752
rect 26146 25880 26202 25936
rect 26054 25336 26110 25392
rect 26514 26968 26570 27024
rect 26698 26288 26754 26344
rect 25962 23044 26018 23080
rect 25962 23024 25964 23044
rect 25964 23024 26016 23044
rect 26016 23024 26018 23044
rect 25594 22616 25650 22672
rect 25778 21564 25780 21584
rect 25780 21564 25832 21584
rect 25832 21564 25834 21584
rect 25778 21528 25834 21564
rect 25778 19352 25834 19408
rect 27710 31084 27712 31104
rect 27712 31084 27764 31104
rect 27764 31084 27766 31104
rect 27710 31048 27766 31084
rect 28446 29572 28502 29608
rect 28446 29552 28448 29572
rect 28448 29552 28500 29572
rect 28500 29552 28502 29572
rect 27802 24656 27858 24712
rect 28262 26424 28318 26480
rect 27710 21548 27766 21584
rect 27710 21528 27712 21548
rect 27712 21528 27764 21548
rect 27764 21528 27766 21548
rect 26882 20032 26938 20088
rect 26054 19624 26110 19680
rect 25594 14900 25596 14920
rect 25596 14900 25648 14920
rect 25648 14900 25650 14920
rect 25594 14864 25650 14900
rect 26054 13932 26110 13968
rect 26054 13912 26056 13932
rect 26056 13912 26108 13932
rect 26108 13912 26110 13932
rect 25318 9036 25374 9072
rect 25318 9016 25320 9036
rect 25320 9016 25372 9036
rect 25372 9016 25374 9036
rect 25410 8336 25466 8392
rect 26238 13388 26294 13424
rect 26238 13368 26240 13388
rect 26240 13368 26292 13388
rect 26292 13368 26294 13388
rect 26146 12860 26148 12880
rect 26148 12860 26200 12880
rect 26200 12860 26202 12880
rect 26146 12824 26202 12860
rect 26422 13368 26478 13424
rect 27434 19488 27490 19544
rect 28262 19372 28318 19408
rect 28262 19352 28264 19372
rect 28264 19352 28316 19372
rect 28316 19352 28318 19372
rect 27710 17740 27766 17776
rect 27710 17720 27712 17740
rect 27712 17720 27764 17740
rect 27764 17720 27766 17740
rect 26606 12824 26662 12880
rect 26054 9016 26110 9072
rect 29550 33088 29606 33144
rect 29090 28600 29146 28656
rect 34940 38650 34996 38652
rect 35020 38650 35076 38652
rect 35100 38650 35156 38652
rect 35180 38650 35236 38652
rect 34940 38598 34986 38650
rect 34986 38598 34996 38650
rect 35020 38598 35050 38650
rect 35050 38598 35062 38650
rect 35062 38598 35076 38650
rect 35100 38598 35114 38650
rect 35114 38598 35126 38650
rect 35126 38598 35156 38650
rect 35180 38598 35190 38650
rect 35190 38598 35236 38650
rect 34940 38596 34996 38598
rect 35020 38596 35076 38598
rect 35100 38596 35156 38598
rect 35180 38596 35236 38598
rect 37646 38820 37702 38856
rect 37646 38800 37648 38820
rect 37648 38800 37700 38820
rect 37700 38800 37702 38820
rect 37922 38800 37978 38856
rect 30194 30640 30250 30696
rect 30378 30096 30434 30152
rect 29826 29588 29828 29608
rect 29828 29588 29880 29608
rect 29880 29588 29882 29608
rect 29826 29552 29882 29588
rect 29918 27920 29974 27976
rect 35600 38106 35656 38108
rect 35680 38106 35736 38108
rect 35760 38106 35816 38108
rect 35840 38106 35896 38108
rect 35600 38054 35646 38106
rect 35646 38054 35656 38106
rect 35680 38054 35710 38106
rect 35710 38054 35722 38106
rect 35722 38054 35736 38106
rect 35760 38054 35774 38106
rect 35774 38054 35786 38106
rect 35786 38054 35816 38106
rect 35840 38054 35850 38106
rect 35850 38054 35896 38106
rect 35600 38052 35656 38054
rect 35680 38052 35736 38054
rect 35760 38052 35816 38054
rect 35840 38052 35896 38054
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 35600 37018 35656 37020
rect 35680 37018 35736 37020
rect 35760 37018 35816 37020
rect 35840 37018 35896 37020
rect 35600 36966 35646 37018
rect 35646 36966 35656 37018
rect 35680 36966 35710 37018
rect 35710 36966 35722 37018
rect 35722 36966 35736 37018
rect 35760 36966 35774 37018
rect 35774 36966 35786 37018
rect 35786 36966 35816 37018
rect 35840 36966 35850 37018
rect 35850 36966 35896 37018
rect 35600 36964 35656 36966
rect 35680 36964 35736 36966
rect 35760 36964 35816 36966
rect 35840 36964 35896 36966
rect 37830 36760 37886 36816
rect 30562 29144 30618 29200
rect 30470 26288 30526 26344
rect 30930 26832 30986 26888
rect 31390 28600 31446 28656
rect 29918 19896 29974 19952
rect 29550 18284 29606 18320
rect 29550 18264 29552 18284
rect 29552 18264 29604 18284
rect 29604 18264 29606 18284
rect 27618 13368 27674 13424
rect 27158 13232 27214 13288
rect 27710 11600 27766 11656
rect 27986 10512 28042 10568
rect 28354 10376 28410 10432
rect 27618 9016 27674 9072
rect 28722 14900 28724 14920
rect 28724 14900 28776 14920
rect 28776 14900 28778 14920
rect 28722 14864 28778 14900
rect 28906 12044 28908 12064
rect 28908 12044 28960 12064
rect 28960 12044 28962 12064
rect 28906 12008 28962 12044
rect 30378 18284 30434 18320
rect 30378 18264 30380 18284
rect 30380 18264 30432 18284
rect 30432 18264 30434 18284
rect 31114 22344 31170 22400
rect 31206 22092 31262 22128
rect 31206 22072 31208 22092
rect 31208 22072 31260 22092
rect 31260 22072 31262 22092
rect 31114 19352 31170 19408
rect 30286 14320 30342 14376
rect 30010 10920 30066 10976
rect 29918 9560 29974 9616
rect 29826 9016 29882 9072
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 35600 35930 35656 35932
rect 35680 35930 35736 35932
rect 35760 35930 35816 35932
rect 35840 35930 35896 35932
rect 35600 35878 35646 35930
rect 35646 35878 35656 35930
rect 35680 35878 35710 35930
rect 35710 35878 35722 35930
rect 35722 35878 35736 35930
rect 35760 35878 35774 35930
rect 35774 35878 35786 35930
rect 35786 35878 35816 35930
rect 35840 35878 35850 35930
rect 35850 35878 35896 35930
rect 35600 35876 35656 35878
rect 35680 35876 35736 35878
rect 35760 35876 35816 35878
rect 35840 35876 35896 35878
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 35600 34842 35656 34844
rect 35680 34842 35736 34844
rect 35760 34842 35816 34844
rect 35840 34842 35896 34844
rect 35600 34790 35646 34842
rect 35646 34790 35656 34842
rect 35680 34790 35710 34842
rect 35710 34790 35722 34842
rect 35722 34790 35736 34842
rect 35760 34790 35774 34842
rect 35774 34790 35786 34842
rect 35786 34790 35816 34842
rect 35840 34790 35850 34842
rect 35850 34790 35896 34842
rect 35600 34788 35656 34790
rect 35680 34788 35736 34790
rect 35760 34788 35816 34790
rect 35840 34788 35896 34790
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 33782 32408 33838 32464
rect 35600 33754 35656 33756
rect 35680 33754 35736 33756
rect 35760 33754 35816 33756
rect 35840 33754 35896 33756
rect 35600 33702 35646 33754
rect 35646 33702 35656 33754
rect 35680 33702 35710 33754
rect 35710 33702 35722 33754
rect 35722 33702 35736 33754
rect 35760 33702 35774 33754
rect 35774 33702 35786 33754
rect 35786 33702 35816 33754
rect 35840 33702 35850 33754
rect 35850 33702 35896 33754
rect 35600 33700 35656 33702
rect 35680 33700 35736 33702
rect 35760 33700 35816 33702
rect 35840 33700 35896 33702
rect 37922 34040 37978 34096
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 35600 32666 35656 32668
rect 35680 32666 35736 32668
rect 35760 32666 35816 32668
rect 35840 32666 35896 32668
rect 35600 32614 35646 32666
rect 35646 32614 35656 32666
rect 35680 32614 35710 32666
rect 35710 32614 35722 32666
rect 35722 32614 35736 32666
rect 35760 32614 35774 32666
rect 35774 32614 35786 32666
rect 35786 32614 35816 32666
rect 35840 32614 35850 32666
rect 35850 32614 35896 32666
rect 35600 32612 35656 32614
rect 35680 32612 35736 32614
rect 35760 32612 35816 32614
rect 35840 32612 35896 32614
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 35600 31578 35656 31580
rect 35680 31578 35736 31580
rect 35760 31578 35816 31580
rect 35840 31578 35896 31580
rect 35600 31526 35646 31578
rect 35646 31526 35656 31578
rect 35680 31526 35710 31578
rect 35710 31526 35722 31578
rect 35722 31526 35736 31578
rect 35760 31526 35774 31578
rect 35774 31526 35786 31578
rect 35786 31526 35816 31578
rect 35840 31526 35850 31578
rect 35850 31526 35896 31578
rect 35600 31524 35656 31526
rect 35680 31524 35736 31526
rect 35760 31524 35816 31526
rect 35840 31524 35896 31526
rect 35600 30490 35656 30492
rect 35680 30490 35736 30492
rect 35760 30490 35816 30492
rect 35840 30490 35896 30492
rect 35600 30438 35646 30490
rect 35646 30438 35656 30490
rect 35680 30438 35710 30490
rect 35710 30438 35722 30490
rect 35722 30438 35736 30490
rect 35760 30438 35774 30490
rect 35774 30438 35786 30490
rect 35786 30438 35816 30490
rect 35840 30438 35850 30490
rect 35850 30438 35896 30490
rect 35600 30436 35656 30438
rect 35680 30436 35736 30438
rect 35760 30436 35816 30438
rect 35840 30436 35896 30438
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 36634 29552 36690 29608
rect 35600 29402 35656 29404
rect 35680 29402 35736 29404
rect 35760 29402 35816 29404
rect 35840 29402 35896 29404
rect 35600 29350 35646 29402
rect 35646 29350 35656 29402
rect 35680 29350 35710 29402
rect 35710 29350 35722 29402
rect 35722 29350 35736 29402
rect 35760 29350 35774 29402
rect 35774 29350 35786 29402
rect 35786 29350 35816 29402
rect 35840 29350 35850 29402
rect 35850 29350 35896 29402
rect 35600 29348 35656 29350
rect 35680 29348 35736 29350
rect 35760 29348 35816 29350
rect 35840 29348 35896 29350
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 35600 28314 35656 28316
rect 35680 28314 35736 28316
rect 35760 28314 35816 28316
rect 35840 28314 35896 28316
rect 35600 28262 35646 28314
rect 35646 28262 35656 28314
rect 35680 28262 35710 28314
rect 35710 28262 35722 28314
rect 35722 28262 35736 28314
rect 35760 28262 35774 28314
rect 35774 28262 35786 28314
rect 35786 28262 35816 28314
rect 35840 28262 35850 28314
rect 35850 28262 35896 28314
rect 35600 28260 35656 28262
rect 35680 28260 35736 28262
rect 35760 28260 35816 28262
rect 35840 28260 35896 28262
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 35600 27226 35656 27228
rect 35680 27226 35736 27228
rect 35760 27226 35816 27228
rect 35840 27226 35896 27228
rect 35600 27174 35646 27226
rect 35646 27174 35656 27226
rect 35680 27174 35710 27226
rect 35710 27174 35722 27226
rect 35722 27174 35736 27226
rect 35760 27174 35774 27226
rect 35774 27174 35786 27226
rect 35786 27174 35816 27226
rect 35840 27174 35850 27226
rect 35850 27174 35896 27226
rect 35600 27172 35656 27174
rect 35680 27172 35736 27174
rect 35760 27172 35816 27174
rect 35840 27172 35896 27174
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 35600 26138 35656 26140
rect 35680 26138 35736 26140
rect 35760 26138 35816 26140
rect 35840 26138 35896 26140
rect 35600 26086 35646 26138
rect 35646 26086 35656 26138
rect 35680 26086 35710 26138
rect 35710 26086 35722 26138
rect 35722 26086 35736 26138
rect 35760 26086 35774 26138
rect 35774 26086 35786 26138
rect 35786 26086 35816 26138
rect 35840 26086 35850 26138
rect 35850 26086 35896 26138
rect 35600 26084 35656 26086
rect 35680 26084 35736 26086
rect 35760 26084 35816 26086
rect 35840 26084 35896 26086
rect 32862 22092 32918 22128
rect 32862 22072 32864 22092
rect 32864 22072 32916 22092
rect 32916 22072 32918 22092
rect 30654 9016 30710 9072
rect 31298 10920 31354 10976
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 35600 25050 35656 25052
rect 35680 25050 35736 25052
rect 35760 25050 35816 25052
rect 35840 25050 35896 25052
rect 35600 24998 35646 25050
rect 35646 24998 35656 25050
rect 35680 24998 35710 25050
rect 35710 24998 35722 25050
rect 35722 24998 35736 25050
rect 35760 24998 35774 25050
rect 35774 24998 35786 25050
rect 35786 24998 35816 25050
rect 35840 24998 35850 25050
rect 35850 24998 35896 25050
rect 35600 24996 35656 24998
rect 35680 24996 35736 24998
rect 35760 24996 35816 24998
rect 35840 24996 35896 24998
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 35600 23962 35656 23964
rect 35680 23962 35736 23964
rect 35760 23962 35816 23964
rect 35840 23962 35896 23964
rect 35600 23910 35646 23962
rect 35646 23910 35656 23962
rect 35680 23910 35710 23962
rect 35710 23910 35722 23962
rect 35722 23910 35736 23962
rect 35760 23910 35774 23962
rect 35774 23910 35786 23962
rect 35786 23910 35816 23962
rect 35840 23910 35850 23962
rect 35850 23910 35896 23962
rect 35600 23908 35656 23910
rect 35680 23908 35736 23910
rect 35760 23908 35816 23910
rect 35840 23908 35896 23910
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 35162 23196 35164 23216
rect 35164 23196 35216 23216
rect 35216 23196 35218 23216
rect 35162 23160 35218 23196
rect 36082 23196 36084 23216
rect 36084 23196 36136 23216
rect 36136 23196 36138 23216
rect 36082 23160 36138 23196
rect 35600 22874 35656 22876
rect 35680 22874 35736 22876
rect 35760 22874 35816 22876
rect 35840 22874 35896 22876
rect 35600 22822 35646 22874
rect 35646 22822 35656 22874
rect 35680 22822 35710 22874
rect 35710 22822 35722 22874
rect 35722 22822 35736 22874
rect 35760 22822 35774 22874
rect 35774 22822 35786 22874
rect 35786 22822 35816 22874
rect 35840 22822 35850 22874
rect 35850 22822 35896 22874
rect 35600 22820 35656 22822
rect 35680 22820 35736 22822
rect 35760 22820 35816 22822
rect 35840 22820 35896 22822
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 35600 21786 35656 21788
rect 35680 21786 35736 21788
rect 35760 21786 35816 21788
rect 35840 21786 35896 21788
rect 35600 21734 35646 21786
rect 35646 21734 35656 21786
rect 35680 21734 35710 21786
rect 35710 21734 35722 21786
rect 35722 21734 35736 21786
rect 35760 21734 35774 21786
rect 35774 21734 35786 21786
rect 35786 21734 35816 21786
rect 35840 21734 35850 21786
rect 35850 21734 35896 21786
rect 35600 21732 35656 21734
rect 35680 21732 35736 21734
rect 35760 21732 35816 21734
rect 35840 21732 35896 21734
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 35070 20984 35126 21040
rect 35714 21020 35716 21040
rect 35716 21020 35768 21040
rect 35768 21020 35770 21040
rect 35714 20984 35770 21020
rect 35600 20698 35656 20700
rect 35680 20698 35736 20700
rect 35760 20698 35816 20700
rect 35840 20698 35896 20700
rect 35600 20646 35646 20698
rect 35646 20646 35656 20698
rect 35680 20646 35710 20698
rect 35710 20646 35722 20698
rect 35722 20646 35736 20698
rect 35760 20646 35774 20698
rect 35774 20646 35786 20698
rect 35786 20646 35816 20698
rect 35840 20646 35850 20698
rect 35850 20646 35896 20698
rect 35600 20644 35656 20646
rect 35680 20644 35736 20646
rect 35760 20644 35816 20646
rect 35840 20644 35896 20646
rect 33598 18264 33654 18320
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 35346 19896 35402 19952
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 35600 19610 35656 19612
rect 35680 19610 35736 19612
rect 35760 19610 35816 19612
rect 35840 19610 35896 19612
rect 35600 19558 35646 19610
rect 35646 19558 35656 19610
rect 35680 19558 35710 19610
rect 35710 19558 35722 19610
rect 35722 19558 35736 19610
rect 35760 19558 35774 19610
rect 35774 19558 35786 19610
rect 35786 19558 35816 19610
rect 35840 19558 35850 19610
rect 35850 19558 35896 19610
rect 35600 19556 35656 19558
rect 35680 19556 35736 19558
rect 35760 19556 35816 19558
rect 35840 19556 35896 19558
rect 36450 19916 36506 19952
rect 36450 19896 36452 19916
rect 36452 19896 36504 19916
rect 36504 19896 36506 19916
rect 37830 22500 37886 22536
rect 37830 22480 37832 22500
rect 37832 22480 37884 22500
rect 37884 22480 37886 22500
rect 36818 21528 36874 21584
rect 35600 18522 35656 18524
rect 35680 18522 35736 18524
rect 35760 18522 35816 18524
rect 35840 18522 35896 18524
rect 35600 18470 35646 18522
rect 35646 18470 35656 18522
rect 35680 18470 35710 18522
rect 35710 18470 35722 18522
rect 35722 18470 35736 18522
rect 35760 18470 35774 18522
rect 35774 18470 35786 18522
rect 35786 18470 35816 18522
rect 35840 18470 35850 18522
rect 35850 18470 35896 18522
rect 35600 18468 35656 18470
rect 35680 18468 35736 18470
rect 35760 18468 35816 18470
rect 35840 18468 35896 18470
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 35600 17434 35656 17436
rect 35680 17434 35736 17436
rect 35760 17434 35816 17436
rect 35840 17434 35896 17436
rect 35600 17382 35646 17434
rect 35646 17382 35656 17434
rect 35680 17382 35710 17434
rect 35710 17382 35722 17434
rect 35722 17382 35736 17434
rect 35760 17382 35774 17434
rect 35774 17382 35786 17434
rect 35786 17382 35816 17434
rect 35840 17382 35850 17434
rect 35850 17382 35896 17434
rect 35600 17380 35656 17382
rect 35680 17380 35736 17382
rect 35760 17380 35816 17382
rect 35840 17380 35896 17382
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 35600 16346 35656 16348
rect 35680 16346 35736 16348
rect 35760 16346 35816 16348
rect 35840 16346 35896 16348
rect 35600 16294 35646 16346
rect 35646 16294 35656 16346
rect 35680 16294 35710 16346
rect 35710 16294 35722 16346
rect 35722 16294 35736 16346
rect 35760 16294 35774 16346
rect 35774 16294 35786 16346
rect 35786 16294 35816 16346
rect 35840 16294 35850 16346
rect 35850 16294 35896 16346
rect 35600 16292 35656 16294
rect 35680 16292 35736 16294
rect 35760 16292 35816 16294
rect 35840 16292 35896 16294
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 35600 15258 35656 15260
rect 35680 15258 35736 15260
rect 35760 15258 35816 15260
rect 35840 15258 35896 15260
rect 35600 15206 35646 15258
rect 35646 15206 35656 15258
rect 35680 15206 35710 15258
rect 35710 15206 35722 15258
rect 35722 15206 35736 15258
rect 35760 15206 35774 15258
rect 35774 15206 35786 15258
rect 35786 15206 35816 15258
rect 35840 15206 35850 15258
rect 35850 15206 35896 15258
rect 35600 15204 35656 15206
rect 35680 15204 35736 15206
rect 35760 15204 35816 15206
rect 35840 15204 35896 15206
rect 35600 14170 35656 14172
rect 35680 14170 35736 14172
rect 35760 14170 35816 14172
rect 35840 14170 35896 14172
rect 35600 14118 35646 14170
rect 35646 14118 35656 14170
rect 35680 14118 35710 14170
rect 35710 14118 35722 14170
rect 35722 14118 35736 14170
rect 35760 14118 35774 14170
rect 35774 14118 35786 14170
rect 35786 14118 35816 14170
rect 35840 14118 35850 14170
rect 35850 14118 35896 14170
rect 35600 14116 35656 14118
rect 35680 14116 35736 14118
rect 35760 14116 35816 14118
rect 35840 14116 35896 14118
rect 35600 13082 35656 13084
rect 35680 13082 35736 13084
rect 35760 13082 35816 13084
rect 35840 13082 35896 13084
rect 35600 13030 35646 13082
rect 35646 13030 35656 13082
rect 35680 13030 35710 13082
rect 35710 13030 35722 13082
rect 35722 13030 35736 13082
rect 35760 13030 35774 13082
rect 35774 13030 35786 13082
rect 35786 13030 35816 13082
rect 35840 13030 35850 13082
rect 35850 13030 35896 13082
rect 35600 13028 35656 13030
rect 35680 13028 35736 13030
rect 35760 13028 35816 13030
rect 35840 13028 35896 13030
rect 35600 11994 35656 11996
rect 35680 11994 35736 11996
rect 35760 11994 35816 11996
rect 35840 11994 35896 11996
rect 35600 11942 35646 11994
rect 35646 11942 35656 11994
rect 35680 11942 35710 11994
rect 35710 11942 35722 11994
rect 35722 11942 35736 11994
rect 35760 11942 35774 11994
rect 35774 11942 35786 11994
rect 35786 11942 35816 11994
rect 35840 11942 35850 11994
rect 35850 11942 35896 11994
rect 35600 11940 35656 11942
rect 35680 11940 35736 11942
rect 35760 11940 35816 11942
rect 35840 11940 35896 11942
rect 35600 10906 35656 10908
rect 35680 10906 35736 10908
rect 35760 10906 35816 10908
rect 35840 10906 35896 10908
rect 35600 10854 35646 10906
rect 35646 10854 35656 10906
rect 35680 10854 35710 10906
rect 35710 10854 35722 10906
rect 35722 10854 35736 10906
rect 35760 10854 35774 10906
rect 35774 10854 35786 10906
rect 35786 10854 35816 10906
rect 35840 10854 35850 10906
rect 35850 10854 35896 10906
rect 35600 10852 35656 10854
rect 35680 10852 35736 10854
rect 35760 10852 35816 10854
rect 35840 10852 35896 10854
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 35600 9818 35656 9820
rect 35680 9818 35736 9820
rect 35760 9818 35816 9820
rect 35840 9818 35896 9820
rect 35600 9766 35646 9818
rect 35646 9766 35656 9818
rect 35680 9766 35710 9818
rect 35710 9766 35722 9818
rect 35722 9766 35736 9818
rect 35760 9766 35774 9818
rect 35774 9766 35786 9818
rect 35786 9766 35816 9818
rect 35840 9766 35850 9818
rect 35850 9766 35896 9818
rect 35600 9764 35656 9766
rect 35680 9764 35736 9766
rect 35760 9764 35816 9766
rect 35840 9764 35896 9766
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 38382 20440 38438 20496
rect 35600 8730 35656 8732
rect 35680 8730 35736 8732
rect 35760 8730 35816 8732
rect 35840 8730 35896 8732
rect 35600 8678 35646 8730
rect 35646 8678 35656 8730
rect 35680 8678 35710 8730
rect 35710 8678 35722 8730
rect 35722 8678 35736 8730
rect 35760 8678 35774 8730
rect 35774 8678 35786 8730
rect 35786 8678 35816 8730
rect 35840 8678 35850 8730
rect 35850 8678 35896 8730
rect 35600 8676 35656 8678
rect 35680 8676 35736 8678
rect 35760 8676 35816 8678
rect 35840 8676 35896 8678
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 35600 7642 35656 7644
rect 35680 7642 35736 7644
rect 35760 7642 35816 7644
rect 35840 7642 35896 7644
rect 35600 7590 35646 7642
rect 35646 7590 35656 7642
rect 35680 7590 35710 7642
rect 35710 7590 35722 7642
rect 35722 7590 35736 7642
rect 35760 7590 35774 7642
rect 35774 7590 35786 7642
rect 35786 7590 35816 7642
rect 35840 7590 35850 7642
rect 35850 7590 35896 7642
rect 35600 7588 35656 7590
rect 35680 7588 35736 7590
rect 35760 7588 35816 7590
rect 35840 7588 35896 7590
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 35600 6554 35656 6556
rect 35680 6554 35736 6556
rect 35760 6554 35816 6556
rect 35840 6554 35896 6556
rect 35600 6502 35646 6554
rect 35646 6502 35656 6554
rect 35680 6502 35710 6554
rect 35710 6502 35722 6554
rect 35722 6502 35736 6554
rect 35760 6502 35774 6554
rect 35774 6502 35786 6554
rect 35786 6502 35816 6554
rect 35840 6502 35850 6554
rect 35850 6502 35896 6554
rect 35600 6500 35656 6502
rect 35680 6500 35736 6502
rect 35760 6500 35816 6502
rect 35840 6500 35896 6502
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 35600 5466 35656 5468
rect 35680 5466 35736 5468
rect 35760 5466 35816 5468
rect 35840 5466 35896 5468
rect 35600 5414 35646 5466
rect 35646 5414 35656 5466
rect 35680 5414 35710 5466
rect 35710 5414 35722 5466
rect 35722 5414 35736 5466
rect 35760 5414 35774 5466
rect 35774 5414 35786 5466
rect 35786 5414 35816 5466
rect 35840 5414 35850 5466
rect 35850 5414 35896 5466
rect 35600 5412 35656 5414
rect 35680 5412 35736 5414
rect 35760 5412 35816 5414
rect 35840 5412 35896 5414
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 35600 4378 35656 4380
rect 35680 4378 35736 4380
rect 35760 4378 35816 4380
rect 35840 4378 35896 4380
rect 35600 4326 35646 4378
rect 35646 4326 35656 4378
rect 35680 4326 35710 4378
rect 35710 4326 35722 4378
rect 35722 4326 35736 4378
rect 35760 4326 35774 4378
rect 35774 4326 35786 4378
rect 35786 4326 35816 4378
rect 35840 4326 35850 4378
rect 35850 4326 35896 4378
rect 35600 4324 35656 4326
rect 35680 4324 35736 4326
rect 35760 4324 35816 4326
rect 35840 4324 35896 4326
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 35600 3290 35656 3292
rect 35680 3290 35736 3292
rect 35760 3290 35816 3292
rect 35840 3290 35896 3292
rect 35600 3238 35646 3290
rect 35646 3238 35656 3290
rect 35680 3238 35710 3290
rect 35710 3238 35722 3290
rect 35722 3238 35736 3290
rect 35760 3238 35774 3290
rect 35774 3238 35786 3290
rect 35786 3238 35816 3290
rect 35840 3238 35850 3290
rect 35850 3238 35896 3290
rect 35600 3236 35656 3238
rect 35680 3236 35736 3238
rect 35760 3236 35816 3238
rect 35840 3236 35896 3238
rect 38382 17720 38438 17776
rect 37830 15680 37886 15736
rect 37922 10920 37978 10976
rect 38290 8916 38292 8936
rect 38292 8916 38344 8936
rect 38344 8916 38346 8936
rect 38290 8880 38346 8916
rect 4880 2202 4936 2204
rect 4960 2202 5016 2204
rect 5040 2202 5096 2204
rect 5120 2202 5176 2204
rect 4880 2150 4926 2202
rect 4926 2150 4936 2202
rect 4960 2150 4990 2202
rect 4990 2150 5002 2202
rect 5002 2150 5016 2202
rect 5040 2150 5054 2202
rect 5054 2150 5066 2202
rect 5066 2150 5096 2202
rect 5120 2150 5130 2202
rect 5130 2150 5176 2202
rect 4880 2148 4936 2150
rect 4960 2148 5016 2150
rect 5040 2148 5096 2150
rect 5120 2148 5176 2150
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 35600 2202 35656 2204
rect 35680 2202 35736 2204
rect 35760 2202 35816 2204
rect 35840 2202 35896 2204
rect 35600 2150 35646 2202
rect 35646 2150 35656 2202
rect 35680 2150 35710 2202
rect 35710 2150 35722 2202
rect 35722 2150 35736 2202
rect 35760 2150 35774 2202
rect 35774 2150 35786 2202
rect 35786 2150 35816 2202
rect 35840 2150 35850 2202
rect 35850 2150 35896 2202
rect 35600 2148 35656 2150
rect 35680 2148 35736 2150
rect 35760 2148 35816 2150
rect 35840 2148 35896 2150
rect 37186 1400 37242 1456
<< metal3 >>
rect 0 39448 800 39568
rect 4870 39200 5186 39201
rect 4870 39136 4876 39200
rect 4940 39136 4956 39200
rect 5020 39136 5036 39200
rect 5100 39136 5116 39200
rect 5180 39136 5186 39200
rect 4870 39135 5186 39136
rect 35590 39200 35906 39201
rect 35590 39136 35596 39200
rect 35660 39136 35676 39200
rect 35740 39136 35756 39200
rect 35820 39136 35836 39200
rect 35900 39136 35906 39200
rect 35590 39135 35906 39136
rect 9806 38796 9812 38860
rect 9876 38858 9882 38860
rect 37641 38858 37707 38861
rect 9876 38856 37707 38858
rect 9876 38800 37646 38856
rect 37702 38800 37707 38856
rect 9876 38798 37707 38800
rect 9876 38796 9882 38798
rect 37641 38795 37707 38798
rect 37917 38858 37983 38861
rect 38618 38858 39418 38888
rect 37917 38856 39418 38858
rect 37917 38800 37922 38856
rect 37978 38800 39418 38856
rect 37917 38798 39418 38800
rect 37917 38795 37983 38798
rect 38618 38768 39418 38798
rect 10358 38660 10364 38724
rect 10428 38722 10434 38724
rect 15561 38722 15627 38725
rect 10428 38720 15627 38722
rect 10428 38664 15566 38720
rect 15622 38664 15627 38720
rect 10428 38662 15627 38664
rect 10428 38660 10434 38662
rect 15561 38659 15627 38662
rect 22369 38722 22435 38725
rect 22870 38722 22876 38724
rect 22369 38720 22876 38722
rect 22369 38664 22374 38720
rect 22430 38664 22876 38720
rect 22369 38662 22876 38664
rect 22369 38659 22435 38662
rect 22870 38660 22876 38662
rect 22940 38660 22946 38724
rect 23974 38660 23980 38724
rect 24044 38722 24050 38724
rect 27061 38722 27127 38725
rect 24044 38720 27127 38722
rect 24044 38664 27066 38720
rect 27122 38664 27127 38720
rect 24044 38662 27127 38664
rect 24044 38660 24050 38662
rect 27061 38659 27127 38662
rect 4210 38656 4526 38657
rect 4210 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4526 38656
rect 4210 38591 4526 38592
rect 34930 38656 35246 38657
rect 34930 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35246 38656
rect 34930 38591 35246 38592
rect 5165 38450 5231 38453
rect 25773 38450 25839 38453
rect 5165 38448 25839 38450
rect 5165 38392 5170 38448
rect 5226 38392 25778 38448
rect 25834 38392 25839 38448
rect 5165 38390 25839 38392
rect 5165 38387 5231 38390
rect 25773 38387 25839 38390
rect 4870 38112 5186 38113
rect 4870 38048 4876 38112
rect 4940 38048 4956 38112
rect 5020 38048 5036 38112
rect 5100 38048 5116 38112
rect 5180 38048 5186 38112
rect 4870 38047 5186 38048
rect 35590 38112 35906 38113
rect 35590 38048 35596 38112
rect 35660 38048 35676 38112
rect 35740 38048 35756 38112
rect 35820 38048 35836 38112
rect 35900 38048 35906 38112
rect 35590 38047 35906 38048
rect 13169 37906 13235 37909
rect 25313 37906 25379 37909
rect 13169 37904 25379 37906
rect 13169 37848 13174 37904
rect 13230 37848 25318 37904
rect 25374 37848 25379 37904
rect 13169 37846 25379 37848
rect 13169 37843 13235 37846
rect 25313 37843 25379 37846
rect 4210 37568 4526 37569
rect 4210 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4526 37568
rect 4210 37503 4526 37504
rect 34930 37568 35246 37569
rect 34930 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35246 37568
rect 34930 37503 35246 37504
rect 22134 37300 22140 37364
rect 22204 37362 22210 37364
rect 22921 37362 22987 37365
rect 22204 37360 22987 37362
rect 22204 37304 22926 37360
rect 22982 37304 22987 37360
rect 22204 37302 22987 37304
rect 22204 37300 22210 37302
rect 22921 37299 22987 37302
rect 25221 37364 25287 37365
rect 25221 37360 25268 37364
rect 25332 37362 25338 37364
rect 25221 37304 25226 37360
rect 25221 37300 25268 37304
rect 25332 37302 25378 37362
rect 25332 37300 25338 37302
rect 27838 37300 27844 37364
rect 27908 37362 27914 37364
rect 27981 37362 28047 37365
rect 27908 37360 28047 37362
rect 27908 37304 27986 37360
rect 28042 37304 28047 37360
rect 27908 37302 28047 37304
rect 27908 37300 27914 37302
rect 25221 37299 25287 37300
rect 27981 37299 28047 37302
rect 4870 37024 5186 37025
rect 4870 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5186 37024
rect 4870 36959 5186 36960
rect 35590 37024 35906 37025
rect 35590 36960 35596 37024
rect 35660 36960 35676 37024
rect 35740 36960 35756 37024
rect 35820 36960 35836 37024
rect 35900 36960 35906 37024
rect 35590 36959 35906 36960
rect 0 36818 800 36848
rect 933 36818 999 36821
rect 0 36816 999 36818
rect 0 36760 938 36816
rect 994 36760 999 36816
rect 0 36758 999 36760
rect 0 36728 800 36758
rect 933 36755 999 36758
rect 37825 36818 37891 36821
rect 38618 36818 39418 36848
rect 37825 36816 39418 36818
rect 37825 36760 37830 36816
rect 37886 36760 39418 36816
rect 37825 36758 39418 36760
rect 37825 36755 37891 36758
rect 38618 36728 39418 36758
rect 4210 36480 4526 36481
rect 4210 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4526 36480
rect 4210 36415 4526 36416
rect 34930 36480 35246 36481
rect 34930 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35246 36480
rect 34930 36415 35246 36416
rect 11513 36138 11579 36141
rect 15561 36138 15627 36141
rect 11513 36136 15627 36138
rect 11513 36080 11518 36136
rect 11574 36080 15566 36136
rect 15622 36080 15627 36136
rect 11513 36078 15627 36080
rect 11513 36075 11579 36078
rect 15561 36075 15627 36078
rect 25589 36138 25655 36141
rect 28809 36138 28875 36141
rect 25589 36136 28875 36138
rect 25589 36080 25594 36136
rect 25650 36080 28814 36136
rect 28870 36080 28875 36136
rect 25589 36078 28875 36080
rect 25589 36075 25655 36078
rect 28809 36075 28875 36078
rect 17401 36002 17467 36005
rect 17534 36002 17540 36004
rect 17401 36000 17540 36002
rect 17401 35944 17406 36000
rect 17462 35944 17540 36000
rect 17401 35942 17540 35944
rect 17401 35939 17467 35942
rect 17534 35940 17540 35942
rect 17604 35940 17610 36004
rect 20161 36002 20227 36005
rect 24945 36004 25011 36005
rect 20294 36002 20300 36004
rect 20161 36000 20300 36002
rect 20161 35944 20166 36000
rect 20222 35944 20300 36000
rect 20161 35942 20300 35944
rect 20161 35939 20227 35942
rect 20294 35940 20300 35942
rect 20364 35940 20370 36004
rect 24894 36002 24900 36004
rect 24854 35942 24900 36002
rect 24964 36000 25011 36004
rect 25006 35944 25011 36000
rect 24894 35940 24900 35942
rect 24964 35940 25011 35944
rect 24945 35939 25011 35940
rect 28441 36002 28507 36005
rect 28942 36002 28948 36004
rect 28441 36000 28948 36002
rect 28441 35944 28446 36000
rect 28502 35944 28948 36000
rect 28441 35942 28948 35944
rect 28441 35939 28507 35942
rect 28942 35940 28948 35942
rect 29012 35940 29018 36004
rect 4870 35936 5186 35937
rect 4870 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5186 35936
rect 4870 35871 5186 35872
rect 35590 35936 35906 35937
rect 35590 35872 35596 35936
rect 35660 35872 35676 35936
rect 35740 35872 35756 35936
rect 35820 35872 35836 35936
rect 35900 35872 35906 35936
rect 35590 35871 35906 35872
rect 25589 35730 25655 35733
rect 26877 35730 26943 35733
rect 25589 35728 26943 35730
rect 25589 35672 25594 35728
rect 25650 35672 26882 35728
rect 26938 35672 26943 35728
rect 25589 35670 26943 35672
rect 25589 35667 25655 35670
rect 26877 35667 26943 35670
rect 25589 35594 25655 35597
rect 26417 35594 26483 35597
rect 25589 35592 26483 35594
rect 25589 35536 25594 35592
rect 25650 35536 26422 35592
rect 26478 35536 26483 35592
rect 25589 35534 26483 35536
rect 25589 35531 25655 35534
rect 26417 35531 26483 35534
rect 4210 35392 4526 35393
rect 4210 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4526 35392
rect 4210 35327 4526 35328
rect 34930 35392 35246 35393
rect 34930 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35246 35392
rect 34930 35327 35246 35328
rect 25865 35186 25931 35189
rect 28349 35186 28415 35189
rect 25865 35184 28415 35186
rect 25865 35128 25870 35184
rect 25926 35128 28354 35184
rect 28410 35128 28415 35184
rect 25865 35126 28415 35128
rect 25865 35123 25931 35126
rect 28349 35123 28415 35126
rect 25129 34914 25195 34917
rect 19290 34912 25195 34914
rect 19290 34856 25134 34912
rect 25190 34856 25195 34912
rect 19290 34854 25195 34856
rect 4870 34848 5186 34849
rect 0 34688 800 34808
rect 4870 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5186 34848
rect 4870 34783 5186 34784
rect 13854 34580 13860 34644
rect 13924 34642 13930 34644
rect 19290 34642 19350 34854
rect 25129 34851 25195 34854
rect 35590 34848 35906 34849
rect 35590 34784 35596 34848
rect 35660 34784 35676 34848
rect 35740 34784 35756 34848
rect 35820 34784 35836 34848
rect 35900 34784 35906 34848
rect 35590 34783 35906 34784
rect 23473 34644 23539 34645
rect 23422 34642 23428 34644
rect 13924 34582 19350 34642
rect 23382 34582 23428 34642
rect 23492 34640 23539 34644
rect 23534 34584 23539 34640
rect 13924 34580 13930 34582
rect 23422 34580 23428 34582
rect 23492 34580 23539 34584
rect 23473 34579 23539 34580
rect 22277 34370 22343 34373
rect 23841 34370 23907 34373
rect 22277 34368 23907 34370
rect 22277 34312 22282 34368
rect 22338 34312 23846 34368
rect 23902 34312 23907 34368
rect 22277 34310 23907 34312
rect 22277 34307 22343 34310
rect 23841 34307 23907 34310
rect 4210 34304 4526 34305
rect 4210 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4526 34304
rect 4210 34239 4526 34240
rect 34930 34304 35246 34305
rect 34930 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35246 34304
rect 34930 34239 35246 34240
rect 19701 34098 19767 34101
rect 22921 34098 22987 34101
rect 19701 34096 22987 34098
rect 19701 34040 19706 34096
rect 19762 34040 22926 34096
rect 22982 34040 22987 34096
rect 19701 34038 22987 34040
rect 19701 34035 19767 34038
rect 22921 34035 22987 34038
rect 37917 34098 37983 34101
rect 38618 34098 39418 34128
rect 37917 34096 39418 34098
rect 37917 34040 37922 34096
rect 37978 34040 39418 34096
rect 37917 34038 39418 34040
rect 37917 34035 37983 34038
rect 38618 34008 39418 34038
rect 15653 33962 15719 33965
rect 20253 33962 20319 33965
rect 20897 33962 20963 33965
rect 15653 33960 20963 33962
rect 15653 33904 15658 33960
rect 15714 33904 20258 33960
rect 20314 33904 20902 33960
rect 20958 33904 20963 33960
rect 15653 33902 20963 33904
rect 15653 33899 15719 33902
rect 20253 33899 20319 33902
rect 20897 33899 20963 33902
rect 15561 33826 15627 33829
rect 23197 33826 23263 33829
rect 15561 33824 23263 33826
rect 15561 33768 15566 33824
rect 15622 33768 23202 33824
rect 23258 33768 23263 33824
rect 15561 33766 23263 33768
rect 15561 33763 15627 33766
rect 23197 33763 23263 33766
rect 4870 33760 5186 33761
rect 4870 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5186 33760
rect 4870 33695 5186 33696
rect 35590 33760 35906 33761
rect 35590 33696 35596 33760
rect 35660 33696 35676 33760
rect 35740 33696 35756 33760
rect 35820 33696 35836 33760
rect 35900 33696 35906 33760
rect 35590 33695 35906 33696
rect 15009 33690 15075 33693
rect 19333 33690 19399 33693
rect 15009 33688 19399 33690
rect 15009 33632 15014 33688
rect 15070 33632 19338 33688
rect 19394 33632 19399 33688
rect 15009 33630 19399 33632
rect 15009 33627 15075 33630
rect 19333 33627 19399 33630
rect 21449 33690 21515 33693
rect 23238 33690 23244 33692
rect 21449 33688 23244 33690
rect 21449 33632 21454 33688
rect 21510 33632 23244 33688
rect 21449 33630 23244 33632
rect 21449 33627 21515 33630
rect 23238 33628 23244 33630
rect 23308 33690 23314 33692
rect 23473 33690 23539 33693
rect 23308 33688 23539 33690
rect 23308 33632 23478 33688
rect 23534 33632 23539 33688
rect 23308 33630 23539 33632
rect 23308 33628 23314 33630
rect 23473 33627 23539 33630
rect 15193 33554 15259 33557
rect 17493 33554 17559 33557
rect 15193 33552 17559 33554
rect 15193 33496 15198 33552
rect 15254 33496 17498 33552
rect 17554 33496 17559 33552
rect 15193 33494 17559 33496
rect 15193 33491 15259 33494
rect 17493 33491 17559 33494
rect 20161 33554 20227 33557
rect 22829 33554 22895 33557
rect 23933 33554 23999 33557
rect 20161 33552 23999 33554
rect 20161 33496 20166 33552
rect 20222 33496 22834 33552
rect 22890 33496 23938 33552
rect 23994 33496 23999 33552
rect 20161 33494 23999 33496
rect 20161 33491 20227 33494
rect 22829 33491 22895 33494
rect 23933 33491 23999 33494
rect 23381 33418 23447 33421
rect 26182 33418 26188 33420
rect 23381 33416 26188 33418
rect 23381 33360 23386 33416
rect 23442 33360 26188 33416
rect 23381 33358 26188 33360
rect 23381 33355 23447 33358
rect 26182 33356 26188 33358
rect 26252 33356 26258 33420
rect 19057 33284 19123 33285
rect 19006 33282 19012 33284
rect 18966 33222 19012 33282
rect 19076 33280 19123 33284
rect 19118 33224 19123 33280
rect 19006 33220 19012 33222
rect 19076 33220 19123 33224
rect 19057 33219 19123 33220
rect 24025 33282 24091 33285
rect 24526 33282 24532 33284
rect 24025 33280 24532 33282
rect 24025 33224 24030 33280
rect 24086 33224 24532 33280
rect 24025 33222 24532 33224
rect 24025 33219 24091 33222
rect 24526 33220 24532 33222
rect 24596 33220 24602 33284
rect 25078 33220 25084 33284
rect 25148 33282 25154 33284
rect 25405 33282 25471 33285
rect 25148 33280 25471 33282
rect 25148 33224 25410 33280
rect 25466 33224 25471 33280
rect 25148 33222 25471 33224
rect 25148 33220 25154 33222
rect 25405 33219 25471 33222
rect 4210 33216 4526 33217
rect 4210 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4526 33216
rect 4210 33151 4526 33152
rect 34930 33216 35246 33217
rect 34930 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35246 33216
rect 34930 33151 35246 33152
rect 17861 33146 17927 33149
rect 17861 33144 17970 33146
rect 17861 33088 17866 33144
rect 17922 33088 17970 33144
rect 17861 33083 17970 33088
rect 19374 33084 19380 33148
rect 19444 33146 19450 33148
rect 19977 33146 20043 33149
rect 19444 33144 20043 33146
rect 19444 33088 19982 33144
rect 20038 33088 20043 33144
rect 19444 33086 20043 33088
rect 19444 33084 19450 33086
rect 19977 33083 20043 33086
rect 23933 33144 23999 33149
rect 23933 33088 23938 33144
rect 23994 33088 23999 33144
rect 23933 33083 23999 33088
rect 28942 33084 28948 33148
rect 29012 33146 29018 33148
rect 29545 33146 29611 33149
rect 29012 33144 29611 33146
rect 29012 33088 29550 33144
rect 29606 33088 29611 33144
rect 29012 33086 29611 33088
rect 29012 33084 29018 33086
rect 29545 33083 29611 33086
rect 17910 33010 17970 33083
rect 23936 33010 23996 33083
rect 17910 32950 23996 33010
rect 12157 32874 12223 32877
rect 20437 32874 20503 32877
rect 12157 32872 20503 32874
rect 12157 32816 12162 32872
rect 12218 32816 20442 32872
rect 20498 32816 20503 32872
rect 12157 32814 20503 32816
rect 12157 32811 12223 32814
rect 20437 32811 20503 32814
rect 4870 32672 5186 32673
rect 4870 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5186 32672
rect 4870 32607 5186 32608
rect 35590 32672 35906 32673
rect 35590 32608 35596 32672
rect 35660 32608 35676 32672
rect 35740 32608 35756 32672
rect 35820 32608 35836 32672
rect 35900 32608 35906 32672
rect 35590 32607 35906 32608
rect 21633 32466 21699 32469
rect 33777 32466 33843 32469
rect 21633 32464 33843 32466
rect 21633 32408 21638 32464
rect 21694 32408 33782 32464
rect 33838 32408 33843 32464
rect 21633 32406 33843 32408
rect 21633 32403 21699 32406
rect 33777 32403 33843 32406
rect 17125 32330 17191 32333
rect 19057 32330 19123 32333
rect 23013 32332 23079 32333
rect 23013 32330 23060 32332
rect 17125 32328 19123 32330
rect 17125 32272 17130 32328
rect 17186 32272 19062 32328
rect 19118 32272 19123 32328
rect 17125 32270 19123 32272
rect 22968 32328 23060 32330
rect 22968 32272 23018 32328
rect 22968 32270 23060 32272
rect 17125 32267 17191 32270
rect 19057 32267 19123 32270
rect 23013 32268 23060 32270
rect 23124 32268 23130 32332
rect 23197 32330 23263 32333
rect 24485 32330 24551 32333
rect 23197 32328 24551 32330
rect 23197 32272 23202 32328
rect 23258 32272 24490 32328
rect 24546 32272 24551 32328
rect 23197 32270 24551 32272
rect 23013 32267 23079 32268
rect 23197 32267 23263 32270
rect 24485 32267 24551 32270
rect 12617 32194 12683 32197
rect 20110 32194 20116 32196
rect 12617 32192 20116 32194
rect 12617 32136 12622 32192
rect 12678 32136 20116 32192
rect 12617 32134 20116 32136
rect 12617 32131 12683 32134
rect 20110 32132 20116 32134
rect 20180 32132 20186 32196
rect 4210 32128 4526 32129
rect 0 31968 800 32088
rect 4210 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4526 32128
rect 4210 32063 4526 32064
rect 34930 32128 35246 32129
rect 34930 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35246 32128
rect 34930 32063 35246 32064
rect 18413 32060 18479 32061
rect 18413 32056 18460 32060
rect 18524 32058 18530 32060
rect 21725 32058 21791 32061
rect 25405 32058 25471 32061
rect 18413 32000 18418 32056
rect 18413 31996 18460 32000
rect 18524 31998 18570 32058
rect 21725 32056 25471 32058
rect 21725 32000 21730 32056
rect 21786 32000 25410 32056
rect 25466 32000 25471 32056
rect 21725 31998 25471 32000
rect 18524 31996 18530 31998
rect 18413 31995 18479 31996
rect 21725 31995 21791 31998
rect 25405 31995 25471 31998
rect 38618 31968 39418 32088
rect 13077 31922 13143 31925
rect 18873 31922 18939 31925
rect 26693 31922 26759 31925
rect 28942 31922 28948 31924
rect 13077 31920 28948 31922
rect 13077 31864 13082 31920
rect 13138 31864 18878 31920
rect 18934 31864 26698 31920
rect 26754 31864 28948 31920
rect 13077 31862 28948 31864
rect 13077 31859 13143 31862
rect 18873 31859 18939 31862
rect 26693 31859 26759 31862
rect 28942 31860 28948 31862
rect 29012 31860 29018 31924
rect 21081 31786 21147 31789
rect 21081 31784 22202 31786
rect 21081 31728 21086 31784
rect 21142 31728 22202 31784
rect 21081 31726 22202 31728
rect 21081 31723 21147 31726
rect 17309 31650 17375 31653
rect 20345 31650 20411 31653
rect 21633 31650 21699 31653
rect 17309 31648 21699 31650
rect 17309 31592 17314 31648
rect 17370 31592 20350 31648
rect 20406 31592 21638 31648
rect 21694 31592 21699 31648
rect 17309 31590 21699 31592
rect 17309 31587 17375 31590
rect 20345 31587 20411 31590
rect 21633 31587 21699 31590
rect 4870 31584 5186 31585
rect 4870 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5186 31584
rect 4870 31519 5186 31520
rect 16297 31514 16363 31517
rect 21541 31514 21607 31517
rect 16297 31512 21607 31514
rect 16297 31456 16302 31512
rect 16358 31456 21546 31512
rect 21602 31456 21607 31512
rect 16297 31454 21607 31456
rect 16297 31451 16363 31454
rect 21541 31451 21607 31454
rect 21725 31378 21791 31381
rect 22142 31378 22202 31726
rect 35590 31584 35906 31585
rect 35590 31520 35596 31584
rect 35660 31520 35676 31584
rect 35740 31520 35756 31584
rect 35820 31520 35836 31584
rect 35900 31520 35906 31584
rect 35590 31519 35906 31520
rect 23381 31380 23447 31381
rect 23381 31378 23428 31380
rect 21725 31376 22202 31378
rect 21725 31320 21730 31376
rect 21786 31320 22202 31376
rect 21725 31318 22202 31320
rect 23336 31376 23428 31378
rect 23336 31320 23386 31376
rect 23336 31318 23428 31320
rect 21725 31315 21791 31318
rect 23381 31316 23428 31318
rect 23492 31316 23498 31380
rect 23381 31315 23447 31316
rect 19333 31242 19399 31245
rect 20713 31242 20779 31245
rect 23749 31242 23815 31245
rect 19333 31240 23815 31242
rect 19333 31184 19338 31240
rect 19394 31184 20718 31240
rect 20774 31184 23754 31240
rect 23810 31184 23815 31240
rect 19333 31182 23815 31184
rect 19333 31179 19399 31182
rect 20713 31179 20779 31182
rect 23749 31179 23815 31182
rect 19977 31106 20043 31109
rect 22277 31106 22343 31109
rect 19977 31104 22343 31106
rect 19977 31048 19982 31104
rect 20038 31048 22282 31104
rect 22338 31048 22343 31104
rect 19977 31046 22343 31048
rect 19977 31043 20043 31046
rect 22277 31043 22343 31046
rect 27705 31106 27771 31109
rect 27838 31106 27844 31108
rect 27705 31104 27844 31106
rect 27705 31048 27710 31104
rect 27766 31048 27844 31104
rect 27705 31046 27844 31048
rect 27705 31043 27771 31046
rect 27838 31044 27844 31046
rect 27908 31044 27914 31108
rect 4210 31040 4526 31041
rect 4210 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4526 31040
rect 4210 30975 4526 30976
rect 34930 31040 35246 31041
rect 34930 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35246 31040
rect 34930 30975 35246 30976
rect 19425 30970 19491 30973
rect 20621 30970 20687 30973
rect 19425 30968 20687 30970
rect 19425 30912 19430 30968
rect 19486 30912 20626 30968
rect 20682 30912 20687 30968
rect 19425 30910 20687 30912
rect 19425 30907 19491 30910
rect 20621 30907 20687 30910
rect 19057 30698 19123 30701
rect 30189 30698 30255 30701
rect 19057 30696 30255 30698
rect 19057 30640 19062 30696
rect 19118 30640 30194 30696
rect 30250 30640 30255 30696
rect 19057 30638 30255 30640
rect 19057 30635 19123 30638
rect 30189 30635 30255 30638
rect 4870 30496 5186 30497
rect 4870 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5186 30496
rect 4870 30431 5186 30432
rect 35590 30496 35906 30497
rect 35590 30432 35596 30496
rect 35660 30432 35676 30496
rect 35740 30432 35756 30496
rect 35820 30432 35836 30496
rect 35900 30432 35906 30496
rect 35590 30431 35906 30432
rect 18321 30428 18387 30429
rect 18270 30426 18276 30428
rect 18230 30366 18276 30426
rect 18340 30424 18387 30428
rect 18382 30368 18387 30424
rect 18270 30364 18276 30366
rect 18340 30364 18387 30368
rect 18321 30363 18387 30364
rect 23381 30426 23447 30429
rect 26693 30428 26759 30429
rect 23974 30426 23980 30428
rect 23381 30424 23980 30426
rect 23381 30368 23386 30424
rect 23442 30368 23980 30424
rect 23381 30366 23980 30368
rect 23381 30363 23447 30366
rect 23974 30364 23980 30366
rect 24044 30364 24050 30428
rect 26693 30424 26740 30428
rect 26804 30426 26810 30428
rect 26693 30368 26698 30424
rect 26693 30364 26740 30368
rect 26804 30366 26850 30426
rect 26804 30364 26810 30366
rect 26693 30363 26759 30364
rect 16665 30290 16731 30293
rect 18137 30290 18203 30293
rect 16665 30288 18203 30290
rect 16665 30232 16670 30288
rect 16726 30232 18142 30288
rect 18198 30232 18203 30288
rect 16665 30230 18203 30232
rect 16665 30227 16731 30230
rect 18137 30227 18203 30230
rect 24025 30290 24091 30293
rect 24894 30290 24900 30292
rect 24025 30288 24900 30290
rect 24025 30232 24030 30288
rect 24086 30232 24900 30288
rect 24025 30230 24900 30232
rect 24025 30227 24091 30230
rect 24894 30228 24900 30230
rect 24964 30228 24970 30292
rect 15653 30154 15719 30157
rect 18413 30154 18479 30157
rect 25865 30154 25931 30157
rect 30373 30154 30439 30157
rect 15653 30152 30439 30154
rect 15653 30096 15658 30152
rect 15714 30096 18418 30152
rect 18474 30096 25870 30152
rect 25926 30096 30378 30152
rect 30434 30096 30439 30152
rect 15653 30094 30439 30096
rect 15653 30091 15719 30094
rect 18413 30091 18479 30094
rect 25865 30091 25931 30094
rect 30373 30091 30439 30094
rect 0 29928 800 30048
rect 19977 30018 20043 30021
rect 24853 30018 24919 30021
rect 19977 30016 24919 30018
rect 19977 29960 19982 30016
rect 20038 29960 24858 30016
rect 24914 29960 24919 30016
rect 19977 29958 24919 29960
rect 19977 29955 20043 29958
rect 24853 29955 24919 29958
rect 25589 30018 25655 30021
rect 26877 30018 26943 30021
rect 25589 30016 26943 30018
rect 25589 29960 25594 30016
rect 25650 29960 26882 30016
rect 26938 29960 26943 30016
rect 25589 29958 26943 29960
rect 25589 29955 25655 29958
rect 26877 29955 26943 29958
rect 4210 29952 4526 29953
rect 4210 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4526 29952
rect 4210 29887 4526 29888
rect 34930 29952 35246 29953
rect 34930 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35246 29952
rect 34930 29887 35246 29888
rect 25773 29882 25839 29885
rect 26601 29882 26667 29885
rect 25773 29880 26667 29882
rect 25773 29824 25778 29880
rect 25834 29824 26606 29880
rect 26662 29824 26667 29880
rect 25773 29822 26667 29824
rect 25773 29819 25839 29822
rect 26601 29819 26667 29822
rect 15193 29746 15259 29749
rect 22277 29746 22343 29749
rect 15193 29744 22343 29746
rect 15193 29688 15198 29744
rect 15254 29688 22282 29744
rect 22338 29688 22343 29744
rect 15193 29686 22343 29688
rect 15193 29683 15259 29686
rect 22277 29683 22343 29686
rect 15837 29610 15903 29613
rect 18873 29610 18939 29613
rect 23289 29610 23355 29613
rect 15837 29608 18939 29610
rect 15837 29552 15842 29608
rect 15898 29552 18878 29608
rect 18934 29552 18939 29608
rect 15837 29550 18939 29552
rect 15837 29547 15903 29550
rect 18873 29547 18939 29550
rect 22326 29608 23355 29610
rect 22326 29552 23294 29608
rect 23350 29552 23355 29608
rect 22326 29550 23355 29552
rect 18413 29474 18479 29477
rect 22326 29474 22386 29550
rect 23289 29547 23355 29550
rect 24577 29610 24643 29613
rect 28441 29610 28507 29613
rect 24577 29608 28507 29610
rect 24577 29552 24582 29608
rect 24638 29552 28446 29608
rect 28502 29552 28507 29608
rect 24577 29550 28507 29552
rect 24577 29547 24643 29550
rect 28441 29547 28507 29550
rect 29821 29610 29887 29613
rect 36629 29610 36695 29613
rect 29821 29608 36695 29610
rect 29821 29552 29826 29608
rect 29882 29552 36634 29608
rect 36690 29552 36695 29608
rect 29821 29550 36695 29552
rect 29821 29547 29887 29550
rect 36629 29547 36695 29550
rect 18413 29472 22386 29474
rect 18413 29416 18418 29472
rect 18474 29416 22386 29472
rect 18413 29414 22386 29416
rect 22461 29474 22527 29477
rect 23105 29474 23171 29477
rect 22461 29472 23171 29474
rect 22461 29416 22466 29472
rect 22522 29416 23110 29472
rect 23166 29416 23171 29472
rect 22461 29414 23171 29416
rect 18413 29411 18479 29414
rect 22461 29411 22527 29414
rect 23105 29411 23171 29414
rect 4870 29408 5186 29409
rect 4870 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5186 29408
rect 4870 29343 5186 29344
rect 35590 29408 35906 29409
rect 35590 29344 35596 29408
rect 35660 29344 35676 29408
rect 35740 29344 35756 29408
rect 35820 29344 35836 29408
rect 35900 29344 35906 29408
rect 35590 29343 35906 29344
rect 8385 29338 8451 29341
rect 19333 29338 19399 29341
rect 8385 29336 19399 29338
rect 8385 29280 8390 29336
rect 8446 29280 19338 29336
rect 19394 29280 19399 29336
rect 8385 29278 19399 29280
rect 8385 29275 8451 29278
rect 19333 29275 19399 29278
rect 20805 29338 20871 29341
rect 24025 29338 24091 29341
rect 20805 29336 24091 29338
rect 20805 29280 20810 29336
rect 20866 29280 24030 29336
rect 24086 29280 24091 29336
rect 20805 29278 24091 29280
rect 20805 29275 20871 29278
rect 24025 29275 24091 29278
rect 38618 29248 39418 29368
rect 18229 29202 18295 29205
rect 20897 29202 20963 29205
rect 30557 29202 30623 29205
rect 18229 29200 30623 29202
rect 18229 29144 18234 29200
rect 18290 29144 20902 29200
rect 20958 29144 30562 29200
rect 30618 29144 30623 29200
rect 18229 29142 30623 29144
rect 18229 29139 18295 29142
rect 20897 29139 20963 29142
rect 30557 29139 30623 29142
rect 5625 29066 5691 29069
rect 9581 29066 9647 29069
rect 5625 29064 9647 29066
rect 5625 29008 5630 29064
rect 5686 29008 9586 29064
rect 9642 29008 9647 29064
rect 5625 29006 9647 29008
rect 5625 29003 5691 29006
rect 9581 29003 9647 29006
rect 12893 29066 12959 29069
rect 13302 29066 13308 29068
rect 12893 29064 13308 29066
rect 12893 29008 12898 29064
rect 12954 29008 13308 29064
rect 12893 29006 13308 29008
rect 12893 29003 12959 29006
rect 13302 29004 13308 29006
rect 13372 29004 13378 29068
rect 16430 29004 16436 29068
rect 16500 29066 16506 29068
rect 18873 29066 18939 29069
rect 16500 29064 18939 29066
rect 16500 29008 18878 29064
rect 18934 29008 18939 29064
rect 16500 29006 18939 29008
rect 16500 29004 16506 29006
rect 18873 29003 18939 29006
rect 21081 29066 21147 29069
rect 23565 29068 23631 29069
rect 23238 29066 23244 29068
rect 21081 29064 23244 29066
rect 21081 29008 21086 29064
rect 21142 29008 23244 29064
rect 21081 29006 23244 29008
rect 21081 29003 21147 29006
rect 23238 29004 23244 29006
rect 23308 29004 23314 29068
rect 23565 29064 23612 29068
rect 23676 29066 23682 29068
rect 23565 29008 23570 29064
rect 23565 29004 23612 29008
rect 23676 29006 23722 29066
rect 23676 29004 23682 29006
rect 24158 29004 24164 29068
rect 24228 29066 24234 29068
rect 24853 29066 24919 29069
rect 24228 29064 24919 29066
rect 24228 29008 24858 29064
rect 24914 29008 24919 29064
rect 24228 29006 24919 29008
rect 24228 29004 24234 29006
rect 23565 29003 23631 29004
rect 24853 29003 24919 29006
rect 25865 29066 25931 29069
rect 26233 29066 26299 29069
rect 25865 29064 26299 29066
rect 25865 29008 25870 29064
rect 25926 29008 26238 29064
rect 26294 29008 26299 29064
rect 25865 29006 26299 29008
rect 25865 29003 25931 29006
rect 26233 29003 26299 29006
rect 4210 28864 4526 28865
rect 4210 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4526 28864
rect 4210 28799 4526 28800
rect 34930 28864 35246 28865
rect 34930 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35246 28864
rect 34930 28799 35246 28800
rect 20253 28660 20319 28661
rect 20253 28658 20300 28660
rect 20172 28656 20300 28658
rect 20364 28658 20370 28660
rect 22737 28658 22803 28661
rect 20364 28656 22803 28658
rect 20172 28600 20258 28656
rect 20364 28600 22742 28656
rect 22798 28600 22803 28656
rect 20172 28598 20300 28600
rect 20253 28596 20300 28598
rect 20364 28598 22803 28600
rect 20364 28596 20370 28598
rect 20253 28595 20319 28596
rect 22737 28595 22803 28598
rect 29085 28658 29151 28661
rect 31385 28658 31451 28661
rect 29085 28656 31451 28658
rect 29085 28600 29090 28656
rect 29146 28600 31390 28656
rect 31446 28600 31451 28656
rect 29085 28598 31451 28600
rect 29085 28595 29151 28598
rect 31385 28595 31451 28598
rect 19609 28522 19675 28525
rect 24853 28522 24919 28525
rect 19609 28520 24919 28522
rect 19609 28464 19614 28520
rect 19670 28464 24858 28520
rect 24914 28464 24919 28520
rect 19609 28462 24919 28464
rect 19609 28459 19675 28462
rect 24853 28459 24919 28462
rect 4870 28320 5186 28321
rect 4870 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5186 28320
rect 4870 28255 5186 28256
rect 35590 28320 35906 28321
rect 35590 28256 35596 28320
rect 35660 28256 35676 28320
rect 35740 28256 35756 28320
rect 35820 28256 35836 28320
rect 35900 28256 35906 28320
rect 35590 28255 35906 28256
rect 19425 28250 19491 28253
rect 19793 28250 19859 28253
rect 19425 28248 19859 28250
rect 19425 28192 19430 28248
rect 19486 28192 19798 28248
rect 19854 28192 19859 28248
rect 19425 28190 19859 28192
rect 19425 28187 19491 28190
rect 19793 28187 19859 28190
rect 11237 28114 11303 28117
rect 17401 28114 17467 28117
rect 11237 28112 17467 28114
rect 11237 28056 11242 28112
rect 11298 28056 17406 28112
rect 17462 28056 17467 28112
rect 11237 28054 17467 28056
rect 11237 28051 11303 28054
rect 17401 28051 17467 28054
rect 19609 28114 19675 28117
rect 26693 28114 26759 28117
rect 19609 28112 26759 28114
rect 19609 28056 19614 28112
rect 19670 28056 26698 28112
rect 26754 28056 26759 28112
rect 19609 28054 26759 28056
rect 19609 28051 19675 28054
rect 26693 28051 26759 28054
rect 19241 27978 19307 27981
rect 20437 27978 20503 27981
rect 21081 27978 21147 27981
rect 19241 27976 21147 27978
rect 19241 27920 19246 27976
rect 19302 27920 20442 27976
rect 20498 27920 21086 27976
rect 21142 27920 21147 27976
rect 19241 27918 21147 27920
rect 19241 27915 19307 27918
rect 20437 27915 20503 27918
rect 21081 27915 21147 27918
rect 22921 27978 22987 27981
rect 23054 27978 23060 27980
rect 22921 27976 23060 27978
rect 22921 27920 22926 27976
rect 22982 27920 23060 27976
rect 22921 27918 23060 27920
rect 22921 27915 22987 27918
rect 23054 27916 23060 27918
rect 23124 27916 23130 27980
rect 28942 27916 28948 27980
rect 29012 27978 29018 27980
rect 29913 27978 29979 27981
rect 29012 27976 29979 27978
rect 29012 27920 29918 27976
rect 29974 27920 29979 27976
rect 29012 27918 29979 27920
rect 29012 27916 29018 27918
rect 29913 27915 29979 27918
rect 22369 27842 22435 27845
rect 24761 27842 24827 27845
rect 22369 27840 24827 27842
rect 22369 27784 22374 27840
rect 22430 27784 24766 27840
rect 24822 27784 24827 27840
rect 22369 27782 24827 27784
rect 22369 27779 22435 27782
rect 24761 27779 24827 27782
rect 4210 27776 4526 27777
rect 4210 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4526 27776
rect 4210 27711 4526 27712
rect 34930 27776 35246 27777
rect 34930 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35246 27776
rect 34930 27711 35246 27712
rect 21909 27708 21975 27709
rect 21909 27704 21956 27708
rect 22020 27706 22026 27708
rect 21909 27648 21914 27704
rect 21909 27644 21956 27648
rect 22020 27646 22066 27706
rect 22020 27644 22026 27646
rect 21909 27643 21975 27644
rect 0 27298 800 27328
rect 4061 27298 4127 27301
rect 0 27296 4127 27298
rect 0 27240 4066 27296
rect 4122 27240 4127 27296
rect 0 27238 4127 27240
rect 0 27208 800 27238
rect 4061 27235 4127 27238
rect 4870 27232 5186 27233
rect 4870 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5186 27232
rect 4870 27167 5186 27168
rect 35590 27232 35906 27233
rect 35590 27168 35596 27232
rect 35660 27168 35676 27232
rect 35740 27168 35756 27232
rect 35820 27168 35836 27232
rect 35900 27168 35906 27232
rect 38618 27208 39418 27328
rect 35590 27167 35906 27168
rect 26509 27026 26575 27029
rect 19014 27024 26575 27026
rect 19014 26968 26514 27024
rect 26570 26968 26575 27024
rect 19014 26966 26575 26968
rect 19014 26893 19074 26966
rect 26509 26963 26575 26966
rect 14733 26890 14799 26893
rect 18965 26890 19074 26893
rect 30925 26890 30991 26893
rect 14733 26888 19074 26890
rect 14733 26832 14738 26888
rect 14794 26832 18970 26888
rect 19026 26832 19074 26888
rect 14733 26830 19074 26832
rect 19290 26888 30991 26890
rect 19290 26832 30930 26888
rect 30986 26832 30991 26888
rect 19290 26830 30991 26832
rect 14733 26827 14799 26830
rect 18965 26827 19031 26830
rect 17125 26754 17191 26757
rect 19290 26754 19350 26830
rect 30925 26827 30991 26830
rect 17125 26752 19350 26754
rect 17125 26696 17130 26752
rect 17186 26696 19350 26752
rect 17125 26694 19350 26696
rect 21909 26754 21975 26757
rect 26233 26754 26299 26757
rect 21909 26752 26299 26754
rect 21909 26696 21914 26752
rect 21970 26696 26238 26752
rect 26294 26696 26299 26752
rect 21909 26694 26299 26696
rect 17125 26691 17191 26694
rect 21909 26691 21975 26694
rect 26233 26691 26299 26694
rect 4210 26688 4526 26689
rect 4210 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4526 26688
rect 4210 26623 4526 26624
rect 34930 26688 35246 26689
rect 34930 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35246 26688
rect 34930 26623 35246 26624
rect 13537 26618 13603 26621
rect 17769 26618 17835 26621
rect 13537 26616 17835 26618
rect 13537 26560 13542 26616
rect 13598 26560 17774 26616
rect 17830 26560 17835 26616
rect 13537 26558 17835 26560
rect 13537 26555 13603 26558
rect 17769 26555 17835 26558
rect 19149 26618 19215 26621
rect 23013 26618 23079 26621
rect 19149 26616 23079 26618
rect 19149 26560 19154 26616
rect 19210 26560 23018 26616
rect 23074 26560 23079 26616
rect 19149 26558 23079 26560
rect 19149 26555 19215 26558
rect 23013 26555 23079 26558
rect 20345 26482 20411 26485
rect 24577 26482 24643 26485
rect 20345 26480 24643 26482
rect 20345 26424 20350 26480
rect 20406 26424 24582 26480
rect 24638 26424 24643 26480
rect 20345 26422 24643 26424
rect 20345 26419 20411 26422
rect 24577 26419 24643 26422
rect 25037 26482 25103 26485
rect 28257 26482 28323 26485
rect 25037 26480 28323 26482
rect 25037 26424 25042 26480
rect 25098 26424 28262 26480
rect 28318 26424 28323 26480
rect 25037 26422 28323 26424
rect 25037 26419 25103 26422
rect 28257 26419 28323 26422
rect 18781 26346 18847 26349
rect 20662 26346 20668 26348
rect 18781 26344 20668 26346
rect 18781 26288 18786 26344
rect 18842 26288 20668 26344
rect 18781 26286 20668 26288
rect 18781 26283 18847 26286
rect 20662 26284 20668 26286
rect 20732 26284 20738 26348
rect 22737 26346 22803 26349
rect 26693 26346 26759 26349
rect 30465 26346 30531 26349
rect 22737 26344 30531 26346
rect 22737 26288 22742 26344
rect 22798 26288 26698 26344
rect 26754 26288 30470 26344
rect 30526 26288 30531 26344
rect 22737 26286 30531 26288
rect 22737 26283 22803 26286
rect 26693 26283 26759 26286
rect 30465 26283 30531 26286
rect 20621 26210 20687 26213
rect 24853 26210 24919 26213
rect 25313 26212 25379 26213
rect 20621 26208 24919 26210
rect 20621 26152 20626 26208
rect 20682 26152 24858 26208
rect 24914 26152 24919 26208
rect 20621 26150 24919 26152
rect 20621 26147 20687 26150
rect 24853 26147 24919 26150
rect 25262 26148 25268 26212
rect 25332 26210 25379 26212
rect 25332 26208 25424 26210
rect 25374 26152 25424 26208
rect 25332 26150 25424 26152
rect 25332 26148 25379 26150
rect 25270 26147 25379 26148
rect 4870 26144 5186 26145
rect 4870 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5186 26144
rect 4870 26079 5186 26080
rect 17585 26074 17651 26077
rect 19149 26074 19215 26077
rect 22829 26074 22895 26077
rect 17585 26072 22895 26074
rect 17585 26016 17590 26072
rect 17646 26016 19154 26072
rect 19210 26016 22834 26072
rect 22890 26016 22895 26072
rect 17585 26014 22895 26016
rect 17585 26011 17651 26014
rect 19149 26011 19215 26014
rect 22829 26011 22895 26014
rect 24025 26074 24091 26077
rect 24158 26074 24164 26076
rect 24025 26072 24164 26074
rect 24025 26016 24030 26072
rect 24086 26016 24164 26072
rect 24025 26014 24164 26016
rect 24025 26011 24091 26014
rect 24158 26012 24164 26014
rect 24228 26012 24234 26076
rect 25037 26074 25103 26077
rect 25270 26074 25330 26147
rect 35590 26144 35906 26145
rect 35590 26080 35596 26144
rect 35660 26080 35676 26144
rect 35740 26080 35756 26144
rect 35820 26080 35836 26144
rect 35900 26080 35906 26144
rect 35590 26079 35906 26080
rect 25037 26072 25330 26074
rect 25037 26016 25042 26072
rect 25098 26016 25330 26072
rect 25037 26014 25330 26016
rect 25037 26011 25103 26014
rect 13905 25938 13971 25941
rect 23105 25938 23171 25941
rect 13905 25936 23171 25938
rect 13905 25880 13910 25936
rect 13966 25880 23110 25936
rect 23166 25880 23171 25936
rect 13905 25878 23171 25880
rect 13905 25875 13971 25878
rect 23105 25875 23171 25878
rect 24301 25938 24367 25941
rect 26141 25938 26207 25941
rect 24301 25936 26207 25938
rect 24301 25880 24306 25936
rect 24362 25880 26146 25936
rect 26202 25880 26207 25936
rect 24301 25878 26207 25880
rect 24301 25875 24367 25878
rect 26141 25875 26207 25878
rect 19333 25802 19399 25805
rect 20069 25802 20135 25805
rect 19333 25800 20135 25802
rect 19333 25744 19338 25800
rect 19394 25744 20074 25800
rect 20130 25744 20135 25800
rect 19333 25742 20135 25744
rect 19333 25739 19399 25742
rect 20069 25739 20135 25742
rect 21449 25802 21515 25805
rect 25313 25802 25379 25805
rect 21449 25800 25379 25802
rect 21449 25744 21454 25800
rect 21510 25744 25318 25800
rect 25374 25744 25379 25800
rect 21449 25742 25379 25744
rect 21449 25739 21515 25742
rect 25313 25739 25379 25742
rect 4210 25600 4526 25601
rect 4210 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4526 25600
rect 4210 25535 4526 25536
rect 34930 25600 35246 25601
rect 34930 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35246 25600
rect 34930 25535 35246 25536
rect 24945 25394 25011 25397
rect 26049 25394 26115 25397
rect 24945 25392 26115 25394
rect 24945 25336 24950 25392
rect 25006 25336 26054 25392
rect 26110 25336 26115 25392
rect 24945 25334 26115 25336
rect 24945 25331 25011 25334
rect 26049 25331 26115 25334
rect 0 25258 800 25288
rect 933 25258 999 25261
rect 0 25256 999 25258
rect 0 25200 938 25256
rect 994 25200 999 25256
rect 0 25198 999 25200
rect 0 25168 800 25198
rect 933 25195 999 25198
rect 38618 25168 39418 25288
rect 12341 25122 12407 25125
rect 19374 25122 19380 25124
rect 12341 25120 19380 25122
rect 12341 25064 12346 25120
rect 12402 25064 19380 25120
rect 12341 25062 19380 25064
rect 12341 25059 12407 25062
rect 19374 25060 19380 25062
rect 19444 25122 19450 25124
rect 20529 25122 20595 25125
rect 19444 25120 20595 25122
rect 19444 25064 20534 25120
rect 20590 25064 20595 25120
rect 19444 25062 20595 25064
rect 19444 25060 19450 25062
rect 20529 25059 20595 25062
rect 4870 25056 5186 25057
rect 4870 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5186 25056
rect 4870 24991 5186 24992
rect 35590 25056 35906 25057
rect 35590 24992 35596 25056
rect 35660 24992 35676 25056
rect 35740 24992 35756 25056
rect 35820 24992 35836 25056
rect 35900 24992 35906 25056
rect 35590 24991 35906 24992
rect 14457 24986 14523 24989
rect 15510 24986 15516 24988
rect 14457 24984 15516 24986
rect 14457 24928 14462 24984
rect 14518 24928 15516 24984
rect 14457 24926 15516 24928
rect 14457 24923 14523 24926
rect 15510 24924 15516 24926
rect 15580 24924 15586 24988
rect 19333 24986 19399 24989
rect 21449 24986 21515 24989
rect 19333 24984 21515 24986
rect 19333 24928 19338 24984
rect 19394 24928 21454 24984
rect 21510 24928 21515 24984
rect 19333 24926 21515 24928
rect 19333 24923 19399 24926
rect 21449 24923 21515 24926
rect 12985 24714 13051 24717
rect 24025 24714 24091 24717
rect 27797 24714 27863 24717
rect 12985 24712 27863 24714
rect 12985 24656 12990 24712
rect 13046 24656 24030 24712
rect 24086 24656 27802 24712
rect 27858 24656 27863 24712
rect 12985 24654 27863 24656
rect 12985 24651 13051 24654
rect 24025 24651 24091 24654
rect 27797 24651 27863 24654
rect 4210 24512 4526 24513
rect 4210 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4526 24512
rect 4210 24447 4526 24448
rect 34930 24512 35246 24513
rect 34930 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35246 24512
rect 34930 24447 35246 24448
rect 9857 24306 9923 24309
rect 22185 24308 22251 24309
rect 22134 24306 22140 24308
rect 9857 24304 22140 24306
rect 22204 24306 22251 24308
rect 22204 24304 22332 24306
rect 9857 24248 9862 24304
rect 9918 24248 22140 24304
rect 22246 24248 22332 24304
rect 9857 24246 22140 24248
rect 9857 24243 9923 24246
rect 22134 24244 22140 24246
rect 22204 24246 22332 24248
rect 22204 24244 22251 24246
rect 22185 24243 22251 24244
rect 16665 24170 16731 24173
rect 17861 24170 17927 24173
rect 16665 24168 17927 24170
rect 16665 24112 16670 24168
rect 16726 24112 17866 24168
rect 17922 24112 17927 24168
rect 16665 24110 17927 24112
rect 16665 24107 16731 24110
rect 17861 24107 17927 24110
rect 4870 23968 5186 23969
rect 4870 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5186 23968
rect 4870 23903 5186 23904
rect 35590 23968 35906 23969
rect 35590 23904 35596 23968
rect 35660 23904 35676 23968
rect 35740 23904 35756 23968
rect 35820 23904 35836 23968
rect 35900 23904 35906 23968
rect 35590 23903 35906 23904
rect 14273 23762 14339 23765
rect 19425 23762 19491 23765
rect 22829 23762 22895 23765
rect 14273 23760 22895 23762
rect 14273 23704 14278 23760
rect 14334 23704 19430 23760
rect 19486 23704 22834 23760
rect 22890 23704 22895 23760
rect 14273 23702 22895 23704
rect 14273 23699 14339 23702
rect 19425 23699 19491 23702
rect 22829 23699 22895 23702
rect 13721 23626 13787 23629
rect 24301 23626 24367 23629
rect 13721 23624 24367 23626
rect 13721 23568 13726 23624
rect 13782 23568 24306 23624
rect 24362 23568 24367 23624
rect 13721 23566 24367 23568
rect 13721 23563 13787 23566
rect 24301 23563 24367 23566
rect 12617 23492 12683 23493
rect 12566 23490 12572 23492
rect 12526 23430 12572 23490
rect 12636 23488 12683 23492
rect 12678 23432 12683 23488
rect 12566 23428 12572 23430
rect 12636 23428 12683 23432
rect 12617 23427 12683 23428
rect 13905 23490 13971 23493
rect 18045 23490 18111 23493
rect 13905 23488 18111 23490
rect 13905 23432 13910 23488
rect 13966 23432 18050 23488
rect 18106 23432 18111 23488
rect 13905 23430 18111 23432
rect 13905 23427 13971 23430
rect 18045 23427 18111 23430
rect 4210 23424 4526 23425
rect 4210 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4526 23424
rect 4210 23359 4526 23360
rect 34930 23424 35246 23425
rect 34930 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35246 23424
rect 34930 23359 35246 23360
rect 0 23128 800 23248
rect 35157 23218 35223 23221
rect 36077 23218 36143 23221
rect 35157 23216 36143 23218
rect 35157 23160 35162 23216
rect 35218 23160 36082 23216
rect 36138 23160 36143 23216
rect 35157 23158 36143 23160
rect 35157 23155 35223 23158
rect 36077 23155 36143 23158
rect 4889 23082 4955 23085
rect 7925 23082 7991 23085
rect 25957 23082 26023 23085
rect 4889 23080 26023 23082
rect 4889 23024 4894 23080
rect 4950 23024 7930 23080
rect 7986 23024 25962 23080
rect 26018 23024 26023 23080
rect 4889 23022 26023 23024
rect 4889 23019 4955 23022
rect 7925 23019 7991 23022
rect 25957 23019 26023 23022
rect 4870 22880 5186 22881
rect 4870 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5186 22880
rect 4870 22815 5186 22816
rect 35590 22880 35906 22881
rect 35590 22816 35596 22880
rect 35660 22816 35676 22880
rect 35740 22816 35756 22880
rect 35820 22816 35836 22880
rect 35900 22816 35906 22880
rect 35590 22815 35906 22816
rect 2957 22674 3023 22677
rect 25589 22674 25655 22677
rect 2957 22672 25655 22674
rect 2957 22616 2962 22672
rect 3018 22616 25594 22672
rect 25650 22616 25655 22672
rect 2957 22614 25655 22616
rect 2957 22611 3023 22614
rect 25589 22611 25655 22614
rect 8201 22538 8267 22541
rect 24761 22538 24827 22541
rect 8201 22536 24827 22538
rect 8201 22480 8206 22536
rect 8262 22480 24766 22536
rect 24822 22480 24827 22536
rect 8201 22478 24827 22480
rect 8201 22475 8267 22478
rect 24761 22475 24827 22478
rect 37825 22538 37891 22541
rect 38618 22538 39418 22568
rect 37825 22536 39418 22538
rect 37825 22480 37830 22536
rect 37886 22480 39418 22536
rect 37825 22478 39418 22480
rect 37825 22475 37891 22478
rect 38618 22448 39418 22478
rect 25313 22402 25379 22405
rect 31109 22402 31175 22405
rect 25313 22400 31175 22402
rect 25313 22344 25318 22400
rect 25374 22344 31114 22400
rect 31170 22344 31175 22400
rect 25313 22342 31175 22344
rect 25313 22339 25379 22342
rect 31109 22339 31175 22342
rect 4210 22336 4526 22337
rect 4210 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4526 22336
rect 4210 22271 4526 22272
rect 34930 22336 35246 22337
rect 34930 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35246 22336
rect 34930 22271 35246 22272
rect 19241 22130 19307 22133
rect 22645 22130 22711 22133
rect 19241 22128 22711 22130
rect 19241 22072 19246 22128
rect 19302 22072 22650 22128
rect 22706 22072 22711 22128
rect 19241 22070 22711 22072
rect 19241 22067 19307 22070
rect 22645 22067 22711 22070
rect 31201 22130 31267 22133
rect 32857 22130 32923 22133
rect 31201 22128 32923 22130
rect 31201 22072 31206 22128
rect 31262 22072 32862 22128
rect 32918 22072 32923 22128
rect 31201 22070 32923 22072
rect 31201 22067 31267 22070
rect 32857 22067 32923 22070
rect 16021 21994 16087 21997
rect 16757 21994 16823 21997
rect 16021 21992 16823 21994
rect 16021 21936 16026 21992
rect 16082 21936 16762 21992
rect 16818 21936 16823 21992
rect 16021 21934 16823 21936
rect 16021 21931 16087 21934
rect 16757 21931 16823 21934
rect 22369 21994 22435 21997
rect 25129 21994 25195 21997
rect 22369 21992 25195 21994
rect 22369 21936 22374 21992
rect 22430 21936 25134 21992
rect 25190 21936 25195 21992
rect 22369 21934 25195 21936
rect 22369 21931 22435 21934
rect 25129 21931 25195 21934
rect 4870 21792 5186 21793
rect 4870 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5186 21792
rect 4870 21727 5186 21728
rect 35590 21792 35906 21793
rect 35590 21728 35596 21792
rect 35660 21728 35676 21792
rect 35740 21728 35756 21792
rect 35820 21728 35836 21792
rect 35900 21728 35906 21792
rect 35590 21727 35906 21728
rect 13905 21724 13971 21725
rect 13854 21722 13860 21724
rect 13814 21662 13860 21722
rect 13924 21720 13971 21724
rect 13966 21664 13971 21720
rect 13854 21660 13860 21662
rect 13924 21660 13971 21664
rect 13905 21659 13971 21660
rect 9673 21586 9739 21589
rect 10317 21588 10383 21589
rect 9806 21586 9812 21588
rect 9673 21584 9812 21586
rect 9673 21528 9678 21584
rect 9734 21528 9812 21584
rect 9673 21526 9812 21528
rect 9673 21523 9739 21526
rect 9806 21524 9812 21526
rect 9876 21524 9882 21588
rect 10317 21586 10364 21588
rect 10272 21584 10364 21586
rect 10272 21528 10322 21584
rect 10272 21526 10364 21528
rect 10317 21524 10364 21526
rect 10428 21524 10434 21588
rect 11881 21586 11947 21589
rect 15561 21586 15627 21589
rect 25773 21586 25839 21589
rect 11881 21584 15627 21586
rect 11881 21528 11886 21584
rect 11942 21528 15566 21584
rect 15622 21528 15627 21584
rect 11881 21526 15627 21528
rect 10317 21523 10383 21524
rect 11881 21523 11947 21526
rect 15561 21523 15627 21526
rect 19290 21584 25839 21586
rect 19290 21528 25778 21584
rect 25834 21528 25839 21584
rect 19290 21526 25839 21528
rect 13537 21450 13603 21453
rect 19290 21450 19350 21526
rect 25773 21523 25839 21526
rect 27705 21586 27771 21589
rect 36813 21586 36879 21589
rect 27705 21584 36879 21586
rect 27705 21528 27710 21584
rect 27766 21528 36818 21584
rect 36874 21528 36879 21584
rect 27705 21526 36879 21528
rect 27705 21523 27771 21526
rect 36813 21523 36879 21526
rect 13537 21448 19350 21450
rect 13537 21392 13542 21448
rect 13598 21392 19350 21448
rect 13537 21390 19350 21392
rect 19793 21450 19859 21453
rect 22185 21450 22251 21453
rect 22829 21452 22895 21453
rect 22829 21450 22876 21452
rect 19793 21448 22251 21450
rect 19793 21392 19798 21448
rect 19854 21392 22190 21448
rect 22246 21392 22251 21448
rect 19793 21390 22251 21392
rect 22784 21448 22876 21450
rect 22784 21392 22834 21448
rect 22784 21390 22876 21392
rect 13537 21387 13603 21390
rect 19793 21387 19859 21390
rect 22185 21387 22251 21390
rect 22829 21388 22876 21390
rect 22940 21388 22946 21452
rect 22829 21387 22895 21388
rect 10041 21314 10107 21317
rect 20161 21314 20227 21317
rect 10041 21312 20227 21314
rect 10041 21256 10046 21312
rect 10102 21256 20166 21312
rect 20222 21256 20227 21312
rect 10041 21254 20227 21256
rect 10041 21251 10107 21254
rect 20161 21251 20227 21254
rect 4210 21248 4526 21249
rect 4210 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4526 21248
rect 4210 21183 4526 21184
rect 34930 21248 35246 21249
rect 34930 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35246 21248
rect 34930 21183 35246 21184
rect 5717 21178 5783 21181
rect 24853 21178 24919 21181
rect 5717 21176 24919 21178
rect 5717 21120 5722 21176
rect 5778 21120 24858 21176
rect 24914 21120 24919 21176
rect 5717 21118 24919 21120
rect 5717 21115 5783 21118
rect 24853 21115 24919 21118
rect 14273 21042 14339 21045
rect 18229 21042 18295 21045
rect 14273 21040 18295 21042
rect 14273 20984 14278 21040
rect 14334 20984 18234 21040
rect 18290 20984 18295 21040
rect 14273 20982 18295 20984
rect 14273 20979 14339 20982
rect 18229 20979 18295 20982
rect 35065 21042 35131 21045
rect 35709 21042 35775 21045
rect 35065 21040 35775 21042
rect 35065 20984 35070 21040
rect 35126 20984 35714 21040
rect 35770 20984 35775 21040
rect 35065 20982 35775 20984
rect 35065 20979 35131 20982
rect 35709 20979 35775 20982
rect 5625 20906 5691 20909
rect 22369 20906 22435 20909
rect 5625 20904 22435 20906
rect 5625 20848 5630 20904
rect 5686 20848 22374 20904
rect 22430 20848 22435 20904
rect 5625 20846 22435 20848
rect 5625 20843 5691 20846
rect 22369 20843 22435 20846
rect 9581 20772 9647 20773
rect 9581 20768 9628 20772
rect 9692 20770 9698 20772
rect 9581 20712 9586 20768
rect 9581 20708 9628 20712
rect 9692 20710 9738 20770
rect 9814 20710 19350 20770
rect 9692 20708 9698 20710
rect 9581 20707 9647 20708
rect 4870 20704 5186 20705
rect 4870 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5186 20704
rect 4870 20639 5186 20640
rect 9814 20637 9874 20710
rect 1485 20634 1551 20637
rect 798 20632 1551 20634
rect 798 20576 1490 20632
rect 1546 20576 1551 20632
rect 798 20574 1551 20576
rect 798 20528 858 20574
rect 1485 20571 1551 20574
rect 9765 20632 9874 20637
rect 9765 20576 9770 20632
rect 9826 20576 9874 20632
rect 9765 20574 9874 20576
rect 12433 20634 12499 20637
rect 15285 20634 15351 20637
rect 12433 20632 15351 20634
rect 12433 20576 12438 20632
rect 12494 20576 15290 20632
rect 15346 20576 15351 20632
rect 12433 20574 15351 20576
rect 9765 20571 9831 20574
rect 12433 20571 12499 20574
rect 15285 20571 15351 20574
rect 15561 20634 15627 20637
rect 16573 20634 16639 20637
rect 15561 20632 16639 20634
rect 15561 20576 15566 20632
rect 15622 20576 16578 20632
rect 16634 20576 16639 20632
rect 15561 20574 16639 20576
rect 15561 20571 15627 20574
rect 16573 20571 16639 20574
rect 17033 20634 17099 20637
rect 18321 20634 18387 20637
rect 17033 20632 18387 20634
rect 17033 20576 17038 20632
rect 17094 20576 18326 20632
rect 18382 20576 18387 20632
rect 17033 20574 18387 20576
rect 19290 20634 19350 20710
rect 35590 20704 35906 20705
rect 35590 20640 35596 20704
rect 35660 20640 35676 20704
rect 35740 20640 35756 20704
rect 35820 20640 35836 20704
rect 35900 20640 35906 20704
rect 35590 20639 35906 20640
rect 23105 20634 23171 20637
rect 19290 20632 23171 20634
rect 19290 20576 23110 20632
rect 23166 20576 23171 20632
rect 19290 20574 23171 20576
rect 17033 20571 17099 20574
rect 18321 20571 18387 20574
rect 23105 20571 23171 20574
rect 25078 20572 25084 20636
rect 25148 20634 25154 20636
rect 25221 20634 25287 20637
rect 25148 20632 25287 20634
rect 25148 20576 25226 20632
rect 25282 20576 25287 20632
rect 25148 20574 25287 20576
rect 25148 20572 25154 20574
rect 25221 20571 25287 20574
rect 0 20438 858 20528
rect 14825 20498 14891 20501
rect 18045 20498 18111 20501
rect 14825 20496 18111 20498
rect 14825 20440 14830 20496
rect 14886 20440 18050 20496
rect 18106 20440 18111 20496
rect 14825 20438 18111 20440
rect 0 20408 800 20438
rect 14825 20435 14891 20438
rect 18045 20435 18111 20438
rect 38377 20498 38443 20501
rect 38618 20498 39418 20528
rect 38377 20496 39418 20498
rect 38377 20440 38382 20496
rect 38438 20440 39418 20496
rect 38377 20438 39418 20440
rect 38377 20435 38443 20438
rect 38618 20408 39418 20438
rect 10133 20362 10199 20365
rect 22001 20362 22067 20365
rect 10133 20360 22067 20362
rect 10133 20304 10138 20360
rect 10194 20304 22006 20360
rect 22062 20304 22067 20360
rect 10133 20302 22067 20304
rect 10133 20299 10199 20302
rect 22001 20299 22067 20302
rect 13629 20226 13695 20229
rect 23473 20226 23539 20229
rect 13629 20224 23539 20226
rect 13629 20168 13634 20224
rect 13690 20168 23478 20224
rect 23534 20168 23539 20224
rect 13629 20166 23539 20168
rect 13629 20163 13695 20166
rect 23473 20163 23539 20166
rect 24393 20226 24459 20229
rect 24945 20226 25011 20229
rect 24393 20224 25011 20226
rect 24393 20168 24398 20224
rect 24454 20168 24950 20224
rect 25006 20168 25011 20224
rect 24393 20166 25011 20168
rect 24393 20163 24459 20166
rect 24945 20163 25011 20166
rect 4210 20160 4526 20161
rect 4210 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4526 20160
rect 4210 20095 4526 20096
rect 34930 20160 35246 20161
rect 34930 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35246 20160
rect 34930 20095 35246 20096
rect 9121 20090 9187 20093
rect 22829 20090 22895 20093
rect 9121 20088 22895 20090
rect 9121 20032 9126 20088
rect 9182 20032 22834 20088
rect 22890 20032 22895 20088
rect 9121 20030 22895 20032
rect 9121 20027 9187 20030
rect 22829 20027 22895 20030
rect 23105 20090 23171 20093
rect 26877 20090 26943 20093
rect 23105 20088 26943 20090
rect 23105 20032 23110 20088
rect 23166 20032 26882 20088
rect 26938 20032 26943 20088
rect 23105 20030 26943 20032
rect 23105 20027 23171 20030
rect 26877 20027 26943 20030
rect 9489 19954 9555 19957
rect 22461 19954 22527 19957
rect 9489 19952 22527 19954
rect 9489 19896 9494 19952
rect 9550 19896 22466 19952
rect 22522 19896 22527 19952
rect 9489 19894 22527 19896
rect 9489 19891 9555 19894
rect 22461 19891 22527 19894
rect 23289 19954 23355 19957
rect 29913 19954 29979 19957
rect 23289 19952 29979 19954
rect 23289 19896 23294 19952
rect 23350 19896 29918 19952
rect 29974 19896 29979 19952
rect 23289 19894 29979 19896
rect 23289 19891 23355 19894
rect 29913 19891 29979 19894
rect 35341 19954 35407 19957
rect 36445 19954 36511 19957
rect 35341 19952 36511 19954
rect 35341 19896 35346 19952
rect 35402 19896 36450 19952
rect 36506 19896 36511 19952
rect 35341 19894 36511 19896
rect 35341 19891 35407 19894
rect 36445 19891 36511 19894
rect 4981 19818 5047 19821
rect 5349 19818 5415 19821
rect 6545 19818 6611 19821
rect 4981 19816 6611 19818
rect 4981 19760 4986 19816
rect 5042 19760 5354 19816
rect 5410 19760 6550 19816
rect 6606 19760 6611 19816
rect 4981 19758 6611 19760
rect 4981 19755 5047 19758
rect 5349 19755 5415 19758
rect 6545 19755 6611 19758
rect 7925 19818 7991 19821
rect 25313 19818 25379 19821
rect 7925 19816 25379 19818
rect 7925 19760 7930 19816
rect 7986 19760 25318 19816
rect 25374 19760 25379 19816
rect 7925 19758 25379 19760
rect 7925 19755 7991 19758
rect 25313 19755 25379 19758
rect 8385 19682 8451 19685
rect 26049 19682 26115 19685
rect 8385 19680 26115 19682
rect 8385 19624 8390 19680
rect 8446 19624 26054 19680
rect 26110 19624 26115 19680
rect 8385 19622 26115 19624
rect 8385 19619 8451 19622
rect 26049 19619 26115 19622
rect 4870 19616 5186 19617
rect 4870 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5186 19616
rect 4870 19551 5186 19552
rect 35590 19616 35906 19617
rect 35590 19552 35596 19616
rect 35660 19552 35676 19616
rect 35740 19552 35756 19616
rect 35820 19552 35836 19616
rect 35900 19552 35906 19616
rect 35590 19551 35906 19552
rect 12525 19546 12591 19549
rect 12893 19546 12959 19549
rect 13537 19546 13603 19549
rect 12525 19544 13603 19546
rect 12525 19488 12530 19544
rect 12586 19488 12898 19544
rect 12954 19488 13542 19544
rect 13598 19488 13603 19544
rect 12525 19486 13603 19488
rect 12525 19483 12591 19486
rect 12893 19483 12959 19486
rect 13537 19483 13603 19486
rect 14549 19546 14615 19549
rect 16021 19546 16087 19549
rect 14549 19544 16087 19546
rect 14549 19488 14554 19544
rect 14610 19488 16026 19544
rect 16082 19488 16087 19544
rect 14549 19486 16087 19488
rect 14549 19483 14615 19486
rect 16021 19483 16087 19486
rect 22461 19546 22527 19549
rect 27429 19546 27495 19549
rect 22461 19544 27495 19546
rect 22461 19488 22466 19544
rect 22522 19488 27434 19544
rect 27490 19488 27495 19544
rect 22461 19486 27495 19488
rect 22461 19483 22527 19486
rect 27429 19483 27495 19486
rect 9029 19410 9095 19413
rect 22369 19412 22435 19413
rect 22318 19410 22324 19412
rect 9029 19408 22324 19410
rect 22388 19410 22435 19412
rect 25773 19410 25839 19413
rect 22388 19408 25839 19410
rect 9029 19352 9034 19408
rect 9090 19352 22324 19408
rect 22430 19352 25778 19408
rect 25834 19352 25839 19408
rect 9029 19350 22324 19352
rect 9029 19347 9095 19350
rect 22318 19348 22324 19350
rect 22388 19350 25839 19352
rect 22388 19348 22435 19350
rect 22369 19347 22435 19348
rect 25773 19347 25839 19350
rect 28257 19410 28323 19413
rect 31109 19410 31175 19413
rect 28257 19408 31175 19410
rect 28257 19352 28262 19408
rect 28318 19352 31114 19408
rect 31170 19352 31175 19408
rect 28257 19350 31175 19352
rect 28257 19347 28323 19350
rect 31109 19347 31175 19350
rect 20110 19212 20116 19276
rect 20180 19274 20186 19276
rect 22369 19274 22435 19277
rect 20180 19272 22435 19274
rect 20180 19216 22374 19272
rect 22430 19216 22435 19272
rect 20180 19214 22435 19216
rect 20180 19212 20186 19214
rect 22369 19211 22435 19214
rect 4210 19072 4526 19073
rect 4210 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4526 19072
rect 4210 19007 4526 19008
rect 34930 19072 35246 19073
rect 34930 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35246 19072
rect 34930 19007 35246 19008
rect 11145 19002 11211 19005
rect 18505 19002 18571 19005
rect 11145 19000 18571 19002
rect 11145 18944 11150 19000
rect 11206 18944 18510 19000
rect 18566 18944 18571 19000
rect 11145 18942 18571 18944
rect 11145 18939 11211 18942
rect 18505 18939 18571 18942
rect 5993 18866 6059 18869
rect 23565 18866 23631 18869
rect 5993 18864 23631 18866
rect 5993 18808 5998 18864
rect 6054 18808 23570 18864
rect 23626 18808 23631 18864
rect 5993 18806 23631 18808
rect 5993 18803 6059 18806
rect 23565 18803 23631 18806
rect 18965 18730 19031 18733
rect 19793 18730 19859 18733
rect 18965 18728 19859 18730
rect 18965 18672 18970 18728
rect 19026 18672 19798 18728
rect 19854 18672 19859 18728
rect 18965 18670 19859 18672
rect 18965 18667 19031 18670
rect 19793 18667 19859 18670
rect 12157 18594 12223 18597
rect 24853 18594 24919 18597
rect 12157 18592 24919 18594
rect 12157 18536 12162 18592
rect 12218 18536 24858 18592
rect 24914 18536 24919 18592
rect 12157 18534 24919 18536
rect 12157 18531 12223 18534
rect 24853 18531 24919 18534
rect 4870 18528 5186 18529
rect 0 18458 800 18488
rect 4870 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5186 18528
rect 4870 18463 5186 18464
rect 35590 18528 35906 18529
rect 35590 18464 35596 18528
rect 35660 18464 35676 18528
rect 35740 18464 35756 18528
rect 35820 18464 35836 18528
rect 35900 18464 35906 18528
rect 35590 18463 35906 18464
rect 933 18458 999 18461
rect 0 18456 999 18458
rect 0 18400 938 18456
rect 994 18400 999 18456
rect 0 18398 999 18400
rect 0 18368 800 18398
rect 933 18395 999 18398
rect 10501 18458 10567 18461
rect 12709 18458 12775 18461
rect 15101 18458 15167 18461
rect 17125 18458 17191 18461
rect 20161 18458 20227 18461
rect 10501 18456 20227 18458
rect 10501 18400 10506 18456
rect 10562 18400 12714 18456
rect 12770 18400 15106 18456
rect 15162 18400 17130 18456
rect 17186 18400 20166 18456
rect 20222 18400 20227 18456
rect 10501 18398 20227 18400
rect 10501 18395 10567 18398
rect 12709 18395 12775 18398
rect 15101 18395 15167 18398
rect 17125 18395 17191 18398
rect 20161 18395 20227 18398
rect 29545 18322 29611 18325
rect 30373 18322 30439 18325
rect 33593 18322 33659 18325
rect 29545 18320 33659 18322
rect 29545 18264 29550 18320
rect 29606 18264 30378 18320
rect 30434 18264 33598 18320
rect 33654 18264 33659 18320
rect 29545 18262 33659 18264
rect 29545 18259 29611 18262
rect 30373 18259 30439 18262
rect 33593 18259 33659 18262
rect 18873 18186 18939 18189
rect 20069 18186 20135 18189
rect 18873 18184 20135 18186
rect 18873 18128 18878 18184
rect 18934 18128 20074 18184
rect 20130 18128 20135 18184
rect 18873 18126 20135 18128
rect 18873 18123 18939 18126
rect 20069 18123 20135 18126
rect 10869 18050 10935 18053
rect 10869 18048 17234 18050
rect 10869 17992 10874 18048
rect 10930 17992 17234 18048
rect 10869 17990 17234 17992
rect 10869 17987 10935 17990
rect 4210 17984 4526 17985
rect 4210 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4526 17984
rect 4210 17919 4526 17920
rect 8937 17914 9003 17917
rect 9806 17914 9812 17916
rect 8937 17912 9812 17914
rect 8937 17856 8942 17912
rect 8998 17856 9812 17912
rect 8937 17854 9812 17856
rect 8937 17851 9003 17854
rect 9806 17852 9812 17854
rect 9876 17852 9882 17916
rect 11697 17914 11763 17917
rect 11881 17914 11947 17917
rect 13353 17914 13419 17917
rect 11697 17912 13419 17914
rect 11697 17856 11702 17912
rect 11758 17856 11886 17912
rect 11942 17856 13358 17912
rect 13414 17856 13419 17912
rect 11697 17854 13419 17856
rect 11697 17851 11763 17854
rect 11881 17851 11947 17854
rect 13353 17851 13419 17854
rect 10869 17778 10935 17781
rect 12249 17778 12315 17781
rect 10869 17776 12315 17778
rect 10869 17720 10874 17776
rect 10930 17720 12254 17776
rect 12310 17720 12315 17776
rect 10869 17718 12315 17720
rect 17174 17778 17234 17990
rect 17534 17988 17540 18052
rect 17604 18050 17610 18052
rect 17604 17990 18522 18050
rect 17604 17988 17610 17990
rect 18229 17916 18295 17917
rect 18229 17912 18276 17916
rect 18340 17914 18346 17916
rect 18462 17914 18522 17990
rect 34930 17984 35246 17985
rect 34930 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35246 17984
rect 34930 17919 35246 17920
rect 18597 17914 18663 17917
rect 18229 17856 18234 17912
rect 18229 17852 18276 17856
rect 18340 17854 18386 17914
rect 18462 17912 18663 17914
rect 18462 17856 18602 17912
rect 18658 17856 18663 17912
rect 18462 17854 18663 17856
rect 18340 17852 18346 17854
rect 18229 17851 18295 17852
rect 18597 17851 18663 17854
rect 21950 17852 21956 17916
rect 22020 17914 22026 17916
rect 22737 17914 22803 17917
rect 22020 17912 22803 17914
rect 22020 17856 22742 17912
rect 22798 17856 22803 17912
rect 22020 17854 22803 17856
rect 22020 17852 22026 17854
rect 22737 17851 22803 17854
rect 23381 17914 23447 17917
rect 23606 17914 23612 17916
rect 23381 17912 23612 17914
rect 23381 17856 23386 17912
rect 23442 17856 23612 17912
rect 23381 17854 23612 17856
rect 23381 17851 23447 17854
rect 23606 17852 23612 17854
rect 23676 17852 23682 17916
rect 27705 17778 27771 17781
rect 17174 17776 27771 17778
rect 17174 17720 27710 17776
rect 27766 17720 27771 17776
rect 17174 17718 27771 17720
rect 10869 17715 10935 17718
rect 12249 17715 12315 17718
rect 27705 17715 27771 17718
rect 38377 17778 38443 17781
rect 38618 17778 39418 17808
rect 38377 17776 39418 17778
rect 38377 17720 38382 17776
rect 38438 17720 39418 17776
rect 38377 17718 39418 17720
rect 38377 17715 38443 17718
rect 38618 17688 39418 17718
rect 11697 17642 11763 17645
rect 12525 17642 12591 17645
rect 11697 17640 12591 17642
rect 11697 17584 11702 17640
rect 11758 17584 12530 17640
rect 12586 17584 12591 17640
rect 11697 17582 12591 17584
rect 11697 17579 11763 17582
rect 12525 17579 12591 17582
rect 23197 17642 23263 17645
rect 26182 17642 26188 17644
rect 23197 17640 26188 17642
rect 23197 17584 23202 17640
rect 23258 17584 26188 17640
rect 23197 17582 26188 17584
rect 23197 17579 23263 17582
rect 26182 17580 26188 17582
rect 26252 17580 26258 17644
rect 16205 17506 16271 17509
rect 16941 17506 17007 17509
rect 24669 17508 24735 17509
rect 24669 17506 24716 17508
rect 16205 17504 17007 17506
rect 16205 17448 16210 17504
rect 16266 17448 16946 17504
rect 17002 17448 17007 17504
rect 16205 17446 17007 17448
rect 24624 17504 24716 17506
rect 24624 17448 24674 17504
rect 24624 17446 24716 17448
rect 16205 17443 16271 17446
rect 16941 17443 17007 17446
rect 24669 17444 24716 17446
rect 24780 17444 24786 17508
rect 24669 17443 24735 17444
rect 4870 17440 5186 17441
rect 4870 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5186 17440
rect 4870 17375 5186 17376
rect 35590 17440 35906 17441
rect 35590 17376 35596 17440
rect 35660 17376 35676 17440
rect 35740 17376 35756 17440
rect 35820 17376 35836 17440
rect 35900 17376 35906 17440
rect 35590 17375 35906 17376
rect 4210 16896 4526 16897
rect 4210 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4526 16896
rect 4210 16831 4526 16832
rect 34930 16896 35246 16897
rect 34930 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35246 16896
rect 34930 16831 35246 16832
rect 4429 16690 4495 16693
rect 7925 16690 7991 16693
rect 4429 16688 7991 16690
rect 4429 16632 4434 16688
rect 4490 16632 7930 16688
rect 7986 16632 7991 16688
rect 4429 16630 7991 16632
rect 4429 16627 4495 16630
rect 7925 16627 7991 16630
rect 14365 16690 14431 16693
rect 16573 16690 16639 16693
rect 17953 16690 18019 16693
rect 14365 16688 18019 16690
rect 14365 16632 14370 16688
rect 14426 16632 16578 16688
rect 16634 16632 17958 16688
rect 18014 16632 18019 16688
rect 14365 16630 18019 16632
rect 14365 16627 14431 16630
rect 16573 16627 16639 16630
rect 17953 16627 18019 16630
rect 24485 16556 24551 16557
rect 24485 16554 24532 16556
rect 24440 16552 24532 16554
rect 24440 16496 24490 16552
rect 24440 16494 24532 16496
rect 24485 16492 24532 16494
rect 24596 16492 24602 16556
rect 24485 16491 24551 16492
rect 4870 16352 5186 16353
rect 4870 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5186 16352
rect 4870 16287 5186 16288
rect 35590 16352 35906 16353
rect 35590 16288 35596 16352
rect 35660 16288 35676 16352
rect 35740 16288 35756 16352
rect 35820 16288 35836 16352
rect 35900 16288 35906 16352
rect 35590 16287 35906 16288
rect 12341 16146 12407 16149
rect 24485 16146 24551 16149
rect 12341 16144 24551 16146
rect 12341 16088 12346 16144
rect 12402 16088 24490 16144
rect 24546 16088 24551 16144
rect 12341 16086 24551 16088
rect 12341 16083 12407 16086
rect 24485 16083 24551 16086
rect 12249 16010 12315 16013
rect 23749 16010 23815 16013
rect 12249 16008 23815 16010
rect 12249 15952 12254 16008
rect 12310 15952 23754 16008
rect 23810 15952 23815 16008
rect 12249 15950 23815 15952
rect 12249 15947 12315 15950
rect 23749 15947 23815 15950
rect 12525 15874 12591 15877
rect 18873 15874 18939 15877
rect 12525 15872 18939 15874
rect 12525 15816 12530 15872
rect 12586 15816 18878 15872
rect 18934 15816 18939 15872
rect 12525 15814 18939 15816
rect 12525 15811 12591 15814
rect 18873 15811 18939 15814
rect 4210 15808 4526 15809
rect 0 15738 800 15768
rect 4210 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4526 15808
rect 4210 15743 4526 15744
rect 34930 15808 35246 15809
rect 34930 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35246 15808
rect 34930 15743 35246 15744
rect 933 15738 999 15741
rect 0 15736 999 15738
rect 0 15680 938 15736
rect 994 15680 999 15736
rect 0 15678 999 15680
rect 0 15648 800 15678
rect 933 15675 999 15678
rect 37825 15738 37891 15741
rect 38618 15738 39418 15768
rect 37825 15736 39418 15738
rect 37825 15680 37830 15736
rect 37886 15680 39418 15736
rect 37825 15678 39418 15680
rect 37825 15675 37891 15678
rect 38618 15648 39418 15678
rect 11421 15466 11487 15469
rect 25129 15466 25195 15469
rect 11421 15464 25195 15466
rect 11421 15408 11426 15464
rect 11482 15408 25134 15464
rect 25190 15408 25195 15464
rect 11421 15406 25195 15408
rect 11421 15403 11487 15406
rect 25129 15403 25195 15406
rect 4870 15264 5186 15265
rect 4870 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5186 15264
rect 4870 15199 5186 15200
rect 35590 15264 35906 15265
rect 35590 15200 35596 15264
rect 35660 15200 35676 15264
rect 35740 15200 35756 15264
rect 35820 15200 35836 15264
rect 35900 15200 35906 15264
rect 35590 15199 35906 15200
rect 25589 14922 25655 14925
rect 28717 14922 28783 14925
rect 25589 14920 28783 14922
rect 25589 14864 25594 14920
rect 25650 14864 28722 14920
rect 28778 14864 28783 14920
rect 25589 14862 28783 14864
rect 25589 14859 25655 14862
rect 28717 14859 28783 14862
rect 4210 14720 4526 14721
rect 4210 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4526 14720
rect 4210 14655 4526 14656
rect 34930 14720 35246 14721
rect 34930 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35246 14720
rect 34930 14655 35246 14656
rect 9581 14378 9647 14381
rect 30281 14378 30347 14381
rect 9581 14376 30347 14378
rect 9581 14320 9586 14376
rect 9642 14320 30286 14376
rect 30342 14320 30347 14376
rect 9581 14318 30347 14320
rect 9581 14315 9647 14318
rect 30281 14315 30347 14318
rect 4870 14176 5186 14177
rect 4870 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5186 14176
rect 4870 14111 5186 14112
rect 35590 14176 35906 14177
rect 35590 14112 35596 14176
rect 35660 14112 35676 14176
rect 35740 14112 35756 14176
rect 35820 14112 35836 14176
rect 35900 14112 35906 14176
rect 35590 14111 35906 14112
rect 24393 13970 24459 13973
rect 26049 13970 26115 13973
rect 24393 13968 26115 13970
rect 24393 13912 24398 13968
rect 24454 13912 26054 13968
rect 26110 13912 26115 13968
rect 24393 13910 26115 13912
rect 24393 13907 24459 13910
rect 26049 13907 26115 13910
rect 0 13698 800 13728
rect 1485 13698 1551 13701
rect 9581 13700 9647 13701
rect 9581 13698 9628 13700
rect 0 13696 1551 13698
rect 0 13640 1490 13696
rect 1546 13640 1551 13696
rect 0 13638 1551 13640
rect 9536 13696 9628 13698
rect 9536 13640 9586 13696
rect 9536 13638 9628 13640
rect 0 13608 800 13638
rect 1485 13635 1551 13638
rect 9581 13636 9628 13638
rect 9692 13636 9698 13700
rect 9581 13635 9647 13636
rect 4210 13632 4526 13633
rect 4210 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4526 13632
rect 4210 13567 4526 13568
rect 34930 13632 35246 13633
rect 34930 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35246 13632
rect 38618 13608 39418 13728
rect 34930 13567 35246 13568
rect 24393 13426 24459 13429
rect 26233 13426 26299 13429
rect 26417 13426 26483 13429
rect 24393 13424 26664 13426
rect 24393 13368 24398 13424
rect 24454 13368 26238 13424
rect 26294 13368 26422 13424
rect 26478 13368 26664 13424
rect 24393 13366 26664 13368
rect 24393 13363 24459 13366
rect 26233 13363 26299 13366
rect 26417 13363 26483 13366
rect 26604 13290 26664 13366
rect 26734 13364 26740 13428
rect 26804 13426 26810 13428
rect 27613 13426 27679 13429
rect 26804 13424 27679 13426
rect 26804 13368 27618 13424
rect 27674 13368 27679 13424
rect 26804 13366 27679 13368
rect 26804 13364 26810 13366
rect 27613 13363 27679 13366
rect 27153 13290 27219 13293
rect 26604 13288 27219 13290
rect 26604 13232 27158 13288
rect 27214 13232 27219 13288
rect 26604 13230 27219 13232
rect 27153 13227 27219 13230
rect 4870 13088 5186 13089
rect 4870 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5186 13088
rect 4870 13023 5186 13024
rect 35590 13088 35906 13089
rect 35590 13024 35596 13088
rect 35660 13024 35676 13088
rect 35740 13024 35756 13088
rect 35820 13024 35836 13088
rect 35900 13024 35906 13088
rect 35590 13023 35906 13024
rect 10225 13018 10291 13021
rect 18689 13018 18755 13021
rect 10225 13016 18755 13018
rect 10225 12960 10230 13016
rect 10286 12960 18694 13016
rect 18750 12960 18755 13016
rect 10225 12958 18755 12960
rect 10225 12955 10291 12958
rect 18689 12955 18755 12958
rect 26141 12882 26207 12885
rect 26601 12882 26667 12885
rect 26141 12880 26667 12882
rect 26141 12824 26146 12880
rect 26202 12824 26606 12880
rect 26662 12824 26667 12880
rect 26141 12822 26667 12824
rect 26141 12819 26207 12822
rect 26601 12819 26667 12822
rect 4210 12544 4526 12545
rect 4210 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4526 12544
rect 4210 12479 4526 12480
rect 34930 12544 35246 12545
rect 34930 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35246 12544
rect 34930 12479 35246 12480
rect 24117 12066 24183 12069
rect 28901 12066 28967 12069
rect 24117 12064 28967 12066
rect 24117 12008 24122 12064
rect 24178 12008 28906 12064
rect 28962 12008 28967 12064
rect 24117 12006 28967 12008
rect 24117 12003 24183 12006
rect 28901 12003 28967 12006
rect 4870 12000 5186 12001
rect 4870 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5186 12000
rect 4870 11935 5186 11936
rect 35590 12000 35906 12001
rect 35590 11936 35596 12000
rect 35660 11936 35676 12000
rect 35740 11936 35756 12000
rect 35820 11936 35836 12000
rect 35900 11936 35906 12000
rect 35590 11935 35906 11936
rect 0 11658 800 11688
rect 933 11658 999 11661
rect 0 11656 999 11658
rect 0 11600 938 11656
rect 994 11600 999 11656
rect 0 11598 999 11600
rect 0 11568 800 11598
rect 933 11595 999 11598
rect 18689 11658 18755 11661
rect 27705 11658 27771 11661
rect 18689 11656 27771 11658
rect 18689 11600 18694 11656
rect 18750 11600 27710 11656
rect 27766 11600 27771 11656
rect 18689 11598 27771 11600
rect 18689 11595 18755 11598
rect 27705 11595 27771 11598
rect 4210 11456 4526 11457
rect 4210 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4526 11456
rect 4210 11391 4526 11392
rect 34930 11456 35246 11457
rect 34930 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35246 11456
rect 34930 11391 35246 11392
rect 16430 10916 16436 10980
rect 16500 10978 16506 10980
rect 18229 10978 18295 10981
rect 16500 10976 18295 10978
rect 16500 10920 18234 10976
rect 18290 10920 18295 10976
rect 16500 10918 18295 10920
rect 16500 10916 16506 10918
rect 18229 10915 18295 10918
rect 20805 10978 20871 10981
rect 22093 10978 22159 10981
rect 22645 10978 22711 10981
rect 20805 10976 22711 10978
rect 20805 10920 20810 10976
rect 20866 10920 22098 10976
rect 22154 10920 22650 10976
rect 22706 10920 22711 10976
rect 20805 10918 22711 10920
rect 20805 10915 20871 10918
rect 22093 10915 22159 10918
rect 22645 10915 22711 10918
rect 30005 10978 30071 10981
rect 31293 10978 31359 10981
rect 30005 10976 31359 10978
rect 30005 10920 30010 10976
rect 30066 10920 31298 10976
rect 31354 10920 31359 10976
rect 30005 10918 31359 10920
rect 30005 10915 30071 10918
rect 31293 10915 31359 10918
rect 37917 10978 37983 10981
rect 38618 10978 39418 11008
rect 37917 10976 39418 10978
rect 37917 10920 37922 10976
rect 37978 10920 39418 10976
rect 37917 10918 39418 10920
rect 37917 10915 37983 10918
rect 4870 10912 5186 10913
rect 4870 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5186 10912
rect 4870 10847 5186 10848
rect 35590 10912 35906 10913
rect 35590 10848 35596 10912
rect 35660 10848 35676 10912
rect 35740 10848 35756 10912
rect 35820 10848 35836 10912
rect 35900 10848 35906 10912
rect 38618 10888 39418 10918
rect 35590 10847 35906 10848
rect 22001 10706 22067 10709
rect 23013 10706 23079 10709
rect 22001 10704 23079 10706
rect 22001 10648 22006 10704
rect 22062 10648 23018 10704
rect 23074 10648 23079 10704
rect 22001 10646 23079 10648
rect 22001 10643 22067 10646
rect 23013 10643 23079 10646
rect 17493 10570 17559 10573
rect 27981 10570 28047 10573
rect 17493 10568 28047 10570
rect 17493 10512 17498 10568
rect 17554 10512 27986 10568
rect 28042 10512 28047 10568
rect 17493 10510 28047 10512
rect 17493 10507 17559 10510
rect 27981 10507 28047 10510
rect 22185 10434 22251 10437
rect 28349 10434 28415 10437
rect 22185 10432 28415 10434
rect 22185 10376 22190 10432
rect 22246 10376 28354 10432
rect 28410 10376 28415 10432
rect 22185 10374 28415 10376
rect 22185 10371 22251 10374
rect 28349 10371 28415 10374
rect 4210 10368 4526 10369
rect 4210 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4526 10368
rect 4210 10303 4526 10304
rect 34930 10368 35246 10369
rect 34930 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35246 10368
rect 34930 10303 35246 10304
rect 20621 10026 20687 10029
rect 21909 10026 21975 10029
rect 20621 10024 21975 10026
rect 20621 9968 20626 10024
rect 20682 9968 21914 10024
rect 21970 9968 21975 10024
rect 20621 9966 21975 9968
rect 20621 9963 20687 9966
rect 21909 9963 21975 9966
rect 4870 9824 5186 9825
rect 4870 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5186 9824
rect 4870 9759 5186 9760
rect 35590 9824 35906 9825
rect 35590 9760 35596 9824
rect 35660 9760 35676 9824
rect 35740 9760 35756 9824
rect 35820 9760 35836 9824
rect 35900 9760 35906 9824
rect 35590 9759 35906 9760
rect 3233 9618 3299 9621
rect 22277 9620 22343 9621
rect 22277 9618 22324 9620
rect 3233 9616 22110 9618
rect 3233 9560 3238 9616
rect 3294 9560 22110 9616
rect 3233 9558 22110 9560
rect 22232 9616 22324 9618
rect 22232 9560 22282 9616
rect 22232 9558 22324 9560
rect 3233 9555 3299 9558
rect 6637 9482 6703 9485
rect 9305 9482 9371 9485
rect 6637 9480 9371 9482
rect 6637 9424 6642 9480
rect 6698 9424 9310 9480
rect 9366 9424 9371 9480
rect 6637 9422 9371 9424
rect 6637 9419 6703 9422
rect 9305 9419 9371 9422
rect 15377 9482 15443 9485
rect 15510 9482 15516 9484
rect 15377 9480 15516 9482
rect 15377 9424 15382 9480
rect 15438 9424 15516 9480
rect 15377 9422 15516 9424
rect 15377 9419 15443 9422
rect 15510 9420 15516 9422
rect 15580 9420 15586 9484
rect 18873 9482 18939 9485
rect 20662 9482 20668 9484
rect 18873 9480 20668 9482
rect 18873 9424 18878 9480
rect 18934 9424 20668 9480
rect 18873 9422 20668 9424
rect 18873 9419 18939 9422
rect 20662 9420 20668 9422
rect 20732 9420 20738 9484
rect 22050 9482 22110 9558
rect 22277 9556 22324 9558
rect 22388 9556 22394 9620
rect 29913 9618 29979 9621
rect 22510 9616 29979 9618
rect 22510 9560 29918 9616
rect 29974 9560 29979 9616
rect 22510 9558 29979 9560
rect 22277 9555 22343 9556
rect 22510 9482 22570 9558
rect 29913 9555 29979 9558
rect 22050 9422 22570 9482
rect 4210 9280 4526 9281
rect 4210 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4526 9280
rect 4210 9215 4526 9216
rect 34930 9280 35246 9281
rect 34930 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35246 9280
rect 34930 9215 35246 9216
rect 9949 9210 10015 9213
rect 13813 9210 13879 9213
rect 17033 9210 17099 9213
rect 9949 9208 17099 9210
rect 9949 9152 9954 9208
rect 10010 9152 13818 9208
rect 13874 9152 17038 9208
rect 17094 9152 17099 9208
rect 9949 9150 17099 9152
rect 9949 9147 10015 9150
rect 13813 9147 13879 9150
rect 17033 9147 17099 9150
rect 22737 9210 22803 9213
rect 22737 9208 24962 9210
rect 22737 9152 22742 9208
rect 22798 9152 24962 9208
rect 22737 9150 24962 9152
rect 22737 9147 22803 9150
rect 4153 9074 4219 9077
rect 22645 9074 22711 9077
rect 24710 9074 24716 9076
rect 4153 9072 24716 9074
rect 4153 9016 4158 9072
rect 4214 9016 22650 9072
rect 22706 9016 24716 9072
rect 4153 9014 24716 9016
rect 4153 9011 4219 9014
rect 22645 9011 22711 9014
rect 24710 9012 24716 9014
rect 24780 9012 24786 9076
rect 24902 9074 24962 9150
rect 25313 9074 25379 9077
rect 26049 9074 26115 9077
rect 27613 9074 27679 9077
rect 24902 9072 27679 9074
rect 24902 9016 25318 9072
rect 25374 9016 26054 9072
rect 26110 9016 27618 9072
rect 27674 9016 27679 9072
rect 24902 9014 27679 9016
rect 25313 9011 25379 9014
rect 26049 9011 26115 9014
rect 27613 9011 27679 9014
rect 29821 9074 29887 9077
rect 30649 9074 30715 9077
rect 29821 9072 30715 9074
rect 29821 9016 29826 9072
rect 29882 9016 30654 9072
rect 30710 9016 30715 9072
rect 29821 9014 30715 9016
rect 29821 9011 29887 9014
rect 30649 9011 30715 9014
rect 0 8938 800 8968
rect 933 8938 999 8941
rect 0 8936 999 8938
rect 0 8880 938 8936
rect 994 8880 999 8936
rect 0 8878 999 8880
rect 0 8848 800 8878
rect 933 8875 999 8878
rect 38285 8938 38351 8941
rect 38618 8938 39418 8968
rect 38285 8936 39418 8938
rect 38285 8880 38290 8936
rect 38346 8880 39418 8936
rect 38285 8878 39418 8880
rect 38285 8875 38351 8878
rect 38618 8848 39418 8878
rect 4870 8736 5186 8737
rect 4870 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5186 8736
rect 4870 8671 5186 8672
rect 35590 8736 35906 8737
rect 35590 8672 35596 8736
rect 35660 8672 35676 8736
rect 35740 8672 35756 8736
rect 35820 8672 35836 8736
rect 35900 8672 35906 8736
rect 35590 8671 35906 8672
rect 18965 8532 19031 8533
rect 18965 8530 19012 8532
rect 18920 8528 19012 8530
rect 18920 8472 18970 8528
rect 18920 8470 19012 8472
rect 18965 8468 19012 8470
rect 19076 8468 19082 8532
rect 18965 8467 19031 8468
rect 21817 8394 21883 8397
rect 23473 8394 23539 8397
rect 25405 8394 25471 8397
rect 21817 8392 25471 8394
rect 21817 8336 21822 8392
rect 21878 8336 23478 8392
rect 23534 8336 25410 8392
rect 25466 8336 25471 8392
rect 21817 8334 25471 8336
rect 21817 8331 21883 8334
rect 23473 8331 23539 8334
rect 25405 8331 25471 8334
rect 4210 8192 4526 8193
rect 4210 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4526 8192
rect 4210 8127 4526 8128
rect 34930 8192 35246 8193
rect 34930 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35246 8192
rect 34930 8127 35246 8128
rect 4870 7648 5186 7649
rect 4870 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5186 7648
rect 4870 7583 5186 7584
rect 35590 7648 35906 7649
rect 35590 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35906 7648
rect 35590 7583 35906 7584
rect 4210 7104 4526 7105
rect 4210 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4526 7104
rect 4210 7039 4526 7040
rect 34930 7104 35246 7105
rect 34930 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35246 7104
rect 34930 7039 35246 7040
rect 0 6898 800 6928
rect 1485 6898 1551 6901
rect 0 6896 1551 6898
rect 0 6840 1490 6896
rect 1546 6840 1551 6896
rect 0 6838 1551 6840
rect 0 6808 800 6838
rect 1485 6835 1551 6838
rect 18229 6898 18295 6901
rect 18454 6898 18460 6900
rect 18229 6896 18460 6898
rect 18229 6840 18234 6896
rect 18290 6840 18460 6896
rect 18229 6838 18460 6840
rect 18229 6835 18295 6838
rect 18454 6836 18460 6838
rect 18524 6836 18530 6900
rect 4870 6560 5186 6561
rect 4870 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5186 6560
rect 4870 6495 5186 6496
rect 35590 6560 35906 6561
rect 35590 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35906 6560
rect 35590 6495 35906 6496
rect 38618 6128 39418 6248
rect 4210 6016 4526 6017
rect 4210 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4526 6016
rect 4210 5951 4526 5952
rect 34930 6016 35246 6017
rect 34930 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35246 6016
rect 34930 5951 35246 5952
rect 4870 5472 5186 5473
rect 4870 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5186 5472
rect 4870 5407 5186 5408
rect 35590 5472 35906 5473
rect 35590 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35906 5472
rect 35590 5407 35906 5408
rect 4210 4928 4526 4929
rect 4210 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4526 4928
rect 4210 4863 4526 4864
rect 34930 4928 35246 4929
rect 34930 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35246 4928
rect 34930 4863 35246 4864
rect 4870 4384 5186 4385
rect 4870 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5186 4384
rect 4870 4319 5186 4320
rect 35590 4384 35906 4385
rect 35590 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35906 4384
rect 35590 4319 35906 4320
rect 0 4178 800 4208
rect 933 4178 999 4181
rect 0 4176 999 4178
rect 0 4120 938 4176
rect 994 4120 999 4176
rect 0 4118 999 4120
rect 0 4088 800 4118
rect 933 4115 999 4118
rect 38618 4088 39418 4208
rect 12525 4044 12591 4045
rect 12525 4040 12572 4044
rect 12636 4042 12642 4044
rect 13169 4042 13235 4045
rect 13302 4042 13308 4044
rect 12525 3984 12530 4040
rect 12525 3980 12572 3984
rect 12636 3982 12682 4042
rect 13169 4040 13308 4042
rect 13169 3984 13174 4040
rect 13230 3984 13308 4040
rect 13169 3982 13308 3984
rect 12636 3980 12642 3982
rect 12525 3979 12591 3980
rect 13169 3979 13235 3982
rect 13302 3980 13308 3982
rect 13372 3980 13378 4044
rect 4210 3840 4526 3841
rect 4210 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4526 3840
rect 4210 3775 4526 3776
rect 34930 3840 35246 3841
rect 34930 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35246 3840
rect 34930 3775 35246 3776
rect 4870 3296 5186 3297
rect 4870 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5186 3296
rect 4870 3231 5186 3232
rect 35590 3296 35906 3297
rect 35590 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35906 3296
rect 35590 3231 35906 3232
rect 4210 2752 4526 2753
rect 4210 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4526 2752
rect 4210 2687 4526 2688
rect 34930 2752 35246 2753
rect 34930 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35246 2752
rect 34930 2687 35246 2688
rect 4870 2208 5186 2209
rect 0 2048 800 2168
rect 4870 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5186 2208
rect 4870 2143 5186 2144
rect 35590 2208 35906 2209
rect 35590 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35906 2208
rect 35590 2143 35906 2144
rect 37181 1458 37247 1461
rect 38618 1458 39418 1488
rect 37181 1456 39418 1458
rect 37181 1400 37186 1456
rect 37242 1400 39418 1456
rect 37181 1398 39418 1400
rect 37181 1395 37247 1398
rect 38618 1368 39418 1398
<< via3 >>
rect 4876 39196 4940 39200
rect 4876 39140 4880 39196
rect 4880 39140 4936 39196
rect 4936 39140 4940 39196
rect 4876 39136 4940 39140
rect 4956 39196 5020 39200
rect 4956 39140 4960 39196
rect 4960 39140 5016 39196
rect 5016 39140 5020 39196
rect 4956 39136 5020 39140
rect 5036 39196 5100 39200
rect 5036 39140 5040 39196
rect 5040 39140 5096 39196
rect 5096 39140 5100 39196
rect 5036 39136 5100 39140
rect 5116 39196 5180 39200
rect 5116 39140 5120 39196
rect 5120 39140 5176 39196
rect 5176 39140 5180 39196
rect 5116 39136 5180 39140
rect 35596 39196 35660 39200
rect 35596 39140 35600 39196
rect 35600 39140 35656 39196
rect 35656 39140 35660 39196
rect 35596 39136 35660 39140
rect 35676 39196 35740 39200
rect 35676 39140 35680 39196
rect 35680 39140 35736 39196
rect 35736 39140 35740 39196
rect 35676 39136 35740 39140
rect 35756 39196 35820 39200
rect 35756 39140 35760 39196
rect 35760 39140 35816 39196
rect 35816 39140 35820 39196
rect 35756 39136 35820 39140
rect 35836 39196 35900 39200
rect 35836 39140 35840 39196
rect 35840 39140 35896 39196
rect 35896 39140 35900 39196
rect 35836 39136 35900 39140
rect 9812 38796 9876 38860
rect 10364 38660 10428 38724
rect 22876 38660 22940 38724
rect 23980 38660 24044 38724
rect 4216 38652 4280 38656
rect 4216 38596 4220 38652
rect 4220 38596 4276 38652
rect 4276 38596 4280 38652
rect 4216 38592 4280 38596
rect 4296 38652 4360 38656
rect 4296 38596 4300 38652
rect 4300 38596 4356 38652
rect 4356 38596 4360 38652
rect 4296 38592 4360 38596
rect 4376 38652 4440 38656
rect 4376 38596 4380 38652
rect 4380 38596 4436 38652
rect 4436 38596 4440 38652
rect 4376 38592 4440 38596
rect 4456 38652 4520 38656
rect 4456 38596 4460 38652
rect 4460 38596 4516 38652
rect 4516 38596 4520 38652
rect 4456 38592 4520 38596
rect 34936 38652 35000 38656
rect 34936 38596 34940 38652
rect 34940 38596 34996 38652
rect 34996 38596 35000 38652
rect 34936 38592 35000 38596
rect 35016 38652 35080 38656
rect 35016 38596 35020 38652
rect 35020 38596 35076 38652
rect 35076 38596 35080 38652
rect 35016 38592 35080 38596
rect 35096 38652 35160 38656
rect 35096 38596 35100 38652
rect 35100 38596 35156 38652
rect 35156 38596 35160 38652
rect 35096 38592 35160 38596
rect 35176 38652 35240 38656
rect 35176 38596 35180 38652
rect 35180 38596 35236 38652
rect 35236 38596 35240 38652
rect 35176 38592 35240 38596
rect 4876 38108 4940 38112
rect 4876 38052 4880 38108
rect 4880 38052 4936 38108
rect 4936 38052 4940 38108
rect 4876 38048 4940 38052
rect 4956 38108 5020 38112
rect 4956 38052 4960 38108
rect 4960 38052 5016 38108
rect 5016 38052 5020 38108
rect 4956 38048 5020 38052
rect 5036 38108 5100 38112
rect 5036 38052 5040 38108
rect 5040 38052 5096 38108
rect 5096 38052 5100 38108
rect 5036 38048 5100 38052
rect 5116 38108 5180 38112
rect 5116 38052 5120 38108
rect 5120 38052 5176 38108
rect 5176 38052 5180 38108
rect 5116 38048 5180 38052
rect 35596 38108 35660 38112
rect 35596 38052 35600 38108
rect 35600 38052 35656 38108
rect 35656 38052 35660 38108
rect 35596 38048 35660 38052
rect 35676 38108 35740 38112
rect 35676 38052 35680 38108
rect 35680 38052 35736 38108
rect 35736 38052 35740 38108
rect 35676 38048 35740 38052
rect 35756 38108 35820 38112
rect 35756 38052 35760 38108
rect 35760 38052 35816 38108
rect 35816 38052 35820 38108
rect 35756 38048 35820 38052
rect 35836 38108 35900 38112
rect 35836 38052 35840 38108
rect 35840 38052 35896 38108
rect 35896 38052 35900 38108
rect 35836 38048 35900 38052
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 22140 37300 22204 37364
rect 25268 37360 25332 37364
rect 25268 37304 25282 37360
rect 25282 37304 25332 37360
rect 25268 37300 25332 37304
rect 27844 37300 27908 37364
rect 4876 37020 4940 37024
rect 4876 36964 4880 37020
rect 4880 36964 4936 37020
rect 4936 36964 4940 37020
rect 4876 36960 4940 36964
rect 4956 37020 5020 37024
rect 4956 36964 4960 37020
rect 4960 36964 5016 37020
rect 5016 36964 5020 37020
rect 4956 36960 5020 36964
rect 5036 37020 5100 37024
rect 5036 36964 5040 37020
rect 5040 36964 5096 37020
rect 5096 36964 5100 37020
rect 5036 36960 5100 36964
rect 5116 37020 5180 37024
rect 5116 36964 5120 37020
rect 5120 36964 5176 37020
rect 5176 36964 5180 37020
rect 5116 36960 5180 36964
rect 35596 37020 35660 37024
rect 35596 36964 35600 37020
rect 35600 36964 35656 37020
rect 35656 36964 35660 37020
rect 35596 36960 35660 36964
rect 35676 37020 35740 37024
rect 35676 36964 35680 37020
rect 35680 36964 35736 37020
rect 35736 36964 35740 37020
rect 35676 36960 35740 36964
rect 35756 37020 35820 37024
rect 35756 36964 35760 37020
rect 35760 36964 35816 37020
rect 35816 36964 35820 37020
rect 35756 36960 35820 36964
rect 35836 37020 35900 37024
rect 35836 36964 35840 37020
rect 35840 36964 35896 37020
rect 35896 36964 35900 37020
rect 35836 36960 35900 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 17540 35940 17604 36004
rect 20300 35940 20364 36004
rect 24900 36000 24964 36004
rect 24900 35944 24950 36000
rect 24950 35944 24964 36000
rect 24900 35940 24964 35944
rect 28948 35940 29012 36004
rect 4876 35932 4940 35936
rect 4876 35876 4880 35932
rect 4880 35876 4936 35932
rect 4936 35876 4940 35932
rect 4876 35872 4940 35876
rect 4956 35932 5020 35936
rect 4956 35876 4960 35932
rect 4960 35876 5016 35932
rect 5016 35876 5020 35932
rect 4956 35872 5020 35876
rect 5036 35932 5100 35936
rect 5036 35876 5040 35932
rect 5040 35876 5096 35932
rect 5096 35876 5100 35932
rect 5036 35872 5100 35876
rect 5116 35932 5180 35936
rect 5116 35876 5120 35932
rect 5120 35876 5176 35932
rect 5176 35876 5180 35932
rect 5116 35872 5180 35876
rect 35596 35932 35660 35936
rect 35596 35876 35600 35932
rect 35600 35876 35656 35932
rect 35656 35876 35660 35932
rect 35596 35872 35660 35876
rect 35676 35932 35740 35936
rect 35676 35876 35680 35932
rect 35680 35876 35736 35932
rect 35736 35876 35740 35932
rect 35676 35872 35740 35876
rect 35756 35932 35820 35936
rect 35756 35876 35760 35932
rect 35760 35876 35816 35932
rect 35816 35876 35820 35932
rect 35756 35872 35820 35876
rect 35836 35932 35900 35936
rect 35836 35876 35840 35932
rect 35840 35876 35896 35932
rect 35896 35876 35900 35932
rect 35836 35872 35900 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 4876 34844 4940 34848
rect 4876 34788 4880 34844
rect 4880 34788 4936 34844
rect 4936 34788 4940 34844
rect 4876 34784 4940 34788
rect 4956 34844 5020 34848
rect 4956 34788 4960 34844
rect 4960 34788 5016 34844
rect 5016 34788 5020 34844
rect 4956 34784 5020 34788
rect 5036 34844 5100 34848
rect 5036 34788 5040 34844
rect 5040 34788 5096 34844
rect 5096 34788 5100 34844
rect 5036 34784 5100 34788
rect 5116 34844 5180 34848
rect 5116 34788 5120 34844
rect 5120 34788 5176 34844
rect 5176 34788 5180 34844
rect 5116 34784 5180 34788
rect 13860 34580 13924 34644
rect 35596 34844 35660 34848
rect 35596 34788 35600 34844
rect 35600 34788 35656 34844
rect 35656 34788 35660 34844
rect 35596 34784 35660 34788
rect 35676 34844 35740 34848
rect 35676 34788 35680 34844
rect 35680 34788 35736 34844
rect 35736 34788 35740 34844
rect 35676 34784 35740 34788
rect 35756 34844 35820 34848
rect 35756 34788 35760 34844
rect 35760 34788 35816 34844
rect 35816 34788 35820 34844
rect 35756 34784 35820 34788
rect 35836 34844 35900 34848
rect 35836 34788 35840 34844
rect 35840 34788 35896 34844
rect 35896 34788 35900 34844
rect 35836 34784 35900 34788
rect 23428 34640 23492 34644
rect 23428 34584 23478 34640
rect 23478 34584 23492 34640
rect 23428 34580 23492 34584
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 4876 33756 4940 33760
rect 4876 33700 4880 33756
rect 4880 33700 4936 33756
rect 4936 33700 4940 33756
rect 4876 33696 4940 33700
rect 4956 33756 5020 33760
rect 4956 33700 4960 33756
rect 4960 33700 5016 33756
rect 5016 33700 5020 33756
rect 4956 33696 5020 33700
rect 5036 33756 5100 33760
rect 5036 33700 5040 33756
rect 5040 33700 5096 33756
rect 5096 33700 5100 33756
rect 5036 33696 5100 33700
rect 5116 33756 5180 33760
rect 5116 33700 5120 33756
rect 5120 33700 5176 33756
rect 5176 33700 5180 33756
rect 5116 33696 5180 33700
rect 35596 33756 35660 33760
rect 35596 33700 35600 33756
rect 35600 33700 35656 33756
rect 35656 33700 35660 33756
rect 35596 33696 35660 33700
rect 35676 33756 35740 33760
rect 35676 33700 35680 33756
rect 35680 33700 35736 33756
rect 35736 33700 35740 33756
rect 35676 33696 35740 33700
rect 35756 33756 35820 33760
rect 35756 33700 35760 33756
rect 35760 33700 35816 33756
rect 35816 33700 35820 33756
rect 35756 33696 35820 33700
rect 35836 33756 35900 33760
rect 35836 33700 35840 33756
rect 35840 33700 35896 33756
rect 35896 33700 35900 33756
rect 35836 33696 35900 33700
rect 23244 33628 23308 33692
rect 26188 33356 26252 33420
rect 19012 33280 19076 33284
rect 19012 33224 19062 33280
rect 19062 33224 19076 33280
rect 19012 33220 19076 33224
rect 24532 33220 24596 33284
rect 25084 33220 25148 33284
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19380 33084 19444 33148
rect 28948 33084 29012 33148
rect 4876 32668 4940 32672
rect 4876 32612 4880 32668
rect 4880 32612 4936 32668
rect 4936 32612 4940 32668
rect 4876 32608 4940 32612
rect 4956 32668 5020 32672
rect 4956 32612 4960 32668
rect 4960 32612 5016 32668
rect 5016 32612 5020 32668
rect 4956 32608 5020 32612
rect 5036 32668 5100 32672
rect 5036 32612 5040 32668
rect 5040 32612 5096 32668
rect 5096 32612 5100 32668
rect 5036 32608 5100 32612
rect 5116 32668 5180 32672
rect 5116 32612 5120 32668
rect 5120 32612 5176 32668
rect 5176 32612 5180 32668
rect 5116 32608 5180 32612
rect 35596 32668 35660 32672
rect 35596 32612 35600 32668
rect 35600 32612 35656 32668
rect 35656 32612 35660 32668
rect 35596 32608 35660 32612
rect 35676 32668 35740 32672
rect 35676 32612 35680 32668
rect 35680 32612 35736 32668
rect 35736 32612 35740 32668
rect 35676 32608 35740 32612
rect 35756 32668 35820 32672
rect 35756 32612 35760 32668
rect 35760 32612 35816 32668
rect 35816 32612 35820 32668
rect 35756 32608 35820 32612
rect 35836 32668 35900 32672
rect 35836 32612 35840 32668
rect 35840 32612 35896 32668
rect 35896 32612 35900 32668
rect 35836 32608 35900 32612
rect 23060 32328 23124 32332
rect 23060 32272 23074 32328
rect 23074 32272 23124 32328
rect 23060 32268 23124 32272
rect 20116 32132 20180 32196
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 18460 32056 18524 32060
rect 18460 32000 18474 32056
rect 18474 32000 18524 32056
rect 18460 31996 18524 32000
rect 28948 31860 29012 31924
rect 4876 31580 4940 31584
rect 4876 31524 4880 31580
rect 4880 31524 4936 31580
rect 4936 31524 4940 31580
rect 4876 31520 4940 31524
rect 4956 31580 5020 31584
rect 4956 31524 4960 31580
rect 4960 31524 5016 31580
rect 5016 31524 5020 31580
rect 4956 31520 5020 31524
rect 5036 31580 5100 31584
rect 5036 31524 5040 31580
rect 5040 31524 5096 31580
rect 5096 31524 5100 31580
rect 5036 31520 5100 31524
rect 5116 31580 5180 31584
rect 5116 31524 5120 31580
rect 5120 31524 5176 31580
rect 5176 31524 5180 31580
rect 5116 31520 5180 31524
rect 35596 31580 35660 31584
rect 35596 31524 35600 31580
rect 35600 31524 35656 31580
rect 35656 31524 35660 31580
rect 35596 31520 35660 31524
rect 35676 31580 35740 31584
rect 35676 31524 35680 31580
rect 35680 31524 35736 31580
rect 35736 31524 35740 31580
rect 35676 31520 35740 31524
rect 35756 31580 35820 31584
rect 35756 31524 35760 31580
rect 35760 31524 35816 31580
rect 35816 31524 35820 31580
rect 35756 31520 35820 31524
rect 35836 31580 35900 31584
rect 35836 31524 35840 31580
rect 35840 31524 35896 31580
rect 35896 31524 35900 31580
rect 35836 31520 35900 31524
rect 23428 31376 23492 31380
rect 23428 31320 23442 31376
rect 23442 31320 23492 31376
rect 23428 31316 23492 31320
rect 27844 31044 27908 31108
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 4876 30492 4940 30496
rect 4876 30436 4880 30492
rect 4880 30436 4936 30492
rect 4936 30436 4940 30492
rect 4876 30432 4940 30436
rect 4956 30492 5020 30496
rect 4956 30436 4960 30492
rect 4960 30436 5016 30492
rect 5016 30436 5020 30492
rect 4956 30432 5020 30436
rect 5036 30492 5100 30496
rect 5036 30436 5040 30492
rect 5040 30436 5096 30492
rect 5096 30436 5100 30492
rect 5036 30432 5100 30436
rect 5116 30492 5180 30496
rect 5116 30436 5120 30492
rect 5120 30436 5176 30492
rect 5176 30436 5180 30492
rect 5116 30432 5180 30436
rect 35596 30492 35660 30496
rect 35596 30436 35600 30492
rect 35600 30436 35656 30492
rect 35656 30436 35660 30492
rect 35596 30432 35660 30436
rect 35676 30492 35740 30496
rect 35676 30436 35680 30492
rect 35680 30436 35736 30492
rect 35736 30436 35740 30492
rect 35676 30432 35740 30436
rect 35756 30492 35820 30496
rect 35756 30436 35760 30492
rect 35760 30436 35816 30492
rect 35816 30436 35820 30492
rect 35756 30432 35820 30436
rect 35836 30492 35900 30496
rect 35836 30436 35840 30492
rect 35840 30436 35896 30492
rect 35896 30436 35900 30492
rect 35836 30432 35900 30436
rect 18276 30424 18340 30428
rect 18276 30368 18326 30424
rect 18326 30368 18340 30424
rect 18276 30364 18340 30368
rect 23980 30364 24044 30428
rect 26740 30424 26804 30428
rect 26740 30368 26754 30424
rect 26754 30368 26804 30424
rect 26740 30364 26804 30368
rect 24900 30228 24964 30292
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 4876 29404 4940 29408
rect 4876 29348 4880 29404
rect 4880 29348 4936 29404
rect 4936 29348 4940 29404
rect 4876 29344 4940 29348
rect 4956 29404 5020 29408
rect 4956 29348 4960 29404
rect 4960 29348 5016 29404
rect 5016 29348 5020 29404
rect 4956 29344 5020 29348
rect 5036 29404 5100 29408
rect 5036 29348 5040 29404
rect 5040 29348 5096 29404
rect 5096 29348 5100 29404
rect 5036 29344 5100 29348
rect 5116 29404 5180 29408
rect 5116 29348 5120 29404
rect 5120 29348 5176 29404
rect 5176 29348 5180 29404
rect 5116 29344 5180 29348
rect 35596 29404 35660 29408
rect 35596 29348 35600 29404
rect 35600 29348 35656 29404
rect 35656 29348 35660 29404
rect 35596 29344 35660 29348
rect 35676 29404 35740 29408
rect 35676 29348 35680 29404
rect 35680 29348 35736 29404
rect 35736 29348 35740 29404
rect 35676 29344 35740 29348
rect 35756 29404 35820 29408
rect 35756 29348 35760 29404
rect 35760 29348 35816 29404
rect 35816 29348 35820 29404
rect 35756 29344 35820 29348
rect 35836 29404 35900 29408
rect 35836 29348 35840 29404
rect 35840 29348 35896 29404
rect 35896 29348 35900 29404
rect 35836 29344 35900 29348
rect 13308 29004 13372 29068
rect 16436 29004 16500 29068
rect 23244 29004 23308 29068
rect 23612 29064 23676 29068
rect 23612 29008 23626 29064
rect 23626 29008 23676 29064
rect 23612 29004 23676 29008
rect 24164 29004 24228 29068
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 20300 28656 20364 28660
rect 20300 28600 20314 28656
rect 20314 28600 20364 28656
rect 20300 28596 20364 28600
rect 4876 28316 4940 28320
rect 4876 28260 4880 28316
rect 4880 28260 4936 28316
rect 4936 28260 4940 28316
rect 4876 28256 4940 28260
rect 4956 28316 5020 28320
rect 4956 28260 4960 28316
rect 4960 28260 5016 28316
rect 5016 28260 5020 28316
rect 4956 28256 5020 28260
rect 5036 28316 5100 28320
rect 5036 28260 5040 28316
rect 5040 28260 5096 28316
rect 5096 28260 5100 28316
rect 5036 28256 5100 28260
rect 5116 28316 5180 28320
rect 5116 28260 5120 28316
rect 5120 28260 5176 28316
rect 5176 28260 5180 28316
rect 5116 28256 5180 28260
rect 35596 28316 35660 28320
rect 35596 28260 35600 28316
rect 35600 28260 35656 28316
rect 35656 28260 35660 28316
rect 35596 28256 35660 28260
rect 35676 28316 35740 28320
rect 35676 28260 35680 28316
rect 35680 28260 35736 28316
rect 35736 28260 35740 28316
rect 35676 28256 35740 28260
rect 35756 28316 35820 28320
rect 35756 28260 35760 28316
rect 35760 28260 35816 28316
rect 35816 28260 35820 28316
rect 35756 28256 35820 28260
rect 35836 28316 35900 28320
rect 35836 28260 35840 28316
rect 35840 28260 35896 28316
rect 35896 28260 35900 28316
rect 35836 28256 35900 28260
rect 23060 27916 23124 27980
rect 28948 27916 29012 27980
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 21956 27704 22020 27708
rect 21956 27648 21970 27704
rect 21970 27648 22020 27704
rect 21956 27644 22020 27648
rect 4876 27228 4940 27232
rect 4876 27172 4880 27228
rect 4880 27172 4936 27228
rect 4936 27172 4940 27228
rect 4876 27168 4940 27172
rect 4956 27228 5020 27232
rect 4956 27172 4960 27228
rect 4960 27172 5016 27228
rect 5016 27172 5020 27228
rect 4956 27168 5020 27172
rect 5036 27228 5100 27232
rect 5036 27172 5040 27228
rect 5040 27172 5096 27228
rect 5096 27172 5100 27228
rect 5036 27168 5100 27172
rect 5116 27228 5180 27232
rect 5116 27172 5120 27228
rect 5120 27172 5176 27228
rect 5176 27172 5180 27228
rect 5116 27168 5180 27172
rect 35596 27228 35660 27232
rect 35596 27172 35600 27228
rect 35600 27172 35656 27228
rect 35656 27172 35660 27228
rect 35596 27168 35660 27172
rect 35676 27228 35740 27232
rect 35676 27172 35680 27228
rect 35680 27172 35736 27228
rect 35736 27172 35740 27228
rect 35676 27168 35740 27172
rect 35756 27228 35820 27232
rect 35756 27172 35760 27228
rect 35760 27172 35816 27228
rect 35816 27172 35820 27228
rect 35756 27168 35820 27172
rect 35836 27228 35900 27232
rect 35836 27172 35840 27228
rect 35840 27172 35896 27228
rect 35896 27172 35900 27228
rect 35836 27168 35900 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 20668 26284 20732 26348
rect 25268 26208 25332 26212
rect 25268 26152 25318 26208
rect 25318 26152 25332 26208
rect 25268 26148 25332 26152
rect 4876 26140 4940 26144
rect 4876 26084 4880 26140
rect 4880 26084 4936 26140
rect 4936 26084 4940 26140
rect 4876 26080 4940 26084
rect 4956 26140 5020 26144
rect 4956 26084 4960 26140
rect 4960 26084 5016 26140
rect 5016 26084 5020 26140
rect 4956 26080 5020 26084
rect 5036 26140 5100 26144
rect 5036 26084 5040 26140
rect 5040 26084 5096 26140
rect 5096 26084 5100 26140
rect 5036 26080 5100 26084
rect 5116 26140 5180 26144
rect 5116 26084 5120 26140
rect 5120 26084 5176 26140
rect 5176 26084 5180 26140
rect 5116 26080 5180 26084
rect 24164 26012 24228 26076
rect 35596 26140 35660 26144
rect 35596 26084 35600 26140
rect 35600 26084 35656 26140
rect 35656 26084 35660 26140
rect 35596 26080 35660 26084
rect 35676 26140 35740 26144
rect 35676 26084 35680 26140
rect 35680 26084 35736 26140
rect 35736 26084 35740 26140
rect 35676 26080 35740 26084
rect 35756 26140 35820 26144
rect 35756 26084 35760 26140
rect 35760 26084 35816 26140
rect 35816 26084 35820 26140
rect 35756 26080 35820 26084
rect 35836 26140 35900 26144
rect 35836 26084 35840 26140
rect 35840 26084 35896 26140
rect 35896 26084 35900 26140
rect 35836 26080 35900 26084
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19380 25060 19444 25124
rect 4876 25052 4940 25056
rect 4876 24996 4880 25052
rect 4880 24996 4936 25052
rect 4936 24996 4940 25052
rect 4876 24992 4940 24996
rect 4956 25052 5020 25056
rect 4956 24996 4960 25052
rect 4960 24996 5016 25052
rect 5016 24996 5020 25052
rect 4956 24992 5020 24996
rect 5036 25052 5100 25056
rect 5036 24996 5040 25052
rect 5040 24996 5096 25052
rect 5096 24996 5100 25052
rect 5036 24992 5100 24996
rect 5116 25052 5180 25056
rect 5116 24996 5120 25052
rect 5120 24996 5176 25052
rect 5176 24996 5180 25052
rect 5116 24992 5180 24996
rect 35596 25052 35660 25056
rect 35596 24996 35600 25052
rect 35600 24996 35656 25052
rect 35656 24996 35660 25052
rect 35596 24992 35660 24996
rect 35676 25052 35740 25056
rect 35676 24996 35680 25052
rect 35680 24996 35736 25052
rect 35736 24996 35740 25052
rect 35676 24992 35740 24996
rect 35756 25052 35820 25056
rect 35756 24996 35760 25052
rect 35760 24996 35816 25052
rect 35816 24996 35820 25052
rect 35756 24992 35820 24996
rect 35836 25052 35900 25056
rect 35836 24996 35840 25052
rect 35840 24996 35896 25052
rect 35896 24996 35900 25052
rect 35836 24992 35900 24996
rect 15516 24924 15580 24988
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 22140 24304 22204 24308
rect 22140 24248 22190 24304
rect 22190 24248 22204 24304
rect 22140 24244 22204 24248
rect 4876 23964 4940 23968
rect 4876 23908 4880 23964
rect 4880 23908 4936 23964
rect 4936 23908 4940 23964
rect 4876 23904 4940 23908
rect 4956 23964 5020 23968
rect 4956 23908 4960 23964
rect 4960 23908 5016 23964
rect 5016 23908 5020 23964
rect 4956 23904 5020 23908
rect 5036 23964 5100 23968
rect 5036 23908 5040 23964
rect 5040 23908 5096 23964
rect 5096 23908 5100 23964
rect 5036 23904 5100 23908
rect 5116 23964 5180 23968
rect 5116 23908 5120 23964
rect 5120 23908 5176 23964
rect 5176 23908 5180 23964
rect 5116 23904 5180 23908
rect 35596 23964 35660 23968
rect 35596 23908 35600 23964
rect 35600 23908 35656 23964
rect 35656 23908 35660 23964
rect 35596 23904 35660 23908
rect 35676 23964 35740 23968
rect 35676 23908 35680 23964
rect 35680 23908 35736 23964
rect 35736 23908 35740 23964
rect 35676 23904 35740 23908
rect 35756 23964 35820 23968
rect 35756 23908 35760 23964
rect 35760 23908 35816 23964
rect 35816 23908 35820 23964
rect 35756 23904 35820 23908
rect 35836 23964 35900 23968
rect 35836 23908 35840 23964
rect 35840 23908 35896 23964
rect 35896 23908 35900 23964
rect 35836 23904 35900 23908
rect 12572 23488 12636 23492
rect 12572 23432 12622 23488
rect 12622 23432 12636 23488
rect 12572 23428 12636 23432
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 4876 22876 4940 22880
rect 4876 22820 4880 22876
rect 4880 22820 4936 22876
rect 4936 22820 4940 22876
rect 4876 22816 4940 22820
rect 4956 22876 5020 22880
rect 4956 22820 4960 22876
rect 4960 22820 5016 22876
rect 5016 22820 5020 22876
rect 4956 22816 5020 22820
rect 5036 22876 5100 22880
rect 5036 22820 5040 22876
rect 5040 22820 5096 22876
rect 5096 22820 5100 22876
rect 5036 22816 5100 22820
rect 5116 22876 5180 22880
rect 5116 22820 5120 22876
rect 5120 22820 5176 22876
rect 5176 22820 5180 22876
rect 5116 22816 5180 22820
rect 35596 22876 35660 22880
rect 35596 22820 35600 22876
rect 35600 22820 35656 22876
rect 35656 22820 35660 22876
rect 35596 22816 35660 22820
rect 35676 22876 35740 22880
rect 35676 22820 35680 22876
rect 35680 22820 35736 22876
rect 35736 22820 35740 22876
rect 35676 22816 35740 22820
rect 35756 22876 35820 22880
rect 35756 22820 35760 22876
rect 35760 22820 35816 22876
rect 35816 22820 35820 22876
rect 35756 22816 35820 22820
rect 35836 22876 35900 22880
rect 35836 22820 35840 22876
rect 35840 22820 35896 22876
rect 35896 22820 35900 22876
rect 35836 22816 35900 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 4876 21788 4940 21792
rect 4876 21732 4880 21788
rect 4880 21732 4936 21788
rect 4936 21732 4940 21788
rect 4876 21728 4940 21732
rect 4956 21788 5020 21792
rect 4956 21732 4960 21788
rect 4960 21732 5016 21788
rect 5016 21732 5020 21788
rect 4956 21728 5020 21732
rect 5036 21788 5100 21792
rect 5036 21732 5040 21788
rect 5040 21732 5096 21788
rect 5096 21732 5100 21788
rect 5036 21728 5100 21732
rect 5116 21788 5180 21792
rect 5116 21732 5120 21788
rect 5120 21732 5176 21788
rect 5176 21732 5180 21788
rect 5116 21728 5180 21732
rect 35596 21788 35660 21792
rect 35596 21732 35600 21788
rect 35600 21732 35656 21788
rect 35656 21732 35660 21788
rect 35596 21728 35660 21732
rect 35676 21788 35740 21792
rect 35676 21732 35680 21788
rect 35680 21732 35736 21788
rect 35736 21732 35740 21788
rect 35676 21728 35740 21732
rect 35756 21788 35820 21792
rect 35756 21732 35760 21788
rect 35760 21732 35816 21788
rect 35816 21732 35820 21788
rect 35756 21728 35820 21732
rect 35836 21788 35900 21792
rect 35836 21732 35840 21788
rect 35840 21732 35896 21788
rect 35896 21732 35900 21788
rect 35836 21728 35900 21732
rect 13860 21720 13924 21724
rect 13860 21664 13910 21720
rect 13910 21664 13924 21720
rect 13860 21660 13924 21664
rect 9812 21524 9876 21588
rect 10364 21584 10428 21588
rect 10364 21528 10378 21584
rect 10378 21528 10428 21584
rect 10364 21524 10428 21528
rect 22876 21448 22940 21452
rect 22876 21392 22890 21448
rect 22890 21392 22940 21448
rect 22876 21388 22940 21392
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 9628 20768 9692 20772
rect 9628 20712 9642 20768
rect 9642 20712 9692 20768
rect 9628 20708 9692 20712
rect 4876 20700 4940 20704
rect 4876 20644 4880 20700
rect 4880 20644 4936 20700
rect 4936 20644 4940 20700
rect 4876 20640 4940 20644
rect 4956 20700 5020 20704
rect 4956 20644 4960 20700
rect 4960 20644 5016 20700
rect 5016 20644 5020 20700
rect 4956 20640 5020 20644
rect 5036 20700 5100 20704
rect 5036 20644 5040 20700
rect 5040 20644 5096 20700
rect 5096 20644 5100 20700
rect 5036 20640 5100 20644
rect 5116 20700 5180 20704
rect 5116 20644 5120 20700
rect 5120 20644 5176 20700
rect 5176 20644 5180 20700
rect 5116 20640 5180 20644
rect 35596 20700 35660 20704
rect 35596 20644 35600 20700
rect 35600 20644 35656 20700
rect 35656 20644 35660 20700
rect 35596 20640 35660 20644
rect 35676 20700 35740 20704
rect 35676 20644 35680 20700
rect 35680 20644 35736 20700
rect 35736 20644 35740 20700
rect 35676 20640 35740 20644
rect 35756 20700 35820 20704
rect 35756 20644 35760 20700
rect 35760 20644 35816 20700
rect 35816 20644 35820 20700
rect 35756 20640 35820 20644
rect 35836 20700 35900 20704
rect 35836 20644 35840 20700
rect 35840 20644 35896 20700
rect 35896 20644 35900 20700
rect 35836 20640 35900 20644
rect 25084 20572 25148 20636
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 4876 19612 4940 19616
rect 4876 19556 4880 19612
rect 4880 19556 4936 19612
rect 4936 19556 4940 19612
rect 4876 19552 4940 19556
rect 4956 19612 5020 19616
rect 4956 19556 4960 19612
rect 4960 19556 5016 19612
rect 5016 19556 5020 19612
rect 4956 19552 5020 19556
rect 5036 19612 5100 19616
rect 5036 19556 5040 19612
rect 5040 19556 5096 19612
rect 5096 19556 5100 19612
rect 5036 19552 5100 19556
rect 5116 19612 5180 19616
rect 5116 19556 5120 19612
rect 5120 19556 5176 19612
rect 5176 19556 5180 19612
rect 5116 19552 5180 19556
rect 35596 19612 35660 19616
rect 35596 19556 35600 19612
rect 35600 19556 35656 19612
rect 35656 19556 35660 19612
rect 35596 19552 35660 19556
rect 35676 19612 35740 19616
rect 35676 19556 35680 19612
rect 35680 19556 35736 19612
rect 35736 19556 35740 19612
rect 35676 19552 35740 19556
rect 35756 19612 35820 19616
rect 35756 19556 35760 19612
rect 35760 19556 35816 19612
rect 35816 19556 35820 19612
rect 35756 19552 35820 19556
rect 35836 19612 35900 19616
rect 35836 19556 35840 19612
rect 35840 19556 35896 19612
rect 35896 19556 35900 19612
rect 35836 19552 35900 19556
rect 22324 19408 22388 19412
rect 22324 19352 22374 19408
rect 22374 19352 22388 19408
rect 22324 19348 22388 19352
rect 20116 19212 20180 19276
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 4876 18524 4940 18528
rect 4876 18468 4880 18524
rect 4880 18468 4936 18524
rect 4936 18468 4940 18524
rect 4876 18464 4940 18468
rect 4956 18524 5020 18528
rect 4956 18468 4960 18524
rect 4960 18468 5016 18524
rect 5016 18468 5020 18524
rect 4956 18464 5020 18468
rect 5036 18524 5100 18528
rect 5036 18468 5040 18524
rect 5040 18468 5096 18524
rect 5096 18468 5100 18524
rect 5036 18464 5100 18468
rect 5116 18524 5180 18528
rect 5116 18468 5120 18524
rect 5120 18468 5176 18524
rect 5176 18468 5180 18524
rect 5116 18464 5180 18468
rect 35596 18524 35660 18528
rect 35596 18468 35600 18524
rect 35600 18468 35656 18524
rect 35656 18468 35660 18524
rect 35596 18464 35660 18468
rect 35676 18524 35740 18528
rect 35676 18468 35680 18524
rect 35680 18468 35736 18524
rect 35736 18468 35740 18524
rect 35676 18464 35740 18468
rect 35756 18524 35820 18528
rect 35756 18468 35760 18524
rect 35760 18468 35816 18524
rect 35816 18468 35820 18524
rect 35756 18464 35820 18468
rect 35836 18524 35900 18528
rect 35836 18468 35840 18524
rect 35840 18468 35896 18524
rect 35896 18468 35900 18524
rect 35836 18464 35900 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 9812 17852 9876 17916
rect 17540 17988 17604 18052
rect 18276 17912 18340 17916
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 18276 17856 18290 17912
rect 18290 17856 18340 17912
rect 18276 17852 18340 17856
rect 21956 17852 22020 17916
rect 23612 17852 23676 17916
rect 26188 17580 26252 17644
rect 24716 17504 24780 17508
rect 24716 17448 24730 17504
rect 24730 17448 24780 17504
rect 24716 17444 24780 17448
rect 4876 17436 4940 17440
rect 4876 17380 4880 17436
rect 4880 17380 4936 17436
rect 4936 17380 4940 17436
rect 4876 17376 4940 17380
rect 4956 17436 5020 17440
rect 4956 17380 4960 17436
rect 4960 17380 5016 17436
rect 5016 17380 5020 17436
rect 4956 17376 5020 17380
rect 5036 17436 5100 17440
rect 5036 17380 5040 17436
rect 5040 17380 5096 17436
rect 5096 17380 5100 17436
rect 5036 17376 5100 17380
rect 5116 17436 5180 17440
rect 5116 17380 5120 17436
rect 5120 17380 5176 17436
rect 5176 17380 5180 17436
rect 5116 17376 5180 17380
rect 35596 17436 35660 17440
rect 35596 17380 35600 17436
rect 35600 17380 35656 17436
rect 35656 17380 35660 17436
rect 35596 17376 35660 17380
rect 35676 17436 35740 17440
rect 35676 17380 35680 17436
rect 35680 17380 35736 17436
rect 35736 17380 35740 17436
rect 35676 17376 35740 17380
rect 35756 17436 35820 17440
rect 35756 17380 35760 17436
rect 35760 17380 35816 17436
rect 35816 17380 35820 17436
rect 35756 17376 35820 17380
rect 35836 17436 35900 17440
rect 35836 17380 35840 17436
rect 35840 17380 35896 17436
rect 35896 17380 35900 17436
rect 35836 17376 35900 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 24532 16552 24596 16556
rect 24532 16496 24546 16552
rect 24546 16496 24596 16552
rect 24532 16492 24596 16496
rect 4876 16348 4940 16352
rect 4876 16292 4880 16348
rect 4880 16292 4936 16348
rect 4936 16292 4940 16348
rect 4876 16288 4940 16292
rect 4956 16348 5020 16352
rect 4956 16292 4960 16348
rect 4960 16292 5016 16348
rect 5016 16292 5020 16348
rect 4956 16288 5020 16292
rect 5036 16348 5100 16352
rect 5036 16292 5040 16348
rect 5040 16292 5096 16348
rect 5096 16292 5100 16348
rect 5036 16288 5100 16292
rect 5116 16348 5180 16352
rect 5116 16292 5120 16348
rect 5120 16292 5176 16348
rect 5176 16292 5180 16348
rect 5116 16288 5180 16292
rect 35596 16348 35660 16352
rect 35596 16292 35600 16348
rect 35600 16292 35656 16348
rect 35656 16292 35660 16348
rect 35596 16288 35660 16292
rect 35676 16348 35740 16352
rect 35676 16292 35680 16348
rect 35680 16292 35736 16348
rect 35736 16292 35740 16348
rect 35676 16288 35740 16292
rect 35756 16348 35820 16352
rect 35756 16292 35760 16348
rect 35760 16292 35816 16348
rect 35816 16292 35820 16348
rect 35756 16288 35820 16292
rect 35836 16348 35900 16352
rect 35836 16292 35840 16348
rect 35840 16292 35896 16348
rect 35896 16292 35900 16348
rect 35836 16288 35900 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 4876 15260 4940 15264
rect 4876 15204 4880 15260
rect 4880 15204 4936 15260
rect 4936 15204 4940 15260
rect 4876 15200 4940 15204
rect 4956 15260 5020 15264
rect 4956 15204 4960 15260
rect 4960 15204 5016 15260
rect 5016 15204 5020 15260
rect 4956 15200 5020 15204
rect 5036 15260 5100 15264
rect 5036 15204 5040 15260
rect 5040 15204 5096 15260
rect 5096 15204 5100 15260
rect 5036 15200 5100 15204
rect 5116 15260 5180 15264
rect 5116 15204 5120 15260
rect 5120 15204 5176 15260
rect 5176 15204 5180 15260
rect 5116 15200 5180 15204
rect 35596 15260 35660 15264
rect 35596 15204 35600 15260
rect 35600 15204 35656 15260
rect 35656 15204 35660 15260
rect 35596 15200 35660 15204
rect 35676 15260 35740 15264
rect 35676 15204 35680 15260
rect 35680 15204 35736 15260
rect 35736 15204 35740 15260
rect 35676 15200 35740 15204
rect 35756 15260 35820 15264
rect 35756 15204 35760 15260
rect 35760 15204 35816 15260
rect 35816 15204 35820 15260
rect 35756 15200 35820 15204
rect 35836 15260 35900 15264
rect 35836 15204 35840 15260
rect 35840 15204 35896 15260
rect 35896 15204 35900 15260
rect 35836 15200 35900 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 4876 14172 4940 14176
rect 4876 14116 4880 14172
rect 4880 14116 4936 14172
rect 4936 14116 4940 14172
rect 4876 14112 4940 14116
rect 4956 14172 5020 14176
rect 4956 14116 4960 14172
rect 4960 14116 5016 14172
rect 5016 14116 5020 14172
rect 4956 14112 5020 14116
rect 5036 14172 5100 14176
rect 5036 14116 5040 14172
rect 5040 14116 5096 14172
rect 5096 14116 5100 14172
rect 5036 14112 5100 14116
rect 5116 14172 5180 14176
rect 5116 14116 5120 14172
rect 5120 14116 5176 14172
rect 5176 14116 5180 14172
rect 5116 14112 5180 14116
rect 35596 14172 35660 14176
rect 35596 14116 35600 14172
rect 35600 14116 35656 14172
rect 35656 14116 35660 14172
rect 35596 14112 35660 14116
rect 35676 14172 35740 14176
rect 35676 14116 35680 14172
rect 35680 14116 35736 14172
rect 35736 14116 35740 14172
rect 35676 14112 35740 14116
rect 35756 14172 35820 14176
rect 35756 14116 35760 14172
rect 35760 14116 35816 14172
rect 35816 14116 35820 14172
rect 35756 14112 35820 14116
rect 35836 14172 35900 14176
rect 35836 14116 35840 14172
rect 35840 14116 35896 14172
rect 35896 14116 35900 14172
rect 35836 14112 35900 14116
rect 9628 13696 9692 13700
rect 9628 13640 9642 13696
rect 9642 13640 9692 13696
rect 9628 13636 9692 13640
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 26740 13364 26804 13428
rect 4876 13084 4940 13088
rect 4876 13028 4880 13084
rect 4880 13028 4936 13084
rect 4936 13028 4940 13084
rect 4876 13024 4940 13028
rect 4956 13084 5020 13088
rect 4956 13028 4960 13084
rect 4960 13028 5016 13084
rect 5016 13028 5020 13084
rect 4956 13024 5020 13028
rect 5036 13084 5100 13088
rect 5036 13028 5040 13084
rect 5040 13028 5096 13084
rect 5096 13028 5100 13084
rect 5036 13024 5100 13028
rect 5116 13084 5180 13088
rect 5116 13028 5120 13084
rect 5120 13028 5176 13084
rect 5176 13028 5180 13084
rect 5116 13024 5180 13028
rect 35596 13084 35660 13088
rect 35596 13028 35600 13084
rect 35600 13028 35656 13084
rect 35656 13028 35660 13084
rect 35596 13024 35660 13028
rect 35676 13084 35740 13088
rect 35676 13028 35680 13084
rect 35680 13028 35736 13084
rect 35736 13028 35740 13084
rect 35676 13024 35740 13028
rect 35756 13084 35820 13088
rect 35756 13028 35760 13084
rect 35760 13028 35816 13084
rect 35816 13028 35820 13084
rect 35756 13024 35820 13028
rect 35836 13084 35900 13088
rect 35836 13028 35840 13084
rect 35840 13028 35896 13084
rect 35896 13028 35900 13084
rect 35836 13024 35900 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 4876 11996 4940 12000
rect 4876 11940 4880 11996
rect 4880 11940 4936 11996
rect 4936 11940 4940 11996
rect 4876 11936 4940 11940
rect 4956 11996 5020 12000
rect 4956 11940 4960 11996
rect 4960 11940 5016 11996
rect 5016 11940 5020 11996
rect 4956 11936 5020 11940
rect 5036 11996 5100 12000
rect 5036 11940 5040 11996
rect 5040 11940 5096 11996
rect 5096 11940 5100 11996
rect 5036 11936 5100 11940
rect 5116 11996 5180 12000
rect 5116 11940 5120 11996
rect 5120 11940 5176 11996
rect 5176 11940 5180 11996
rect 5116 11936 5180 11940
rect 35596 11996 35660 12000
rect 35596 11940 35600 11996
rect 35600 11940 35656 11996
rect 35656 11940 35660 11996
rect 35596 11936 35660 11940
rect 35676 11996 35740 12000
rect 35676 11940 35680 11996
rect 35680 11940 35736 11996
rect 35736 11940 35740 11996
rect 35676 11936 35740 11940
rect 35756 11996 35820 12000
rect 35756 11940 35760 11996
rect 35760 11940 35816 11996
rect 35816 11940 35820 11996
rect 35756 11936 35820 11940
rect 35836 11996 35900 12000
rect 35836 11940 35840 11996
rect 35840 11940 35896 11996
rect 35896 11940 35900 11996
rect 35836 11936 35900 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 16436 10916 16500 10980
rect 4876 10908 4940 10912
rect 4876 10852 4880 10908
rect 4880 10852 4936 10908
rect 4936 10852 4940 10908
rect 4876 10848 4940 10852
rect 4956 10908 5020 10912
rect 4956 10852 4960 10908
rect 4960 10852 5016 10908
rect 5016 10852 5020 10908
rect 4956 10848 5020 10852
rect 5036 10908 5100 10912
rect 5036 10852 5040 10908
rect 5040 10852 5096 10908
rect 5096 10852 5100 10908
rect 5036 10848 5100 10852
rect 5116 10908 5180 10912
rect 5116 10852 5120 10908
rect 5120 10852 5176 10908
rect 5176 10852 5180 10908
rect 5116 10848 5180 10852
rect 35596 10908 35660 10912
rect 35596 10852 35600 10908
rect 35600 10852 35656 10908
rect 35656 10852 35660 10908
rect 35596 10848 35660 10852
rect 35676 10908 35740 10912
rect 35676 10852 35680 10908
rect 35680 10852 35736 10908
rect 35736 10852 35740 10908
rect 35676 10848 35740 10852
rect 35756 10908 35820 10912
rect 35756 10852 35760 10908
rect 35760 10852 35816 10908
rect 35816 10852 35820 10908
rect 35756 10848 35820 10852
rect 35836 10908 35900 10912
rect 35836 10852 35840 10908
rect 35840 10852 35896 10908
rect 35896 10852 35900 10908
rect 35836 10848 35900 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 4876 9820 4940 9824
rect 4876 9764 4880 9820
rect 4880 9764 4936 9820
rect 4936 9764 4940 9820
rect 4876 9760 4940 9764
rect 4956 9820 5020 9824
rect 4956 9764 4960 9820
rect 4960 9764 5016 9820
rect 5016 9764 5020 9820
rect 4956 9760 5020 9764
rect 5036 9820 5100 9824
rect 5036 9764 5040 9820
rect 5040 9764 5096 9820
rect 5096 9764 5100 9820
rect 5036 9760 5100 9764
rect 5116 9820 5180 9824
rect 5116 9764 5120 9820
rect 5120 9764 5176 9820
rect 5176 9764 5180 9820
rect 5116 9760 5180 9764
rect 35596 9820 35660 9824
rect 35596 9764 35600 9820
rect 35600 9764 35656 9820
rect 35656 9764 35660 9820
rect 35596 9760 35660 9764
rect 35676 9820 35740 9824
rect 35676 9764 35680 9820
rect 35680 9764 35736 9820
rect 35736 9764 35740 9820
rect 35676 9760 35740 9764
rect 35756 9820 35820 9824
rect 35756 9764 35760 9820
rect 35760 9764 35816 9820
rect 35816 9764 35820 9820
rect 35756 9760 35820 9764
rect 35836 9820 35900 9824
rect 35836 9764 35840 9820
rect 35840 9764 35896 9820
rect 35896 9764 35900 9820
rect 35836 9760 35900 9764
rect 22324 9616 22388 9620
rect 22324 9560 22338 9616
rect 22338 9560 22388 9616
rect 15516 9420 15580 9484
rect 20668 9420 20732 9484
rect 22324 9556 22388 9560
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 24716 9012 24780 9076
rect 4876 8732 4940 8736
rect 4876 8676 4880 8732
rect 4880 8676 4936 8732
rect 4936 8676 4940 8732
rect 4876 8672 4940 8676
rect 4956 8732 5020 8736
rect 4956 8676 4960 8732
rect 4960 8676 5016 8732
rect 5016 8676 5020 8732
rect 4956 8672 5020 8676
rect 5036 8732 5100 8736
rect 5036 8676 5040 8732
rect 5040 8676 5096 8732
rect 5096 8676 5100 8732
rect 5036 8672 5100 8676
rect 5116 8732 5180 8736
rect 5116 8676 5120 8732
rect 5120 8676 5176 8732
rect 5176 8676 5180 8732
rect 5116 8672 5180 8676
rect 35596 8732 35660 8736
rect 35596 8676 35600 8732
rect 35600 8676 35656 8732
rect 35656 8676 35660 8732
rect 35596 8672 35660 8676
rect 35676 8732 35740 8736
rect 35676 8676 35680 8732
rect 35680 8676 35736 8732
rect 35736 8676 35740 8732
rect 35676 8672 35740 8676
rect 35756 8732 35820 8736
rect 35756 8676 35760 8732
rect 35760 8676 35816 8732
rect 35816 8676 35820 8732
rect 35756 8672 35820 8676
rect 35836 8732 35900 8736
rect 35836 8676 35840 8732
rect 35840 8676 35896 8732
rect 35896 8676 35900 8732
rect 35836 8672 35900 8676
rect 19012 8528 19076 8532
rect 19012 8472 19026 8528
rect 19026 8472 19076 8528
rect 19012 8468 19076 8472
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 4876 7644 4940 7648
rect 4876 7588 4880 7644
rect 4880 7588 4936 7644
rect 4936 7588 4940 7644
rect 4876 7584 4940 7588
rect 4956 7644 5020 7648
rect 4956 7588 4960 7644
rect 4960 7588 5016 7644
rect 5016 7588 5020 7644
rect 4956 7584 5020 7588
rect 5036 7644 5100 7648
rect 5036 7588 5040 7644
rect 5040 7588 5096 7644
rect 5096 7588 5100 7644
rect 5036 7584 5100 7588
rect 5116 7644 5180 7648
rect 5116 7588 5120 7644
rect 5120 7588 5176 7644
rect 5176 7588 5180 7644
rect 5116 7584 5180 7588
rect 35596 7644 35660 7648
rect 35596 7588 35600 7644
rect 35600 7588 35656 7644
rect 35656 7588 35660 7644
rect 35596 7584 35660 7588
rect 35676 7644 35740 7648
rect 35676 7588 35680 7644
rect 35680 7588 35736 7644
rect 35736 7588 35740 7644
rect 35676 7584 35740 7588
rect 35756 7644 35820 7648
rect 35756 7588 35760 7644
rect 35760 7588 35816 7644
rect 35816 7588 35820 7644
rect 35756 7584 35820 7588
rect 35836 7644 35900 7648
rect 35836 7588 35840 7644
rect 35840 7588 35896 7644
rect 35896 7588 35900 7644
rect 35836 7584 35900 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 18460 6836 18524 6900
rect 4876 6556 4940 6560
rect 4876 6500 4880 6556
rect 4880 6500 4936 6556
rect 4936 6500 4940 6556
rect 4876 6496 4940 6500
rect 4956 6556 5020 6560
rect 4956 6500 4960 6556
rect 4960 6500 5016 6556
rect 5016 6500 5020 6556
rect 4956 6496 5020 6500
rect 5036 6556 5100 6560
rect 5036 6500 5040 6556
rect 5040 6500 5096 6556
rect 5096 6500 5100 6556
rect 5036 6496 5100 6500
rect 5116 6556 5180 6560
rect 5116 6500 5120 6556
rect 5120 6500 5176 6556
rect 5176 6500 5180 6556
rect 5116 6496 5180 6500
rect 35596 6556 35660 6560
rect 35596 6500 35600 6556
rect 35600 6500 35656 6556
rect 35656 6500 35660 6556
rect 35596 6496 35660 6500
rect 35676 6556 35740 6560
rect 35676 6500 35680 6556
rect 35680 6500 35736 6556
rect 35736 6500 35740 6556
rect 35676 6496 35740 6500
rect 35756 6556 35820 6560
rect 35756 6500 35760 6556
rect 35760 6500 35816 6556
rect 35816 6500 35820 6556
rect 35756 6496 35820 6500
rect 35836 6556 35900 6560
rect 35836 6500 35840 6556
rect 35840 6500 35896 6556
rect 35896 6500 35900 6556
rect 35836 6496 35900 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 4876 5468 4940 5472
rect 4876 5412 4880 5468
rect 4880 5412 4936 5468
rect 4936 5412 4940 5468
rect 4876 5408 4940 5412
rect 4956 5468 5020 5472
rect 4956 5412 4960 5468
rect 4960 5412 5016 5468
rect 5016 5412 5020 5468
rect 4956 5408 5020 5412
rect 5036 5468 5100 5472
rect 5036 5412 5040 5468
rect 5040 5412 5096 5468
rect 5096 5412 5100 5468
rect 5036 5408 5100 5412
rect 5116 5468 5180 5472
rect 5116 5412 5120 5468
rect 5120 5412 5176 5468
rect 5176 5412 5180 5468
rect 5116 5408 5180 5412
rect 35596 5468 35660 5472
rect 35596 5412 35600 5468
rect 35600 5412 35656 5468
rect 35656 5412 35660 5468
rect 35596 5408 35660 5412
rect 35676 5468 35740 5472
rect 35676 5412 35680 5468
rect 35680 5412 35736 5468
rect 35736 5412 35740 5468
rect 35676 5408 35740 5412
rect 35756 5468 35820 5472
rect 35756 5412 35760 5468
rect 35760 5412 35816 5468
rect 35816 5412 35820 5468
rect 35756 5408 35820 5412
rect 35836 5468 35900 5472
rect 35836 5412 35840 5468
rect 35840 5412 35896 5468
rect 35896 5412 35900 5468
rect 35836 5408 35900 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 4876 4380 4940 4384
rect 4876 4324 4880 4380
rect 4880 4324 4936 4380
rect 4936 4324 4940 4380
rect 4876 4320 4940 4324
rect 4956 4380 5020 4384
rect 4956 4324 4960 4380
rect 4960 4324 5016 4380
rect 5016 4324 5020 4380
rect 4956 4320 5020 4324
rect 5036 4380 5100 4384
rect 5036 4324 5040 4380
rect 5040 4324 5096 4380
rect 5096 4324 5100 4380
rect 5036 4320 5100 4324
rect 5116 4380 5180 4384
rect 5116 4324 5120 4380
rect 5120 4324 5176 4380
rect 5176 4324 5180 4380
rect 5116 4320 5180 4324
rect 35596 4380 35660 4384
rect 35596 4324 35600 4380
rect 35600 4324 35656 4380
rect 35656 4324 35660 4380
rect 35596 4320 35660 4324
rect 35676 4380 35740 4384
rect 35676 4324 35680 4380
rect 35680 4324 35736 4380
rect 35736 4324 35740 4380
rect 35676 4320 35740 4324
rect 35756 4380 35820 4384
rect 35756 4324 35760 4380
rect 35760 4324 35816 4380
rect 35816 4324 35820 4380
rect 35756 4320 35820 4324
rect 35836 4380 35900 4384
rect 35836 4324 35840 4380
rect 35840 4324 35896 4380
rect 35896 4324 35900 4380
rect 35836 4320 35900 4324
rect 12572 4040 12636 4044
rect 12572 3984 12586 4040
rect 12586 3984 12636 4040
rect 12572 3980 12636 3984
rect 13308 3980 13372 4044
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 4876 3292 4940 3296
rect 4876 3236 4880 3292
rect 4880 3236 4936 3292
rect 4936 3236 4940 3292
rect 4876 3232 4940 3236
rect 4956 3292 5020 3296
rect 4956 3236 4960 3292
rect 4960 3236 5016 3292
rect 5016 3236 5020 3292
rect 4956 3232 5020 3236
rect 5036 3292 5100 3296
rect 5036 3236 5040 3292
rect 5040 3236 5096 3292
rect 5096 3236 5100 3292
rect 5036 3232 5100 3236
rect 5116 3292 5180 3296
rect 5116 3236 5120 3292
rect 5120 3236 5176 3292
rect 5176 3236 5180 3292
rect 5116 3232 5180 3236
rect 35596 3292 35660 3296
rect 35596 3236 35600 3292
rect 35600 3236 35656 3292
rect 35656 3236 35660 3292
rect 35596 3232 35660 3236
rect 35676 3292 35740 3296
rect 35676 3236 35680 3292
rect 35680 3236 35736 3292
rect 35736 3236 35740 3292
rect 35676 3232 35740 3236
rect 35756 3292 35820 3296
rect 35756 3236 35760 3292
rect 35760 3236 35816 3292
rect 35816 3236 35820 3292
rect 35756 3232 35820 3236
rect 35836 3292 35900 3296
rect 35836 3236 35840 3292
rect 35840 3236 35896 3292
rect 35896 3236 35900 3292
rect 35836 3232 35900 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 4876 2204 4940 2208
rect 4876 2148 4880 2204
rect 4880 2148 4936 2204
rect 4936 2148 4940 2204
rect 4876 2144 4940 2148
rect 4956 2204 5020 2208
rect 4956 2148 4960 2204
rect 4960 2148 5016 2204
rect 5016 2148 5020 2204
rect 4956 2144 5020 2148
rect 5036 2204 5100 2208
rect 5036 2148 5040 2204
rect 5040 2148 5096 2204
rect 5096 2148 5100 2204
rect 5036 2144 5100 2148
rect 5116 2204 5180 2208
rect 5116 2148 5120 2204
rect 5120 2148 5176 2204
rect 5176 2148 5180 2204
rect 5116 2144 5180 2148
rect 35596 2204 35660 2208
rect 35596 2148 35600 2204
rect 35600 2148 35656 2204
rect 35656 2148 35660 2204
rect 35596 2144 35660 2148
rect 35676 2204 35740 2208
rect 35676 2148 35680 2204
rect 35680 2148 35736 2204
rect 35736 2148 35740 2204
rect 35676 2144 35740 2148
rect 35756 2204 35820 2208
rect 35756 2148 35760 2204
rect 35760 2148 35816 2204
rect 35816 2148 35820 2204
rect 35756 2144 35820 2148
rect 35836 2204 35900 2208
rect 35836 2148 35840 2204
rect 35840 2148 35896 2204
rect 35896 2148 35900 2204
rect 35836 2144 35900 2148
<< metal4 >>
rect 4208 38656 4528 39216
rect 4208 38592 4216 38656
rect 4280 38592 4296 38656
rect 4360 38592 4376 38656
rect 4440 38592 4456 38656
rect 4520 38592 4528 38656
rect 4208 37568 4528 38592
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36260 4528 36416
rect 4208 36024 4250 36260
rect 4486 36024 4528 36260
rect 4208 35392 4528 36024
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5624 4528 5952
rect 4208 5388 4250 5624
rect 4486 5388 4528 5624
rect 4208 4928 4528 5388
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 4868 39200 5188 39216
rect 4868 39136 4876 39200
rect 4940 39136 4956 39200
rect 5020 39136 5036 39200
rect 5100 39136 5116 39200
rect 5180 39136 5188 39200
rect 4868 38112 5188 39136
rect 9811 38860 9877 38861
rect 9811 38796 9812 38860
rect 9876 38796 9877 38860
rect 9811 38795 9877 38796
rect 4868 38048 4876 38112
rect 4940 38048 4956 38112
rect 5020 38048 5036 38112
rect 5100 38048 5116 38112
rect 5180 38048 5188 38112
rect 4868 37024 5188 38048
rect 4868 36960 4876 37024
rect 4940 36960 4956 37024
rect 5020 36960 5036 37024
rect 5100 36960 5116 37024
rect 5180 36960 5188 37024
rect 4868 36920 5188 36960
rect 4868 36684 4910 36920
rect 5146 36684 5188 36920
rect 4868 35936 5188 36684
rect 4868 35872 4876 35936
rect 4940 35872 4956 35936
rect 5020 35872 5036 35936
rect 5100 35872 5116 35936
rect 5180 35872 5188 35936
rect 4868 34848 5188 35872
rect 4868 34784 4876 34848
rect 4940 34784 4956 34848
rect 5020 34784 5036 34848
rect 5100 34784 5116 34848
rect 5180 34784 5188 34848
rect 4868 33760 5188 34784
rect 4868 33696 4876 33760
rect 4940 33696 4956 33760
rect 5020 33696 5036 33760
rect 5100 33696 5116 33760
rect 5180 33696 5188 33760
rect 4868 32672 5188 33696
rect 4868 32608 4876 32672
rect 4940 32608 4956 32672
rect 5020 32608 5036 32672
rect 5100 32608 5116 32672
rect 5180 32608 5188 32672
rect 4868 31584 5188 32608
rect 4868 31520 4876 31584
rect 4940 31520 4956 31584
rect 5020 31520 5036 31584
rect 5100 31520 5116 31584
rect 5180 31520 5188 31584
rect 4868 30496 5188 31520
rect 4868 30432 4876 30496
rect 4940 30432 4956 30496
rect 5020 30432 5036 30496
rect 5100 30432 5116 30496
rect 5180 30432 5188 30496
rect 4868 29408 5188 30432
rect 4868 29344 4876 29408
rect 4940 29344 4956 29408
rect 5020 29344 5036 29408
rect 5100 29344 5116 29408
rect 5180 29344 5188 29408
rect 4868 28320 5188 29344
rect 4868 28256 4876 28320
rect 4940 28256 4956 28320
rect 5020 28256 5036 28320
rect 5100 28256 5116 28320
rect 5180 28256 5188 28320
rect 4868 27232 5188 28256
rect 4868 27168 4876 27232
rect 4940 27168 4956 27232
rect 5020 27168 5036 27232
rect 5100 27168 5116 27232
rect 5180 27168 5188 27232
rect 4868 26144 5188 27168
rect 4868 26080 4876 26144
rect 4940 26080 4956 26144
rect 5020 26080 5036 26144
rect 5100 26080 5116 26144
rect 5180 26080 5188 26144
rect 4868 25056 5188 26080
rect 4868 24992 4876 25056
rect 4940 24992 4956 25056
rect 5020 24992 5036 25056
rect 5100 24992 5116 25056
rect 5180 24992 5188 25056
rect 4868 23968 5188 24992
rect 4868 23904 4876 23968
rect 4940 23904 4956 23968
rect 5020 23904 5036 23968
rect 5100 23904 5116 23968
rect 5180 23904 5188 23968
rect 4868 22880 5188 23904
rect 4868 22816 4876 22880
rect 4940 22816 4956 22880
rect 5020 22816 5036 22880
rect 5100 22816 5116 22880
rect 5180 22816 5188 22880
rect 4868 21792 5188 22816
rect 4868 21728 4876 21792
rect 4940 21728 4956 21792
rect 5020 21728 5036 21792
rect 5100 21728 5116 21792
rect 5180 21728 5188 21792
rect 4868 20704 5188 21728
rect 9814 21589 9874 38795
rect 10363 38724 10429 38725
rect 10363 38660 10364 38724
rect 10428 38660 10429 38724
rect 10363 38659 10429 38660
rect 22875 38724 22941 38725
rect 22875 38660 22876 38724
rect 22940 38660 22941 38724
rect 22875 38659 22941 38660
rect 23979 38724 24045 38725
rect 23979 38660 23980 38724
rect 24044 38660 24045 38724
rect 23979 38659 24045 38660
rect 10366 21589 10426 38659
rect 22139 37364 22205 37365
rect 22139 37300 22140 37364
rect 22204 37300 22205 37364
rect 22139 37299 22205 37300
rect 17539 36004 17605 36005
rect 17539 35940 17540 36004
rect 17604 35940 17605 36004
rect 17539 35939 17605 35940
rect 20299 36004 20365 36005
rect 20299 35940 20300 36004
rect 20364 35940 20365 36004
rect 20299 35939 20365 35940
rect 13859 34644 13925 34645
rect 13859 34580 13860 34644
rect 13924 34580 13925 34644
rect 13859 34579 13925 34580
rect 13307 29068 13373 29069
rect 13307 29004 13308 29068
rect 13372 29004 13373 29068
rect 13307 29003 13373 29004
rect 12571 23492 12637 23493
rect 12571 23428 12572 23492
rect 12636 23428 12637 23492
rect 12571 23427 12637 23428
rect 9811 21588 9877 21589
rect 9811 21524 9812 21588
rect 9876 21524 9877 21588
rect 9811 21523 9877 21524
rect 10363 21588 10429 21589
rect 10363 21524 10364 21588
rect 10428 21524 10429 21588
rect 10363 21523 10429 21524
rect 9627 20772 9693 20773
rect 9627 20708 9628 20772
rect 9692 20708 9693 20772
rect 9627 20707 9693 20708
rect 4868 20640 4876 20704
rect 4940 20640 4956 20704
rect 5020 20640 5036 20704
rect 5100 20640 5116 20704
rect 5180 20640 5188 20704
rect 4868 19616 5188 20640
rect 4868 19552 4876 19616
rect 4940 19552 4956 19616
rect 5020 19552 5036 19616
rect 5100 19552 5116 19616
rect 5180 19552 5188 19616
rect 4868 18528 5188 19552
rect 4868 18464 4876 18528
rect 4940 18464 4956 18528
rect 5020 18464 5036 18528
rect 5100 18464 5116 18528
rect 5180 18464 5188 18528
rect 4868 17440 5188 18464
rect 4868 17376 4876 17440
rect 4940 17376 4956 17440
rect 5020 17376 5036 17440
rect 5100 17376 5116 17440
rect 5180 17376 5188 17440
rect 4868 16352 5188 17376
rect 4868 16288 4876 16352
rect 4940 16288 4956 16352
rect 5020 16288 5036 16352
rect 5100 16288 5116 16352
rect 5180 16288 5188 16352
rect 4868 15264 5188 16288
rect 4868 15200 4876 15264
rect 4940 15200 4956 15264
rect 5020 15200 5036 15264
rect 5100 15200 5116 15264
rect 5180 15200 5188 15264
rect 4868 14176 5188 15200
rect 4868 14112 4876 14176
rect 4940 14112 4956 14176
rect 5020 14112 5036 14176
rect 5100 14112 5116 14176
rect 5180 14112 5188 14176
rect 4868 13088 5188 14112
rect 9630 13701 9690 20707
rect 9814 17917 9874 21523
rect 9811 17916 9877 17917
rect 9811 17852 9812 17916
rect 9876 17852 9877 17916
rect 9811 17851 9877 17852
rect 9627 13700 9693 13701
rect 9627 13636 9628 13700
rect 9692 13636 9693 13700
rect 9627 13635 9693 13636
rect 4868 13024 4876 13088
rect 4940 13024 4956 13088
rect 5020 13024 5036 13088
rect 5100 13024 5116 13088
rect 5180 13024 5188 13088
rect 4868 12000 5188 13024
rect 4868 11936 4876 12000
rect 4940 11936 4956 12000
rect 5020 11936 5036 12000
rect 5100 11936 5116 12000
rect 5180 11936 5188 12000
rect 4868 10912 5188 11936
rect 4868 10848 4876 10912
rect 4940 10848 4956 10912
rect 5020 10848 5036 10912
rect 5100 10848 5116 10912
rect 5180 10848 5188 10912
rect 4868 9824 5188 10848
rect 4868 9760 4876 9824
rect 4940 9760 4956 9824
rect 5020 9760 5036 9824
rect 5100 9760 5116 9824
rect 5180 9760 5188 9824
rect 4868 8736 5188 9760
rect 4868 8672 4876 8736
rect 4940 8672 4956 8736
rect 5020 8672 5036 8736
rect 5100 8672 5116 8736
rect 5180 8672 5188 8736
rect 4868 7648 5188 8672
rect 4868 7584 4876 7648
rect 4940 7584 4956 7648
rect 5020 7584 5036 7648
rect 5100 7584 5116 7648
rect 5180 7584 5188 7648
rect 4868 6560 5188 7584
rect 4868 6496 4876 6560
rect 4940 6496 4956 6560
rect 5020 6496 5036 6560
rect 5100 6496 5116 6560
rect 5180 6496 5188 6560
rect 4868 6284 5188 6496
rect 4868 6048 4910 6284
rect 5146 6048 5188 6284
rect 4868 5472 5188 6048
rect 4868 5408 4876 5472
rect 4940 5408 4956 5472
rect 5020 5408 5036 5472
rect 5100 5408 5116 5472
rect 5180 5408 5188 5472
rect 4868 4384 5188 5408
rect 4868 4320 4876 4384
rect 4940 4320 4956 4384
rect 5020 4320 5036 4384
rect 5100 4320 5116 4384
rect 5180 4320 5188 4384
rect 4868 3296 5188 4320
rect 12574 4045 12634 23427
rect 13310 4045 13370 29003
rect 13862 21725 13922 34579
rect 16435 29068 16501 29069
rect 16435 29004 16436 29068
rect 16500 29004 16501 29068
rect 16435 29003 16501 29004
rect 15515 24988 15581 24989
rect 15515 24924 15516 24988
rect 15580 24924 15581 24988
rect 15515 24923 15581 24924
rect 13859 21724 13925 21725
rect 13859 21660 13860 21724
rect 13924 21660 13925 21724
rect 13859 21659 13925 21660
rect 15518 9485 15578 24923
rect 16438 10981 16498 29003
rect 17542 18053 17602 35939
rect 19011 33284 19077 33285
rect 19011 33220 19012 33284
rect 19076 33220 19077 33284
rect 19011 33219 19077 33220
rect 18459 32060 18525 32061
rect 18459 31996 18460 32060
rect 18524 31996 18525 32060
rect 18459 31995 18525 31996
rect 18275 30428 18341 30429
rect 18275 30364 18276 30428
rect 18340 30364 18341 30428
rect 18275 30363 18341 30364
rect 17539 18052 17605 18053
rect 17539 17988 17540 18052
rect 17604 17988 17605 18052
rect 17539 17987 17605 17988
rect 18278 17917 18338 30363
rect 18275 17916 18341 17917
rect 18275 17852 18276 17916
rect 18340 17852 18341 17916
rect 18275 17851 18341 17852
rect 16435 10980 16501 10981
rect 16435 10916 16436 10980
rect 16500 10916 16501 10980
rect 16435 10915 16501 10916
rect 15515 9484 15581 9485
rect 15515 9420 15516 9484
rect 15580 9420 15581 9484
rect 15515 9419 15581 9420
rect 18462 6901 18522 31995
rect 19014 8533 19074 33219
rect 19379 33148 19445 33149
rect 19379 33084 19380 33148
rect 19444 33084 19445 33148
rect 19379 33083 19445 33084
rect 19382 25125 19442 33083
rect 20115 32196 20181 32197
rect 20115 32132 20116 32196
rect 20180 32132 20181 32196
rect 20115 32131 20181 32132
rect 19379 25124 19445 25125
rect 19379 25060 19380 25124
rect 19444 25060 19445 25124
rect 19379 25059 19445 25060
rect 20118 19277 20178 32131
rect 20302 28661 20362 35939
rect 20299 28660 20365 28661
rect 20299 28596 20300 28660
rect 20364 28596 20365 28660
rect 20299 28595 20365 28596
rect 21955 27708 22021 27709
rect 21955 27644 21956 27708
rect 22020 27644 22021 27708
rect 21955 27643 22021 27644
rect 20667 26348 20733 26349
rect 20667 26284 20668 26348
rect 20732 26284 20733 26348
rect 20667 26283 20733 26284
rect 20115 19276 20181 19277
rect 20115 19212 20116 19276
rect 20180 19212 20181 19276
rect 20115 19211 20181 19212
rect 20670 9485 20730 26283
rect 21958 17917 22018 27643
rect 22142 24309 22202 37299
rect 22139 24308 22205 24309
rect 22139 24244 22140 24308
rect 22204 24244 22205 24308
rect 22139 24243 22205 24244
rect 22878 21453 22938 38659
rect 23427 34644 23493 34645
rect 23427 34580 23428 34644
rect 23492 34580 23493 34644
rect 23427 34579 23493 34580
rect 23243 33692 23309 33693
rect 23243 33628 23244 33692
rect 23308 33628 23309 33692
rect 23243 33627 23309 33628
rect 23059 32332 23125 32333
rect 23059 32268 23060 32332
rect 23124 32268 23125 32332
rect 23059 32267 23125 32268
rect 23062 27981 23122 32267
rect 23246 29069 23306 33627
rect 23430 31381 23490 34579
rect 23427 31380 23493 31381
rect 23427 31316 23428 31380
rect 23492 31316 23493 31380
rect 23427 31315 23493 31316
rect 23982 30429 24042 38659
rect 34928 38656 35248 39216
rect 34928 38592 34936 38656
rect 35000 38592 35016 38656
rect 35080 38592 35096 38656
rect 35160 38592 35176 38656
rect 35240 38592 35248 38656
rect 34928 37568 35248 38592
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 25267 37364 25333 37365
rect 25267 37300 25268 37364
rect 25332 37300 25333 37364
rect 25267 37299 25333 37300
rect 27843 37364 27909 37365
rect 27843 37300 27844 37364
rect 27908 37300 27909 37364
rect 27843 37299 27909 37300
rect 24899 36004 24965 36005
rect 24899 35940 24900 36004
rect 24964 35940 24965 36004
rect 24899 35939 24965 35940
rect 24531 33284 24597 33285
rect 24531 33220 24532 33284
rect 24596 33220 24597 33284
rect 24531 33219 24597 33220
rect 23979 30428 24045 30429
rect 23979 30364 23980 30428
rect 24044 30364 24045 30428
rect 23979 30363 24045 30364
rect 23243 29068 23309 29069
rect 23243 29004 23244 29068
rect 23308 29004 23309 29068
rect 23243 29003 23309 29004
rect 23611 29068 23677 29069
rect 23611 29004 23612 29068
rect 23676 29004 23677 29068
rect 23611 29003 23677 29004
rect 24163 29068 24229 29069
rect 24163 29004 24164 29068
rect 24228 29004 24229 29068
rect 24163 29003 24229 29004
rect 23059 27980 23125 27981
rect 23059 27916 23060 27980
rect 23124 27916 23125 27980
rect 23059 27915 23125 27916
rect 22875 21452 22941 21453
rect 22875 21388 22876 21452
rect 22940 21388 22941 21452
rect 22875 21387 22941 21388
rect 22323 19412 22389 19413
rect 22323 19348 22324 19412
rect 22388 19348 22389 19412
rect 22323 19347 22389 19348
rect 21955 17916 22021 17917
rect 21955 17852 21956 17916
rect 22020 17852 22021 17916
rect 21955 17851 22021 17852
rect 22326 9621 22386 19347
rect 23614 17917 23674 29003
rect 24166 26077 24226 29003
rect 24163 26076 24229 26077
rect 24163 26012 24164 26076
rect 24228 26012 24229 26076
rect 24163 26011 24229 26012
rect 23611 17916 23677 17917
rect 23611 17852 23612 17916
rect 23676 17852 23677 17916
rect 23611 17851 23677 17852
rect 24534 16557 24594 33219
rect 24902 30293 24962 35939
rect 25083 33284 25149 33285
rect 25083 33220 25084 33284
rect 25148 33220 25149 33284
rect 25083 33219 25149 33220
rect 24899 30292 24965 30293
rect 24899 30228 24900 30292
rect 24964 30228 24965 30292
rect 24899 30227 24965 30228
rect 25086 20637 25146 33219
rect 25270 26213 25330 37299
rect 26187 33420 26253 33421
rect 26187 33356 26188 33420
rect 26252 33356 26253 33420
rect 26187 33355 26253 33356
rect 25267 26212 25333 26213
rect 25267 26148 25268 26212
rect 25332 26148 25333 26212
rect 25267 26147 25333 26148
rect 25083 20636 25149 20637
rect 25083 20572 25084 20636
rect 25148 20572 25149 20636
rect 25083 20571 25149 20572
rect 26190 17645 26250 33355
rect 27846 31109 27906 37299
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36260 35248 36416
rect 34928 36024 34970 36260
rect 35206 36024 35248 36260
rect 28947 36004 29013 36005
rect 28947 35940 28948 36004
rect 29012 35940 29013 36004
rect 28947 35939 29013 35940
rect 28950 33149 29010 35939
rect 34928 35392 35248 36024
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 28947 33148 29013 33149
rect 28947 33084 28948 33148
rect 29012 33084 29013 33148
rect 28947 33083 29013 33084
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 28947 31924 29013 31925
rect 28947 31860 28948 31924
rect 29012 31860 29013 31924
rect 28947 31859 29013 31860
rect 27843 31108 27909 31109
rect 27843 31044 27844 31108
rect 27908 31044 27909 31108
rect 27843 31043 27909 31044
rect 26739 30428 26805 30429
rect 26739 30364 26740 30428
rect 26804 30364 26805 30428
rect 26739 30363 26805 30364
rect 26187 17644 26253 17645
rect 26187 17580 26188 17644
rect 26252 17580 26253 17644
rect 26187 17579 26253 17580
rect 24715 17508 24781 17509
rect 24715 17444 24716 17508
rect 24780 17444 24781 17508
rect 24715 17443 24781 17444
rect 24531 16556 24597 16557
rect 24531 16492 24532 16556
rect 24596 16492 24597 16556
rect 24531 16491 24597 16492
rect 22323 9620 22389 9621
rect 22323 9556 22324 9620
rect 22388 9556 22389 9620
rect 22323 9555 22389 9556
rect 20667 9484 20733 9485
rect 20667 9420 20668 9484
rect 20732 9420 20733 9484
rect 20667 9419 20733 9420
rect 24718 9077 24778 17443
rect 26742 13429 26802 30363
rect 28950 27981 29010 31859
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 28947 27980 29013 27981
rect 28947 27916 28948 27980
rect 29012 27916 29013 27980
rect 28947 27915 29013 27916
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 26739 13428 26805 13429
rect 26739 13364 26740 13428
rect 26804 13364 26805 13428
rect 26739 13363 26805 13364
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 24715 9076 24781 9077
rect 24715 9012 24716 9076
rect 24780 9012 24781 9076
rect 24715 9011 24781 9012
rect 19011 8532 19077 8533
rect 19011 8468 19012 8532
rect 19076 8468 19077 8532
rect 19011 8467 19077 8468
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 18459 6900 18525 6901
rect 18459 6836 18460 6900
rect 18524 6836 18525 6900
rect 18459 6835 18525 6836
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5624 35248 5952
rect 34928 5388 34970 5624
rect 35206 5388 35248 5624
rect 34928 4928 35248 5388
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 12571 4044 12637 4045
rect 12571 3980 12572 4044
rect 12636 3980 12637 4044
rect 12571 3979 12637 3980
rect 13307 4044 13373 4045
rect 13307 3980 13308 4044
rect 13372 3980 13373 4044
rect 13307 3979 13373 3980
rect 4868 3232 4876 3296
rect 4940 3232 4956 3296
rect 5020 3232 5036 3296
rect 5100 3232 5116 3296
rect 5180 3232 5188 3296
rect 4868 2208 5188 3232
rect 4868 2144 4876 2208
rect 4940 2144 4956 2208
rect 5020 2144 5036 2208
rect 5100 2144 5116 2208
rect 5180 2144 5188 2208
rect 4868 2128 5188 2144
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 35588 39200 35908 39216
rect 35588 39136 35596 39200
rect 35660 39136 35676 39200
rect 35740 39136 35756 39200
rect 35820 39136 35836 39200
rect 35900 39136 35908 39200
rect 35588 38112 35908 39136
rect 35588 38048 35596 38112
rect 35660 38048 35676 38112
rect 35740 38048 35756 38112
rect 35820 38048 35836 38112
rect 35900 38048 35908 38112
rect 35588 37024 35908 38048
rect 35588 36960 35596 37024
rect 35660 36960 35676 37024
rect 35740 36960 35756 37024
rect 35820 36960 35836 37024
rect 35900 36960 35908 37024
rect 35588 36920 35908 36960
rect 35588 36684 35630 36920
rect 35866 36684 35908 36920
rect 35588 35936 35908 36684
rect 35588 35872 35596 35936
rect 35660 35872 35676 35936
rect 35740 35872 35756 35936
rect 35820 35872 35836 35936
rect 35900 35872 35908 35936
rect 35588 34848 35908 35872
rect 35588 34784 35596 34848
rect 35660 34784 35676 34848
rect 35740 34784 35756 34848
rect 35820 34784 35836 34848
rect 35900 34784 35908 34848
rect 35588 33760 35908 34784
rect 35588 33696 35596 33760
rect 35660 33696 35676 33760
rect 35740 33696 35756 33760
rect 35820 33696 35836 33760
rect 35900 33696 35908 33760
rect 35588 32672 35908 33696
rect 35588 32608 35596 32672
rect 35660 32608 35676 32672
rect 35740 32608 35756 32672
rect 35820 32608 35836 32672
rect 35900 32608 35908 32672
rect 35588 31584 35908 32608
rect 35588 31520 35596 31584
rect 35660 31520 35676 31584
rect 35740 31520 35756 31584
rect 35820 31520 35836 31584
rect 35900 31520 35908 31584
rect 35588 30496 35908 31520
rect 35588 30432 35596 30496
rect 35660 30432 35676 30496
rect 35740 30432 35756 30496
rect 35820 30432 35836 30496
rect 35900 30432 35908 30496
rect 35588 29408 35908 30432
rect 35588 29344 35596 29408
rect 35660 29344 35676 29408
rect 35740 29344 35756 29408
rect 35820 29344 35836 29408
rect 35900 29344 35908 29408
rect 35588 28320 35908 29344
rect 35588 28256 35596 28320
rect 35660 28256 35676 28320
rect 35740 28256 35756 28320
rect 35820 28256 35836 28320
rect 35900 28256 35908 28320
rect 35588 27232 35908 28256
rect 35588 27168 35596 27232
rect 35660 27168 35676 27232
rect 35740 27168 35756 27232
rect 35820 27168 35836 27232
rect 35900 27168 35908 27232
rect 35588 26144 35908 27168
rect 35588 26080 35596 26144
rect 35660 26080 35676 26144
rect 35740 26080 35756 26144
rect 35820 26080 35836 26144
rect 35900 26080 35908 26144
rect 35588 25056 35908 26080
rect 35588 24992 35596 25056
rect 35660 24992 35676 25056
rect 35740 24992 35756 25056
rect 35820 24992 35836 25056
rect 35900 24992 35908 25056
rect 35588 23968 35908 24992
rect 35588 23904 35596 23968
rect 35660 23904 35676 23968
rect 35740 23904 35756 23968
rect 35820 23904 35836 23968
rect 35900 23904 35908 23968
rect 35588 22880 35908 23904
rect 35588 22816 35596 22880
rect 35660 22816 35676 22880
rect 35740 22816 35756 22880
rect 35820 22816 35836 22880
rect 35900 22816 35908 22880
rect 35588 21792 35908 22816
rect 35588 21728 35596 21792
rect 35660 21728 35676 21792
rect 35740 21728 35756 21792
rect 35820 21728 35836 21792
rect 35900 21728 35908 21792
rect 35588 20704 35908 21728
rect 35588 20640 35596 20704
rect 35660 20640 35676 20704
rect 35740 20640 35756 20704
rect 35820 20640 35836 20704
rect 35900 20640 35908 20704
rect 35588 19616 35908 20640
rect 35588 19552 35596 19616
rect 35660 19552 35676 19616
rect 35740 19552 35756 19616
rect 35820 19552 35836 19616
rect 35900 19552 35908 19616
rect 35588 18528 35908 19552
rect 35588 18464 35596 18528
rect 35660 18464 35676 18528
rect 35740 18464 35756 18528
rect 35820 18464 35836 18528
rect 35900 18464 35908 18528
rect 35588 17440 35908 18464
rect 35588 17376 35596 17440
rect 35660 17376 35676 17440
rect 35740 17376 35756 17440
rect 35820 17376 35836 17440
rect 35900 17376 35908 17440
rect 35588 16352 35908 17376
rect 35588 16288 35596 16352
rect 35660 16288 35676 16352
rect 35740 16288 35756 16352
rect 35820 16288 35836 16352
rect 35900 16288 35908 16352
rect 35588 15264 35908 16288
rect 35588 15200 35596 15264
rect 35660 15200 35676 15264
rect 35740 15200 35756 15264
rect 35820 15200 35836 15264
rect 35900 15200 35908 15264
rect 35588 14176 35908 15200
rect 35588 14112 35596 14176
rect 35660 14112 35676 14176
rect 35740 14112 35756 14176
rect 35820 14112 35836 14176
rect 35900 14112 35908 14176
rect 35588 13088 35908 14112
rect 35588 13024 35596 13088
rect 35660 13024 35676 13088
rect 35740 13024 35756 13088
rect 35820 13024 35836 13088
rect 35900 13024 35908 13088
rect 35588 12000 35908 13024
rect 35588 11936 35596 12000
rect 35660 11936 35676 12000
rect 35740 11936 35756 12000
rect 35820 11936 35836 12000
rect 35900 11936 35908 12000
rect 35588 10912 35908 11936
rect 35588 10848 35596 10912
rect 35660 10848 35676 10912
rect 35740 10848 35756 10912
rect 35820 10848 35836 10912
rect 35900 10848 35908 10912
rect 35588 9824 35908 10848
rect 35588 9760 35596 9824
rect 35660 9760 35676 9824
rect 35740 9760 35756 9824
rect 35820 9760 35836 9824
rect 35900 9760 35908 9824
rect 35588 8736 35908 9760
rect 35588 8672 35596 8736
rect 35660 8672 35676 8736
rect 35740 8672 35756 8736
rect 35820 8672 35836 8736
rect 35900 8672 35908 8736
rect 35588 7648 35908 8672
rect 35588 7584 35596 7648
rect 35660 7584 35676 7648
rect 35740 7584 35756 7648
rect 35820 7584 35836 7648
rect 35900 7584 35908 7648
rect 35588 6560 35908 7584
rect 35588 6496 35596 6560
rect 35660 6496 35676 6560
rect 35740 6496 35756 6560
rect 35820 6496 35836 6560
rect 35900 6496 35908 6560
rect 35588 6284 35908 6496
rect 35588 6048 35630 6284
rect 35866 6048 35908 6284
rect 35588 5472 35908 6048
rect 35588 5408 35596 5472
rect 35660 5408 35676 5472
rect 35740 5408 35756 5472
rect 35820 5408 35836 5472
rect 35900 5408 35908 5472
rect 35588 4384 35908 5408
rect 35588 4320 35596 4384
rect 35660 4320 35676 4384
rect 35740 4320 35756 4384
rect 35820 4320 35836 4384
rect 35900 4320 35908 4384
rect 35588 3296 35908 4320
rect 35588 3232 35596 3296
rect 35660 3232 35676 3296
rect 35740 3232 35756 3296
rect 35820 3232 35836 3296
rect 35900 3232 35908 3296
rect 35588 2208 35908 3232
rect 35588 2144 35596 2208
rect 35660 2144 35676 2208
rect 35740 2144 35756 2208
rect 35820 2144 35836 2208
rect 35900 2144 35908 2208
rect 35588 2128 35908 2144
<< via4 >>
rect 4250 36024 4486 36260
rect 4250 5388 4486 5624
rect 4910 36684 5146 36920
rect 4910 6048 5146 6284
rect 34970 36024 35206 36260
rect 34970 5388 35206 5624
rect 35630 36684 35866 36920
rect 35630 6048 35866 6284
<< metal5 >>
rect 1056 36920 38320 36962
rect 1056 36684 4910 36920
rect 5146 36684 35630 36920
rect 35866 36684 38320 36920
rect 1056 36642 38320 36684
rect 1056 36260 38320 36302
rect 1056 36024 4250 36260
rect 4486 36024 34970 36260
rect 35206 36024 38320 36260
rect 1056 35982 38320 36024
rect 1056 6284 38320 6326
rect 1056 6048 4910 6284
rect 5146 6048 35630 6284
rect 35866 6048 38320 6284
rect 1056 6006 38320 6048
rect 1056 5624 38320 5666
rect 1056 5388 4250 5624
rect 4486 5388 34970 5624
rect 35206 5388 38320 5624
rect 1056 5346 38320 5388
use sky130_fd_sc_hd__inv_2  _1275_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 20332 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_8  _1276_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13156 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__inv_2  _1277_
timestamp 1688980957
transform 1 0 17388 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1278_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20332 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  _1279_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14168 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _1280_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13248 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_8  _1281_
timestamp 1688980957
transform 1 0 16836 0 -1 13056
box -38 -48 1050 592
use sky130_fd_sc_hd__or2_1  _1282_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14996 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _1283_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15272 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1284_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12696 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _1285_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 14812 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_8  _1286_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13708 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_8  _1287_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22724 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__o21a_2  _1288_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 22172 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2b_4  _1289_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15364 0 -1 14144
box -38 -48 1050 592
use sky130_fd_sc_hd__a21boi_1  _1290_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15456 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1291_
timestamp 1688980957
transform -1 0 16468 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_4  _1292_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 2062 592
use sky130_fd_sc_hd__nand3b_2  _1293_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 14904 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and3b_1  _1294_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14260 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_4  _1295_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15824 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__and2b_1  _1296_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 14536 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1297_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 16100 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _1298_
timestamp 1688980957
transform 1 0 18768 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and4bb_4  _1299_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 18768 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__or4bb_1  _1300_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15088 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__o221ai_4  _1301_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_8  _1302_
timestamp 1688980957
transform -1 0 16468 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__a221oi_2  _1303_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 16928 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1304_
timestamp 1688980957
transform 1 0 20700 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _1305_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1306_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 21252 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1307_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 20884 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _1308_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20424 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _1309_
timestamp 1688980957
transform 1 0 20792 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1310_
timestamp 1688980957
transform -1 0 14536 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_8  _1311_
timestamp 1688980957
transform -1 0 14260 0 -1 23936
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_8  _1312_
timestamp 1688980957
transform 1 0 23000 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__nand2_1  _1313_
timestamp 1688980957
transform -1 0 18216 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1314_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17020 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1315_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12052 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _1316_
timestamp 1688980957
transform 1 0 12512 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1317_
timestamp 1688980957
transform 1 0 15364 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and3b_1  _1318_
timestamp 1688980957
transform 1 0 16100 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1319_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 17296 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1320_
timestamp 1688980957
transform 1 0 16560 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o311a_4  _1321_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 18308 0 -1 15232
box -38 -48 1602 592
use sky130_fd_sc_hd__o211a_1  _1322_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20240 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _1323_
timestamp 1688980957
transform -1 0 20056 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__or4bb_1  _1324_
timestamp 1688980957
transform 1 0 18676 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__nand2b_1  _1325_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19504 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1326_
timestamp 1688980957
transform 1 0 18768 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1327_
timestamp 1688980957
transform 1 0 17756 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _1328_
timestamp 1688980957
transform 1 0 16652 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_4  _1329_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 -1 18496
box -38 -48 2062 592
use sky130_fd_sc_hd__o211a_1  _1330_
timestamp 1688980957
transform -1 0 18676 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_4  _1331_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 19780 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_8  _1332_
timestamp 1688980957
transform 1 0 18216 0 -1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_4  _1333_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 28796 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_2  _1334_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15640 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_8  _1335_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12420 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__or3_4  _1336_
timestamp 1688980957
transform -1 0 14904 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _1337_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15364 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__a22o_4  _1338_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14720 0 1 22848
box -38 -48 1326 592
use sky130_fd_sc_hd__and2_1  _1339_
timestamp 1688980957
transform 1 0 12880 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_8  _1340_
timestamp 1688980957
transform 1 0 13984 0 -1 35904
box -38 -48 1050 592
use sky130_fd_sc_hd__o2bb2a_2  _1341_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15180 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_4  _1342_
timestamp 1688980957
transform 1 0 14168 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__and3_1  _1343_
timestamp 1688980957
transform 1 0 13524 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_8  _1344_
timestamp 1688980957
transform 1 0 15364 0 -1 25024
box -38 -48 1050 592
use sky130_fd_sc_hd__a221o_1  _1345_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27232 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1346_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 28520 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1347_
timestamp 1688980957
transform -1 0 30268 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1348_
timestamp 1688980957
transform 1 0 29900 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_2  _1349_
timestamp 1688980957
transform 1 0 18492 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_8  _1350_
timestamp 1688980957
transform 1 0 19228 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__or2_2  _1351_
timestamp 1688980957
transform 1 0 16100 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1352_
timestamp 1688980957
transform -1 0 19044 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or3b_4  _1353_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19964 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1354_
timestamp 1688980957
transform -1 0 12328 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o2111ai_4  _1355_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16836 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__a21o_4  _1356_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16192 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _1357_
timestamp 1688980957
transform 1 0 17296 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1358_
timestamp 1688980957
transform -1 0 20424 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1359_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 19872 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_4  _1360_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18860 0 -1 21760
box -38 -48 1326 592
use sky130_fd_sc_hd__nand2_8  _1361_
timestamp 1688980957
transform 1 0 19228 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_8  _1362_
timestamp 1688980957
transform 1 0 16100 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__o22ai_4  _1363_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 20700 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_8  _1364_
timestamp 1688980957
transform 1 0 20884 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__a21oi_4  _1365_
timestamp 1688980957
transform -1 0 18124 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_4  _1366_
timestamp 1688980957
transform -1 0 20056 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1367_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24840 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_8  _1368_
timestamp 1688980957
transform 1 0 20700 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__a211o_1  _1369_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 26772 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1370_
timestamp 1688980957
transform 1 0 26036 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1371_
timestamp 1688980957
transform 1 0 25668 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1372_
timestamp 1688980957
transform -1 0 30728 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1373_
timestamp 1688980957
transform -1 0 29900 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1374_
timestamp 1688980957
transform -1 0 30452 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1375_
timestamp 1688980957
transform 1 0 29624 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1376_
timestamp 1688980957
transform 1 0 30268 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1377_
timestamp 1688980957
transform -1 0 32016 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_2  _1378_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 32108 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1379_
timestamp 1688980957
transform 1 0 25668 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1380_
timestamp 1688980957
transform 1 0 26220 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1381_
timestamp 1688980957
transform 1 0 25484 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _1382_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25760 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _1383_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 36064 0 -1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__a221o_1  _1384_
timestamp 1688980957
transform 1 0 30360 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1385_
timestamp 1688980957
transform -1 0 32016 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1386_
timestamp 1688980957
transform -1 0 33672 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1387_
timestamp 1688980957
transform 1 0 25392 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1388_
timestamp 1688980957
transform 1 0 26036 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1389_
timestamp 1688980957
transform -1 0 26680 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1390_
timestamp 1688980957
transform 1 0 26956 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1391_
timestamp 1688980957
transform -1 0 36616 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1392_
timestamp 1688980957
transform 1 0 36616 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1393_
timestamp 1688980957
transform -1 0 37076 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1394_
timestamp 1688980957
transform 1 0 36616 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1395_
timestamp 1688980957
transform 1 0 30452 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1396_
timestamp 1688980957
transform -1 0 32016 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_4  _1397_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 33672 0 -1 32640
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_1  _1398_
timestamp 1688980957
transform 1 0 21804 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1399_
timestamp 1688980957
transform -1 0 26680 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1400_
timestamp 1688980957
transform 1 0 25392 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1401_
timestamp 1688980957
transform 1 0 24840 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1402_
timestamp 1688980957
transform 1 0 25024 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1403_
timestamp 1688980957
transform -1 0 33672 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1404_
timestamp 1688980957
transform 1 0 27140 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1405_
timestamp 1688980957
transform -1 0 28980 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1406_
timestamp 1688980957
transform -1 0 30728 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1407_
timestamp 1688980957
transform -1 0 25944 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1408_
timestamp 1688980957
transform 1 0 24748 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1409_
timestamp 1688980957
transform -1 0 25300 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1410_
timestamp 1688980957
transform 1 0 25024 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1411_
timestamp 1688980957
transform 1 0 31004 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1412_
timestamp 1688980957
transform 1 0 31004 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1413_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 31464 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1414_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16284 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _1415_
timestamp 1688980957
transform -1 0 18584 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1416_
timestamp 1688980957
transform 1 0 17296 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _1417_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17756 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__and4_4  _1418_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15088 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a31oi_4  _1419_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17296 0 1 22848
box -38 -48 1602 592
use sky130_fd_sc_hd__o211a_2  _1420_
timestamp 1688980957
transform -1 0 17572 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1421_
timestamp 1688980957
transform -1 0 23460 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_2  _1422_
timestamp 1688980957
transform 1 0 15732 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1423_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 17756 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_2  _1424_
timestamp 1688980957
transform -1 0 17112 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _1425_
timestamp 1688980957
transform 1 0 20700 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1426_
timestamp 1688980957
transform 1 0 21896 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _1427_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19872 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_4  _1428_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 17940 0 -1 25024
box -38 -48 1326 592
use sky130_fd_sc_hd__nor4_1  _1429_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15640 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1430_
timestamp 1688980957
transform 1 0 22632 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _1431_
timestamp 1688980957
transform 1 0 21344 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o32a_2  _1432_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22540 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _1433_
timestamp 1688980957
transform 1 0 11684 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1434_
timestamp 1688980957
transform 1 0 11500 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _1435_
timestamp 1688980957
transform 1 0 12236 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1436_
timestamp 1688980957
transform 1 0 18400 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _1437_
timestamp 1688980957
transform 1 0 19228 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_4  _1438_
timestamp 1688980957
transform 1 0 22080 0 -1 18496
box -38 -48 1602 592
use sky130_fd_sc_hd__nand2_1  _1439_
timestamp 1688980957
transform -1 0 18860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _1440_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18400 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and3_4  _1441_
timestamp 1688980957
transform 1 0 18308 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_2  _1442_
timestamp 1688980957
transform -1 0 17572 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and3_2  _1443_
timestamp 1688980957
transform 1 0 16652 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1444_
timestamp 1688980957
transform 1 0 24380 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and3_4  _1445_
timestamp 1688980957
transform 1 0 18308 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _1446_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16928 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1447_
timestamp 1688980957
transform 1 0 23184 0 1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1448_
timestamp 1688980957
transform 1 0 23736 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1449_
timestamp 1688980957
transform 1 0 17848 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _1450_
timestamp 1688980957
transform 1 0 20424 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _1451_
timestamp 1688980957
transform 1 0 17296 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1452_
timestamp 1688980957
transform 1 0 21804 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1453_
timestamp 1688980957
transform 1 0 23368 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _1454_
timestamp 1688980957
transform 1 0 24472 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1455_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 25668 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1456_
timestamp 1688980957
transform 1 0 20148 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1457_
timestamp 1688980957
transform 1 0 20976 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1458_
timestamp 1688980957
transform 1 0 20332 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_4  _1459_
timestamp 1688980957
transform 1 0 25208 0 -1 31552
box -38 -48 1602 592
use sky130_fd_sc_hd__nand2_1  _1460_
timestamp 1688980957
transform 1 0 28244 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1461_
timestamp 1688980957
transform -1 0 32384 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1462_
timestamp 1688980957
transform -1 0 32844 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1463_
timestamp 1688980957
transform 1 0 32844 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and4_1  _1464_
timestamp 1688980957
transform 1 0 14076 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1465_
timestamp 1688980957
transform 1 0 13524 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _1466_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14168 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1467_
timestamp 1688980957
transform -1 0 15732 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1468_
timestamp 1688980957
transform -1 0 15088 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _1469_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14260 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1470_
timestamp 1688980957
transform 1 0 12236 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1471_
timestamp 1688980957
transform 1 0 12420 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_2  _1472_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13248 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _1473_
timestamp 1688980957
transform 1 0 17940 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__and3_2  _1474_
timestamp 1688980957
transform -1 0 21528 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1475_
timestamp 1688980957
transform -1 0 17296 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1476_
timestamp 1688980957
transform 1 0 16652 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1477_
timestamp 1688980957
transform 1 0 16008 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1478_
timestamp 1688980957
transform 1 0 16836 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1479_
timestamp 1688980957
transform 1 0 16100 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1480_
timestamp 1688980957
transform 1 0 17664 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1481_
timestamp 1688980957
transform -1 0 19228 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1482_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 16100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1483_
timestamp 1688980957
transform 1 0 16652 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1484_
timestamp 1688980957
transform -1 0 18124 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or2_2  _1485_
timestamp 1688980957
transform -1 0 18492 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_2  _1486_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 18952 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _1487_
timestamp 1688980957
transform -1 0 18216 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_4  _1488_
timestamp 1688980957
transform -1 0 19504 0 -1 9792
box -38 -48 1326 592
use sky130_fd_sc_hd__nor2_1  _1489_
timestamp 1688980957
transform -1 0 25208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and4_1  _1490_
timestamp 1688980957
transform -1 0 17296 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1491_
timestamp 1688980957
transform 1 0 16560 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1492_
timestamp 1688980957
transform 1 0 16100 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1493_
timestamp 1688980957
transform 1 0 17388 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1494_
timestamp 1688980957
transform 1 0 15916 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1495_
timestamp 1688980957
transform 1 0 17664 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1496_
timestamp 1688980957
transform 1 0 18492 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _1497_
timestamp 1688980957
transform -1 0 15916 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1498_
timestamp 1688980957
transform 1 0 16652 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1499_
timestamp 1688980957
transform 1 0 18124 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a311o_1  _1500_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 18952 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1501_
timestamp 1688980957
transform -1 0 18768 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__and4_1  _1502_
timestamp 1688980957
transform 1 0 13340 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1503_
timestamp 1688980957
transform 1 0 13064 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _1504_
timestamp 1688980957
transform 1 0 14076 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1505_
timestamp 1688980957
transform -1 0 16376 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1506_
timestamp 1688980957
transform -1 0 15732 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o32a_1  _1507_
timestamp 1688980957
transform 1 0 14076 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1508_
timestamp 1688980957
transform 1 0 11592 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1509_
timestamp 1688980957
transform 1 0 11500 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1510_
timestamp 1688980957
transform 1 0 13248 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1511_
timestamp 1688980957
transform 1 0 17572 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1512_
timestamp 1688980957
transform 1 0 19228 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1513_
timestamp 1688980957
transform 1 0 28980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1514_
timestamp 1688980957
transform 1 0 13984 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1515_
timestamp 1688980957
transform 1 0 13156 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _1516_
timestamp 1688980957
transform -1 0 15180 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1517_
timestamp 1688980957
transform -1 0 20516 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1518_
timestamp 1688980957
transform 1 0 18400 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _1519_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 19596 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1520_
timestamp 1688980957
transform 1 0 20700 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1521_
timestamp 1688980957
transform -1 0 12236 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1522_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11592 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _1523_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 19964 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_4  _1524_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 20700 0 -1 33728
box -38 -48 1694 592
use sky130_fd_sc_hd__or2_1  _1525_
timestamp 1688980957
transform 1 0 18860 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1526_
timestamp 1688980957
transform -1 0 18032 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1527_
timestamp 1688980957
transform -1 0 18768 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a22oi_1  _1528_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19780 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1529_
timestamp 1688980957
transform -1 0 17480 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1530_
timestamp 1688980957
transform 1 0 15364 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1531_
timestamp 1688980957
transform -1 0 16744 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a2111oi_1  _1532_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16652 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _1533_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18676 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__and3_1  _1534_
timestamp 1688980957
transform 1 0 17204 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1535_
timestamp 1688980957
transform 1 0 17664 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a211oi_1  _1536_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18308 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_2  _1537_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18308 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1538_
timestamp 1688980957
transform 1 0 18032 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1539_
timestamp 1688980957
transform 1 0 19320 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1540_
timestamp 1688980957
transform 1 0 18308 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_1  _1541_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17572 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _1542_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18400 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1543_
timestamp 1688980957
transform -1 0 22816 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1544_
timestamp 1688980957
transform 1 0 21068 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1545_
timestamp 1688980957
transform 1 0 22172 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1546_
timestamp 1688980957
transform 1 0 20240 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1547_
timestamp 1688980957
transform 1 0 20792 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1548_
timestamp 1688980957
transform -1 0 23920 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1549_
timestamp 1688980957
transform 1 0 22264 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1550_
timestamp 1688980957
transform 1 0 20424 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1551_
timestamp 1688980957
transform -1 0 21804 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1552_
timestamp 1688980957
transform 1 0 20516 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _1553_
timestamp 1688980957
transform -1 0 22172 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__and4_1  _1554_
timestamp 1688980957
transform 1 0 18492 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1555_
timestamp 1688980957
transform -1 0 19872 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o2111a_1  _1556_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20056 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__o2111a_1  _1557_
timestamp 1688980957
transform 1 0 19228 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__o2111a_1  _1558_
timestamp 1688980957
transform 1 0 19504 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a2111o_1  _1559_
timestamp 1688980957
transform 1 0 18676 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a2111o_1  _1560_
timestamp 1688980957
transform 1 0 18308 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_1  _1561_
timestamp 1688980957
transform -1 0 13524 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1562_
timestamp 1688980957
transform 1 0 12144 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1563_
timestamp 1688980957
transform 1 0 12788 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1564_
timestamp 1688980957
transform 1 0 18216 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1565_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19320 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1566_
timestamp 1688980957
transform 1 0 19504 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1567_
timestamp 1688980957
transform -1 0 20056 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1568_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _1569_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 20700 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1570_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1571_
timestamp 1688980957
transform -1 0 23736 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1572_
timestamp 1688980957
transform 1 0 20608 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1573_
timestamp 1688980957
transform 1 0 21804 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1574_
timestamp 1688980957
transform -1 0 23460 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_1  _1575_
timestamp 1688980957
transform -1 0 23276 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1576_
timestamp 1688980957
transform 1 0 20792 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1577_
timestamp 1688980957
transform 1 0 20700 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_4  _1578_
timestamp 1688980957
transform 1 0 21804 0 -1 28288
box -38 -48 1326 592
use sky130_fd_sc_hd__nand2_2  _1579_
timestamp 1688980957
transform 1 0 26404 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1580_
timestamp 1688980957
transform -1 0 24380 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1581_
timestamp 1688980957
transform -1 0 25024 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1582_
timestamp 1688980957
transform 1 0 23460 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1583_
timestamp 1688980957
transform 1 0 22724 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1584_
timestamp 1688980957
transform 1 0 23184 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a2111o_1  _1585_
timestamp 1688980957
transform -1 0 24564 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__a21o_1  _1586_
timestamp 1688980957
transform 1 0 23368 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1587_
timestamp 1688980957
transform 1 0 19044 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1588_
timestamp 1688980957
transform -1 0 20148 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1589_
timestamp 1688980957
transform 1 0 20148 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1590_
timestamp 1688980957
transform -1 0 20148 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1591_
timestamp 1688980957
transform 1 0 22816 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1592_
timestamp 1688980957
transform 1 0 28704 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1593_
timestamp 1688980957
transform 1 0 28796 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1594_
timestamp 1688980957
transform 1 0 31832 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o311a_1  _1595_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 30268 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1596_
timestamp 1688980957
transform -1 0 24196 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__and4_1  _1597_
timestamp 1688980957
transform 1 0 20792 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1598_
timestamp 1688980957
transform 1 0 21896 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1599_
timestamp 1688980957
transform 1 0 22816 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_1  _1600_
timestamp 1688980957
transform -1 0 24012 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1601_
timestamp 1688980957
transform 1 0 23184 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1602_
timestamp 1688980957
transform 1 0 23368 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_2  _1603_
timestamp 1688980957
transform -1 0 24196 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_4  _1604_
timestamp 1688980957
transform 1 0 24380 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__or3_1  _1605_
timestamp 1688980957
transform -1 0 24840 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1606_
timestamp 1688980957
transform 1 0 23644 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1607_
timestamp 1688980957
transform 1 0 23276 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1608_
timestamp 1688980957
transform 1 0 24012 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1609_
timestamp 1688980957
transform 1 0 23368 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1610_
timestamp 1688980957
transform 1 0 23552 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1611_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 24472 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1612_
timestamp 1688980957
transform 1 0 23552 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1613_
timestamp 1688980957
transform 1 0 20976 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1614_
timestamp 1688980957
transform 1 0 21896 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_1  _1615_
timestamp 1688980957
transform -1 0 23184 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_2  _1616_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 24012 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_4  _1617_
timestamp 1688980957
transform 1 0 24104 0 -1 16320
box -38 -48 2062 592
use sky130_fd_sc_hd__a22oi_1  _1618_
timestamp 1688980957
transform -1 0 14812 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__and4_1  _1619_
timestamp 1688980957
transform 1 0 13340 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_1  _1620_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14260 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a221oi_1  _1621_
timestamp 1688980957
transform 1 0 15272 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1622_
timestamp 1688980957
transform 1 0 13248 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1623_
timestamp 1688980957
transform 1 0 13524 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1624_
timestamp 1688980957
transform -1 0 13432 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1625_
timestamp 1688980957
transform 1 0 11224 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_2  _1626_
timestamp 1688980957
transform 1 0 11868 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_2  _1627_
timestamp 1688980957
transform 1 0 26128 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1628_
timestamp 1688980957
transform -1 0 19136 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1629_
timestamp 1688980957
transform -1 0 18768 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1630_
timestamp 1688980957
transform 1 0 15916 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1631_
timestamp 1688980957
transform 1 0 16652 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1632_
timestamp 1688980957
transform 1 0 17204 0 -1 38080
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1633_
timestamp 1688980957
transform 1 0 17480 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _1634_
timestamp 1688980957
transform 1 0 17756 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1635_
timestamp 1688980957
transform 1 0 18308 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1636_
timestamp 1688980957
transform 1 0 15916 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1637_
timestamp 1688980957
transform 1 0 16744 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1638_
timestamp 1688980957
transform 1 0 18216 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_4  _1639_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 19136 0 1 16320
box -38 -48 1602 592
use sky130_fd_sc_hd__xnor2_2  _1640_
timestamp 1688980957
transform 1 0 29532 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _1641_
timestamp 1688980957
transform -1 0 30636 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1642_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 31372 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1643_
timestamp 1688980957
transform 1 0 25944 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1644_
timestamp 1688980957
transform 1 0 26036 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o31a_1  _1645_
timestamp 1688980957
transform -1 0 27600 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _1646_
timestamp 1688980957
transform 1 0 30176 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _1647_
timestamp 1688980957
transform -1 0 30636 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1648_
timestamp 1688980957
transform -1 0 33212 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1649_
timestamp 1688980957
transform 1 0 31188 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1650_
timestamp 1688980957
transform -1 0 31648 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1651_
timestamp 1688980957
transform -1 0 33028 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1652_
timestamp 1688980957
transform 1 0 37260 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1653_
timestamp 1688980957
transform 1 0 36064 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1654_
timestamp 1688980957
transform 1 0 35420 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1655_
timestamp 1688980957
transform 1 0 34684 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1656_
timestamp 1688980957
transform 1 0 36156 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1657_
timestamp 1688980957
transform 1 0 35144 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1658_
timestamp 1688980957
transform 1 0 29532 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1659_
timestamp 1688980957
transform -1 0 32016 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1660_
timestamp 1688980957
transform -1 0 32844 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1661_
timestamp 1688980957
transform -1 0 26588 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1662_
timestamp 1688980957
transform -1 0 26680 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1663_
timestamp 1688980957
transform -1 0 27692 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1664_
timestamp 1688980957
transform 1 0 27692 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1665_
timestamp 1688980957
transform 1 0 33028 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1666_
timestamp 1688980957
transform 1 0 33580 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1667_
timestamp 1688980957
transform -1 0 34132 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1668_
timestamp 1688980957
transform 1 0 34132 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1669_
timestamp 1688980957
transform 1 0 30360 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1670_
timestamp 1688980957
transform 1 0 31096 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_2  _1671_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 31096 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1672_
timestamp 1688980957
transform -1 0 26404 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1673_
timestamp 1688980957
transform -1 0 26128 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1674_
timestamp 1688980957
transform -1 0 26864 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1675_
timestamp 1688980957
transform 1 0 27048 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1676_
timestamp 1688980957
transform -1 0 31648 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1677_
timestamp 1688980957
transform 1 0 32108 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1678_
timestamp 1688980957
transform 1 0 32200 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1679_
timestamp 1688980957
transform 1 0 32844 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1680_
timestamp 1688980957
transform -1 0 33580 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1681_
timestamp 1688980957
transform 1 0 32568 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _1682_
timestamp 1688980957
transform 1 0 32200 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1683_
timestamp 1688980957
transform -1 0 31004 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1684_
timestamp 1688980957
transform 1 0 29624 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1685_
timestamp 1688980957
transform 1 0 30360 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1686_
timestamp 1688980957
transform 1 0 29532 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1687_
timestamp 1688980957
transform 1 0 25484 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1688_
timestamp 1688980957
transform 1 0 25484 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1689_
timestamp 1688980957
transform -1 0 26036 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1690_
timestamp 1688980957
transform 1 0 25760 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1691_
timestamp 1688980957
transform 1 0 28980 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1692_
timestamp 1688980957
transform 1 0 28888 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1693_
timestamp 1688980957
transform 1 0 29716 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1694_
timestamp 1688980957
transform 1 0 29992 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1695_
timestamp 1688980957
transform 1 0 30176 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1696_
timestamp 1688980957
transform 1 0 20332 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a221o_1  _1697_
timestamp 1688980957
transform 1 0 19596 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1698_
timestamp 1688980957
transform 1 0 20332 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1699_
timestamp 1688980957
transform 1 0 20240 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_4  _1700_
timestamp 1688980957
transform 1 0 20976 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__and3b_2  _1701_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19228 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1702_
timestamp 1688980957
transform -1 0 20608 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1703_
timestamp 1688980957
transform 1 0 19688 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_4  _1704_
timestamp 1688980957
transform 1 0 19688 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__o211ai_4  _1705_
timestamp 1688980957
transform 1 0 20148 0 1 14144
box -38 -48 1602 592
use sky130_fd_sc_hd__nand2_8  _1706_
timestamp 1688980957
transform -1 0 23276 0 1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__nor2_2  _1707_
timestamp 1688980957
transform 1 0 27876 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__o31ai_2  _1708_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30176 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__inv_2  _1709_
timestamp 1688980957
transform 1 0 35144 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1710_
timestamp 1688980957
transform 1 0 33856 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1711_
timestamp 1688980957
transform 1 0 34684 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1712_
timestamp 1688980957
transform 1 0 32016 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1713_
timestamp 1688980957
transform -1 0 29164 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_4  _1714_
timestamp 1688980957
transform 1 0 21160 0 1 4352
box -38 -48 2062 592
use sky130_fd_sc_hd__o211a_1  _1715_
timestamp 1688980957
transform -1 0 18860 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _1716_
timestamp 1688980957
transform 1 0 20240 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _1717_
timestamp 1688980957
transform -1 0 21712 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1718_
timestamp 1688980957
transform 1 0 26404 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1719_
timestamp 1688980957
transform 1 0 25576 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _1720_
timestamp 1688980957
transform -1 0 26680 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1721_
timestamp 1688980957
transform -1 0 29440 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1722_
timestamp 1688980957
transform -1 0 29900 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1723_
timestamp 1688980957
transform 1 0 25208 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1724_
timestamp 1688980957
transform 1 0 25484 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1725_
timestamp 1688980957
transform 1 0 25208 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _1726_
timestamp 1688980957
transform 1 0 26404 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1727_
timestamp 1688980957
transform -1 0 27324 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1728_
timestamp 1688980957
transform 1 0 27692 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nand4_2  _1729_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22908 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1730_
timestamp 1688980957
transform -1 0 27968 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1731_
timestamp 1688980957
transform 1 0 26956 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1732_
timestamp 1688980957
transform -1 0 26036 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1733_
timestamp 1688980957
transform -1 0 26864 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1734_
timestamp 1688980957
transform 1 0 26220 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1735_
timestamp 1688980957
transform -1 0 25944 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a41o_1  _1736_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29256 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _1737_
timestamp 1688980957
transform 1 0 32108 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _1738_
timestamp 1688980957
transform 1 0 33304 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1739_
timestamp 1688980957
transform -1 0 34684 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1740_
timestamp 1688980957
transform 1 0 34960 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1741_
timestamp 1688980957
transform -1 0 36156 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1742_
timestamp 1688980957
transform 1 0 35512 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1743_
timestamp 1688980957
transform 1 0 31648 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1744_
timestamp 1688980957
transform -1 0 33580 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1745_
timestamp 1688980957
transform 1 0 32844 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1746_
timestamp 1688980957
transform 1 0 29716 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1747_
timestamp 1688980957
transform 1 0 29532 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1748_
timestamp 1688980957
transform 1 0 21804 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  _1749_
timestamp 1688980957
transform 1 0 22540 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _1750_
timestamp 1688980957
transform 1 0 30084 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__o22ai_4  _1751_
timestamp 1688980957
transform 1 0 30268 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2_1  _1752_
timestamp 1688980957
transform 1 0 29072 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1753_
timestamp 1688980957
transform 1 0 30544 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1754_
timestamp 1688980957
transform 1 0 31004 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1755_
timestamp 1688980957
transform 1 0 31464 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1756_
timestamp 1688980957
transform 1 0 29348 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1757_
timestamp 1688980957
transform 1 0 29900 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1758_
timestamp 1688980957
transform -1 0 33028 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1759_
timestamp 1688980957
transform -1 0 33672 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1760_
timestamp 1688980957
transform -1 0 33304 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1761_
timestamp 1688980957
transform 1 0 29532 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1762_
timestamp 1688980957
transform 1 0 31648 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1763_
timestamp 1688980957
transform 1 0 25208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1764_
timestamp 1688980957
transform 1 0 19780 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1765_
timestamp 1688980957
transform 1 0 19504 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1766_
timestamp 1688980957
transform -1 0 20332 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1767_
timestamp 1688980957
transform 1 0 19596 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1768_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 19964 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1769_
timestamp 1688980957
transform -1 0 25576 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1770_
timestamp 1688980957
transform -1 0 28980 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1771_
timestamp 1688980957
transform -1 0 27140 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1772_
timestamp 1688980957
transform 1 0 30912 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1773_
timestamp 1688980957
transform 1 0 32108 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1774_
timestamp 1688980957
transform -1 0 33396 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1775_
timestamp 1688980957
transform -1 0 32844 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _1776_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 33580 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1777_
timestamp 1688980957
transform -1 0 34132 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _1778_
timestamp 1688980957
transform -1 0 33488 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_2  _1779_
timestamp 1688980957
transform 1 0 20884 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_2  _1780_
timestamp 1688980957
transform -1 0 21436 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1781_
timestamp 1688980957
transform -1 0 29072 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1782_
timestamp 1688980957
transform -1 0 32568 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1783_
timestamp 1688980957
transform -1 0 33028 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or3_2  _1784_
timestamp 1688980957
transform 1 0 28888 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1785_
timestamp 1688980957
transform 1 0 28888 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1786_
timestamp 1688980957
transform -1 0 29348 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1787_
timestamp 1688980957
transform -1 0 29072 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1788_
timestamp 1688980957
transform 1 0 30452 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1789_
timestamp 1688980957
transform 1 0 32568 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1790_
timestamp 1688980957
transform -1 0 30176 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1791_
timestamp 1688980957
transform -1 0 32752 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1792_
timestamp 1688980957
transform 1 0 29532 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1793_
timestamp 1688980957
transform 1 0 29992 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _1794_
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _1795_
timestamp 1688980957
transform 1 0 18952 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1796_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20056 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nand3b_1  _1797_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19780 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1798_
timestamp 1688980957
transform 1 0 20792 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1799_
timestamp 1688980957
transform 1 0 21528 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1800_
timestamp 1688980957
transform 1 0 22172 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1801_
timestamp 1688980957
transform 1 0 25576 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1802_
timestamp 1688980957
transform 1 0 26956 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1803_
timestamp 1688980957
transform 1 0 28060 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_2  _1804_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 31924 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1805_
timestamp 1688980957
transform -1 0 31464 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1806_
timestamp 1688980957
transform -1 0 29808 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _1807_
timestamp 1688980957
transform -1 0 21528 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  _1808_
timestamp 1688980957
transform 1 0 22172 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__a2111oi_1  _1809_
timestamp 1688980957
transform 1 0 28060 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1810_
timestamp 1688980957
transform -1 0 28796 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1811_
timestamp 1688980957
transform 1 0 30268 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _1812_
timestamp 1688980957
transform 1 0 32108 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1813_
timestamp 1688980957
transform -1 0 30912 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1814_
timestamp 1688980957
transform 1 0 27968 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1815_
timestamp 1688980957
transform -1 0 27876 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1816_
timestamp 1688980957
transform 1 0 20424 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and2_2  _1817_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21896 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1818_
timestamp 1688980957
transform -1 0 23828 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1819_
timestamp 1688980957
transform 1 0 22448 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_2  _1820_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 20608 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1821_
timestamp 1688980957
transform -1 0 23276 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1822_
timestamp 1688980957
transform 1 0 22356 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_4  _1823_
timestamp 1688980957
transform 1 0 33028 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__a31o_1  _1824_
timestamp 1688980957
transform -1 0 23552 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_4  _1825_
timestamp 1688980957
transform 1 0 21804 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1826_
timestamp 1688980957
transform 1 0 26312 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1827_
timestamp 1688980957
transform 1 0 25392 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1828_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21068 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1829_
timestamp 1688980957
transform -1 0 21804 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1830_
timestamp 1688980957
transform 1 0 19504 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1831_
timestamp 1688980957
transform 1 0 24840 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1832_
timestamp 1688980957
transform 1 0 23460 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _1833_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25208 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1834_
timestamp 1688980957
transform 1 0 24932 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1835_
timestamp 1688980957
transform -1 0 24932 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1836_
timestamp 1688980957
transform -1 0 25392 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1837_
timestamp 1688980957
transform -1 0 27508 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1838_
timestamp 1688980957
transform -1 0 29348 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_2  _1839_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27508 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _1840_
timestamp 1688980957
transform -1 0 25024 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1841_
timestamp 1688980957
transform 1 0 25668 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1842_
timestamp 1688980957
transform -1 0 19596 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1843_
timestamp 1688980957
transform -1 0 20608 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1844_
timestamp 1688980957
transform 1 0 20148 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_2  _1845_
timestamp 1688980957
transform 1 0 20608 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1846_
timestamp 1688980957
transform -1 0 19964 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1847_
timestamp 1688980957
transform -1 0 20240 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _1848_
timestamp 1688980957
transform 1 0 20516 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_4  _1849_
timestamp 1688980957
transform 1 0 22264 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__a221o_2  _1850_
timestamp 1688980957
transform 1 0 21344 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_1  _1851_
timestamp 1688980957
transform -1 0 14812 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1852_
timestamp 1688980957
transform -1 0 16560 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1853_
timestamp 1688980957
transform 1 0 14812 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1854_
timestamp 1688980957
transform 1 0 16744 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1855_
timestamp 1688980957
transform -1 0 16376 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _1856_
timestamp 1688980957
transform 1 0 15456 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or3b_1  _1857_
timestamp 1688980957
transform 1 0 14168 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _1858_
timestamp 1688980957
transform 1 0 15640 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o21bai_4  _1859_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22908 0 1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__nor2_4  _1860_
timestamp 1688980957
transform -1 0 25576 0 1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1861_
timestamp 1688980957
transform -1 0 33856 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1862_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 34132 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _1863_
timestamp 1688980957
transform -1 0 33212 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _1864_
timestamp 1688980957
transform -1 0 33212 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_2  _1865_
timestamp 1688980957
transform 1 0 28152 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1866_
timestamp 1688980957
transform 1 0 32108 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1867_
timestamp 1688980957
transform 1 0 31464 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1868_
timestamp 1688980957
transform 1 0 24380 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1869_
timestamp 1688980957
transform 1 0 30176 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1870_
timestamp 1688980957
transform 1 0 30636 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_4  _1871_
timestamp 1688980957
transform 1 0 23552 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_2  _1872_
timestamp 1688980957
transform 1 0 23276 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1873_
timestamp 1688980957
transform 1 0 26036 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1874_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25944 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1875_
timestamp 1688980957
transform -1 0 26956 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _1876_
timestamp 1688980957
transform -1 0 27508 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1877_
timestamp 1688980957
transform 1 0 30176 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _1878_
timestamp 1688980957
transform -1 0 32016 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1879_
timestamp 1688980957
transform -1 0 31464 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1880_
timestamp 1688980957
transform 1 0 30728 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_2  _1881_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 30728 0 1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _1882_
timestamp 1688980957
transform -1 0 27876 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1883_
timestamp 1688980957
transform -1 0 27416 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1884_
timestamp 1688980957
transform 1 0 26588 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1885_
timestamp 1688980957
transform -1 0 26864 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1886_
timestamp 1688980957
transform 1 0 31464 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _1887_
timestamp 1688980957
transform 1 0 31096 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1888_
timestamp 1688980957
transform 1 0 32384 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1889_
timestamp 1688980957
transform 1 0 25392 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _1890_
timestamp 1688980957
transform 1 0 26864 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _1891_
timestamp 1688980957
transform -1 0 26864 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _1892_
timestamp 1688980957
transform -1 0 27692 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1893_
timestamp 1688980957
transform 1 0 30084 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__or2_1  _1894_
timestamp 1688980957
transform 1 0 32844 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1895_
timestamp 1688980957
transform -1 0 28704 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _1896_
timestamp 1688980957
transform -1 0 33028 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1897_
timestamp 1688980957
transform 1 0 32384 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_4  _1898_
timestamp 1688980957
transform -1 0 32016 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _1899_
timestamp 1688980957
transform 1 0 33120 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1900_
timestamp 1688980957
transform -1 0 33764 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1901_
timestamp 1688980957
transform -1 0 32384 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1902_
timestamp 1688980957
transform 1 0 32292 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _1903_
timestamp 1688980957
transform -1 0 32200 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1904_
timestamp 1688980957
transform 1 0 32476 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1905_
timestamp 1688980957
transform 1 0 32476 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1906_
timestamp 1688980957
transform 1 0 27968 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1907_
timestamp 1688980957
transform 1 0 30084 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1908_
timestamp 1688980957
transform -1 0 29900 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_1  _1909_
timestamp 1688980957
transform 1 0 30912 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1910_
timestamp 1688980957
transform 1 0 30268 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1911_
timestamp 1688980957
transform -1 0 30360 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1912_
timestamp 1688980957
transform 1 0 30084 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1913_
timestamp 1688980957
transform 1 0 23828 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1914_
timestamp 1688980957
transform -1 0 23828 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1915_
timestamp 1688980957
transform 1 0 21528 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1916_
timestamp 1688980957
transform -1 0 24380 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1917_
timestamp 1688980957
transform 1 0 25944 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1918_
timestamp 1688980957
transform 1 0 27600 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o221a_1  _1919_
timestamp 1688980957
transform 1 0 26772 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1920_
timestamp 1688980957
transform 1 0 24380 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1921_
timestamp 1688980957
transform -1 0 27692 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__o211a_1  _1922_
timestamp 1688980957
transform -1 0 28888 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o221ai_2  _1923_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 29900 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__o211a_1  _1924_
timestamp 1688980957
transform 1 0 31464 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__a211o_4  _1925_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30728 0 -1 7616
box -38 -48 1326 592
use sky130_fd_sc_hd__mux2_1  _1926_
timestamp 1688980957
transform 1 0 34684 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1927_
timestamp 1688980957
transform -1 0 34040 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1928_
timestamp 1688980957
transform 1 0 33028 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1929_
timestamp 1688980957
transform 1 0 28612 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1930_
timestamp 1688980957
transform 1 0 34224 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1931_
timestamp 1688980957
transform -1 0 34592 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1932_
timestamp 1688980957
transform 1 0 26128 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1933_
timestamp 1688980957
transform 1 0 27140 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1934_
timestamp 1688980957
transform -1 0 27968 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _1935_
timestamp 1688980957
transform -1 0 28060 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1936_
timestamp 1688980957
transform -1 0 28060 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1937_
timestamp 1688980957
transform 1 0 27600 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__o22a_1  _1938_
timestamp 1688980957
transform -1 0 25852 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _1939_
timestamp 1688980957
transform -1 0 26588 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o221a_1  _1940_
timestamp 1688980957
transform 1 0 26956 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_1  _1941_
timestamp 1688980957
transform 1 0 26956 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a221o_1  _1942_
timestamp 1688980957
transform 1 0 27508 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1943_
timestamp 1688980957
transform -1 0 27876 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _1944_
timestamp 1688980957
transform 1 0 27876 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_2  _1945_
timestamp 1688980957
transform -1 0 28888 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _1946_
timestamp 1688980957
transform -1 0 36800 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _1947_
timestamp 1688980957
transform 1 0 35420 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _1948_
timestamp 1688980957
transform -1 0 35696 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_2  _1949_
timestamp 1688980957
transform -1 0 35420 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _1950_
timestamp 1688980957
transform 1 0 27232 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1951_
timestamp 1688980957
transform -1 0 34592 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1952_
timestamp 1688980957
transform -1 0 34868 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1953_
timestamp 1688980957
transform 1 0 22356 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1954_
timestamp 1688980957
transform 1 0 23000 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1955_
timestamp 1688980957
transform -1 0 23552 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _1956_
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _1957_
timestamp 1688980957
transform 1 0 19964 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1958_
timestamp 1688980957
transform 1 0 20884 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1959_
timestamp 1688980957
transform 1 0 25392 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1960_
timestamp 1688980957
transform -1 0 19044 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1961_
timestamp 1688980957
transform 1 0 24380 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _1962_
timestamp 1688980957
transform 1 0 25392 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1963_
timestamp 1688980957
transform -1 0 25392 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__or4b_1  _1964_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 25668 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _1965_
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _1966_
timestamp 1688980957
transform 1 0 23368 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__o2bb2a_4  _1967_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 23920 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__nand2_1  _1968_
timestamp 1688980957
transform 1 0 35788 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1969_
timestamp 1688980957
transform 1 0 35512 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _1970_
timestamp 1688980957
transform 1 0 36340 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_2  _1971_
timestamp 1688980957
transform 1 0 34776 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1972_
timestamp 1688980957
transform -1 0 25760 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1973_
timestamp 1688980957
transform 1 0 24840 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1974_
timestamp 1688980957
transform -1 0 34868 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1975_
timestamp 1688980957
transform -1 0 34960 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1976_
timestamp 1688980957
transform 1 0 20608 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1977_
timestamp 1688980957
transform 1 0 21896 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1978_
timestamp 1688980957
transform 1 0 19688 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1979_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19872 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o22a_1  _1980_
timestamp 1688980957
transform -1 0 22448 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1981_
timestamp 1688980957
transform 1 0 19688 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1982_
timestamp 1688980957
transform 1 0 20056 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _1983_
timestamp 1688980957
transform -1 0 22908 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1984_
timestamp 1688980957
transform 1 0 22908 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _1985_
timestamp 1688980957
transform 1 0 23000 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__o211ai_1  _1986_
timestamp 1688980957
transform 1 0 21804 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a221o_1  _1987_
timestamp 1688980957
transform 1 0 22540 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_4  _1988_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 22356 0 1 7616
box -38 -48 1326 592
use sky130_fd_sc_hd__a21oi_1  _1989_
timestamp 1688980957
transform -1 0 33212 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _1990_
timestamp 1688980957
transform -1 0 34776 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _1991_
timestamp 1688980957
transform 1 0 34684 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_2  _1992_
timestamp 1688980957
transform -1 0 35420 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1993_
timestamp 1688980957
transform -1 0 33764 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1994_
timestamp 1688980957
transform 1 0 27232 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _1995_
timestamp 1688980957
transform -1 0 34684 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1996_
timestamp 1688980957
transform -1 0 34960 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1997_
timestamp 1688980957
transform -1 0 21712 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1998_
timestamp 1688980957
transform -1 0 20884 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1999_
timestamp 1688980957
transform -1 0 20516 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2000_
timestamp 1688980957
transform 1 0 21620 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_1  _2001_
timestamp 1688980957
transform 1 0 20884 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _2002_
timestamp 1688980957
transform 1 0 22724 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _2003_
timestamp 1688980957
transform 1 0 22448 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _2004_
timestamp 1688980957
transform 1 0 21988 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2005_
timestamp 1688980957
transform 1 0 24564 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2006_
timestamp 1688980957
transform 1 0 21344 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _2007_
timestamp 1688980957
transform 1 0 22264 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_2  _2008_
timestamp 1688980957
transform 1 0 21804 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2009_
timestamp 1688980957
transform -1 0 30544 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2010_
timestamp 1688980957
transform -1 0 32568 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2011_
timestamp 1688980957
transform 1 0 31648 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _2012_
timestamp 1688980957
transform -1 0 32844 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _2013_
timestamp 1688980957
transform 1 0 32844 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2014_
timestamp 1688980957
transform -1 0 27048 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2015_
timestamp 1688980957
transform -1 0 29164 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2016_
timestamp 1688980957
transform -1 0 28888 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _2017_
timestamp 1688980957
transform 1 0 23092 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _2018_
timestamp 1688980957
transform 1 0 27600 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2019_
timestamp 1688980957
transform 1 0 29164 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2020_
timestamp 1688980957
transform -1 0 29072 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2021_
timestamp 1688980957
transform 1 0 27324 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2022_
timestamp 1688980957
transform -1 0 26864 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2023_
timestamp 1688980957
transform 1 0 28060 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2024_
timestamp 1688980957
transform 1 0 28060 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2025_
timestamp 1688980957
transform 1 0 29532 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2026_
timestamp 1688980957
transform -1 0 29348 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2027_
timestamp 1688980957
transform -1 0 28336 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2028_
timestamp 1688980957
transform 1 0 28336 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2029_
timestamp 1688980957
transform -1 0 30360 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2030_
timestamp 1688980957
transform 1 0 29808 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2031_
timestamp 1688980957
transform 1 0 28428 0 1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2032_
timestamp 1688980957
transform -1 0 28152 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2033_
timestamp 1688980957
transform 1 0 27784 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2034_
timestamp 1688980957
transform 1 0 27968 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _2035_
timestamp 1688980957
transform -1 0 13984 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_4  _2036_
timestamp 1688980957
transform -1 0 14904 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__and4_2  _2037_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13248 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_2  _2038_
timestamp 1688980957
transform 1 0 14904 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _2039_
timestamp 1688980957
transform 1 0 24288 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2040_
timestamp 1688980957
transform -1 0 23092 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2041_
timestamp 1688980957
transform 1 0 21988 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _2042_
timestamp 1688980957
transform -1 0 22632 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _2043_
timestamp 1688980957
transform 1 0 22172 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_4  _2044_
timestamp 1688980957
transform 1 0 22632 0 -1 23936
box -38 -48 1326 592
use sky130_fd_sc_hd__mux2_1  _2045_
timestamp 1688980957
transform 1 0 19412 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2046_
timestamp 1688980957
transform -1 0 19688 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2047_
timestamp 1688980957
transform 1 0 9568 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2048_
timestamp 1688980957
transform 1 0 10212 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2049_
timestamp 1688980957
transform 1 0 9752 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2050_
timestamp 1688980957
transform -1 0 9752 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2051_
timestamp 1688980957
transform -1 0 10212 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2052_
timestamp 1688980957
transform 1 0 9660 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2053_
timestamp 1688980957
transform -1 0 10396 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2054_
timestamp 1688980957
transform 1 0 8740 0 -1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2055_
timestamp 1688980957
transform -1 0 8556 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2056_
timestamp 1688980957
transform 1 0 9200 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2057_
timestamp 1688980957
transform 1 0 10120 0 -1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2058_
timestamp 1688980957
transform 1 0 9844 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2059_
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2060_
timestamp 1688980957
transform 1 0 11500 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2061_
timestamp 1688980957
transform 1 0 10580 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2062_
timestamp 1688980957
transform 1 0 8740 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2063_
timestamp 1688980957
transform 1 0 9476 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2064_
timestamp 1688980957
transform 1 0 9568 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2065_
timestamp 1688980957
transform 1 0 9844 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2066_
timestamp 1688980957
transform 1 0 11960 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2067_
timestamp 1688980957
transform 1 0 10580 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2068_
timestamp 1688980957
transform -1 0 24012 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _2069_
timestamp 1688980957
transform -1 0 26312 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _2070_
timestamp 1688980957
transform 1 0 22540 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_4  _2071_
timestamp 1688980957
transform -1 0 25392 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2072_
timestamp 1688980957
transform -1 0 31372 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2073_
timestamp 1688980957
transform 1 0 31004 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2074_
timestamp 1688980957
transform 1 0 26036 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2075_
timestamp 1688980957
transform 1 0 26220 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2076_
timestamp 1688980957
transform -1 0 28980 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2077_
timestamp 1688980957
transform 1 0 28980 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2078_
timestamp 1688980957
transform -1 0 33028 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2079_
timestamp 1688980957
transform 1 0 32844 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2080_
timestamp 1688980957
transform -1 0 33856 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2081_
timestamp 1688980957
transform -1 0 34132 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2082_
timestamp 1688980957
transform 1 0 33212 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2083_
timestamp 1688980957
transform -1 0 33396 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2084_
timestamp 1688980957
transform -1 0 33764 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2085_
timestamp 1688980957
transform 1 0 33304 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2086_
timestamp 1688980957
transform -1 0 26864 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2087_
timestamp 1688980957
transform 1 0 26956 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _2088_
timestamp 1688980957
transform 1 0 23276 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  _2089_
timestamp 1688980957
transform 1 0 21988 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2090_
timestamp 1688980957
transform -1 0 21528 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2091_
timestamp 1688980957
transform -1 0 12328 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2092_
timestamp 1688980957
transform -1 0 12328 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2093_
timestamp 1688980957
transform 1 0 5428 0 -1 33728
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2094_
timestamp 1688980957
transform 1 0 5428 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2095_
timestamp 1688980957
transform 1 0 6348 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2096_
timestamp 1688980957
transform 1 0 4600 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2097_
timestamp 1688980957
transform 1 0 7820 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2098_
timestamp 1688980957
transform 1 0 6440 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2099_
timestamp 1688980957
transform 1 0 11592 0 1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2100_
timestamp 1688980957
transform 1 0 10212 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2101_
timestamp 1688980957
transform 1 0 7268 0 -1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2102_
timestamp 1688980957
transform 1 0 6532 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2103_
timestamp 1688980957
transform 1 0 9292 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2104_
timestamp 1688980957
transform 1 0 9016 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _2105_
timestamp 1688980957
transform -1 0 24288 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__o21ai_4  _2106_
timestamp 1688980957
transform 1 0 23092 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  _2107_
timestamp 1688980957
transform 1 0 32568 0 1 35904
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2108_
timestamp 1688980957
transform -1 0 32292 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2109_
timestamp 1688980957
transform -1 0 28152 0 1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2110_
timestamp 1688980957
transform 1 0 28152 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2111_
timestamp 1688980957
transform -1 0 31280 0 -1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2112_
timestamp 1688980957
transform -1 0 31188 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2113_
timestamp 1688980957
transform -1 0 34592 0 1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2114_
timestamp 1688980957
transform -1 0 34500 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2115_
timestamp 1688980957
transform -1 0 35512 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2116_
timestamp 1688980957
transform 1 0 35236 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2117_
timestamp 1688980957
transform 1 0 32108 0 -1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2118_
timestamp 1688980957
transform 1 0 31464 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2119_
timestamp 1688980957
transform 1 0 31188 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2120_
timestamp 1688980957
transform 1 0 31188 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2121_
timestamp 1688980957
transform 1 0 26956 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2122_
timestamp 1688980957
transform 1 0 25944 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_8  _2123_
timestamp 1688980957
transform -1 0 23092 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _2124_
timestamp 1688980957
transform 1 0 22356 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2125_
timestamp 1688980957
transform 1 0 20884 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2126_
timestamp 1688980957
transform 1 0 9292 0 -1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2127_
timestamp 1688980957
transform -1 0 8556 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2128_
timestamp 1688980957
transform 1 0 6256 0 1 32640
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2129_
timestamp 1688980957
transform 1 0 4968 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2130_
timestamp 1688980957
transform 1 0 5428 0 1 29376
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2131_
timestamp 1688980957
transform 1 0 4508 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2132_
timestamp 1688980957
transform 1 0 8924 0 1 30464
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2133_
timestamp 1688980957
transform 1 0 8280 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2134_
timestamp 1688980957
transform 1 0 9568 0 -1 28288
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2135_
timestamp 1688980957
transform 1 0 8280 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2136_
timestamp 1688980957
transform 1 0 7912 0 -1 34816
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2137_
timestamp 1688980957
transform 1 0 7636 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2138_
timestamp 1688980957
transform 1 0 9200 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2139_
timestamp 1688980957
transform 1 0 7912 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2140_
timestamp 1688980957
transform -1 0 24656 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2141_
timestamp 1688980957
transform 1 0 24012 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2142_
timestamp 1688980957
transform 1 0 11500 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _2143_
timestamp 1688980957
transform 1 0 18308 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2144_
timestamp 1688980957
transform -1 0 18308 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2145_
timestamp 1688980957
transform 1 0 17664 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _2146_
timestamp 1688980957
transform 1 0 17480 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a2bb2o_1  _2147_
timestamp 1688980957
transform 1 0 15272 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a211oi_4  _2148_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 25760 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__a31o_2  _2149_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12236 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2150_
timestamp 1688980957
transform 1 0 6900 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2151_
timestamp 1688980957
transform 1 0 5428 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2152_
timestamp 1688980957
transform 1 0 8556 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or4_1  _2153_
timestamp 1688980957
transform -1 0 25392 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _2154_
timestamp 1688980957
transform 1 0 24104 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _2155_
timestamp 1688980957
transform 1 0 23828 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _2156_
timestamp 1688980957
transform 1 0 22172 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_1  _2157_
timestamp 1688980957
transform 1 0 22816 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__or4_2  _2158_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 24012 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2159_
timestamp 1688980957
transform -1 0 10488 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2160_
timestamp 1688980957
transform 1 0 9476 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _2161_
timestamp 1688980957
transform -1 0 9936 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2162_
timestamp 1688980957
transform -1 0 7912 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2163_
timestamp 1688980957
transform -1 0 7360 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2164_
timestamp 1688980957
transform -1 0 8096 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _2165_
timestamp 1688980957
transform 1 0 31740 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_2  _2166_
timestamp 1688980957
transform 1 0 29440 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2167_
timestamp 1688980957
transform -1 0 30360 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _2168_
timestamp 1688980957
transform 1 0 29992 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _2169_
timestamp 1688980957
transform 1 0 23184 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2170_
timestamp 1688980957
transform 1 0 24104 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2171_
timestamp 1688980957
transform 1 0 23828 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _2172_
timestamp 1688980957
transform 1 0 24104 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2173_
timestamp 1688980957
transform 1 0 24748 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2174_
timestamp 1688980957
transform 1 0 33028 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _2175_
timestamp 1688980957
transform 1 0 33488 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_1  _2176_
timestamp 1688980957
transform 1 0 33488 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2177_
timestamp 1688980957
transform -1 0 24656 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2178_
timestamp 1688980957
transform 1 0 33856 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2179_
timestamp 1688980957
transform 1 0 34500 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2180_
timestamp 1688980957
transform -1 0 35972 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2181_
timestamp 1688980957
transform 1 0 32936 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2182_
timestamp 1688980957
transform -1 0 34132 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2183_
timestamp 1688980957
transform 1 0 33764 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _2184_
timestamp 1688980957
transform 1 0 34408 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2185_
timestamp 1688980957
transform 1 0 34868 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o221a_1  _2186_
timestamp 1688980957
transform 1 0 28244 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _2187_
timestamp 1688980957
transform 1 0 30912 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o221a_1  _2188_
timestamp 1688980957
transform 1 0 31188 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2189_
timestamp 1688980957
transform 1 0 32844 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2190_
timestamp 1688980957
transform 1 0 33764 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2191_
timestamp 1688980957
transform 1 0 34684 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2192_
timestamp 1688980957
transform -1 0 35236 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2193_
timestamp 1688980957
transform 1 0 34960 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _2194_
timestamp 1688980957
transform 1 0 35420 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2195_
timestamp 1688980957
transform -1 0 34592 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o221ai_4  _2196_
timestamp 1688980957
transform 1 0 28152 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__a21oi_1  _2197_
timestamp 1688980957
transform -1 0 28336 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2198_
timestamp 1688980957
transform -1 0 28796 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _2199_
timestamp 1688980957
transform 1 0 22172 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2200_
timestamp 1688980957
transform 1 0 23368 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _2201_
timestamp 1688980957
transform 1 0 24380 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2202_
timestamp 1688980957
transform 1 0 25024 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2203_
timestamp 1688980957
transform 1 0 25668 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2204_
timestamp 1688980957
transform 1 0 26036 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2205_
timestamp 1688980957
transform 1 0 26864 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2206_
timestamp 1688980957
transform 1 0 27968 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o31ai_4  _2207_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 29256 0 1 17408
box -38 -48 1602 592
use sky130_fd_sc_hd__mux2_1  _2208_
timestamp 1688980957
transform 1 0 9384 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2209_
timestamp 1688980957
transform 1 0 8004 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2210_
timestamp 1688980957
transform 1 0 7728 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2211_
timestamp 1688980957
transform -1 0 8556 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _2212_
timestamp 1688980957
transform 1 0 7636 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2213_
timestamp 1688980957
transform 1 0 30452 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2214_
timestamp 1688980957
transform -1 0 30268 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2215_
timestamp 1688980957
transform 1 0 29072 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__o21ai_1  _2216_
timestamp 1688980957
transform 1 0 23460 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _2217_
timestamp 1688980957
transform -1 0 23460 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2218_
timestamp 1688980957
transform -1 0 24564 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o2111a_1  _2219_
timestamp 1688980957
transform 1 0 29532 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _2220_
timestamp 1688980957
transform -1 0 30268 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _2221_
timestamp 1688980957
transform -1 0 28980 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2222_
timestamp 1688980957
transform 1 0 28428 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _2223_
timestamp 1688980957
transform 1 0 29532 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__o311a_1  _2224_
timestamp 1688980957
transform -1 0 29716 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_2  _2225_
timestamp 1688980957
transform 1 0 28980 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2226_
timestamp 1688980957
transform -1 0 12236 0 1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2227_
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2228_
timestamp 1688980957
transform 1 0 11040 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2229_
timestamp 1688980957
transform 1 0 12328 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _2230_
timestamp 1688980957
transform -1 0 12328 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__or3b_1  _2231_
timestamp 1688980957
transform -1 0 12972 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _2232_
timestamp 1688980957
transform 1 0 12236 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2233_
timestamp 1688980957
transform -1 0 9936 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2234_
timestamp 1688980957
transform -1 0 15088 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _2235_
timestamp 1688980957
transform -1 0 16928 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_2  _2236_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 15548 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__or3_4  _2237_
timestamp 1688980957
transform -1 0 14628 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__nor3_1  _2238_
timestamp 1688980957
transform 1 0 9016 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2239_
timestamp 1688980957
transform -1 0 10120 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _2240_
timestamp 1688980957
transform 1 0 9384 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2241_
timestamp 1688980957
transform -1 0 10304 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_2  _2242_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 13248 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _2243_
timestamp 1688980957
transform -1 0 13616 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2244_
timestamp 1688980957
transform 1 0 8464 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _2245_
timestamp 1688980957
transform 1 0 8372 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2246_
timestamp 1688980957
transform -1 0 8832 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2247_
timestamp 1688980957
transform 1 0 8924 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _2248_
timestamp 1688980957
transform -1 0 9660 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2249_
timestamp 1688980957
transform -1 0 9108 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _2250_
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2251_
timestamp 1688980957
transform 1 0 7912 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _2252_
timestamp 1688980957
transform -1 0 8740 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _2253_
timestamp 1688980957
transform -1 0 8648 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2254_
timestamp 1688980957
transform -1 0 10396 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a211o_1  _2255_
timestamp 1688980957
transform -1 0 8004 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2256_
timestamp 1688980957
transform -1 0 9752 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_2  _2257_
timestamp 1688980957
transform 1 0 7452 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__and4bb_1  _2258_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8924 0 -1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__o21ai_1  _2259_
timestamp 1688980957
transform 1 0 7452 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _2260_
timestamp 1688980957
transform -1 0 10212 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2261_
timestamp 1688980957
transform 1 0 8280 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and4b_1  _2262_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7820 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _2263_
timestamp 1688980957
transform -1 0 9568 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2264_
timestamp 1688980957
transform -1 0 9200 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _2265_
timestamp 1688980957
transform 1 0 10120 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2266_
timestamp 1688980957
transform -1 0 14352 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2267_
timestamp 1688980957
transform -1 0 14628 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__buf_6  _2268_
timestamp 1688980957
transform 1 0 14352 0 -1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__inv_6  _2269_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7728 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2270_
timestamp 1688980957
transform 1 0 13432 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2271_
timestamp 1688980957
transform 1 0 15548 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2272_
timestamp 1688980957
transform 1 0 15364 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2273_
timestamp 1688980957
transform 1 0 16008 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__buf_6  _2274_
timestamp 1688980957
transform 1 0 16652 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2275_
timestamp 1688980957
transform -1 0 15548 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2276_
timestamp 1688980957
transform 1 0 14904 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2277_
timestamp 1688980957
transform 1 0 35604 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2278_
timestamp 1688980957
transform -1 0 36984 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2279_
timestamp 1688980957
transform 1 0 36708 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__buf_1  _2280_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 36892 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2281_
timestamp 1688980957
transform -1 0 12972 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2282_
timestamp 1688980957
transform -1 0 8832 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2283_
timestamp 1688980957
transform -1 0 13064 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2284_
timestamp 1688980957
transform 1 0 12328 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2285_
timestamp 1688980957
transform -1 0 13340 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2286_
timestamp 1688980957
transform 1 0 12972 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2287_
timestamp 1688980957
transform -1 0 13156 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2288_
timestamp 1688980957
transform 1 0 1748 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2289_
timestamp 1688980957
transform 1 0 36616 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2290_
timestamp 1688980957
transform -1 0 37628 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__a21boi_4  _2291_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 14352 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__and2_1  _2292_
timestamp 1688980957
transform 1 0 1656 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2293_
timestamp 1688980957
transform 1 0 2024 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2294_
timestamp 1688980957
transform 1 0 10488 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2295_
timestamp 1688980957
transform -1 0 12972 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _2296_
timestamp 1688980957
transform -1 0 14812 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2297_
timestamp 1688980957
transform 1 0 5796 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2298_
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2299_
timestamp 1688980957
transform -1 0 5060 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2300_
timestamp 1688980957
transform 1 0 3864 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2301_
timestamp 1688980957
transform 1 0 7176 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2302_
timestamp 1688980957
transform -1 0 17572 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2303_
timestamp 1688980957
transform 1 0 2760 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2304_
timestamp 1688980957
transform 1 0 2944 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2305_
timestamp 1688980957
transform 1 0 3864 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2306_
timestamp 1688980957
transform -1 0 9660 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2307_
timestamp 1688980957
transform 1 0 3036 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2308_
timestamp 1688980957
transform 1 0 2944 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2309_
timestamp 1688980957
transform 1 0 5704 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2310_
timestamp 1688980957
transform -1 0 23000 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2311_
timestamp 1688980957
transform 1 0 17388 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2312_
timestamp 1688980957
transform -1 0 17664 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2313_
timestamp 1688980957
transform -1 0 17480 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2314_
timestamp 1688980957
transform 1 0 2668 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2315_
timestamp 1688980957
transform 1 0 1564 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2316_
timestamp 1688980957
transform 1 0 1748 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2317_
timestamp 1688980957
transform 1 0 2760 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _2318_
timestamp 1688980957
transform 1 0 2208 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2319_
timestamp 1688980957
transform 1 0 5244 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2320_
timestamp 1688980957
transform -1 0 22908 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2321_
timestamp 1688980957
transform 1 0 7820 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2322_
timestamp 1688980957
transform -1 0 25392 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2323_
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2324_
timestamp 1688980957
transform -1 0 13064 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2325_
timestamp 1688980957
transform 1 0 4968 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _2326_
timestamp 1688980957
transform 1 0 5428 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_1  _2327_
timestamp 1688980957
transform -1 0 6348 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _2328_
timestamp 1688980957
transform 1 0 2116 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2329_
timestamp 1688980957
transform 1 0 2208 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _2330_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 27416 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _2331_
timestamp 1688980957
transform 1 0 27692 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2332_
timestamp 1688980957
transform -1 0 25300 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2333_
timestamp 1688980957
transform 1 0 18308 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2334_
timestamp 1688980957
transform -1 0 25392 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2335_
timestamp 1688980957
transform 1 0 1748 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2336_
timestamp 1688980957
transform 1 0 27232 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2337_
timestamp 1688980957
transform -1 0 37444 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2338_
timestamp 1688980957
transform -1 0 25852 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2339_
timestamp 1688980957
transform 1 0 19780 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2340_
timestamp 1688980957
transform 1 0 27508 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2341_
timestamp 1688980957
transform -1 0 34960 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2342_
timestamp 1688980957
transform 1 0 27968 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2343_
timestamp 1688980957
transform -1 0 32292 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2344_
timestamp 1688980957
transform -1 0 26220 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2345_
timestamp 1688980957
transform 1 0 4968 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2346_
timestamp 1688980957
transform -1 0 25760 0 -1 38080
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _2347_
timestamp 1688980957
transform 1 0 12328 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2348_
timestamp 1688980957
transform 1 0 14352 0 1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2349_
timestamp 1688980957
transform -1 0 14628 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2350_
timestamp 1688980957
transform 1 0 8188 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2351_
timestamp 1688980957
transform 1 0 9108 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2352_
timestamp 1688980957
transform 1 0 7360 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2353_
timestamp 1688980957
transform 1 0 6440 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2354_
timestamp 1688980957
transform 1 0 7084 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2355_
timestamp 1688980957
transform 1 0 6624 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2356_
timestamp 1688980957
transform 1 0 6624 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2357_
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2358_
timestamp 1688980957
transform 1 0 6440 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2359_
timestamp 1688980957
transform 1 0 4968 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2360_
timestamp 1688980957
transform 1 0 9384 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_1  _2361_
timestamp 1688980957
transform 1 0 7176 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2362_
timestamp 1688980957
transform 1 0 6900 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2363_
timestamp 1688980957
transform 1 0 8924 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2364_
timestamp 1688980957
transform 1 0 8004 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2365_
timestamp 1688980957
transform 1 0 6900 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2366_
timestamp 1688980957
transform 1 0 6532 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2367_
timestamp 1688980957
transform 1 0 6532 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2368_
timestamp 1688980957
transform -1 0 6256 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2369_
timestamp 1688980957
transform 1 0 7176 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2370_
timestamp 1688980957
transform 1 0 6992 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__or3_1  _2371_
timestamp 1688980957
transform -1 0 13984 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _2372_
timestamp 1688980957
transform -1 0 13156 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2373_
timestamp 1688980957
transform 1 0 11500 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2374_
timestamp 1688980957
transform -1 0 10948 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2375_
timestamp 1688980957
transform -1 0 13524 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2376_
timestamp 1688980957
transform 1 0 13892 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2377_
timestamp 1688980957
transform 1 0 15088 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2378_
timestamp 1688980957
transform -1 0 14996 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2379_
timestamp 1688980957
transform 1 0 12420 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2380_
timestamp 1688980957
transform -1 0 12236 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2381_
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2382_
timestamp 1688980957
transform 1 0 10304 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2383_
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2384_
timestamp 1688980957
transform -1 0 13984 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2385_
timestamp 1688980957
transform 1 0 11776 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2386_
timestamp 1688980957
transform -1 0 11684 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2387_
timestamp 1688980957
transform -1 0 13616 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2388_
timestamp 1688980957
transform 1 0 13616 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2389_
timestamp 1688980957
transform 1 0 9108 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2390_
timestamp 1688980957
transform 1 0 8556 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2391_
timestamp 1688980957
transform 1 0 15364 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2392_
timestamp 1688980957
transform -1 0 15732 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2393_
timestamp 1688980957
transform -1 0 16008 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2394_
timestamp 1688980957
transform 1 0 16008 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2395_
timestamp 1688980957
transform 1 0 12972 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2396_
timestamp 1688980957
transform -1 0 13432 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2397_
timestamp 1688980957
transform 1 0 10304 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2398_
timestamp 1688980957
transform -1 0 10028 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2399_
timestamp 1688980957
transform 1 0 15548 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2400_
timestamp 1688980957
transform -1 0 15824 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2401_
timestamp 1688980957
transform 1 0 10304 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2402_
timestamp 1688980957
transform 1 0 10028 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2403_
timestamp 1688980957
transform 1 0 9752 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2404_
timestamp 1688980957
transform 1 0 9476 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _2405_
timestamp 1688980957
transform 1 0 16192 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _2406_
timestamp 1688980957
transform -1 0 30452 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2407__8
timestamp 1688980957
transform 1 0 10488 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2408__9
timestamp 1688980957
transform -1 0 7360 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2409__10
timestamp 1688980957
transform -1 0 6992 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2410__11
timestamp 1688980957
transform -1 0 4600 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2411__12
timestamp 1688980957
transform -1 0 6164 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2412__13
timestamp 1688980957
transform 1 0 3956 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2413__14
timestamp 1688980957
transform -1 0 9200 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2414__15
timestamp 1688980957
transform 1 0 4508 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2415__16
timestamp 1688980957
transform -1 0 7636 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2416__17
timestamp 1688980957
transform 1 0 6624 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2417__18
timestamp 1688980957
transform -1 0 8372 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2418__19
timestamp 1688980957
transform -1 0 8188 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2419__20
timestamp 1688980957
transform -1 0 4232 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2420__21
timestamp 1688980957
transform 1 0 4048 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2421__22
timestamp 1688980957
transform 1 0 8556 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2422__23
timestamp 1688980957
transform 1 0 20148 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2423__24
timestamp 1688980957
transform -1 0 25944 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2424__25
timestamp 1688980957
transform 1 0 30360 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2425__26
timestamp 1688980957
transform 1 0 30728 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _2426_
timestamp 1688980957
transform -1 0 34040 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2427__27
timestamp 1688980957
transform 1 0 34960 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2428__28
timestamp 1688980957
transform -1 0 35052 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2429__29
timestamp 1688980957
transform -1 0 31556 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2430__30
timestamp 1688980957
transform -1 0 27784 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2431__31
timestamp 1688980957
transform -1 0 32660 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2432__32
timestamp 1688980957
transform -1 0 9200 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2433__33
timestamp 1688980957
transform 1 0 5704 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2434__34
timestamp 1688980957
transform 1 0 9476 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2435__35
timestamp 1688980957
transform 1 0 5612 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2436__36
timestamp 1688980957
transform -1 0 4416 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2437__37
timestamp 1688980957
transform 1 0 4692 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2438__38
timestamp 1688980957
transform -1 0 13432 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2439__39
timestamp 1688980957
transform 1 0 21528 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2440__40
timestamp 1688980957
transform 1 0 25484 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2441__41
timestamp 1688980957
transform -1 0 33028 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2442__42
timestamp 1688980957
transform -1 0 33764 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2443__43
timestamp 1688980957
transform -1 0 34960 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2444__44
timestamp 1688980957
transform -1 0 32016 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2445__45
timestamp 1688980957
transform -1 0 27968 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _2446_
timestamp 1688980957
transform -1 0 27048 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2447__46
timestamp 1688980957
transform 1 0 25024 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2448__47
timestamp 1688980957
transform 1 0 29624 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2449__48
timestamp 1688980957
transform -1 0 10488 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2450__49
timestamp 1688980957
transform -1 0 9568 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2451__50
timestamp 1688980957
transform 1 0 9936 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2452__51
timestamp 1688980957
transform 1 0 9200 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2453__52
timestamp 1688980957
transform 1 0 8556 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2454__53
timestamp 1688980957
transform 1 0 8556 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2455__54
timestamp 1688980957
transform 1 0 9016 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2456__55
timestamp 1688980957
transform 1 0 18860 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2457__56
timestamp 1688980957
transform -1 0 27968 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2458__57
timestamp 1688980957
transform -1 0 28980 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2459__58
timestamp 1688980957
transform 1 0 29532 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2460__59
timestamp 1688980957
transform -1 0 27508 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2461__60
timestamp 1688980957
transform -1 0 29440 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2462__61
timestamp 1688980957
transform -1 0 28060 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2463__62
timestamp 1688980957
transform -1 0 27784 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2464__63
timestamp 1688980957
transform 1 0 29532 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2465__64
timestamp 1688980957
transform -1 0 29256 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2466__1
timestamp 1688980957
transform 1 0 34316 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2467__2
timestamp 1688980957
transform 1 0 35144 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2468__3
timestamp 1688980957
transform -1 0 35144 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2469__4
timestamp 1688980957
transform -1 0 35144 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2470__5
timestamp 1688980957
transform -1 0 30544 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2471__6
timestamp 1688980957
transform -1 0 27324 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2472__7
timestamp 1688980957
transform 1 0 34316 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2473_
timestamp 1688980957
transform 1 0 17480 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _2474_
timestamp 1688980957
transform 1 0 18676 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2475_
timestamp 1688980957
transform -1 0 10672 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2476_
timestamp 1688980957
transform -1 0 19136 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2477_
timestamp 1688980957
transform 1 0 10120 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2478_
timestamp 1688980957
transform -1 0 11408 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2479_
timestamp 1688980957
transform -1 0 12972 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2480_
timestamp 1688980957
transform -1 0 12512 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2481_
timestamp 1688980957
transform -1 0 13248 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2482_
timestamp 1688980957
transform -1 0 11316 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2483_
timestamp 1688980957
transform -1 0 12236 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2484_
timestamp 1688980957
transform 1 0 11316 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2485_
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2486_
timestamp 1688980957
transform -1 0 12604 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__or4b_1  _2487_
timestamp 1688980957
transform -1 0 13064 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__o41a_1  _2488_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 12328 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__o21ai_2  _2489_
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _2490_
timestamp 1688980957
transform 1 0 11500 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__and3b_1  _2491_
timestamp 1688980957
transform -1 0 12052 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2492_
timestamp 1688980957
transform 1 0 10304 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__o211a_1  _2493_
timestamp 1688980957
transform 1 0 16008 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or3_2  _2494_
timestamp 1688980957
transform -1 0 12696 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_4  _2495_
timestamp 1688980957
transform -1 0 11040 0 1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__mux2_1  _2496_
timestamp 1688980957
transform 1 0 9660 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_8  _2497_
timestamp 1688980957
transform -1 0 14812 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__mux2_1  _2498_
timestamp 1688980957
transform 1 0 8004 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2499_
timestamp 1688980957
transform 1 0 7636 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2500_
timestamp 1688980957
transform 1 0 17572 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2501_
timestamp 1688980957
transform -1 0 17572 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_1  _2502_
timestamp 1688980957
transform -1 0 6992 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2503_
timestamp 1688980957
transform 1 0 6072 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2504_
timestamp 1688980957
transform 1 0 5152 0 -1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2505_
timestamp 1688980957
transform 1 0 4692 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2506_
timestamp 1688980957
transform 1 0 14904 0 1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_1  _2507_
timestamp 1688980957
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2508_
timestamp 1688980957
transform -1 0 6808 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2509_
timestamp 1688980957
transform 1 0 5612 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2510_
timestamp 1688980957
transform 1 0 5060 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2511_
timestamp 1688980957
transform 1 0 3772 0 -1 8704
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2512_
timestamp 1688980957
transform 1 0 3220 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2513_
timestamp 1688980957
transform 1 0 13064 0 -1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2514_
timestamp 1688980957
transform -1 0 6164 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2515_
timestamp 1688980957
transform -1 0 6256 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2516_
timestamp 1688980957
transform -1 0 6256 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2517_
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2518_
timestamp 1688980957
transform 1 0 5152 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2519_
timestamp 1688980957
transform 1 0 4600 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2520_
timestamp 1688980957
transform 1 0 10580 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _2521_
timestamp 1688980957
transform 1 0 3128 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2522_
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2523_
timestamp 1688980957
transform 1 0 2300 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2524_
timestamp 1688980957
transform 1 0 1748 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2525_
timestamp 1688980957
transform 1 0 22172 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__mux2_1  _2526_
timestamp 1688980957
transform 1 0 17572 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__and3_1  _2527_
timestamp 1688980957
transform -1 0 4232 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2528_
timestamp 1688980957
transform 1 0 4232 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2529_
timestamp 1688980957
transform 1 0 4416 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2530_
timestamp 1688980957
transform 1 0 3588 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2531_
timestamp 1688980957
transform 1 0 2576 0 1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2532_
timestamp 1688980957
transform 1 0 1932 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2533_
timestamp 1688980957
transform 1 0 10948 0 1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2534_
timestamp 1688980957
transform 1 0 4508 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2535_
timestamp 1688980957
transform -1 0 3680 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2536_
timestamp 1688980957
transform 1 0 4048 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2537_
timestamp 1688980957
transform 1 0 3680 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2538_
timestamp 1688980957
transform 1 0 2484 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2539_
timestamp 1688980957
transform 1 0 1932 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _2540_
timestamp 1688980957
transform 1 0 11868 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_1  _2541_
timestamp 1688980957
transform 1 0 4416 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2542_
timestamp 1688980957
transform 1 0 5152 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__mux2_1  _2543_
timestamp 1688980957
transform 1 0 4508 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2544_
timestamp 1688980957
transform 1 0 4232 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2545_
timestamp 1688980957
transform -1 0 4324 0 -1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2546_
timestamp 1688980957
transform 1 0 4508 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2547_
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_2  _2548_
timestamp 1688980957
transform -1 0 10672 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_1  _2549_
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2550_
timestamp 1688980957
transform 1 0 2300 0 1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2551_
timestamp 1688980957
transform 1 0 2024 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2552_
timestamp 1688980957
transform 1 0 3312 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2553_
timestamp 1688980957
transform 1 0 3772 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2554_
timestamp 1688980957
transform 1 0 3496 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _2555_
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2556_
timestamp 1688980957
transform 1 0 2392 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2557_
timestamp 1688980957
transform 1 0 1748 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2558_
timestamp 1688980957
transform 1 0 3864 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2559_
timestamp 1688980957
transform -1 0 3864 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _2560_
timestamp 1688980957
transform 1 0 2944 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2561_
timestamp 1688980957
transform 1 0 2300 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2562_
timestamp 1688980957
transform 1 0 1748 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2563_
timestamp 1688980957
transform 1 0 3772 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2564_
timestamp 1688980957
transform 1 0 4232 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2565_
timestamp 1688980957
transform -1 0 4416 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a32o_1  _2566_
timestamp 1688980957
transform 1 0 4048 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2567_
timestamp 1688980957
transform 1 0 3220 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2568_
timestamp 1688980957
transform 1 0 1748 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2569_
timestamp 1688980957
transform 1 0 6716 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2570_
timestamp 1688980957
transform 1 0 7728 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _2571_
timestamp 1688980957
transform 1 0 6992 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2572_
timestamp 1688980957
transform 1 0 6348 0 -1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2573_
timestamp 1688980957
transform 1 0 5704 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2574_
timestamp 1688980957
transform -1 0 6716 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2575_
timestamp 1688980957
transform -1 0 5704 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2576_
timestamp 1688980957
transform 1 0 5704 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_1  _2577_
timestamp 1688980957
transform 1 0 4968 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2578_
timestamp 1688980957
transform 1 0 4324 0 -1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2579_
timestamp 1688980957
transform 1 0 3864 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2580_
timestamp 1688980957
transform -1 0 5796 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2581_
timestamp 1688980957
transform -1 0 5520 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _2582_
timestamp 1688980957
transform 1 0 4232 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__mux2_1  _2583_
timestamp 1688980957
transform 1 0 3772 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2584_
timestamp 1688980957
transform 1 0 2852 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2585_
timestamp 1688980957
transform 1 0 4508 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2586_
timestamp 1688980957
transform -1 0 6624 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__mux2_1  _2587_
timestamp 1688980957
transform 1 0 5152 0 1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _2588_
timestamp 1688980957
transform 1 0 4692 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_1  _2589_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14168 0 1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2590_
timestamp 1688980957
transform 1 0 6900 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2591_
timestamp 1688980957
transform 1 0 8004 0 -1 4352
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2592_
timestamp 1688980957
transform 1 0 5060 0 1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2593_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6164 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2594_
timestamp 1688980957
transform 1 0 5612 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2595_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4324 0 1 13056
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2596_
timestamp 1688980957
transform 1 0 6532 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2597_
timestamp 1688980957
transform 1 0 7544 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2598_
timestamp 1688980957
transform 1 0 6072 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2599_
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2600_
timestamp 1688980957
transform 1 0 6624 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2601_
timestamp 1688980957
transform 1 0 10948 0 1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2602_
timestamp 1688980957
transform 1 0 11868 0 1 15232
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_1  _2603_
timestamp 1688980957
transform 1 0 15088 0 1 11968
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2604_
timestamp 1688980957
transform 1 0 12236 0 -1 11968
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2605_
timestamp 1688980957
transform 1 0 9844 0 1 14144
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2606_
timestamp 1688980957
transform 1 0 13892 0 -1 10880
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2607_
timestamp 1688980957
transform 1 0 11684 0 1 9792
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2608_
timestamp 1688980957
transform 1 0 13156 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2609_
timestamp 1688980957
transform 1 0 8280 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2610_
timestamp 1688980957
transform 1 0 15456 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2611_
timestamp 1688980957
transform 1 0 15732 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2612_
timestamp 1688980957
transform 1 0 13432 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2613_
timestamp 1688980957
transform 1 0 10028 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2614_
timestamp 1688980957
transform 1 0 15824 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2615_
timestamp 1688980957
transform 1 0 9752 0 1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2616_
timestamp 1688980957
transform 1 0 9108 0 1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_4  _2617_
timestamp 1688980957
transform 1 0 10764 0 1 22848
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2618_
timestamp 1688980957
transform 1 0 6992 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2619_
timestamp 1688980957
transform 1 0 6624 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2620_
timestamp 1688980957
transform 1 0 4232 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2621_
timestamp 1688980957
transform 1 0 6164 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2622_
timestamp 1688980957
transform 1 0 4232 0 1 31552
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2623_
timestamp 1688980957
transform 1 0 8648 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2624_
timestamp 1688980957
transform 1 0 4784 0 1 26112
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2625_
timestamp 1688980957
transform 1 0 7268 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2626_
timestamp 1688980957
transform 1 0 6900 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2627_
timestamp 1688980957
transform 1 0 7636 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2628_
timestamp 1688980957
transform 1 0 7820 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2629_
timestamp 1688980957
transform 1 0 3864 0 -1 29376
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2630_
timestamp 1688980957
transform 1 0 4324 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2631_
timestamp 1688980957
transform 1 0 8924 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2632_
timestamp 1688980957
transform 1 0 20424 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2633_
timestamp 1688980957
transform 1 0 25576 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2634_
timestamp 1688980957
transform 1 0 30636 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2635_
timestamp 1688980957
transform 1 0 31004 0 1 26112
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2636_
timestamp 1688980957
transform 1 0 34500 0 -1 31552
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2637_
timestamp 1688980957
transform 1 0 34684 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2638_
timestamp 1688980957
transform 1 0 31188 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2639_
timestamp 1688980957
transform 1 0 27416 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2640_
timestamp 1688980957
transform 1 0 32292 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2641_
timestamp 1688980957
transform 1 0 8648 0 -1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2642_
timestamp 1688980957
transform 1 0 5980 0 1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2643_
timestamp 1688980957
transform 1 0 9752 0 1 27200
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2644_
timestamp 1688980957
transform 1 0 5888 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2645_
timestamp 1688980957
transform 1 0 4048 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2646_
timestamp 1688980957
transform 1 0 4968 0 1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2647_
timestamp 1688980957
transform -1 0 13156 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2648_
timestamp 1688980957
transform 1 0 21804 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2649_
timestamp 1688980957
transform 1 0 25760 0 1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2650_
timestamp 1688980957
transform 1 0 32660 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2651_
timestamp 1688980957
transform 1 0 33396 0 -1 27200
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2652_
timestamp 1688980957
transform -1 0 34500 0 -1 31552
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2653_
timestamp 1688980957
transform 1 0 31740 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2654_
timestamp 1688980957
transform 1 0 27508 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2655_
timestamp 1688980957
transform 1 0 25300 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2656_
timestamp 1688980957
transform 1 0 29900 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2657_
timestamp 1688980957
transform 1 0 10120 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2658_
timestamp 1688980957
transform 1 0 9200 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2659_
timestamp 1688980957
transform 1 0 10212 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2660_
timestamp 1688980957
transform 1 0 9476 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2661_
timestamp 1688980957
transform 1 0 8924 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2662_
timestamp 1688980957
transform 1 0 8924 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2663_
timestamp 1688980957
transform 1 0 9292 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2664_
timestamp 1688980957
transform 1 0 19228 0 1 38080
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2665_
timestamp 1688980957
transform 1 0 27508 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2666_
timestamp 1688980957
transform 1 0 28612 0 -1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2667_
timestamp 1688980957
transform 1 0 29440 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2668_
timestamp 1688980957
transform 1 0 27232 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2669_
timestamp 1688980957
transform 1 0 29164 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2670_
timestamp 1688980957
transform 1 0 27692 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2671_
timestamp 1688980957
transform 1 0 27232 0 1 38080
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2672_
timestamp 1688980957
transform 1 0 29072 0 -1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_4  _2673_
timestamp 1688980957
transform 1 0 28888 0 -1 25024
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2674_
timestamp 1688980957
transform 1 0 34684 0 1 32640
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2675_
timestamp 1688980957
transform 1 0 34960 0 1 26112
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2676_
timestamp 1688980957
transform 1 0 34776 0 1 29376
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2677_
timestamp 1688980957
transform 1 0 34684 0 1 25024
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2678_
timestamp 1688980957
transform 1 0 29900 0 -1 31552
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2679_
timestamp 1688980957
transform 1 0 26956 0 -1 33728
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_4  _2680_
timestamp 1688980957
transform 1 0 34684 0 1 33728
box -38 -48 2154 592
use sky130_fd_sc_hd__dfrtp_2  _2681_
timestamp 1688980957
transform 1 0 6900 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2682_
timestamp 1688980957
transform 1 0 4232 0 1 6528
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2683_
timestamp 1688980957
transform 1 0 2576 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2684_
timestamp 1688980957
transform 1 0 4048 0 -1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2685_
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2686_
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2687_
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2688_
timestamp 1688980957
transform 1 0 3956 0 1 17408
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2689_
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2690_
timestamp 1688980957
transform 1 0 1380 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2691_
timestamp 1688980957
transform 1 0 1380 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2692_
timestamp 1688980957
transform 1 0 1380 0 -1 21760
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2693_
timestamp 1688980957
transform 1 0 5244 0 1 23936
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2694_
timestamp 1688980957
transform 1 0 3312 0 -1 26112
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2695_
timestamp 1688980957
transform 1 0 1840 0 1 25024
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2696_
timestamp 1688980957
transform 1 0 4140 0 -1 19584
box -38 -48 1878 592
use sky130_fd_sc_hd__dfstp_1  _2697_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 17572 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2698_
timestamp 1688980957
transform 1 0 13432 0 -1 5440
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_2  _2699_
timestamp 1688980957
transform 1 0 10672 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _2700_
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_1  _2701_
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__dfrtp_1  _2702_
timestamp 1688980957
transform 1 0 9384 0 -1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0514_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30912 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0515_
timestamp 1688980957
transform -1 0 19136 0 1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0516_
timestamp 1688980957
transform -1 0 21344 0 -1 32640
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0__0517_
timestamp 1688980957
transform -1 0 21344 0 1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_clk
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0514_
timestamp 1688980957
transform 1 0 31188 0 1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0515_
timestamp 1688980957
transform -1 0 11408 0 -1 29376
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0516_
timestamp 1688980957
transform -1 0 14812 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_0__f__0517_
timestamp 1688980957
transform -1 0 14812 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0514_
timestamp 1688980957
transform -1 0 30452 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0515_
timestamp 1688980957
transform 1 0 20792 0 1 28288
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0516_
timestamp 1688980957
transform 1 0 23368 0 -1 31552
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_1_1__f__0517_
timestamp 1688980957
transform 1 0 23368 0 -1 30464
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_0__f_clk
timestamp 1688980957
transform 1 0 7820 0 -1 8704
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_1__f_clk
timestamp 1688980957
transform 1 0 10396 0 1 7616
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_2__f_clk
timestamp 1688980957
transform -1 0 4416 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_2_3__f_clk
timestamp 1688980957
transform 1 0 9476 0 -1 18496
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_6  fanout57
timestamp 1688980957
transform 1 0 7820 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__buf_8  fanout58
timestamp 1688980957
transform -1 0 3404 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  fanout59
timestamp 1688980957
transform -1 0 9200 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_4  fanout60
timestamp 1688980957
transform 1 0 7176 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  fanout61
timestamp 1688980957
transform -1 0 8832 0 -1 36992
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_8  fanout62
timestamp 1688980957
transform 1 0 28336 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_6  fanout63
timestamp 1688980957
transform 1 0 20240 0 -1 38080
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1932 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_16 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2576 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_29 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_37
timestamp 1688980957
transform 1 0 4508 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_49 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5612 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_55
timestamp 1688980957
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_57
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_65
timestamp 1688980957
transform 1 0 7084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_77 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8188 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_83
timestamp 1688980957
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_97 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_105
timestamp 1688980957
transform 1 0 10764 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_125 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12604 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_135
timestamp 1688980957
transform 1 0 13524 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 1688980957
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_149
timestamp 1688980957
transform 1 0 14812 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_156
timestamp 1688980957
transform 1 0 15456 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_169
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_177
timestamp 1688980957
transform 1 0 17388 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_184
timestamp 1688980957
transform 1 0 18032 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_197
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_205
timestamp 1688980957
transform 1 0 19964 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_217
timestamp 1688980957
transform 1 0 21068 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_223
timestamp 1688980957
transform 1 0 21620 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_225
timestamp 1688980957
transform 1 0 21804 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_237
timestamp 1688980957
transform 1 0 22908 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_249
timestamp 1688980957
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_265
timestamp 1688980957
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1688980957
transform 1 0 26588 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_287
timestamp 1688980957
transform 1 0 27508 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_299
timestamp 1688980957
transform 1 0 28612 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_307
timestamp 1688980957
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_321
timestamp 1688980957
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_333
timestamp 1688980957
transform 1 0 31740 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_337
timestamp 1688980957
transform 1 0 32108 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_349
timestamp 1688980957
transform 1 0 33212 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_361
timestamp 1688980957
transform 1 0 34316 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_365
timestamp 1688980957
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_377
timestamp 1688980957
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_389
timestamp 1688980957
transform 1 0 36892 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_393
timestamp 1688980957
transform 1 0 37260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_399
timestamp 1688980957
transform 1 0 37812 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_10
timestamp 1688980957
transform 1 0 2024 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_121
timestamp 1688980957
transform 1 0 12236 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_132
timestamp 1688980957
transform 1 0 13248 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_144
timestamp 1688980957
transform 1 0 14352 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_153
timestamp 1688980957
transform 1 0 15180 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_165
timestamp 1688980957
transform 1 0 16284 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_178
timestamp 1688980957
transform 1 0 17480 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_190
timestamp 1688980957
transform 1 0 18584 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_202
timestamp 1688980957
transform 1 0 19688 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_206
timestamp 1688980957
transform 1 0 20056 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_218
timestamp 1688980957
transform 1 0 21160 0 -1 3264
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1688980957
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1688980957
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1688980957
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1688980957
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1688980957
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1688980957
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1688980957
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 1688980957
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_329
timestamp 1688980957
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 1688980957
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_337
timestamp 1688980957
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_349
timestamp 1688980957
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_361
timestamp 1688980957
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_373
timestamp 1688980957
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_385
timestamp 1688980957
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_391
timestamp 1688980957
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_393
timestamp 1688980957
transform 1 0 37260 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1688980957
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1688980957
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1688980957
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1688980957
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1688980957
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1688980957
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1688980957
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_245
timestamp 1688980957
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_251
timestamp 1688980957
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1688980957
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1688980957
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 1688980957
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 1688980957
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1688980957
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1688980957
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1688980957
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_333
timestamp 1688980957
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_345
timestamp 1688980957
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_357
timestamp 1688980957
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_363
timestamp 1688980957
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_365
timestamp 1688980957
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_377
timestamp 1688980957
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_389
timestamp 1688980957
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_95
timestamp 1688980957
transform 1 0 9844 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_107
timestamp 1688980957
transform 1 0 10948 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_143
timestamp 1688980957
transform 1 0 14260 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_147
timestamp 1688980957
transform 1 0 14628 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_159
timestamp 1688980957
transform 1 0 15732 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1688980957
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1688980957
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1688980957
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1688980957
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1688980957
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1688980957
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_249
timestamp 1688980957
transform 1 0 24012 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_257
timestamp 1688980957
transform 1 0 24748 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_265
timestamp 1688980957
transform 1 0 25484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_277
timestamp 1688980957
transform 1 0 26588 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_281
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_289
timestamp 1688980957
transform 1 0 27692 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1688980957
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1688980957
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1688980957
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_329
timestamp 1688980957
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_335
timestamp 1688980957
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1688980957
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1688980957
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_361
timestamp 1688980957
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_373
timestamp 1688980957
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_385
timestamp 1688980957
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_391
timestamp 1688980957
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_393
timestamp 1688980957
transform 1 0 37260 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_9
timestamp 1688980957
transform 1 0 1932 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_21
timestamp 1688980957
transform 1 0 3036 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_93
timestamp 1688980957
transform 1 0 9660 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_100
timestamp 1688980957
transform 1 0 10304 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_125
timestamp 1688980957
transform 1 0 12604 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_137
timestamp 1688980957
transform 1 0 13708 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_169
timestamp 1688980957
transform 1 0 16652 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_181
timestamp 1688980957
transform 1 0 17756 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_193
timestamp 1688980957
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_204
timestamp 1688980957
transform 1 0 19872 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_210
timestamp 1688980957
transform 1 0 20424 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_244
timestamp 1688980957
transform 1 0 23552 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1688980957
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1688980957
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_318
timestamp 1688980957
transform 1 0 30360 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_330
timestamp 1688980957
transform 1 0 31464 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_342
timestamp 1688980957
transform 1 0 32568 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_354
timestamp 1688980957
transform 1 0 33672 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_362
timestamp 1688980957
transform 1 0 34408 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_365
timestamp 1688980957
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_377
timestamp 1688980957
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_389
timestamp 1688980957
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_61
timestamp 1688980957
transform 1 0 6716 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_73
timestamp 1688980957
transform 1 0 7820 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_85
timestamp 1688980957
transform 1 0 8924 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_101
timestamp 1688980957
transform 1 0 10396 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_110
timestamp 1688980957
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_154
timestamp 1688980957
transform 1 0 15272 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_158
timestamp 1688980957
transform 1 0 15640 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1688980957
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_177
timestamp 1688980957
transform 1 0 17388 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_189
timestamp 1688980957
transform 1 0 18492 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_197
timestamp 1688980957
transform 1 0 19228 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_206
timestamp 1688980957
transform 1 0 20056 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_214
timestamp 1688980957
transform 1 0 20792 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_220
timestamp 1688980957
transform 1 0 21344 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_241
timestamp 1688980957
transform 1 0 23276 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_246
timestamp 1688980957
transform 1 0 23736 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_258
timestamp 1688980957
transform 1 0 24840 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_270
timestamp 1688980957
transform 1 0 25944 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_278
timestamp 1688980957
transform 1 0 26680 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_292
timestamp 1688980957
transform 1 0 27968 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_331
timestamp 1688980957
transform 1 0 31556 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 1688980957
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1688980957
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 1688980957
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_361
timestamp 1688980957
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_373
timestamp 1688980957
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_385
timestamp 1688980957
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_391
timestamp 1688980957
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_393
timestamp 1688980957
transform 1 0 37260 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_106
timestamp 1688980957
transform 1 0 10856 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_129
timestamp 1688980957
transform 1 0 12972 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_133
timestamp 1688980957
transform 1 0 13340 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_179
timestamp 1688980957
transform 1 0 17572 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_191
timestamp 1688980957
transform 1 0 18676 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1688980957
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_205
timestamp 1688980957
transform 1 0 19964 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_213
timestamp 1688980957
transform 1 0 20700 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_225
timestamp 1688980957
transform 1 0 21804 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_248
timestamp 1688980957
transform 1 0 23920 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_261
timestamp 1688980957
transform 1 0 25116 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_273
timestamp 1688980957
transform 1 0 26220 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_285
timestamp 1688980957
transform 1 0 27324 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_297
timestamp 1688980957
transform 1 0 28428 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_305
timestamp 1688980957
transform 1 0 29164 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_320
timestamp 1688980957
transform 1 0 30544 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_340
timestamp 1688980957
transform 1 0 32384 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_352
timestamp 1688980957
transform 1 0 33488 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_365
timestamp 1688980957
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_377
timestamp 1688980957
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_389
timestamp 1688980957
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_42
timestamp 1688980957
transform 1 0 4968 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_54
timestamp 1688980957
transform 1 0 6072 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_65
timestamp 1688980957
transform 1 0 7084 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_94
timestamp 1688980957
transform 1 0 9752 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_98
timestamp 1688980957
transform 1 0 10120 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_110
timestamp 1688980957
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_130
timestamp 1688980957
transform 1 0 13064 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_160
timestamp 1688980957
transform 1 0 15824 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_181
timestamp 1688980957
transform 1 0 17756 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_198
timestamp 1688980957
transform 1 0 19320 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1688980957
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1688980957
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1688980957
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_239
timestamp 1688980957
transform 1 0 23092 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_247
timestamp 1688980957
transform 1 0 23828 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_254
timestamp 1688980957
transform 1 0 24472 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_262
timestamp 1688980957
transform 1 0 25208 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_267
timestamp 1688980957
transform 1 0 25668 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1688980957
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_281
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_296
timestamp 1688980957
transform 1 0 28336 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_308
timestamp 1688980957
transform 1 0 29440 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_320
timestamp 1688980957
transform 1 0 30544 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_332
timestamp 1688980957
transform 1 0 31648 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_337
timestamp 1688980957
transform 1 0 32108 0 -1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_345
timestamp 1688980957
transform 1 0 32844 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_357
timestamp 1688980957
transform 1 0 33948 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_369
timestamp 1688980957
transform 1 0 35052 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_381
timestamp 1688980957
transform 1 0 36156 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_389
timestamp 1688980957
transform 1 0 36892 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_393
timestamp 1688980957
transform 1 0 37260 0 -1 6528
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_33
timestamp 1688980957
transform 1 0 4140 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_54
timestamp 1688980957
transform 1 0 6072 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_66
timestamp 1688980957
transform 1 0 7176 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_78
timestamp 1688980957
transform 1 0 8280 0 1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_88
timestamp 1688980957
transform 1 0 9200 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_100
timestamp 1688980957
transform 1 0 10304 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_112
timestamp 1688980957
transform 1 0 11408 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_120
timestamp 1688980957
transform 1 0 12144 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_129
timestamp 1688980957
transform 1 0 12972 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_137
timestamp 1688980957
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_145
timestamp 1688980957
transform 1 0 14444 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_154
timestamp 1688980957
transform 1 0 15272 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_176
timestamp 1688980957
transform 1 0 17296 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_193
timestamp 1688980957
transform 1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_203
timestamp 1688980957
transform 1 0 19780 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_211
timestamp 1688980957
transform 1 0 20516 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_217
timestamp 1688980957
transform 1 0 21068 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_224
timestamp 1688980957
transform 1 0 21712 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_236
timestamp 1688980957
transform 1 0 22816 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_248
timestamp 1688980957
transform 1 0 23920 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_268
timestamp 1688980957
transform 1 0 25760 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_278
timestamp 1688980957
transform 1 0 26680 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_285
timestamp 1688980957
transform 1 0 27324 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_302
timestamp 1688980957
transform 1 0 28888 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_309
timestamp 1688980957
transform 1 0 29532 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_325
timestamp 1688980957
transform 1 0 31004 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_329
timestamp 1688980957
transform 1 0 31372 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_338
timestamp 1688980957
transform 1 0 32200 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_354
timestamp 1688980957
transform 1 0 33672 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_362
timestamp 1688980957
transform 1 0 34408 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_365
timestamp 1688980957
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_377
timestamp 1688980957
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_389
timestamp 1688980957
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_7
timestamp 1688980957
transform 1 0 1748 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_36
timestamp 1688980957
transform 1 0 4416 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_53
timestamp 1688980957
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_64
timestamp 1688980957
transform 1 0 6992 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_70
timestamp 1688980957
transform 1 0 7544 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_74
timestamp 1688980957
transform 1 0 7912 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_86
timestamp 1688980957
transform 1 0 9016 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_110
timestamp 1688980957
transform 1 0 11224 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_133
timestamp 1688980957
transform 1 0 13340 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_137
timestamp 1688980957
transform 1 0 13708 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_152
timestamp 1688980957
transform 1 0 15088 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_159
timestamp 1688980957
transform 1 0 15732 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1688980957
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_184
timestamp 1688980957
transform 1 0 18032 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_192
timestamp 1688980957
transform 1 0 18768 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_199
timestamp 1688980957
transform 1 0 19412 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_210
timestamp 1688980957
transform 1 0 20424 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_219
timestamp 1688980957
transform 1 0 21252 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1688980957
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_232
timestamp 1688980957
transform 1 0 22448 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_241
timestamp 1688980957
transform 1 0 23276 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_267
timestamp 1688980957
transform 1 0 25668 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_278
timestamp 1688980957
transform 1 0 26680 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_281
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_287
timestamp 1688980957
transform 1 0 27508 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_318
timestamp 1688980957
transform 1 0 30360 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_337
timestamp 1688980957
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_349
timestamp 1688980957
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_361
timestamp 1688980957
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_373
timestamp 1688980957
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_385
timestamp 1688980957
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_391
timestamp 1688980957
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_393
timestamp 1688980957
transform 1 0 37260 0 -1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_52
timestamp 1688980957
transform 1 0 5888 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_96
timestamp 1688980957
transform 1 0 9936 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_100
timestamp 1688980957
transform 1 0 10304 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_153
timestamp 1688980957
transform 1 0 15180 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_164
timestamp 1688980957
transform 1 0 16192 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_172
timestamp 1688980957
transform 1 0 16928 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_182
timestamp 1688980957
transform 1 0 17848 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_194
timestamp 1688980957
transform 1 0 18952 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_197
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_201
timestamp 1688980957
transform 1 0 19596 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_205
timestamp 1688980957
transform 1 0 19964 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1688980957
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_221
timestamp 1688980957
transform 1 0 21436 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 1688980957
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1688980957
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1688980957
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 1688980957
transform 1 0 26588 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_289
timestamp 1688980957
transform 1 0 27692 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 1688980957
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1688980957
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_309
timestamp 1688980957
transform 1 0 29532 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_313
timestamp 1688980957
transform 1 0 29900 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_323
timestamp 1688980957
transform 1 0 30820 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_335
timestamp 1688980957
transform 1 0 31924 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_347
timestamp 1688980957
transform 1 0 33028 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_359
timestamp 1688980957
transform 1 0 34132 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_363
timestamp 1688980957
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_365
timestamp 1688980957
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_377
timestamp 1688980957
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_389
timestamp 1688980957
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_15
timestamp 1688980957
transform 1 0 2484 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_26
timestamp 1688980957
transform 1 0 3496 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_38
timestamp 1688980957
transform 1 0 4600 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_42
timestamp 1688980957
transform 1 0 4968 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_62
timestamp 1688980957
transform 1 0 6808 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_70
timestamp 1688980957
transform 1 0 7544 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1688980957
transform 1 0 10764 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_154
timestamp 1688980957
transform 1 0 15272 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_166
timestamp 1688980957
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_180
timestamp 1688980957
transform 1 0 17664 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_195
timestamp 1688980957
transform 1 0 19044 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_199
timestamp 1688980957
transform 1 0 19412 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_204
timestamp 1688980957
transform 1 0 19872 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_216
timestamp 1688980957
transform 1 0 20976 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_225
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_231
timestamp 1688980957
transform 1 0 22356 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_237
timestamp 1688980957
transform 1 0 22908 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_246
timestamp 1688980957
transform 1 0 23736 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_254
timestamp 1688980957
transform 1 0 24472 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_264
timestamp 1688980957
transform 1 0 25392 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_276
timestamp 1688980957
transform 1 0 26496 0 -1 8704
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_290
timestamp 1688980957
transform 1 0 27784 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_308
timestamp 1688980957
transform 1 0 29440 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_320
timestamp 1688980957
transform 1 0 30544 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_326
timestamp 1688980957
transform 1 0 31096 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_335
timestamp 1688980957
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_337
timestamp 1688980957
transform 1 0 32108 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_343
timestamp 1688980957
transform 1 0 32660 0 -1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_351
timestamp 1688980957
transform 1 0 33396 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_363
timestamp 1688980957
transform 1 0 34500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_375
timestamp 1688980957
transform 1 0 35604 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_387
timestamp 1688980957
transform 1 0 36708 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_391
timestamp 1688980957
transform 1 0 37076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_393
timestamp 1688980957
transform 1 0 37260 0 -1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_9
timestamp 1688980957
transform 1 0 1932 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_21
timestamp 1688980957
transform 1 0 3036 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_43
timestamp 1688980957
transform 1 0 5060 0 1 8704
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_56
timestamp 1688980957
transform 1 0 6256 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_68
timestamp 1688980957
transform 1 0 7360 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_74
timestamp 1688980957
transform 1 0 7912 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_93
timestamp 1688980957
transform 1 0 9660 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_114
timestamp 1688980957
transform 1 0 11592 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_138
timestamp 1688980957
transform 1 0 13800 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_149
timestamp 1688980957
transform 1 0 14812 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_179
timestamp 1688980957
transform 1 0 17572 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_192
timestamp 1688980957
transform 1 0 18768 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_206
timestamp 1688980957
transform 1 0 20056 0 1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_216
timestamp 1688980957
transform 1 0 20976 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_228
timestamp 1688980957
transform 1 0 22080 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_245
timestamp 1688980957
transform 1 0 23644 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_250
timestamp 1688980957
transform 1 0 24104 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_261
timestamp 1688980957
transform 1 0 25116 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_277
timestamp 1688980957
transform 1 0 26588 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_293
timestamp 1688980957
transform 1 0 28060 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_319
timestamp 1688980957
transform 1 0 30452 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_325
timestamp 1688980957
transform 1 0 31004 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_339
timestamp 1688980957
transform 1 0 32292 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_353
timestamp 1688980957
transform 1 0 33580 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_361
timestamp 1688980957
transform 1 0 34316 0 1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_365
timestamp 1688980957
transform 1 0 34684 0 1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_377
timestamp 1688980957
transform 1 0 35788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_389
timestamp 1688980957
transform 1 0 36892 0 1 8704
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_15
timestamp 1688980957
transform 1 0 2484 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_19
timestamp 1688980957
transform 1 0 2852 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_28
timestamp 1688980957
transform 1 0 3680 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_40
timestamp 1688980957
transform 1 0 4784 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_52
timestamp 1688980957
transform 1 0 5888 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_65
timestamp 1688980957
transform 1 0 7084 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_79
timestamp 1688980957
transform 1 0 8372 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_83
timestamp 1688980957
transform 1 0 8740 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_95
timestamp 1688980957
transform 1 0 9844 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_109
timestamp 1688980957
transform 1 0 11132 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_125
timestamp 1688980957
transform 1 0 12604 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_129
timestamp 1688980957
transform 1 0 12972 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_139
timestamp 1688980957
transform 1 0 13892 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_151
timestamp 1688980957
transform 1 0 14996 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_165
timestamp 1688980957
transform 1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_178
timestamp 1688980957
transform 1 0 17480 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_200
timestamp 1688980957
transform 1 0 19504 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_208
timestamp 1688980957
transform 1 0 20240 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_220
timestamp 1688980957
transform 1 0 21344 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_225
timestamp 1688980957
transform 1 0 21804 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_231
timestamp 1688980957
transform 1 0 22356 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_240
timestamp 1688980957
transform 1 0 23184 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_248
timestamp 1688980957
transform 1 0 23920 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_260
timestamp 1688980957
transform 1 0 25024 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_268
timestamp 1688980957
transform 1 0 25760 0 -1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_289
timestamp 1688980957
transform 1 0 27692 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_306
timestamp 1688980957
transform 1 0 29256 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_316
timestamp 1688980957
transform 1 0 30176 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_344
timestamp 1688980957
transform 1 0 32752 0 -1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_350
timestamp 1688980957
transform 1 0 33304 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_362
timestamp 1688980957
transform 1 0 34408 0 -1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_374
timestamp 1688980957
transform 1 0 35512 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_386
timestamp 1688980957
transform 1 0 36616 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_393
timestamp 1688980957
transform 1 0 37260 0 -1 9792
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_3
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_15
timestamp 1688980957
transform 1 0 2484 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_23
timestamp 1688980957
transform 1 0 3220 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1688980957
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_37
timestamp 1688980957
transform 1 0 4508 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_41
timestamp 1688980957
transform 1 0 4876 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_56
timestamp 1688980957
transform 1 0 6256 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_68
timestamp 1688980957
transform 1 0 7360 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_81
timestamp 1688980957
transform 1 0 8556 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_92
timestamp 1688980957
transform 1 0 9568 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_14_104
timestamp 1688980957
transform 1 0 10672 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_138
timestamp 1688980957
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_153
timestamp 1688980957
transform 1 0 15180 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_165
timestamp 1688980957
transform 1 0 16284 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_177
timestamp 1688980957
transform 1 0 17388 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_192
timestamp 1688980957
transform 1 0 18768 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_203
timestamp 1688980957
transform 1 0 19780 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_207
timestamp 1688980957
transform 1 0 20148 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_227
timestamp 1688980957
transform 1 0 21988 0 1 9792
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_235
timestamp 1688980957
transform 1 0 22724 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_247
timestamp 1688980957
transform 1 0 23828 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_251
timestamp 1688980957
transform 1 0 24196 0 1 9792
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_253
timestamp 1688980957
transform 1 0 24380 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_265
timestamp 1688980957
transform 1 0 25484 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_277
timestamp 1688980957
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_289
timestamp 1688980957
transform 1 0 27692 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_14_305
timestamp 1688980957
transform 1 0 29164 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_309
timestamp 1688980957
transform 1 0 29532 0 1 9792
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_324
timestamp 1688980957
transform 1 0 30912 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_336
timestamp 1688980957
transform 1 0 32016 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_345
timestamp 1688980957
transform 1 0 32844 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_351
timestamp 1688980957
transform 1 0 33396 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_360
timestamp 1688980957
transform 1 0 34224 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_365
timestamp 1688980957
transform 1 0 34684 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_377
timestamp 1688980957
transform 1 0 35788 0 1 9792
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_389
timestamp 1688980957
transform 1 0 36892 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_3
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_10
timestamp 1688980957
transform 1 0 2024 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_29
timestamp 1688980957
transform 1 0 3772 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_52
timestamp 1688980957
transform 1 0 5888 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_71
timestamp 1688980957
transform 1 0 7636 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_79
timestamp 1688980957
transform 1 0 8372 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_93
timestamp 1688980957
transform 1 0 9660 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_101
timestamp 1688980957
transform 1 0 10396 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_113
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_125
timestamp 1688980957
transform 1 0 12604 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_137
timestamp 1688980957
transform 1 0 13708 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_162
timestamp 1688980957
transform 1 0 16008 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_169
timestamp 1688980957
transform 1 0 16652 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_179
timestamp 1688980957
transform 1 0 17572 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_202
timestamp 1688980957
transform 1 0 19688 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_209
timestamp 1688980957
transform 1 0 20332 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_213
timestamp 1688980957
transform 1 0 20700 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_233
timestamp 1688980957
transform 1 0 22540 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_243
timestamp 1688980957
transform 1 0 23460 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_256
timestamp 1688980957
transform 1 0 24656 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_268
timestamp 1688980957
transform 1 0 25760 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_289
timestamp 1688980957
transform 1 0 27692 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_293
timestamp 1688980957
transform 1 0 28060 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_304
timestamp 1688980957
transform 1 0 29072 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_316
timestamp 1688980957
transform 1 0 30176 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_320
timestamp 1688980957
transform 1 0 30544 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_332
timestamp 1688980957
transform 1 0 31648 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_347
timestamp 1688980957
transform 1 0 33028 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_351
timestamp 1688980957
transform 1 0 33396 0 -1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_370
timestamp 1688980957
transform 1 0 35144 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_382
timestamp 1688980957
transform 1 0 36248 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_390
timestamp 1688980957
transform 1 0 36984 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_393
timestamp 1688980957
transform 1 0 37260 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_23
timestamp 1688980957
transform 1 0 3220 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_27
timestamp 1688980957
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_38
timestamp 1688980957
transform 1 0 4600 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_55
timestamp 1688980957
transform 1 0 6164 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_67
timestamp 1688980957
transform 1 0 7268 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_82
timestamp 1688980957
transform 1 0 8648 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_92
timestamp 1688980957
transform 1 0 9568 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_117
timestamp 1688980957
transform 1 0 11868 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_132
timestamp 1688980957
transform 1 0 13248 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_136
timestamp 1688980957
transform 1 0 13616 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_150
timestamp 1688980957
transform 1 0 14904 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_156
timestamp 1688980957
transform 1 0 15456 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_180
timestamp 1688980957
transform 1 0 17664 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_193
timestamp 1688980957
transform 1 0 18860 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_209
timestamp 1688980957
transform 1 0 20332 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_217
timestamp 1688980957
transform 1 0 21068 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_233
timestamp 1688980957
transform 1 0 22540 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_241
timestamp 1688980957
transform 1 0 23276 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_247
timestamp 1688980957
transform 1 0 23828 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_251
timestamp 1688980957
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_253
timestamp 1688980957
transform 1 0 24380 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_261
timestamp 1688980957
transform 1 0 25116 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_267
timestamp 1688980957
transform 1 0 25668 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_298
timestamp 1688980957
transform 1 0 28520 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_309
timestamp 1688980957
transform 1 0 29532 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_313
timestamp 1688980957
transform 1 0 29900 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_321
timestamp 1688980957
transform 1 0 30636 0 1 10880
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_350
timestamp 1688980957
transform 1 0 33304 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_362
timestamp 1688980957
transform 1 0 34408 0 1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_365
timestamp 1688980957
transform 1 0 34684 0 1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_377
timestamp 1688980957
transform 1 0 35788 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_389
timestamp 1688980957
transform 1 0 36892 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_7
timestamp 1688980957
transform 1 0 1748 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_19
timestamp 1688980957
transform 1 0 2852 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_31
timestamp 1688980957
transform 1 0 3956 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_43
timestamp 1688980957
transform 1 0 5060 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_55
timestamp 1688980957
transform 1 0 6164 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1688980957
transform 1 0 7452 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 1688980957
transform 1 0 8556 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_93
timestamp 1688980957
transform 1 0 9660 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_99
timestamp 1688980957
transform 1 0 10212 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_109
timestamp 1688980957
transform 1 0 11132 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_113
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_117
timestamp 1688980957
transform 1 0 11868 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_144
timestamp 1688980957
transform 1 0 14352 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_156
timestamp 1688980957
transform 1 0 15456 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_166
timestamp 1688980957
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_169
timestamp 1688980957
transform 1 0 16652 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_181
timestamp 1688980957
transform 1 0 17756 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_189
timestamp 1688980957
transform 1 0 18492 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_193
timestamp 1688980957
transform 1 0 18860 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_205
timestamp 1688980957
transform 1 0 19964 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_217
timestamp 1688980957
transform 1 0 21068 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_223
timestamp 1688980957
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_225
timestamp 1688980957
transform 1 0 21804 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_237
timestamp 1688980957
transform 1 0 22908 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_248
timestamp 1688980957
transform 1 0 23920 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_261
timestamp 1688980957
transform 1 0 25116 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_273
timestamp 1688980957
transform 1 0 26220 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_279
timestamp 1688980957
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_292
timestamp 1688980957
transform 1 0 27968 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_304
timestamp 1688980957
transform 1 0 29072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_314
timestamp 1688980957
transform 1 0 29992 0 -1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_324
timestamp 1688980957
transform 1 0 30912 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_337
timestamp 1688980957
transform 1 0 32108 0 -1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_345
timestamp 1688980957
transform 1 0 32844 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_357
timestamp 1688980957
transform 1 0 33948 0 -1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_369
timestamp 1688980957
transform 1 0 35052 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_381
timestamp 1688980957
transform 1 0 36156 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_389
timestamp 1688980957
transform 1 0 36892 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_17_393
timestamp 1688980957
transform 1 0 37260 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_3
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_12
timestamp 1688980957
transform 1 0 2208 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_25
timestamp 1688980957
transform 1 0 3404 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_38
timestamp 1688980957
transform 1 0 4600 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_50
timestamp 1688980957
transform 1 0 5704 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_67
timestamp 1688980957
transform 1 0 7268 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_83
timestamp 1688980957
transform 1 0 8740 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_85
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_93
timestamp 1688980957
transform 1 0 9660 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_99
timestamp 1688980957
transform 1 0 10212 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_111
timestamp 1688980957
transform 1 0 11316 0 1 11968
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_122
timestamp 1688980957
transform 1 0 12328 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_134
timestamp 1688980957
transform 1 0 13432 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_141
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_147
timestamp 1688980957
transform 1 0 14628 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_151
timestamp 1688980957
transform 1 0 14996 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_172
timestamp 1688980957
transform 1 0 16928 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_178
timestamp 1688980957
transform 1 0 17480 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_195
timestamp 1688980957
transform 1 0 19044 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_197
timestamp 1688980957
transform 1 0 19228 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_202
timestamp 1688980957
transform 1 0 19688 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_214
timestamp 1688980957
transform 1 0 20792 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_227
timestamp 1688980957
transform 1 0 21988 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_235
timestamp 1688980957
transform 1 0 22724 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_247
timestamp 1688980957
transform 1 0 23828 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_251
timestamp 1688980957
transform 1 0 24196 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_253
timestamp 1688980957
transform 1 0 24380 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_261
timestamp 1688980957
transform 1 0 25116 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_271
timestamp 1688980957
transform 1 0 26036 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_281
timestamp 1688980957
transform 1 0 26956 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_293
timestamp 1688980957
transform 1 0 28060 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_305
timestamp 1688980957
transform 1 0 29164 0 1 11968
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_321
timestamp 1688980957
transform 1 0 30636 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_333
timestamp 1688980957
transform 1 0 31740 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_345
timestamp 1688980957
transform 1 0 32844 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_356
timestamp 1688980957
transform 1 0 33856 0 1 11968
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_365
timestamp 1688980957
transform 1 0 34684 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_377
timestamp 1688980957
transform 1 0 35788 0 1 11968
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_389
timestamp 1688980957
transform 1 0 36892 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_23
timestamp 1688980957
transform 1 0 3220 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_39
timestamp 1688980957
transform 1 0 4692 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_45
timestamp 1688980957
transform 1 0 5244 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_104
timestamp 1688980957
transform 1 0 10672 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_113
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_119
timestamp 1688980957
transform 1 0 12052 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_161
timestamp 1688980957
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 1688980957
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_169
timestamp 1688980957
transform 1 0 16652 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_182
timestamp 1688980957
transform 1 0 17848 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_194
timestamp 1688980957
transform 1 0 18952 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_212
timestamp 1688980957
transform 1 0 20608 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_216
timestamp 1688980957
transform 1 0 20976 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_234
timestamp 1688980957
transform 1 0 22632 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_246
timestamp 1688980957
transform 1 0 23736 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_263
timestamp 1688980957
transform 1 0 25300 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_271
timestamp 1688980957
transform 1 0 26036 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_281
timestamp 1688980957
transform 1 0 26956 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_293
timestamp 1688980957
transform 1 0 28060 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_301
timestamp 1688980957
transform 1 0 28796 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_308
timestamp 1688980957
transform 1 0 29440 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_316
timestamp 1688980957
transform 1 0 30176 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_326
timestamp 1688980957
transform 1 0 31096 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_335
timestamp 1688980957
transform 1 0 31924 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_342
timestamp 1688980957
transform 1 0 32568 0 -1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_349
timestamp 1688980957
transform 1 0 33212 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_361
timestamp 1688980957
transform 1 0 34316 0 -1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_373
timestamp 1688980957
transform 1 0 35420 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_385
timestamp 1688980957
transform 1 0 36524 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_391
timestamp 1688980957
transform 1 0 37076 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_393
timestamp 1688980957
transform 1 0 37260 0 -1 13056
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_3
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_15
timestamp 1688980957
transform 1 0 2484 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_27
timestamp 1688980957
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_29
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_58
timestamp 1688980957
transform 1 0 6440 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_68
timestamp 1688980957
transform 1 0 7360 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_80
timestamp 1688980957
transform 1 0 8464 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_85
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_139
timestamp 1688980957
transform 1 0 13892 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_141
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_149
timestamp 1688980957
transform 1 0 14812 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_156
timestamp 1688980957
transform 1 0 15456 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_164
timestamp 1688980957
transform 1 0 16192 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_172
timestamp 1688980957
transform 1 0 16928 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_180
timestamp 1688980957
transform 1 0 17664 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_184
timestamp 1688980957
transform 1 0 18032 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_197
timestamp 1688980957
transform 1 0 19228 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_201
timestamp 1688980957
transform 1 0 19596 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_215
timestamp 1688980957
transform 1 0 20884 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_225
timestamp 1688980957
transform 1 0 21804 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_246
timestamp 1688980957
transform 1 0 23736 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_258
timestamp 1688980957
transform 1 0 24840 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_266
timestamp 1688980957
transform 1 0 25576 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_287
timestamp 1688980957
transform 1 0 27508 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_301
timestamp 1688980957
transform 1 0 28796 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_307
timestamp 1688980957
transform 1 0 29348 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_312
timestamp 1688980957
transform 1 0 29808 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_324
timestamp 1688980957
transform 1 0 30912 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_336
timestamp 1688980957
transform 1 0 32016 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_340
timestamp 1688980957
transform 1 0 32384 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_359
timestamp 1688980957
transform 1 0 34132 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_363
timestamp 1688980957
transform 1 0 34500 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_365
timestamp 1688980957
transform 1 0 34684 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_377
timestamp 1688980957
transform 1 0 35788 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_389
timestamp 1688980957
transform 1 0 36892 0 1 13056
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_12
timestamp 1688980957
transform 1 0 2208 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_24
timestamp 1688980957
transform 1 0 3312 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_36
timestamp 1688980957
transform 1 0 4416 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_48
timestamp 1688980957
transform 1 0 5520 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_69
timestamp 1688980957
transform 1 0 7452 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_77
timestamp 1688980957
transform 1 0 8188 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_83
timestamp 1688980957
transform 1 0 8740 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_95
timestamp 1688980957
transform 1 0 9844 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_107
timestamp 1688980957
transform 1 0 10948 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1688980957
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_113
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_125
timestamp 1688980957
transform 1 0 12604 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_137
timestamp 1688980957
transform 1 0 13708 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_143
timestamp 1688980957
transform 1 0 14260 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 1688980957
transform 1 0 16468 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_176
timestamp 1688980957
transform 1 0 17296 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_186
timestamp 1688980957
transform 1 0 18216 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_198
timestamp 1688980957
transform 1 0 19320 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_223
timestamp 1688980957
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_225
timestamp 1688980957
transform 1 0 21804 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_281
timestamp 1688980957
transform 1 0 26956 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_285
timestamp 1688980957
transform 1 0 27324 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_307
timestamp 1688980957
transform 1 0 29348 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_315
timestamp 1688980957
transform 1 0 30084 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_325
timestamp 1688980957
transform 1 0 31004 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_337
timestamp 1688980957
transform 1 0 32108 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_343
timestamp 1688980957
transform 1 0 32660 0 -1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_350
timestamp 1688980957
transform 1 0 33304 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_362
timestamp 1688980957
transform 1 0 34408 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_374
timestamp 1688980957
transform 1 0 35512 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_386
timestamp 1688980957
transform 1 0 36616 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_393
timestamp 1688980957
transform 1 0 37260 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_23
timestamp 1688980957
transform 1 0 3220 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1688980957
transform 1 0 3588 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_29
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_35
timestamp 1688980957
transform 1 0 4324 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_47
timestamp 1688980957
transform 1 0 5428 0 1 14144
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_70
timestamp 1688980957
transform 1 0 7544 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_82
timestamp 1688980957
transform 1 0 8648 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_93
timestamp 1688980957
transform 1 0 9660 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_118
timestamp 1688980957
transform 1 0 11960 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_135
timestamp 1688980957
transform 1 0 13524 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_139
timestamp 1688980957
transform 1 0 13892 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_153
timestamp 1688980957
transform 1 0 15180 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_160
timestamp 1688980957
transform 1 0 15824 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_171
timestamp 1688980957
transform 1 0 16836 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_179
timestamp 1688980957
transform 1 0 17572 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_186
timestamp 1688980957
transform 1 0 18216 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_194
timestamp 1688980957
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_205
timestamp 1688980957
transform 1 0 19964 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_224
timestamp 1688980957
transform 1 0 21712 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_247
timestamp 1688980957
transform 1 0 23828 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_251
timestamp 1688980957
transform 1 0 24196 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_253
timestamp 1688980957
transform 1 0 24380 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_265
timestamp 1688980957
transform 1 0 25484 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_277
timestamp 1688980957
transform 1 0 26588 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_289
timestamp 1688980957
transform 1 0 27692 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_301
timestamp 1688980957
transform 1 0 28796 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_307
timestamp 1688980957
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_309
timestamp 1688980957
transform 1 0 29532 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_315
timestamp 1688980957
transform 1 0 30084 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_326
timestamp 1688980957
transform 1 0 31096 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_336
timestamp 1688980957
transform 1 0 32016 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_348
timestamp 1688980957
transform 1 0 33120 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_360
timestamp 1688980957
transform 1 0 34224 0 1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_365
timestamp 1688980957
transform 1 0 34684 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_377
timestamp 1688980957
transform 1 0 35788 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_389
timestamp 1688980957
transform 1 0 36892 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_3
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_24
timestamp 1688980957
transform 1 0 3312 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_42
timestamp 1688980957
transform 1 0 4968 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_54
timestamp 1688980957
transform 1 0 6072 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_57
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_63
timestamp 1688980957
transform 1 0 6900 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_95
timestamp 1688980957
transform 1 0 9844 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_99
timestamp 1688980957
transform 1 0 10212 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_103
timestamp 1688980957
transform 1 0 10580 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1688980957
transform 1 0 11316 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_122
timestamp 1688980957
transform 1 0 12328 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_153
timestamp 1688980957
transform 1 0 15180 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_160
timestamp 1688980957
transform 1 0 15824 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_169
timestamp 1688980957
transform 1 0 16652 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_187
timestamp 1688980957
transform 1 0 18308 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_203
timestamp 1688980957
transform 1 0 19780 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_212
timestamp 1688980957
transform 1 0 20608 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_230
timestamp 1688980957
transform 1 0 22264 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_242
timestamp 1688980957
transform 1 0 23368 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_254
timestamp 1688980957
transform 1 0 24472 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_262
timestamp 1688980957
transform 1 0 25208 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_271
timestamp 1688980957
transform 1 0 26036 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_279
timestamp 1688980957
transform 1 0 26772 0 -1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_304
timestamp 1688980957
transform 1 0 29072 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_316
timestamp 1688980957
transform 1 0 30176 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_320
timestamp 1688980957
transform 1 0 30544 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_327
timestamp 1688980957
transform 1 0 31188 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_335
timestamp 1688980957
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_337
timestamp 1688980957
transform 1 0 32108 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_352
timestamp 1688980957
transform 1 0 33488 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_362
timestamp 1688980957
transform 1 0 34408 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_374
timestamp 1688980957
transform 1 0 35512 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_386
timestamp 1688980957
transform 1 0 36616 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_393
timestamp 1688980957
transform 1 0 37260 0 -1 15232
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_9
timestamp 1688980957
transform 1 0 1932 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_21
timestamp 1688980957
transform 1 0 3036 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_27
timestamp 1688980957
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_43
timestamp 1688980957
transform 1 0 5060 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_76
timestamp 1688980957
transform 1 0 8096 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_105
timestamp 1688980957
transform 1 0 10764 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_116
timestamp 1688980957
transform 1 0 11776 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_141
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_149
timestamp 1688980957
transform 1 0 14812 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_155
timestamp 1688980957
transform 1 0 15364 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_166
timestamp 1688980957
transform 1 0 16376 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_178
timestamp 1688980957
transform 1 0 17480 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_216
timestamp 1688980957
transform 1 0 20976 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_228
timestamp 1688980957
transform 1 0 22080 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_236
timestamp 1688980957
transform 1 0 22816 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_247
timestamp 1688980957
transform 1 0 23828 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_251
timestamp 1688980957
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_267
timestamp 1688980957
transform 1 0 25668 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_279
timestamp 1688980957
transform 1 0 26772 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_283
timestamp 1688980957
transform 1 0 27140 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_291
timestamp 1688980957
transform 1 0 27876 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_301
timestamp 1688980957
transform 1 0 28796 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_307
timestamp 1688980957
transform 1 0 29348 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_322
timestamp 1688980957
transform 1 0 30728 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_335
timestamp 1688980957
transform 1 0 31924 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_352
timestamp 1688980957
transform 1 0 33488 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_379
timestamp 1688980957
transform 1 0 35972 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_391
timestamp 1688980957
transform 1 0 37076 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_399
timestamp 1688980957
transform 1 0 37812 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_23
timestamp 1688980957
transform 1 0 3220 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_29
timestamp 1688980957
transform 1 0 3772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_35
timestamp 1688980957
transform 1 0 4324 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_43
timestamp 1688980957
transform 1 0 5060 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_53
timestamp 1688980957
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_57
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_69
timestamp 1688980957
transform 1 0 7452 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_81
timestamp 1688980957
transform 1 0 8556 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_89
timestamp 1688980957
transform 1 0 9292 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_103
timestamp 1688980957
transform 1 0 10580 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_111
timestamp 1688980957
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_113
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_126
timestamp 1688980957
transform 1 0 12696 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_138
timestamp 1688980957
transform 1 0 13800 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_149
timestamp 1688980957
transform 1 0 14812 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_161
timestamp 1688980957
transform 1 0 15916 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_167
timestamp 1688980957
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_176
timestamp 1688980957
transform 1 0 17296 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_197
timestamp 1688980957
transform 1 0 19228 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_205
timestamp 1688980957
transform 1 0 19964 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_214
timestamp 1688980957
transform 1 0 20792 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_222
timestamp 1688980957
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_225
timestamp 1688980957
transform 1 0 21804 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_233
timestamp 1688980957
transform 1 0 22540 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_243
timestamp 1688980957
transform 1 0 23460 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_249
timestamp 1688980957
transform 1 0 24012 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_277
timestamp 1688980957
transform 1 0 26588 0 -1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_288
timestamp 1688980957
transform 1 0 27600 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_300
timestamp 1688980957
transform 1 0 28704 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_312
timestamp 1688980957
transform 1 0 29808 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_318
timestamp 1688980957
transform 1 0 30360 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_330
timestamp 1688980957
transform 1 0 31464 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_337
timestamp 1688980957
transform 1 0 32108 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_349
timestamp 1688980957
transform 1 0 33212 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_361
timestamp 1688980957
transform 1 0 34316 0 -1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_371
timestamp 1688980957
transform 1 0 35236 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_383
timestamp 1688980957
transform 1 0 36340 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_391
timestamp 1688980957
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_393
timestamp 1688980957
transform 1 0 37260 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_3
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_22
timestamp 1688980957
transform 1 0 3128 0 1 16320
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_40
timestamp 1688980957
transform 1 0 4784 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_52
timestamp 1688980957
transform 1 0 5888 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_64
timestamp 1688980957
transform 1 0 6992 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_76
timestamp 1688980957
transform 1 0 8096 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_85
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_107
timestamp 1688980957
transform 1 0 10948 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_119
timestamp 1688980957
transform 1 0 12052 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_131
timestamp 1688980957
transform 1 0 13156 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_139
timestamp 1688980957
transform 1 0 13892 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_176
timestamp 1688980957
transform 1 0 17296 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_197
timestamp 1688980957
transform 1 0 19228 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_205
timestamp 1688980957
transform 1 0 19964 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_238
timestamp 1688980957
transform 1 0 23000 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_249
timestamp 1688980957
transform 1 0 24012 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_253
timestamp 1688980957
transform 1 0 24380 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_261
timestamp 1688980957
transform 1 0 25116 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_267
timestamp 1688980957
transform 1 0 25668 0 1 16320
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_276
timestamp 1688980957
transform 1 0 26496 0 1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_288
timestamp 1688980957
transform 1 0 27600 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_300
timestamp 1688980957
transform 1 0 28704 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_309
timestamp 1688980957
transform 1 0 29532 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_313
timestamp 1688980957
transform 1 0 29900 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_317
timestamp 1688980957
transform 1 0 30268 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_323
timestamp 1688980957
transform 1 0 30820 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_330
timestamp 1688980957
transform 1 0 31464 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_336
timestamp 1688980957
transform 1 0 32016 0 1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_342
timestamp 1688980957
transform 1 0 32568 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_354
timestamp 1688980957
transform 1 0 33672 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_365
timestamp 1688980957
transform 1 0 34684 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_378
timestamp 1688980957
transform 1 0 35880 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_390
timestamp 1688980957
transform 1 0 36984 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_398
timestamp 1688980957
transform 1 0 37720 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_3
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_15
timestamp 1688980957
transform 1 0 2484 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_26
timestamp 1688980957
transform 1 0 3496 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_46
timestamp 1688980957
transform 1 0 5336 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_55
timestamp 1688980957
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_62
timestamp 1688980957
transform 1 0 6808 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_72
timestamp 1688980957
transform 1 0 7728 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_84
timestamp 1688980957
transform 1 0 8832 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_90
timestamp 1688980957
transform 1 0 9384 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_104
timestamp 1688980957
transform 1 0 10672 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_113
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_117
timestamp 1688980957
transform 1 0 11868 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_124
timestamp 1688980957
transform 1 0 12512 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_136
timestamp 1688980957
transform 1 0 13616 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_146
timestamp 1688980957
transform 1 0 14536 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_158
timestamp 1688980957
transform 1 0 15640 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_166
timestamp 1688980957
transform 1 0 16376 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_174
timestamp 1688980957
transform 1 0 17112 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_186
timestamp 1688980957
transform 1 0 18216 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_198
timestamp 1688980957
transform 1 0 19320 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_217
timestamp 1688980957
transform 1 0 21068 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_223
timestamp 1688980957
transform 1 0 21620 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_225
timestamp 1688980957
transform 1 0 21804 0 -1 17408
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_245
timestamp 1688980957
transform 1 0 23644 0 -1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_257
timestamp 1688980957
transform 1 0 24748 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_269
timestamp 1688980957
transform 1 0 25852 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_277
timestamp 1688980957
transform 1 0 26588 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_281
timestamp 1688980957
transform 1 0 26956 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_289
timestamp 1688980957
transform 1 0 27692 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_301
timestamp 1688980957
transform 1 0 28796 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_310
timestamp 1688980957
transform 1 0 29624 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_322
timestamp 1688980957
transform 1 0 30728 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_330
timestamp 1688980957
transform 1 0 31464 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_337
timestamp 1688980957
transform 1 0 32108 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_350
timestamp 1688980957
transform 1 0 33304 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_354
timestamp 1688980957
transform 1 0 33672 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_360
timestamp 1688980957
transform 1 0 34224 0 -1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_371
timestamp 1688980957
transform 1 0 35236 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_383
timestamp 1688980957
transform 1 0 36340 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_391
timestamp 1688980957
transform 1 0 37076 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_393
timestamp 1688980957
transform 1 0 37260 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_3
timestamp 1688980957
transform 1 0 1380 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_13
timestamp 1688980957
transform 1 0 2300 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_19
timestamp 1688980957
transform 1 0 2852 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_29
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_51
timestamp 1688980957
transform 1 0 5796 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_78
timestamp 1688980957
transform 1 0 8280 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_94
timestamp 1688980957
transform 1 0 9752 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_132
timestamp 1688980957
transform 1 0 13248 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_141
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_151
timestamp 1688980957
transform 1 0 14996 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_170
timestamp 1688980957
transform 1 0 16744 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_176
timestamp 1688980957
transform 1 0 17296 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_191
timestamp 1688980957
transform 1 0 18676 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_195
timestamp 1688980957
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_197
timestamp 1688980957
transform 1 0 19228 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_214
timestamp 1688980957
transform 1 0 20792 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_226
timestamp 1688980957
transform 1 0 21896 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_238
timestamp 1688980957
transform 1 0 23000 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_249
timestamp 1688980957
transform 1 0 24012 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_267
timestamp 1688980957
transform 1 0 25668 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_278
timestamp 1688980957
transform 1 0 26680 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_287
timestamp 1688980957
transform 1 0 27508 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_306
timestamp 1688980957
transform 1 0 29256 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_320
timestamp 1688980957
transform 1 0 30544 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_326
timestamp 1688980957
transform 1 0 31096 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_330
timestamp 1688980957
transform 1 0 31464 0 1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_339
timestamp 1688980957
transform 1 0 32292 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_351
timestamp 1688980957
transform 1 0 33396 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_359
timestamp 1688980957
transform 1 0 34132 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_363
timestamp 1688980957
transform 1 0 34500 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_365
timestamp 1688980957
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_377
timestamp 1688980957
transform 1 0 35788 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_389
timestamp 1688980957
transform 1 0 36892 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_3
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_36
timestamp 1688980957
transform 1 0 4416 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_48
timestamp 1688980957
transform 1 0 5520 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_57
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_69
timestamp 1688980957
transform 1 0 7452 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 1688980957
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_125
timestamp 1688980957
transform 1 0 12604 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_137
timestamp 1688980957
transform 1 0 13708 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_153
timestamp 1688980957
transform 1 0 15180 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_163
timestamp 1688980957
transform 1 0 16100 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_167
timestamp 1688980957
transform 1 0 16468 0 -1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_205
timestamp 1688980957
transform 1 0 19964 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_217
timestamp 1688980957
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_223
timestamp 1688980957
transform 1 0 21620 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_225
timestamp 1688980957
transform 1 0 21804 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_245
timestamp 1688980957
transform 1 0 23644 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_257
timestamp 1688980957
transform 1 0 24748 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_274
timestamp 1688980957
transform 1 0 26312 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_281
timestamp 1688980957
transform 1 0 26956 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_289
timestamp 1688980957
transform 1 0 27692 0 -1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_295
timestamp 1688980957
transform 1 0 28244 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_307
timestamp 1688980957
transform 1 0 29348 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_313
timestamp 1688980957
transform 1 0 29900 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_324
timestamp 1688980957
transform 1 0 30912 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_335
timestamp 1688980957
transform 1 0 31924 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_349
timestamp 1688980957
transform 1 0 33212 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_373
timestamp 1688980957
transform 1 0 35420 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_385
timestamp 1688980957
transform 1 0 36524 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_393
timestamp 1688980957
transform 1 0 37260 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_9
timestamp 1688980957
transform 1 0 1932 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_26
timestamp 1688980957
transform 1 0 3496 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_29
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_37
timestamp 1688980957
transform 1 0 4508 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_42
timestamp 1688980957
transform 1 0 4968 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_48
timestamp 1688980957
transform 1 0 5520 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_57
timestamp 1688980957
transform 1 0 6348 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_69
timestamp 1688980957
transform 1 0 7452 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_81
timestamp 1688980957
transform 1 0 8556 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_85
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_97
timestamp 1688980957
transform 1 0 10028 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_109
timestamp 1688980957
transform 1 0 11132 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_121
timestamp 1688980957
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_133
timestamp 1688980957
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 1688980957
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_141
timestamp 1688980957
transform 1 0 14076 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_147
timestamp 1688980957
transform 1 0 14628 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_159
timestamp 1688980957
transform 1 0 15732 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_171
timestamp 1688980957
transform 1 0 16836 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_177
timestamp 1688980957
transform 1 0 17388 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_191
timestamp 1688980957
transform 1 0 18676 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp 1688980957
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_204
timestamp 1688980957
transform 1 0 19872 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_219
timestamp 1688980957
transform 1 0 21252 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_235
timestamp 1688980957
transform 1 0 22724 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_247
timestamp 1688980957
transform 1 0 23828 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_251
timestamp 1688980957
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_253
timestamp 1688980957
transform 1 0 24380 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_265
timestamp 1688980957
transform 1 0 25484 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_277
timestamp 1688980957
transform 1 0 26588 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_289
timestamp 1688980957
transform 1 0 27692 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_301
timestamp 1688980957
transform 1 0 28796 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_307
timestamp 1688980957
transform 1 0 29348 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_309
timestamp 1688980957
transform 1 0 29532 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_321
timestamp 1688980957
transform 1 0 30636 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_328
timestamp 1688980957
transform 1 0 31280 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_332
timestamp 1688980957
transform 1 0 31648 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_347
timestamp 1688980957
transform 1 0 33028 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_351
timestamp 1688980957
transform 1 0 33396 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_355
timestamp 1688980957
transform 1 0 33764 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_363
timestamp 1688980957
transform 1 0 34500 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_369
timestamp 1688980957
transform 1 0 35052 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_381
timestamp 1688980957
transform 1 0 36156 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_392
timestamp 1688980957
transform 1 0 37168 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_400
timestamp 1688980957
transform 1 0 37904 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_23
timestamp 1688980957
transform 1 0 3220 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_31
timestamp 1688980957
transform 1 0 3956 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_53
timestamp 1688980957
transform 1 0 5980 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_57
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_63
timestamp 1688980957
transform 1 0 6900 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_67
timestamp 1688980957
transform 1 0 7268 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_82
timestamp 1688980957
transform 1 0 8648 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_95
timestamp 1688980957
transform 1 0 9844 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_107
timestamp 1688980957
transform 1 0 10948 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_136
timestamp 1688980957
transform 1 0 13616 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_140
timestamp 1688980957
transform 1 0 13984 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_150
timestamp 1688980957
transform 1 0 14904 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_162
timestamp 1688980957
transform 1 0 16008 0 -1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_190
timestamp 1688980957
transform 1 0 18584 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_205
timestamp 1688980957
transform 1 0 19964 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_217
timestamp 1688980957
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_223
timestamp 1688980957
transform 1 0 21620 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_225
timestamp 1688980957
transform 1 0 21804 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_253
timestamp 1688980957
transform 1 0 24380 0 -1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_265
timestamp 1688980957
transform 1 0 25484 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_277
timestamp 1688980957
transform 1 0 26588 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_281
timestamp 1688980957
transform 1 0 26956 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_296
timestamp 1688980957
transform 1 0 28336 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_302
timestamp 1688980957
transform 1 0 28888 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_317
timestamp 1688980957
transform 1 0 30268 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_329
timestamp 1688980957
transform 1 0 31372 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_335
timestamp 1688980957
transform 1 0 31924 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_337
timestamp 1688980957
transform 1 0 32108 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_345
timestamp 1688980957
transform 1 0 32844 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_349
timestamp 1688980957
transform 1 0 33212 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_368
timestamp 1688980957
transform 1 0 34960 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_376
timestamp 1688980957
transform 1 0 35696 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_380
timestamp 1688980957
transform 1 0 36064 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_393
timestamp 1688980957
transform 1 0 37260 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_3
timestamp 1688980957
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_10
timestamp 1688980957
transform 1 0 2024 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_25
timestamp 1688980957
transform 1 0 3404 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_81
timestamp 1688980957
transform 1 0 8556 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_85
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_102
timestamp 1688980957
transform 1 0 10488 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_110
timestamp 1688980957
transform 1 0 11224 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_122
timestamp 1688980957
transform 1 0 12328 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_150
timestamp 1688980957
transform 1 0 14904 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_161
timestamp 1688980957
transform 1 0 15916 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 1688980957
transform 1 0 19044 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_197
timestamp 1688980957
transform 1 0 19228 0 1 19584
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_216
timestamp 1688980957
transform 1 0 20976 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_228
timestamp 1688980957
transform 1 0 22080 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_256
timestamp 1688980957
transform 1 0 24656 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_282
timestamp 1688980957
transform 1 0 27048 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_294
timestamp 1688980957
transform 1 0 28152 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_306
timestamp 1688980957
transform 1 0 29256 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_316
timestamp 1688980957
transform 1 0 30176 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_340
timestamp 1688980957
transform 1 0 32384 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_348
timestamp 1688980957
transform 1 0 33120 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_354
timestamp 1688980957
transform 1 0 33672 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_362
timestamp 1688980957
transform 1 0 34408 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_365
timestamp 1688980957
transform 1 0 34684 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_389
timestamp 1688980957
transform 1 0 36892 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_3
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_11
timestamp 1688980957
transform 1 0 2116 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_23
timestamp 1688980957
transform 1 0 3220 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_32
timestamp 1688980957
transform 1 0 4048 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_44
timestamp 1688980957
transform 1 0 5152 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_57
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_65
timestamp 1688980957
transform 1 0 7084 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_75
timestamp 1688980957
transform 1 0 8004 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_87
timestamp 1688980957
transform 1 0 9108 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_99
timestamp 1688980957
transform 1 0 10212 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_111
timestamp 1688980957
transform 1 0 11316 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_120
timestamp 1688980957
transform 1 0 12144 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_132
timestamp 1688980957
transform 1 0 13248 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_140
timestamp 1688980957
transform 1 0 13984 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_150
timestamp 1688980957
transform 1 0 14904 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_162
timestamp 1688980957
transform 1 0 16008 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_169
timestamp 1688980957
transform 1 0 16652 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_177
timestamp 1688980957
transform 1 0 17388 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_200
timestamp 1688980957
transform 1 0 19504 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_221
timestamp 1688980957
transform 1 0 21436 0 -1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_225
timestamp 1688980957
transform 1 0 21804 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_237
timestamp 1688980957
transform 1 0 22908 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_249
timestamp 1688980957
transform 1 0 24012 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_257
timestamp 1688980957
transform 1 0 24748 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_264
timestamp 1688980957
transform 1 0 25392 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_275
timestamp 1688980957
transform 1 0 26404 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_279
timestamp 1688980957
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_281
timestamp 1688980957
transform 1 0 26956 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_291
timestamp 1688980957
transform 1 0 27876 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_299
timestamp 1688980957
transform 1 0 28612 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_305
timestamp 1688980957
transform 1 0 29164 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_326
timestamp 1688980957
transform 1 0 31096 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_334
timestamp 1688980957
transform 1 0 31832 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_337
timestamp 1688980957
transform 1 0 32108 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_345
timestamp 1688980957
transform 1 0 32844 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_353
timestamp 1688980957
transform 1 0 33580 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_365
timestamp 1688980957
transform 1 0 34684 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_380
timestamp 1688980957
transform 1 0 36064 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_393
timestamp 1688980957
transform 1 0 37260 0 -1 20672
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_9
timestamp 1688980957
transform 1 0 1932 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_21
timestamp 1688980957
transform 1 0 3036 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1688980957
transform 1 0 3588 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_36
timestamp 1688980957
transform 1 0 4416 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_44
timestamp 1688980957
transform 1 0 5152 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_50
timestamp 1688980957
transform 1 0 5704 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_62
timestamp 1688980957
transform 1 0 6808 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_75
timestamp 1688980957
transform 1 0 8004 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_83
timestamp 1688980957
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_99
timestamp 1688980957
transform 1 0 10212 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_111
timestamp 1688980957
transform 1 0 11316 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_123
timestamp 1688980957
transform 1 0 12420 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_135
timestamp 1688980957
transform 1 0 13524 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_139
timestamp 1688980957
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_167
timestamp 1688980957
transform 1 0 16468 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_179
timestamp 1688980957
transform 1 0 17572 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_187
timestamp 1688980957
transform 1 0 18308 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_197
timestamp 1688980957
transform 1 0 19228 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_201
timestamp 1688980957
transform 1 0 19596 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_210
timestamp 1688980957
transform 1 0 20424 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_237
timestamp 1688980957
transform 1 0 22908 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_249
timestamp 1688980957
transform 1 0 24012 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_253
timestamp 1688980957
transform 1 0 24380 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_257
timestamp 1688980957
transform 1 0 24748 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_264
timestamp 1688980957
transform 1 0 25392 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_276
timestamp 1688980957
transform 1 0 26496 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_291
timestamp 1688980957
transform 1 0 27876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_303
timestamp 1688980957
transform 1 0 28980 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_307
timestamp 1688980957
transform 1 0 29348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_309
timestamp 1688980957
transform 1 0 29532 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_315
timestamp 1688980957
transform 1 0 30084 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_322
timestamp 1688980957
transform 1 0 30728 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_334
timestamp 1688980957
transform 1 0 31832 0 1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_346
timestamp 1688980957
transform 1 0 32936 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_358
timestamp 1688980957
transform 1 0 34040 0 1 20672
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_376
timestamp 1688980957
transform 1 0 35696 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_388
timestamp 1688980957
transform 1 0 36800 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_40
timestamp 1688980957
transform 1 0 4784 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 1688980957
transform 1 0 6164 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_57
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_80
timestamp 1688980957
transform 1 0 8464 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_86
timestamp 1688980957
transform 1 0 9016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_101
timestamp 1688980957
transform 1 0 10396 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_109
timestamp 1688980957
transform 1 0 11132 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_122
timestamp 1688980957
transform 1 0 12328 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_128
timestamp 1688980957
transform 1 0 12880 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_144
timestamp 1688980957
transform 1 0 14352 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_148
timestamp 1688980957
transform 1 0 14720 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_158
timestamp 1688980957
transform 1 0 15640 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_166
timestamp 1688980957
transform 1 0 16376 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_169
timestamp 1688980957
transform 1 0 16652 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_175
timestamp 1688980957
transform 1 0 17204 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_190
timestamp 1688980957
transform 1 0 18584 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_210
timestamp 1688980957
transform 1 0 20424 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_222
timestamp 1688980957
transform 1 0 21528 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_225
timestamp 1688980957
transform 1 0 21804 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_233
timestamp 1688980957
transform 1 0 22540 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_245
timestamp 1688980957
transform 1 0 23644 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_257
timestamp 1688980957
transform 1 0 24748 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_268
timestamp 1688980957
transform 1 0 25760 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_281
timestamp 1688980957
transform 1 0 26956 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_285
timestamp 1688980957
transform 1 0 27324 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_290
timestamp 1688980957
transform 1 0 27784 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_302
timestamp 1688980957
transform 1 0 28888 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_310
timestamp 1688980957
transform 1 0 29624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_315
timestamp 1688980957
transform 1 0 30084 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_321
timestamp 1688980957
transform 1 0 30636 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_325
timestamp 1688980957
transform 1 0 31004 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_333
timestamp 1688980957
transform 1 0 31740 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_337
timestamp 1688980957
transform 1 0 32108 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_346
timestamp 1688980957
transform 1 0 32936 0 -1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_358
timestamp 1688980957
transform 1 0 34040 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_388
timestamp 1688980957
transform 1 0 36800 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_393
timestamp 1688980957
transform 1 0 37260 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_3
timestamp 1688980957
transform 1 0 1380 0 1 21760
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_10
timestamp 1688980957
transform 1 0 2024 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_22
timestamp 1688980957
transform 1 0 3128 0 1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_37
timestamp 1688980957
transform 1 0 4508 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_49
timestamp 1688980957
transform 1 0 5612 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_61
timestamp 1688980957
transform 1 0 6716 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_69
timestamp 1688980957
transform 1 0 7452 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_79
timestamp 1688980957
transform 1 0 8372 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_83
timestamp 1688980957
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_85
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_89
timestamp 1688980957
transform 1 0 9292 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_102
timestamp 1688980957
transform 1 0 10488 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_110
timestamp 1688980957
transform 1 0 11224 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_128
timestamp 1688980957
transform 1 0 12880 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_141
timestamp 1688980957
transform 1 0 14076 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_181
timestamp 1688980957
transform 1 0 17756 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_193
timestamp 1688980957
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_213
timestamp 1688980957
transform 1 0 20700 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_225
timestamp 1688980957
transform 1 0 21804 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_236
timestamp 1688980957
transform 1 0 22816 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_253
timestamp 1688980957
transform 1 0 24380 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_264
timestamp 1688980957
transform 1 0 25392 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_276
timestamp 1688980957
transform 1 0 26496 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_306
timestamp 1688980957
transform 1 0 29256 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_331
timestamp 1688980957
transform 1 0 31556 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_352
timestamp 1688980957
transform 1 0 33488 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_381
timestamp 1688980957
transform 1 0 36156 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_385
timestamp 1688980957
transform 1 0 36524 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_391
timestamp 1688980957
transform 1 0 37076 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_399
timestamp 1688980957
transform 1 0 37812 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_3
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_15
timestamp 1688980957
transform 1 0 2484 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_21
timestamp 1688980957
transform 1 0 3036 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_33
timestamp 1688980957
transform 1 0 4140 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_41
timestamp 1688980957
transform 1 0 4876 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_51
timestamp 1688980957
transform 1 0 5796 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_55
timestamp 1688980957
transform 1 0 6164 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_62
timestamp 1688980957
transform 1 0 6808 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_70
timestamp 1688980957
transform 1 0 7544 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_78
timestamp 1688980957
transform 1 0 8280 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_90
timestamp 1688980957
transform 1 0 9384 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_97
timestamp 1688980957
transform 1 0 10028 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_105
timestamp 1688980957
transform 1 0 10764 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_111
timestamp 1688980957
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_130
timestamp 1688980957
transform 1 0 13064 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_162
timestamp 1688980957
transform 1 0 16008 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_169
timestamp 1688980957
transform 1 0 16652 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_185
timestamp 1688980957
transform 1 0 18124 0 -1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_197
timestamp 1688980957
transform 1 0 19228 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_215
timestamp 1688980957
transform 1 0 20884 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_223
timestamp 1688980957
transform 1 0 21620 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_225
timestamp 1688980957
transform 1 0 21804 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_255
timestamp 1688980957
transform 1 0 24564 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_263
timestamp 1688980957
transform 1 0 25300 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_269
timestamp 1688980957
transform 1 0 25852 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_277
timestamp 1688980957
transform 1 0 26588 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_294
timestamp 1688980957
transform 1 0 28152 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_306
timestamp 1688980957
transform 1 0 29256 0 -1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_322
timestamp 1688980957
transform 1 0 30728 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_334
timestamp 1688980957
transform 1 0 31832 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_340
timestamp 1688980957
transform 1 0 32384 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_355
timestamp 1688980957
transform 1 0 33764 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_367
timestamp 1688980957
transform 1 0 34868 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_374
timestamp 1688980957
transform 1 0 35512 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_391
timestamp 1688980957
transform 1 0 37076 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_396
timestamp 1688980957
transform 1 0 37536 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_3
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_10
timestamp 1688980957
transform 1 0 2024 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_29
timestamp 1688980957
transform 1 0 3772 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_33
timestamp 1688980957
transform 1 0 4140 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_77
timestamp 1688980957
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 1688980957
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_85
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_96
timestamp 1688980957
transform 1 0 9936 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_128
timestamp 1688980957
transform 1 0 12880 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_146
timestamp 1688980957
transform 1 0 14536 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_162
timestamp 1688980957
transform 1 0 16008 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_193
timestamp 1688980957
transform 1 0 18860 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_197
timestamp 1688980957
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_209
timestamp 1688980957
transform 1 0 20332 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_215
timestamp 1688980957
transform 1 0 20884 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_229
timestamp 1688980957
transform 1 0 22172 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_249
timestamp 1688980957
transform 1 0 24012 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_253
timestamp 1688980957
transform 1 0 24380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_266
timestamp 1688980957
transform 1 0 25576 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_274
timestamp 1688980957
transform 1 0 26312 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_286
timestamp 1688980957
transform 1 0 27416 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_298
timestamp 1688980957
transform 1 0 28520 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_306
timestamp 1688980957
transform 1 0 29256 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_309
timestamp 1688980957
transform 1 0 29532 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_315
timestamp 1688980957
transform 1 0 30084 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_327
timestamp 1688980957
transform 1 0 31188 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_350
timestamp 1688980957
transform 1 0 33304 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_362
timestamp 1688980957
transform 1 0 34408 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_384
timestamp 1688980957
transform 1 0 36432 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_396
timestamp 1688980957
transform 1 0 37536 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_400
timestamp 1688980957
transform 1 0 37904 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_3
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_15
timestamp 1688980957
transform 1 0 2484 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_27
timestamp 1688980957
transform 1 0 3588 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_39
timestamp 1688980957
transform 1 0 4692 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_50
timestamp 1688980957
transform 1 0 5704 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_66
timestamp 1688980957
transform 1 0 7176 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_78
timestamp 1688980957
transform 1 0 8280 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_111
timestamp 1688980957
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_113
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_125
timestamp 1688980957
transform 1 0 12604 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_131
timestamp 1688980957
transform 1 0 13156 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_157
timestamp 1688980957
transform 1 0 15548 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_163
timestamp 1688980957
transform 1 0 16100 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_167
timestamp 1688980957
transform 1 0 16468 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_169
timestamp 1688980957
transform 1 0 16652 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_173
timestamp 1688980957
transform 1 0 17020 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_190
timestamp 1688980957
transform 1 0 18584 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_209
timestamp 1688980957
transform 1 0 20332 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_213
timestamp 1688980957
transform 1 0 20700 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_220
timestamp 1688980957
transform 1 0 21344 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_225
timestamp 1688980957
transform 1 0 21804 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_248
timestamp 1688980957
transform 1 0 23920 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_274
timestamp 1688980957
transform 1 0 26312 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_281
timestamp 1688980957
transform 1 0 26956 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_305
timestamp 1688980957
transform 1 0 29164 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_317
timestamp 1688980957
transform 1 0 30268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_39_329
timestamp 1688980957
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_335
timestamp 1688980957
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_340
timestamp 1688980957
transform 1 0 32384 0 -1 23936
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_351
timestamp 1688980957
transform 1 0 33396 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_363
timestamp 1688980957
transform 1 0 34500 0 -1 23936
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_380
timestamp 1688980957
transform 1 0 36064 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_393
timestamp 1688980957
transform 1 0 37260 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_3
timestamp 1688980957
transform 1 0 1380 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_10
timestamp 1688980957
transform 1 0 2024 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_22
timestamp 1688980957
transform 1 0 3128 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_38
timestamp 1688980957
transform 1 0 4600 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_44
timestamp 1688980957
transform 1 0 5152 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_65
timestamp 1688980957
transform 1 0 7084 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_73
timestamp 1688980957
transform 1 0 7820 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_77
timestamp 1688980957
transform 1 0 8188 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_83
timestamp 1688980957
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_88
timestamp 1688980957
transform 1 0 9200 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_100
timestamp 1688980957
transform 1 0 10304 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_112
timestamp 1688980957
transform 1 0 11408 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_124
timestamp 1688980957
transform 1 0 12512 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_130
timestamp 1688980957
transform 1 0 13064 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_134
timestamp 1688980957
transform 1 0 13432 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_141
timestamp 1688980957
transform 1 0 14076 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_155
timestamp 1688980957
transform 1 0 15364 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_167
timestamp 1688980957
transform 1 0 16468 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_179
timestamp 1688980957
transform 1 0 17572 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_215
timestamp 1688980957
transform 1 0 20884 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_253
timestamp 1688980957
transform 1 0 24380 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_264
timestamp 1688980957
transform 1 0 25392 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_287
timestamp 1688980957
transform 1 0 27508 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_291
timestamp 1688980957
transform 1 0 27876 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_301
timestamp 1688980957
transform 1 0 28796 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_307
timestamp 1688980957
transform 1 0 29348 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_317
timestamp 1688980957
transform 1 0 30268 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_341
timestamp 1688980957
transform 1 0 32476 0 1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_365
timestamp 1688980957
transform 1 0 34684 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_377
timestamp 1688980957
transform 1 0 35788 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_389
timestamp 1688980957
transform 1 0 36892 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_24
timestamp 1688980957
transform 1 0 3312 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_32
timestamp 1688980957
transform 1 0 4048 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_44
timestamp 1688980957
transform 1 0 5152 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_53
timestamp 1688980957
transform 1 0 5980 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_57
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_65
timestamp 1688980957
transform 1 0 7084 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_97
timestamp 1688980957
transform 1 0 10028 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_102
timestamp 1688980957
transform 1 0 10488 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_106
timestamp 1688980957
transform 1 0 10856 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_113
timestamp 1688980957
transform 1 0 11500 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_119
timestamp 1688980957
transform 1 0 12052 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_132
timestamp 1688980957
transform 1 0 13248 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_140
timestamp 1688980957
transform 1 0 13984 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_166
timestamp 1688980957
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_183
timestamp 1688980957
transform 1 0 17940 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_196
timestamp 1688980957
transform 1 0 19136 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_208
timestamp 1688980957
transform 1 0 20240 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_216
timestamp 1688980957
transform 1 0 20976 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_225
timestamp 1688980957
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_237
timestamp 1688980957
transform 1 0 22908 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_254
timestamp 1688980957
transform 1 0 24472 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_266
timestamp 1688980957
transform 1 0 25576 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_273
timestamp 1688980957
transform 1 0 26220 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_279
timestamp 1688980957
transform 1 0 26772 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_290
timestamp 1688980957
transform 1 0 27784 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_298
timestamp 1688980957
transform 1 0 28520 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_325
timestamp 1688980957
transform 1 0 31004 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_337
timestamp 1688980957
transform 1 0 32108 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_345
timestamp 1688980957
transform 1 0 32844 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_353
timestamp 1688980957
transform 1 0 33580 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_359
timestamp 1688980957
transform 1 0 34132 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_369
timestamp 1688980957
transform 1 0 35052 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_381
timestamp 1688980957
transform 1 0 36156 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_389
timestamp 1688980957
transform 1 0 36892 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_393
timestamp 1688980957
transform 1 0 37260 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_3
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_7
timestamp 1688980957
transform 1 0 1748 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_29
timestamp 1688980957
transform 1 0 3772 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_33
timestamp 1688980957
transform 1 0 4140 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_45
timestamp 1688980957
transform 1 0 5244 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_57
timestamp 1688980957
transform 1 0 6348 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_65
timestamp 1688980957
transform 1 0 7084 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_71
timestamp 1688980957
transform 1 0 7636 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_83
timestamp 1688980957
transform 1 0 8740 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_85
timestamp 1688980957
transform 1 0 8924 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_135
timestamp 1688980957
transform 1 0 13524 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_139
timestamp 1688980957
transform 1 0 13892 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_141
timestamp 1688980957
transform 1 0 14076 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_145
timestamp 1688980957
transform 1 0 14444 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_152
timestamp 1688980957
transform 1 0 15088 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_160
timestamp 1688980957
transform 1 0 15824 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_165
timestamp 1688980957
transform 1 0 16284 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_178
timestamp 1688980957
transform 1 0 17480 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_186
timestamp 1688980957
transform 1 0 18216 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_197
timestamp 1688980957
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_209
timestamp 1688980957
transform 1 0 20332 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_225
timestamp 1688980957
transform 1 0 21804 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_237
timestamp 1688980957
transform 1 0 22908 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_250
timestamp 1688980957
transform 1 0 24104 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_253
timestamp 1688980957
transform 1 0 24380 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_264
timestamp 1688980957
transform 1 0 25392 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_276
timestamp 1688980957
transform 1 0 26496 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_282
timestamp 1688980957
transform 1 0 27048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_291
timestamp 1688980957
transform 1 0 27876 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_306
timestamp 1688980957
transform 1 0 29256 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_309
timestamp 1688980957
transform 1 0 29532 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_313
timestamp 1688980957
transform 1 0 29900 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_322
timestamp 1688980957
transform 1 0 30728 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_334
timestamp 1688980957
transform 1 0 31832 0 1 25024
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_346
timestamp 1688980957
transform 1 0 32936 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_358
timestamp 1688980957
transform 1 0 34040 0 1 25024
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_388
timestamp 1688980957
transform 1 0 36800 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_400
timestamp 1688980957
transform 1 0 37904 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_9
timestamp 1688980957
transform 1 0 1932 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_17
timestamp 1688980957
transform 1 0 2668 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_22
timestamp 1688980957
transform 1 0 3128 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_44
timestamp 1688980957
transform 1 0 5152 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_50
timestamp 1688980957
transform 1 0 5704 0 -1 26112
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_57
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_69
timestamp 1688980957
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_81
timestamp 1688980957
transform 1 0 8556 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_103
timestamp 1688980957
transform 1 0 10580 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_111
timestamp 1688980957
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_113
timestamp 1688980957
transform 1 0 11500 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_125
timestamp 1688980957
transform 1 0 12604 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_137
timestamp 1688980957
transform 1 0 13708 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_149
timestamp 1688980957
transform 1 0 14812 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_161
timestamp 1688980957
transform 1 0 15916 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_167
timestamp 1688980957
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_169
timestamp 1688980957
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_181
timestamp 1688980957
transform 1 0 17756 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_204
timestamp 1688980957
transform 1 0 19872 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_217
timestamp 1688980957
transform 1 0 21068 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_223
timestamp 1688980957
transform 1 0 21620 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_225
timestamp 1688980957
transform 1 0 21804 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_229
timestamp 1688980957
transform 1 0 22172 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_253
timestamp 1688980957
transform 1 0 24380 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_278
timestamp 1688980957
transform 1 0 26680 0 -1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_281
timestamp 1688980957
transform 1 0 26956 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_293
timestamp 1688980957
transform 1 0 28060 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_305
timestamp 1688980957
transform 1 0 29164 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_317
timestamp 1688980957
transform 1 0 30268 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_329
timestamp 1688980957
transform 1 0 31372 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_354
timestamp 1688980957
transform 1 0 33672 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_373
timestamp 1688980957
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_385
timestamp 1688980957
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_391
timestamp 1688980957
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_393
timestamp 1688980957
transform 1 0 37260 0 -1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_3
timestamp 1688980957
transform 1 0 1380 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_15
timestamp 1688980957
transform 1 0 2484 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_27
timestamp 1688980957
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_29
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_88
timestamp 1688980957
transform 1 0 9200 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_100
timestamp 1688980957
transform 1 0 10304 0 1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_112
timestamp 1688980957
transform 1 0 11408 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_124
timestamp 1688980957
transform 1 0 12512 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_141
timestamp 1688980957
transform 1 0 14076 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_159
timestamp 1688980957
transform 1 0 15732 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_167
timestamp 1688980957
transform 1 0 16468 0 1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_178
timestamp 1688980957
transform 1 0 17480 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_190
timestamp 1688980957
transform 1 0 18584 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_197
timestamp 1688980957
transform 1 0 19228 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_205
timestamp 1688980957
transform 1 0 19964 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_213
timestamp 1688980957
transform 1 0 20700 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_221
timestamp 1688980957
transform 1 0 21436 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_233
timestamp 1688980957
transform 1 0 22540 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_241
timestamp 1688980957
transform 1 0 23276 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_248
timestamp 1688980957
transform 1 0 23920 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_253
timestamp 1688980957
transform 1 0 24380 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_261
timestamp 1688980957
transform 1 0 25116 0 1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_278
timestamp 1688980957
transform 1 0 26680 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_299
timestamp 1688980957
transform 1 0 28612 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_307
timestamp 1688980957
transform 1 0 29348 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_318
timestamp 1688980957
transform 1 0 30360 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_348
timestamp 1688980957
transform 1 0 33120 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_358
timestamp 1688980957
transform 1 0 34040 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_391
timestamp 1688980957
transform 1 0 37076 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_399
timestamp 1688980957
transform 1 0 37812 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_3
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_15
timestamp 1688980957
transform 1 0 2484 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_27
timestamp 1688980957
transform 1 0 3588 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_39
timestamp 1688980957
transform 1 0 4692 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_51
timestamp 1688980957
transform 1 0 5796 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1688980957
transform 1 0 6164 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_57
timestamp 1688980957
transform 1 0 6348 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_81
timestamp 1688980957
transform 1 0 8556 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_93
timestamp 1688980957
transform 1 0 9660 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_102
timestamp 1688980957
transform 1 0 10488 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_110
timestamp 1688980957
transform 1 0 11224 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_113
timestamp 1688980957
transform 1 0 11500 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_129
timestamp 1688980957
transform 1 0 12972 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_141
timestamp 1688980957
transform 1 0 14076 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_151
timestamp 1688980957
transform 1 0 14996 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_155
timestamp 1688980957
transform 1 0 15364 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_160
timestamp 1688980957
transform 1 0 15824 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_176
timestamp 1688980957
transform 1 0 17296 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_185
timestamp 1688980957
transform 1 0 18124 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_191
timestamp 1688980957
transform 1 0 18676 0 -1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_197
timestamp 1688980957
transform 1 0 19228 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_209
timestamp 1688980957
transform 1 0 20332 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_221
timestamp 1688980957
transform 1 0 21436 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_225
timestamp 1688980957
transform 1 0 21804 0 -1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_236
timestamp 1688980957
transform 1 0 22816 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_248
timestamp 1688980957
transform 1 0 23920 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_260
timestamp 1688980957
transform 1 0 25024 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_268
timestamp 1688980957
transform 1 0 25760 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_284
timestamp 1688980957
transform 1 0 27232 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_329
timestamp 1688980957
transform 1 0 31372 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_333
timestamp 1688980957
transform 1 0 31740 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_337
timestamp 1688980957
transform 1 0 32108 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_345
timestamp 1688980957
transform 1 0 32844 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_374
timestamp 1688980957
transform 1 0 35512 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_45_386
timestamp 1688980957
transform 1 0 36616 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_393
timestamp 1688980957
transform 1 0 37260 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_3
timestamp 1688980957
transform 1 0 1380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_15
timestamp 1688980957
transform 1 0 2484 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1688980957
transform 1 0 3588 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_29
timestamp 1688980957
transform 1 0 3772 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_37
timestamp 1688980957
transform 1 0 4508 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_41
timestamp 1688980957
transform 1 0 4876 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_53
timestamp 1688980957
transform 1 0 5980 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_64
timestamp 1688980957
transform 1 0 6992 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_76
timestamp 1688980957
transform 1 0 8096 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_81
timestamp 1688980957
transform 1 0 8556 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_85
timestamp 1688980957
transform 1 0 8924 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_123
timestamp 1688980957
transform 1 0 12420 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_133
timestamp 1688980957
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_139
timestamp 1688980957
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_148
timestamp 1688980957
transform 1 0 14720 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_156
timestamp 1688980957
transform 1 0 15456 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_163
timestamp 1688980957
transform 1 0 16100 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_194
timestamp 1688980957
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_197
timestamp 1688980957
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_209
timestamp 1688980957
transform 1 0 20332 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_221
timestamp 1688980957
transform 1 0 21436 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_233
timestamp 1688980957
transform 1 0 22540 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_247
timestamp 1688980957
transform 1 0 23828 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_251
timestamp 1688980957
transform 1 0 24196 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_253
timestamp 1688980957
transform 1 0 24380 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_295
timestamp 1688980957
transform 1 0 28244 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_307
timestamp 1688980957
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_315
timestamp 1688980957
transform 1 0 30084 0 1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_326
timestamp 1688980957
transform 1 0 31096 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_338
timestamp 1688980957
transform 1 0 32200 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_350
timestamp 1688980957
transform 1 0 33304 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_358
timestamp 1688980957
transform 1 0 34040 0 1 27200
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_365
timestamp 1688980957
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_377
timestamp 1688980957
transform 1 0 35788 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_389
timestamp 1688980957
transform 1 0 36892 0 1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_3
timestamp 1688980957
transform 1 0 1380 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_15
timestamp 1688980957
transform 1 0 2484 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_27
timestamp 1688980957
transform 1 0 3588 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_31
timestamp 1688980957
transform 1 0 3956 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_53
timestamp 1688980957
transform 1 0 5980 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_66
timestamp 1688980957
transform 1 0 7176 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_70
timestamp 1688980957
transform 1 0 7544 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_101
timestamp 1688980957
transform 1 0 10396 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_106
timestamp 1688980957
transform 1 0 10856 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_122
timestamp 1688980957
transform 1 0 12328 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_130
timestamp 1688980957
transform 1 0 13064 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_134
timestamp 1688980957
transform 1 0 13432 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_151
timestamp 1688980957
transform 1 0 14996 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_163
timestamp 1688980957
transform 1 0 16100 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_167
timestamp 1688980957
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_177
timestamp 1688980957
transform 1 0 17388 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_189
timestamp 1688980957
transform 1 0 18492 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_222
timestamp 1688980957
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_255
timestamp 1688980957
transform 1 0 24564 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_267
timestamp 1688980957
transform 1 0 25668 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_279
timestamp 1688980957
transform 1 0 26772 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_281
timestamp 1688980957
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_293
timestamp 1688980957
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_305
timestamp 1688980957
transform 1 0 29164 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_317
timestamp 1688980957
transform 1 0 30268 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_329
timestamp 1688980957
transform 1 0 31372 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_337
timestamp 1688980957
transform 1 0 32108 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_347
timestamp 1688980957
transform 1 0 33028 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_359
timestamp 1688980957
transform 1 0 34132 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_363
timestamp 1688980957
transform 1 0 34500 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_369
timestamp 1688980957
transform 1 0 35052 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_381
timestamp 1688980957
transform 1 0 36156 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_389
timestamp 1688980957
transform 1 0 36892 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_393
timestamp 1688980957
transform 1 0 37260 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_397
timestamp 1688980957
transform 1 0 37628 0 -1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_3
timestamp 1688980957
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_15
timestamp 1688980957
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_27
timestamp 1688980957
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_29
timestamp 1688980957
transform 1 0 3772 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_36
timestamp 1688980957
transform 1 0 4416 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_40
timestamp 1688980957
transform 1 0 4784 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_79
timestamp 1688980957
transform 1 0 8372 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_83
timestamp 1688980957
transform 1 0 8740 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_85
timestamp 1688980957
transform 1 0 8924 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_93
timestamp 1688980957
transform 1 0 9660 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_119
timestamp 1688980957
transform 1 0 12052 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_131
timestamp 1688980957
transform 1 0 13156 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_139
timestamp 1688980957
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_141
timestamp 1688980957
transform 1 0 14076 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_153
timestamp 1688980957
transform 1 0 15180 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_161
timestamp 1688980957
transform 1 0 15916 0 1 28288
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_170
timestamp 1688980957
transform 1 0 16744 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_182
timestamp 1688980957
transform 1 0 17848 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_194
timestamp 1688980957
transform 1 0 18952 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_197
timestamp 1688980957
transform 1 0 19228 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_207
timestamp 1688980957
transform 1 0 20148 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_213
timestamp 1688980957
transform 1 0 20700 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_234
timestamp 1688980957
transform 1 0 22632 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_246
timestamp 1688980957
transform 1 0 23736 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_260
timestamp 1688980957
transform 1 0 25024 0 1 28288
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_275
timestamp 1688980957
transform 1 0 26404 0 1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_287
timestamp 1688980957
transform 1 0 27508 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_299
timestamp 1688980957
transform 1 0 28612 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_303
timestamp 1688980957
transform 1 0 28980 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_307
timestamp 1688980957
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_332
timestamp 1688980957
transform 1 0 31648 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_354
timestamp 1688980957
transform 1 0 33672 0 1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_386
timestamp 1688980957
transform 1 0 36616 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_398
timestamp 1688980957
transform 1 0 37720 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_3
timestamp 1688980957
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_15
timestamp 1688980957
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_27
timestamp 1688980957
transform 1 0 3588 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_53
timestamp 1688980957
transform 1 0 5980 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_57
timestamp 1688980957
transform 1 0 6348 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_68
timestamp 1688980957
transform 1 0 7360 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_79
timestamp 1688980957
transform 1 0 8372 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_113
timestamp 1688980957
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_125
timestamp 1688980957
transform 1 0 12604 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_133
timestamp 1688980957
transform 1 0 13340 0 -1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_145
timestamp 1688980957
transform 1 0 14444 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_157
timestamp 1688980957
transform 1 0 15548 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_165
timestamp 1688980957
transform 1 0 16284 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_169
timestamp 1688980957
transform 1 0 16652 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_181
timestamp 1688980957
transform 1 0 17756 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_194
timestamp 1688980957
transform 1 0 18952 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_206
timestamp 1688980957
transform 1 0 20056 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_212
timestamp 1688980957
transform 1 0 20608 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_220
timestamp 1688980957
transform 1 0 21344 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_241
timestamp 1688980957
transform 1 0 23276 0 -1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_250
timestamp 1688980957
transform 1 0 24104 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_262
timestamp 1688980957
transform 1 0 25208 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_281
timestamp 1688980957
transform 1 0 26956 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_326
timestamp 1688980957
transform 1 0 31096 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_348
timestamp 1688980957
transform 1 0 33120 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_360
timestamp 1688980957
transform 1 0 34224 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_370
timestamp 1688980957
transform 1 0 35144 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_382
timestamp 1688980957
transform 1 0 36248 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_391
timestamp 1688980957
transform 1 0 37076 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_393
timestamp 1688980957
transform 1 0 37260 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_3
timestamp 1688980957
transform 1 0 1380 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_15
timestamp 1688980957
transform 1 0 2484 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 1688980957
transform 1 0 3588 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_29
timestamp 1688980957
transform 1 0 3772 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_34
timestamp 1688980957
transform 1 0 4232 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_46
timestamp 1688980957
transform 1 0 5336 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_56
timestamp 1688980957
transform 1 0 6256 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_68
timestamp 1688980957
transform 1 0 7360 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_76
timestamp 1688980957
transform 1 0 8096 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_106
timestamp 1688980957
transform 1 0 10856 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_118
timestamp 1688980957
transform 1 0 11960 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_129
timestamp 1688980957
transform 1 0 12972 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_139
timestamp 1688980957
transform 1 0 13892 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_149
timestamp 1688980957
transform 1 0 14812 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_166
timestamp 1688980957
transform 1 0 16376 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_176
timestamp 1688980957
transform 1 0 17296 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_184
timestamp 1688980957
transform 1 0 18032 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_194
timestamp 1688980957
transform 1 0 18952 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_197
timestamp 1688980957
transform 1 0 19228 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_209
timestamp 1688980957
transform 1 0 20332 0 1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_219
timestamp 1688980957
transform 1 0 21252 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_231
timestamp 1688980957
transform 1 0 22356 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_243
timestamp 1688980957
transform 1 0 23460 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_250
timestamp 1688980957
transform 1 0 24104 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_258
timestamp 1688980957
transform 1 0 24840 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_264
timestamp 1688980957
transform 1 0 25392 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_280
timestamp 1688980957
transform 1 0 26864 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_299
timestamp 1688980957
transform 1 0 28612 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_325
timestamp 1688980957
transform 1 0 31004 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_347
timestamp 1688980957
transform 1 0 33028 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_365
timestamp 1688980957
transform 1 0 34684 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_389
timestamp 1688980957
transform 1 0 36892 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_3
timestamp 1688980957
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_15
timestamp 1688980957
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_27
timestamp 1688980957
transform 1 0 3588 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_33
timestamp 1688980957
transform 1 0 4140 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_55
timestamp 1688980957
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_57
timestamp 1688980957
transform 1 0 6348 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_76
timestamp 1688980957
transform 1 0 8096 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_80
timestamp 1688980957
transform 1 0 8464 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_84
timestamp 1688980957
transform 1 0 8832 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_96
timestamp 1688980957
transform 1 0 9936 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_108
timestamp 1688980957
transform 1 0 11040 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_113
timestamp 1688980957
transform 1 0 11500 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_122
timestamp 1688980957
transform 1 0 12328 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_128
timestamp 1688980957
transform 1 0 12880 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_149
timestamp 1688980957
transform 1 0 14812 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_161
timestamp 1688980957
transform 1 0 15916 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_167
timestamp 1688980957
transform 1 0 16468 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_169
timestamp 1688980957
transform 1 0 16652 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_177
timestamp 1688980957
transform 1 0 17388 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_193
timestamp 1688980957
transform 1 0 18860 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_201
timestamp 1688980957
transform 1 0 19596 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_216
timestamp 1688980957
transform 1 0 20976 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_225
timestamp 1688980957
transform 1 0 21804 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_237
timestamp 1688980957
transform 1 0 22908 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_241
timestamp 1688980957
transform 1 0 23276 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_262
timestamp 1688980957
transform 1 0 25208 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_266
timestamp 1688980957
transform 1 0 25576 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_274
timestamp 1688980957
transform 1 0 26312 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_281
timestamp 1688980957
transform 1 0 26956 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_51_293
timestamp 1688980957
transform 1 0 28060 0 -1 30464
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_319
timestamp 1688980957
transform 1 0 30452 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_331
timestamp 1688980957
transform 1 0 31556 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_335
timestamp 1688980957
transform 1 0 31924 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_345
timestamp 1688980957
transform 1 0 32844 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_357
timestamp 1688980957
transform 1 0 33948 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_369
timestamp 1688980957
transform 1 0 35052 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_381
timestamp 1688980957
transform 1 0 36156 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_389
timestamp 1688980957
transform 1 0 36892 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_393
timestamp 1688980957
transform 1 0 37260 0 -1 30464
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_3
timestamp 1688980957
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_15
timestamp 1688980957
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_27
timestamp 1688980957
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_29
timestamp 1688980957
transform 1 0 3772 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_38
timestamp 1688980957
transform 1 0 4600 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_46
timestamp 1688980957
transform 1 0 5336 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_82
timestamp 1688980957
transform 1 0 8648 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_94
timestamp 1688980957
transform 1 0 9752 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_106
timestamp 1688980957
transform 1 0 10856 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_118
timestamp 1688980957
transform 1 0 11960 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_130
timestamp 1688980957
transform 1 0 13064 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_150
timestamp 1688980957
transform 1 0 14904 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_162
timestamp 1688980957
transform 1 0 16008 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_225
timestamp 1688980957
transform 1 0 21804 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_237
timestamp 1688980957
transform 1 0 22908 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_249
timestamp 1688980957
transform 1 0 24012 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_253
timestamp 1688980957
transform 1 0 24380 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_259
timestamp 1688980957
transform 1 0 24932 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_278
timestamp 1688980957
transform 1 0 26680 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_290
timestamp 1688980957
transform 1 0 27784 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_302
timestamp 1688980957
transform 1 0 28888 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_309
timestamp 1688980957
transform 1 0 29532 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_344
timestamp 1688980957
transform 1 0 32752 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_359
timestamp 1688980957
transform 1 0 34132 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_363
timestamp 1688980957
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_374
timestamp 1688980957
transform 1 0 35512 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_386
timestamp 1688980957
transform 1 0 36616 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_398
timestamp 1688980957
transform 1 0 37720 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_3
timestamp 1688980957
transform 1 0 1380 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_15
timestamp 1688980957
transform 1 0 2484 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_27
timestamp 1688980957
transform 1 0 3588 0 -1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_39
timestamp 1688980957
transform 1 0 4692 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_51
timestamp 1688980957
transform 1 0 5796 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_55
timestamp 1688980957
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_57
timestamp 1688980957
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_69
timestamp 1688980957
transform 1 0 7452 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_94
timestamp 1688980957
transform 1 0 9752 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_107
timestamp 1688980957
transform 1 0 10948 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_111
timestamp 1688980957
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_120
timestamp 1688980957
transform 1 0 12144 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_128
timestamp 1688980957
transform 1 0 12880 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_149
timestamp 1688980957
transform 1 0 14812 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_184
timestamp 1688980957
transform 1 0 18032 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_193
timestamp 1688980957
transform 1 0 18860 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_206
timestamp 1688980957
transform 1 0 20056 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_223
timestamp 1688980957
transform 1 0 21620 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_232
timestamp 1688980957
transform 1 0 22448 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_279
timestamp 1688980957
transform 1 0 26772 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_337
timestamp 1688980957
transform 1 0 32108 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_386
timestamp 1688980957
transform 1 0 36616 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_393
timestamp 1688980957
transform 1 0 37260 0 -1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_3
timestamp 1688980957
transform 1 0 1380 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_15
timestamp 1688980957
transform 1 0 2484 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_27
timestamp 1688980957
transform 1 0 3588 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_29
timestamp 1688980957
transform 1 0 3772 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_57
timestamp 1688980957
transform 1 0 6348 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_77
timestamp 1688980957
transform 1 0 8188 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_81
timestamp 1688980957
transform 1 0 8556 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_85
timestamp 1688980957
transform 1 0 8924 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_111
timestamp 1688980957
transform 1 0 11316 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_123
timestamp 1688980957
transform 1 0 12420 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_129
timestamp 1688980957
transform 1 0 12972 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_137
timestamp 1688980957
transform 1 0 13708 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_141
timestamp 1688980957
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_153
timestamp 1688980957
transform 1 0 15180 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_165
timestamp 1688980957
transform 1 0 16284 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_177
timestamp 1688980957
transform 1 0 17388 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_189
timestamp 1688980957
transform 1 0 18492 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_197
timestamp 1688980957
transform 1 0 19228 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_220
timestamp 1688980957
transform 1 0 21344 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_250
timestamp 1688980957
transform 1 0 24104 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_267
timestamp 1688980957
transform 1 0 25668 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_277
timestamp 1688980957
transform 1 0 26588 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_282
timestamp 1688980957
transform 1 0 27048 0 1 31552
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_296
timestamp 1688980957
transform 1 0 28336 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_320
timestamp 1688980957
transform 1 0 30544 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_328
timestamp 1688980957
transform 1 0 31280 0 1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_336
timestamp 1688980957
transform 1 0 32016 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_348
timestamp 1688980957
transform 1 0 33120 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_360
timestamp 1688980957
transform 1 0 34224 0 1 31552
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_374
timestamp 1688980957
transform 1 0 35512 0 1 31552
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_386
timestamp 1688980957
transform 1 0 36616 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_398
timestamp 1688980957
transform 1 0 37720 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_3
timestamp 1688980957
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_15
timestamp 1688980957
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_27
timestamp 1688980957
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_39
timestamp 1688980957
transform 1 0 4692 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_45
timestamp 1688980957
transform 1 0 5244 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_53
timestamp 1688980957
transform 1 0 5980 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_57
timestamp 1688980957
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_69
timestamp 1688980957
transform 1 0 7452 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_81
timestamp 1688980957
transform 1 0 8556 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_93
timestamp 1688980957
transform 1 0 9660 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_105
timestamp 1688980957
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_111
timestamp 1688980957
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_120
timestamp 1688980957
transform 1 0 12144 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_126
timestamp 1688980957
transform 1 0 12696 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_138
timestamp 1688980957
transform 1 0 13800 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_150
timestamp 1688980957
transform 1 0 14904 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_162
timestamp 1688980957
transform 1 0 16008 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_175
timestamp 1688980957
transform 1 0 17204 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_182
timestamp 1688980957
transform 1 0 17848 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_186
timestamp 1688980957
transform 1 0 18216 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_195
timestamp 1688980957
transform 1 0 19044 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_199
timestamp 1688980957
transform 1 0 19412 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_220
timestamp 1688980957
transform 1 0 21344 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_231
timestamp 1688980957
transform 1 0 22356 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_235
timestamp 1688980957
transform 1 0 22724 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_243
timestamp 1688980957
transform 1 0 23460 0 -1 32640
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_253
timestamp 1688980957
transform 1 0 24380 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_265
timestamp 1688980957
transform 1 0 25484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_277
timestamp 1688980957
transform 1 0 26588 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_281
timestamp 1688980957
transform 1 0 26956 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_292
timestamp 1688980957
transform 1 0 27968 0 -1 32640
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_306
timestamp 1688980957
transform 1 0 29256 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_318
timestamp 1688980957
transform 1 0 30360 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_331
timestamp 1688980957
transform 1 0 31556 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_335
timestamp 1688980957
transform 1 0 31924 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_354
timestamp 1688980957
transform 1 0 33672 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_366
timestamp 1688980957
transform 1 0 34776 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_374
timestamp 1688980957
transform 1 0 35512 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_380
timestamp 1688980957
transform 1 0 36064 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_393
timestamp 1688980957
transform 1 0 37260 0 -1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_3
timestamp 1688980957
transform 1 0 1380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_15
timestamp 1688980957
transform 1 0 2484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_27
timestamp 1688980957
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_29
timestamp 1688980957
transform 1 0 3772 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_65
timestamp 1688980957
transform 1 0 7084 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_81
timestamp 1688980957
transform 1 0 8556 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_85
timestamp 1688980957
transform 1 0 8924 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_89
timestamp 1688980957
transform 1 0 9292 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_99
timestamp 1688980957
transform 1 0 10212 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_111
timestamp 1688980957
transform 1 0 11316 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_123
timestamp 1688980957
transform 1 0 12420 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_135
timestamp 1688980957
transform 1 0 13524 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_139
timestamp 1688980957
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_141
timestamp 1688980957
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_153
timestamp 1688980957
transform 1 0 15180 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_161
timestamp 1688980957
transform 1 0 15916 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_179
timestamp 1688980957
transform 1 0 17572 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_193
timestamp 1688980957
transform 1 0 18860 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_197
timestamp 1688980957
transform 1 0 19228 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_205
timestamp 1688980957
transform 1 0 19964 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_214
timestamp 1688980957
transform 1 0 20792 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_231
timestamp 1688980957
transform 1 0 22356 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_239
timestamp 1688980957
transform 1 0 23092 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_245
timestamp 1688980957
transform 1 0 23644 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_251
timestamp 1688980957
transform 1 0 24196 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_253
timestamp 1688980957
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_265
timestamp 1688980957
transform 1 0 25484 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_286
timestamp 1688980957
transform 1 0 27416 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_309
timestamp 1688980957
transform 1 0 29532 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_315
timestamp 1688980957
transform 1 0 30084 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_319
timestamp 1688980957
transform 1 0 30452 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_323
timestamp 1688980957
transform 1 0 30820 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_348
timestamp 1688980957
transform 1 0 33120 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_360
timestamp 1688980957
transform 1 0 34224 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_388
timestamp 1688980957
transform 1 0 36800 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_400
timestamp 1688980957
transform 1 0 37904 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_3
timestamp 1688980957
transform 1 0 1380 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_15
timestamp 1688980957
transform 1 0 2484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_27
timestamp 1688980957
transform 1 0 3588 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_39
timestamp 1688980957
transform 1 0 4692 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_57
timestamp 1688980957
transform 1 0 6348 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_63
timestamp 1688980957
transform 1 0 6900 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_106
timestamp 1688980957
transform 1 0 10856 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_113
timestamp 1688980957
transform 1 0 11500 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_125
timestamp 1688980957
transform 1 0 12604 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_137
timestamp 1688980957
transform 1 0 13708 0 -1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_147
timestamp 1688980957
transform 1 0 14628 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_159
timestamp 1688980957
transform 1 0 15732 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_167
timestamp 1688980957
transform 1 0 16468 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_169
timestamp 1688980957
transform 1 0 16652 0 -1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_180
timestamp 1688980957
transform 1 0 17664 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_192
timestamp 1688980957
transform 1 0 18768 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_222
timestamp 1688980957
transform 1 0 21528 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_228
timestamp 1688980957
transform 1 0 22080 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_240
timestamp 1688980957
transform 1 0 23184 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_251
timestamp 1688980957
transform 1 0 24196 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_257
timestamp 1688980957
transform 1 0 24748 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_265
timestamp 1688980957
transform 1 0 25484 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_304
timestamp 1688980957
transform 1 0 29072 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_316
timestamp 1688980957
transform 1 0 30176 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_328
timestamp 1688980957
transform 1 0 31280 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_337
timestamp 1688980957
transform 1 0 32108 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_345
timestamp 1688980957
transform 1 0 32844 0 -1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_368
timestamp 1688980957
transform 1 0 34960 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_380
timestamp 1688980957
transform 1 0 36064 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_386
timestamp 1688980957
transform 1 0 36616 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_390
timestamp 1688980957
transform 1 0 36984 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_393
timestamp 1688980957
transform 1 0 37260 0 -1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_3
timestamp 1688980957
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_15
timestamp 1688980957
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_27
timestamp 1688980957
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_29
timestamp 1688980957
transform 1 0 3772 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_37
timestamp 1688980957
transform 1 0 4508 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_63
timestamp 1688980957
transform 1 0 6900 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_68
timestamp 1688980957
transform 1 0 7360 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_80
timestamp 1688980957
transform 1 0 8464 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_96
timestamp 1688980957
transform 1 0 9936 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_108
timestamp 1688980957
transform 1 0 11040 0 1 33728
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_118
timestamp 1688980957
transform 1 0 11960 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_130
timestamp 1688980957
transform 1 0 13064 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_138
timestamp 1688980957
transform 1 0 13800 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_141
timestamp 1688980957
transform 1 0 14076 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_153
timestamp 1688980957
transform 1 0 15180 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_170
timestamp 1688980957
transform 1 0 16744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_178
timestamp 1688980957
transform 1 0 17480 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_195
timestamp 1688980957
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_201
timestamp 1688980957
transform 1 0 19596 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_211
timestamp 1688980957
transform 1 0 20516 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_229
timestamp 1688980957
transform 1 0 22172 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_248
timestamp 1688980957
transform 1 0 23920 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_253
timestamp 1688980957
transform 1 0 24380 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_261
timestamp 1688980957
transform 1 0 25116 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_278
timestamp 1688980957
transform 1 0 26680 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_285
timestamp 1688980957
transform 1 0 27324 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_294
timestamp 1688980957
transform 1 0 28152 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_306
timestamp 1688980957
transform 1 0 29256 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_309
timestamp 1688980957
transform 1 0 29532 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_317
timestamp 1688980957
transform 1 0 30268 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_327
timestamp 1688980957
transform 1 0 31188 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_336
timestamp 1688980957
transform 1 0 32016 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_348
timestamp 1688980957
transform 1 0 33120 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_359
timestamp 1688980957
transform 1 0 34132 0 1 33728
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_388
timestamp 1688980957
transform 1 0 36800 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_400
timestamp 1688980957
transform 1 0 37904 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_3
timestamp 1688980957
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_15
timestamp 1688980957
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_27
timestamp 1688980957
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_39
timestamp 1688980957
transform 1 0 4692 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_50
timestamp 1688980957
transform 1 0 5704 0 -1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_57
timestamp 1688980957
transform 1 0 6348 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_69
timestamp 1688980957
transform 1 0 7452 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_83
timestamp 1688980957
transform 1 0 8740 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_95
timestamp 1688980957
transform 1 0 9844 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_107
timestamp 1688980957
transform 1 0 10948 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_111
timestamp 1688980957
transform 1 0 11316 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_121
timestamp 1688980957
transform 1 0 12236 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_133
timestamp 1688980957
transform 1 0 13340 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_145
timestamp 1688980957
transform 1 0 14444 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_157
timestamp 1688980957
transform 1 0 15548 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_165
timestamp 1688980957
transform 1 0 16284 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_177
timestamp 1688980957
transform 1 0 17388 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_189
timestamp 1688980957
transform 1 0 18492 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_201
timestamp 1688980957
transform 1 0 19596 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_213
timestamp 1688980957
transform 1 0 20700 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_221
timestamp 1688980957
transform 1 0 21436 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_225
timestamp 1688980957
transform 1 0 21804 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_234
timestamp 1688980957
transform 1 0 22632 0 -1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_249
timestamp 1688980957
transform 1 0 24012 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_261
timestamp 1688980957
transform 1 0 25116 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_273
timestamp 1688980957
transform 1 0 26220 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_279
timestamp 1688980957
transform 1 0 26772 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_281
timestamp 1688980957
transform 1 0 26956 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_293
timestamp 1688980957
transform 1 0 28060 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_320
timestamp 1688980957
transform 1 0 30544 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_326
timestamp 1688980957
transform 1 0 31096 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_337
timestamp 1688980957
transform 1 0 32108 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_345
timestamp 1688980957
transform 1 0 32844 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_355
timestamp 1688980957
transform 1 0 33764 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_367
timestamp 1688980957
transform 1 0 34868 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_379
timestamp 1688980957
transform 1 0 35972 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_391
timestamp 1688980957
transform 1 0 37076 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_393
timestamp 1688980957
transform 1 0 37260 0 -1 34816
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_3
timestamp 1688980957
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_15
timestamp 1688980957
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_27
timestamp 1688980957
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_29
timestamp 1688980957
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_41
timestamp 1688980957
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_53
timestamp 1688980957
transform 1 0 5980 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_59
timestamp 1688980957
transform 1 0 6532 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_85
timestamp 1688980957
transform 1 0 8924 0 1 34816
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_100
timestamp 1688980957
transform 1 0 10304 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_112
timestamp 1688980957
transform 1 0 11408 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_124
timestamp 1688980957
transform 1 0 12512 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_136
timestamp 1688980957
transform 1 0 13616 0 1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_141
timestamp 1688980957
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_153
timestamp 1688980957
transform 1 0 15180 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_165
timestamp 1688980957
transform 1 0 16284 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_173
timestamp 1688980957
transform 1 0 17020 0 1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_179
timestamp 1688980957
transform 1 0 17572 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_191
timestamp 1688980957
transform 1 0 18676 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_195
timestamp 1688980957
transform 1 0 19044 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_197
timestamp 1688980957
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_209
timestamp 1688980957
transform 1 0 20332 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_221
timestamp 1688980957
transform 1 0 21436 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_233
timestamp 1688980957
transform 1 0 22540 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_249
timestamp 1688980957
transform 1 0 24012 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_253
timestamp 1688980957
transform 1 0 24380 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_261
timestamp 1688980957
transform 1 0 25116 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_279
timestamp 1688980957
transform 1 0 26772 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_297
timestamp 1688980957
transform 1 0 28428 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_303
timestamp 1688980957
transform 1 0 28980 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_307
timestamp 1688980957
transform 1 0 29348 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_309
timestamp 1688980957
transform 1 0 29532 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_317
timestamp 1688980957
transform 1 0 30268 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_342
timestamp 1688980957
transform 1 0 32568 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_365
timestamp 1688980957
transform 1 0 34684 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_377
timestamp 1688980957
transform 1 0 35788 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_389
timestamp 1688980957
transform 1 0 36892 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_3
timestamp 1688980957
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_15
timestamp 1688980957
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_27
timestamp 1688980957
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_39
timestamp 1688980957
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_51
timestamp 1688980957
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_55
timestamp 1688980957
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_57
timestamp 1688980957
transform 1 0 6348 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_62
timestamp 1688980957
transform 1 0 6808 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_66
timestamp 1688980957
transform 1 0 7176 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_109
timestamp 1688980957
transform 1 0 11132 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_113
timestamp 1688980957
transform 1 0 11500 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_125
timestamp 1688980957
transform 1 0 12604 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_151
timestamp 1688980957
transform 1 0 14996 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_163
timestamp 1688980957
transform 1 0 16100 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_167
timestamp 1688980957
transform 1 0 16468 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_169
timestamp 1688980957
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_181
timestamp 1688980957
transform 1 0 17756 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_189
timestamp 1688980957
transform 1 0 18492 0 -1 35904
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_199
timestamp 1688980957
transform 1 0 19412 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_211
timestamp 1688980957
transform 1 0 20516 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_221
timestamp 1688980957
transform 1 0 21436 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_225
timestamp 1688980957
transform 1 0 21804 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_234
timestamp 1688980957
transform 1 0 22632 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_251
timestamp 1688980957
transform 1 0 24196 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_257
timestamp 1688980957
transform 1 0 24748 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_279
timestamp 1688980957
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_281
timestamp 1688980957
transform 1 0 26956 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_285
timestamp 1688980957
transform 1 0 27324 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_307
timestamp 1688980957
transform 1 0 29348 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_324
timestamp 1688980957
transform 1 0 30912 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_330
timestamp 1688980957
transform 1 0 31464 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_337
timestamp 1688980957
transform 1 0 32108 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_343
timestamp 1688980957
transform 1 0 32660 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_347
timestamp 1688980957
transform 1 0 33028 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_353
timestamp 1688980957
transform 1 0 33580 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_365
timestamp 1688980957
transform 1 0 34684 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_377
timestamp 1688980957
transform 1 0 35788 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_389
timestamp 1688980957
transform 1 0 36892 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_393
timestamp 1688980957
transform 1 0 37260 0 -1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_3
timestamp 1688980957
transform 1 0 1380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_15
timestamp 1688980957
transform 1 0 2484 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_27
timestamp 1688980957
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_29
timestamp 1688980957
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_41
timestamp 1688980957
transform 1 0 4876 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_49
timestamp 1688980957
transform 1 0 5612 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_74
timestamp 1688980957
transform 1 0 7912 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_82
timestamp 1688980957
transform 1 0 8648 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_85
timestamp 1688980957
transform 1 0 8924 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_95
timestamp 1688980957
transform 1 0 9844 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_107
timestamp 1688980957
transform 1 0 10948 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_134
timestamp 1688980957
transform 1 0 13432 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_141
timestamp 1688980957
transform 1 0 14076 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_150
timestamp 1688980957
transform 1 0 14904 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_168
timestamp 1688980957
transform 1 0 16560 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_185
timestamp 1688980957
transform 1 0 18124 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_192
timestamp 1688980957
transform 1 0 18768 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_197
timestamp 1688980957
transform 1 0 19228 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_209
timestamp 1688980957
transform 1 0 20332 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_221
timestamp 1688980957
transform 1 0 21436 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_233
timestamp 1688980957
transform 1 0 22540 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_241
timestamp 1688980957
transform 1 0 23276 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_251
timestamp 1688980957
transform 1 0 24196 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_253
timestamp 1688980957
transform 1 0 24380 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_272
timestamp 1688980957
transform 1 0 26128 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_292
timestamp 1688980957
transform 1 0 27968 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_309
timestamp 1688980957
transform 1 0 29532 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_321
timestamp 1688980957
transform 1 0 30636 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_333
timestamp 1688980957
transform 1 0 31740 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_339
timestamp 1688980957
transform 1 0 32292 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_351
timestamp 1688980957
transform 1 0 33396 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_363
timestamp 1688980957
transform 1 0 34500 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_365
timestamp 1688980957
transform 1 0 34684 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_377
timestamp 1688980957
transform 1 0 35788 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_389
timestamp 1688980957
transform 1 0 36892 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_3
timestamp 1688980957
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_15
timestamp 1688980957
transform 1 0 2484 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_27
timestamp 1688980957
transform 1 0 3588 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_39
timestamp 1688980957
transform 1 0 4692 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_51
timestamp 1688980957
transform 1 0 5796 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_55
timestamp 1688980957
transform 1 0 6164 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_57
timestamp 1688980957
transform 1 0 6348 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_65
timestamp 1688980957
transform 1 0 7084 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_72
timestamp 1688980957
transform 1 0 7728 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_84
timestamp 1688980957
transform 1 0 8832 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_88
timestamp 1688980957
transform 1 0 9200 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_98
timestamp 1688980957
transform 1 0 10120 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_110
timestamp 1688980957
transform 1 0 11224 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_113
timestamp 1688980957
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_125
timestamp 1688980957
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_137
timestamp 1688980957
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_149
timestamp 1688980957
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_161
timestamp 1688980957
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_167
timestamp 1688980957
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_169
timestamp 1688980957
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_181
timestamp 1688980957
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_193
timestamp 1688980957
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_205
timestamp 1688980957
transform 1 0 19964 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_213
timestamp 1688980957
transform 1 0 20700 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_218
timestamp 1688980957
transform 1 0 21160 0 -1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_225
timestamp 1688980957
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_237
timestamp 1688980957
transform 1 0 22908 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_250
timestamp 1688980957
transform 1 0 24104 0 -1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_260
timestamp 1688980957
transform 1 0 25024 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_272
timestamp 1688980957
transform 1 0 26128 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_281
timestamp 1688980957
transform 1 0 26956 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_290
timestamp 1688980957
transform 1 0 27784 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_298
timestamp 1688980957
transform 1 0 28520 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_304
timestamp 1688980957
transform 1 0 29072 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_314
timestamp 1688980957
transform 1 0 29992 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63_329
timestamp 1688980957
transform 1 0 31372 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_335
timestamp 1688980957
transform 1 0 31924 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_337
timestamp 1688980957
transform 1 0 32108 0 -1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_360
timestamp 1688980957
transform 1 0 34224 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_372
timestamp 1688980957
transform 1 0 35328 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_384
timestamp 1688980957
transform 1 0 36432 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_393
timestamp 1688980957
transform 1 0 37260 0 -1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_7
timestamp 1688980957
transform 1 0 1748 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_19
timestamp 1688980957
transform 1 0 2852 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_27
timestamp 1688980957
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_29
timestamp 1688980957
transform 1 0 3772 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_41
timestamp 1688980957
transform 1 0 4876 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_53
timestamp 1688980957
transform 1 0 5980 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_65
timestamp 1688980957
transform 1 0 7084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_77
timestamp 1688980957
transform 1 0 8188 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_106
timestamp 1688980957
transform 1 0 10856 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_118
timestamp 1688980957
transform 1 0 11960 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_130
timestamp 1688980957
transform 1 0 13064 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_138
timestamp 1688980957
transform 1 0 13800 0 1 36992
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_141
timestamp 1688980957
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_153
timestamp 1688980957
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_165
timestamp 1688980957
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_177
timestamp 1688980957
transform 1 0 17388 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_192
timestamp 1688980957
transform 1 0 18768 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_197
timestamp 1688980957
transform 1 0 19228 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_205
timestamp 1688980957
transform 1 0 19964 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_240
timestamp 1688980957
transform 1 0 23184 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_248
timestamp 1688980957
transform 1 0 23920 0 1 36992
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_253
timestamp 1688980957
transform 1 0 24380 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_265
timestamp 1688980957
transform 1 0 25484 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_280
timestamp 1688980957
transform 1 0 26864 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_284
timestamp 1688980957
transform 1 0 27232 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_294
timestamp 1688980957
transform 1 0 28152 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_306
timestamp 1688980957
transform 1 0 29256 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_309
timestamp 1688980957
transform 1 0 29532 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_334
timestamp 1688980957
transform 1 0 31832 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_343
timestamp 1688980957
transform 1 0 32660 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_355
timestamp 1688980957
transform 1 0 33764 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_363
timestamp 1688980957
transform 1 0 34500 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_365
timestamp 1688980957
transform 1 0 34684 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_377
timestamp 1688980957
transform 1 0 35788 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_389
timestamp 1688980957
transform 1 0 36892 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_3
timestamp 1688980957
transform 1 0 1380 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_15
timestamp 1688980957
transform 1 0 2484 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_27
timestamp 1688980957
transform 1 0 3588 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_39
timestamp 1688980957
transform 1 0 4692 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_51
timestamp 1688980957
transform 1 0 5796 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_55
timestamp 1688980957
transform 1 0 6164 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_57
timestamp 1688980957
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_69
timestamp 1688980957
transform 1 0 7452 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_81
timestamp 1688980957
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_93
timestamp 1688980957
transform 1 0 9660 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_97
timestamp 1688980957
transform 1 0 10028 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_108
timestamp 1688980957
transform 1 0 11040 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_125
timestamp 1688980957
transform 1 0 12604 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_131
timestamp 1688980957
transform 1 0 13156 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_149
timestamp 1688980957
transform 1 0 14812 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_174
timestamp 1688980957
transform 1 0 17112 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_182
timestamp 1688980957
transform 1 0 17848 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_194
timestamp 1688980957
transform 1 0 18952 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_198
timestamp 1688980957
transform 1 0 19320 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_217
timestamp 1688980957
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_223
timestamp 1688980957
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_225
timestamp 1688980957
transform 1 0 21804 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_236
timestamp 1688980957
transform 1 0 22816 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_254
timestamp 1688980957
transform 1 0 24472 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_276
timestamp 1688980957
transform 1 0 26496 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_281
timestamp 1688980957
transform 1 0 26956 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_297
timestamp 1688980957
transform 1 0 28428 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_328
timestamp 1688980957
transform 1 0 31280 0 -1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_337
timestamp 1688980957
transform 1 0 32108 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_349
timestamp 1688980957
transform 1 0 33212 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_361
timestamp 1688980957
transform 1 0 34316 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_373
timestamp 1688980957
transform 1 0 35420 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_385
timestamp 1688980957
transform 1 0 36524 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_391
timestamp 1688980957
transform 1 0 37076 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_393
timestamp 1688980957
transform 1 0 37260 0 -1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_3
timestamp 1688980957
transform 1 0 1380 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_15
timestamp 1688980957
transform 1 0 2484 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_27
timestamp 1688980957
transform 1 0 3588 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_29
timestamp 1688980957
transform 1 0 3772 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_41
timestamp 1688980957
transform 1 0 4876 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_45
timestamp 1688980957
transform 1 0 5244 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_57
timestamp 1688980957
transform 1 0 6348 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_69
timestamp 1688980957
transform 1 0 7452 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_85
timestamp 1688980957
transform 1 0 8924 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_110
timestamp 1688980957
transform 1 0 11224 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_134
timestamp 1688980957
transform 1 0 13432 0 1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_141
timestamp 1688980957
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_153
timestamp 1688980957
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_165
timestamp 1688980957
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_177
timestamp 1688980957
transform 1 0 17388 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_185
timestamp 1688980957
transform 1 0 18124 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_190
timestamp 1688980957
transform 1 0 18584 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_217
timestamp 1688980957
transform 1 0 21068 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_245
timestamp 1688980957
transform 1 0 23644 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_251
timestamp 1688980957
transform 1 0 24196 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_253
timestamp 1688980957
transform 1 0 24380 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_259
timestamp 1688980957
transform 1 0 24932 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_307
timestamp 1688980957
transform 1 0 29348 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_312
timestamp 1688980957
transform 1 0 29808 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_324
timestamp 1688980957
transform 1 0 30912 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_339
timestamp 1688980957
transform 1 0 32292 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_351
timestamp 1688980957
transform 1 0 33396 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_363
timestamp 1688980957
transform 1 0 34500 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_368
timestamp 1688980957
transform 1 0 34960 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_380
timestamp 1688980957
transform 1 0 36064 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_392
timestamp 1688980957
transform 1 0 37168 0 1 38080
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_9
timestamp 1688980957
transform 1 0 1932 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_21
timestamp 1688980957
transform 1 0 3036 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_27
timestamp 1688980957
transform 1 0 3588 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_29
timestamp 1688980957
transform 1 0 3772 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_37
timestamp 1688980957
transform 1 0 4508 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_44
timestamp 1688980957
transform 1 0 5152 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_57
timestamp 1688980957
transform 1 0 6348 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_69
timestamp 1688980957
transform 1 0 7452 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_81
timestamp 1688980957
transform 1 0 8556 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_85
timestamp 1688980957
transform 1 0 8924 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_93
timestamp 1688980957
transform 1 0 9660 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_105
timestamp 1688980957
transform 1 0 10764 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_111
timestamp 1688980957
transform 1 0 11316 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_122
timestamp 1688980957
transform 1 0 12328 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_128
timestamp 1688980957
transform 1 0 12880 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_133
timestamp 1688980957
transform 1 0 13340 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_139
timestamp 1688980957
transform 1 0 13892 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_141
timestamp 1688980957
transform 1 0 14076 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_153
timestamp 1688980957
transform 1 0 15180 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_161
timestamp 1688980957
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_167
timestamp 1688980957
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_169
timestamp 1688980957
transform 1 0 16652 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_177
timestamp 1688980957
transform 1 0 17388 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_184
timestamp 1688980957
transform 1 0 18032 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_197
timestamp 1688980957
transform 1 0 19228 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_202
timestamp 1688980957
transform 1 0 19688 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_216
timestamp 1688980957
transform 1 0 20976 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_225
timestamp 1688980957
transform 1 0 21804 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_233
timestamp 1688980957
transform 1 0 22540 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_245
timestamp 1688980957
transform 1 0 23644 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_251
timestamp 1688980957
transform 1 0 24196 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_253
timestamp 1688980957
transform 1 0 24380 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_265
timestamp 1688980957
transform 1 0 25484 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_277
timestamp 1688980957
transform 1 0 26588 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_290
timestamp 1688980957
transform 1 0 27784 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_302
timestamp 1688980957
transform 1 0 28888 0 -1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_309
timestamp 1688980957
transform 1 0 29532 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_321
timestamp 1688980957
transform 1 0 30636 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_329
timestamp 1688980957
transform 1 0 31372 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_335
timestamp 1688980957
transform 1 0 31924 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_337
timestamp 1688980957
transform 1 0 32108 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_345
timestamp 1688980957
transform 1 0 32844 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_352
timestamp 1688980957
transform 1 0 33488 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_365
timestamp 1688980957
transform 1 0 34684 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_373
timestamp 1688980957
transform 1 0 35420 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_380
timestamp 1688980957
transform 1 0 36064 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_393
timestamp 1688980957
transform 1 0 37260 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_399
timestamp 1688980957
transform 1 0 37812 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8188 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1688980957
transform 1 0 10488 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1688980957
transform -1 0 10396 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1688980957
transform -1 0 9476 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold5
timestamp 1688980957
transform -1 0 13524 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold6
timestamp 1688980957
transform -1 0 15272 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold7
timestamp 1688980957
transform 1 0 15732 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold8
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold9
timestamp 1688980957
transform -1 0 9660 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold10
timestamp 1688980957
transform -1 0 8372 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold11
timestamp 1688980957
transform 1 0 6716 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold12
timestamp 1688980957
transform 1 0 6532 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold13
timestamp 1688980957
transform -1 0 11316 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold14
timestamp 1688980957
transform -1 0 12696 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__buf_4  input1
timestamp 1688980957
transform -1 0 37996 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input4
timestamp 1688980957
transform -1 0 31372 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input5
timestamp 1688980957
transform -1 0 11408 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1688980957
transform 1 0 8464 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1688980957
transform -1 0 15916 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input8
timestamp 1688980957
transform 1 0 37444 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input9
timestamp 1688980957
transform 1 0 37444 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input10 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20056 0 -1 39168
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1688980957
transform 1 0 1380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  max_cap47
timestamp 1688980957
transform -1 0 6256 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  max_cap48
timestamp 1688980957
transform -1 0 23460 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  max_cap49
timestamp 1688980957
transform 1 0 22816 0 -1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  max_cap52
timestamp 1688980957
transform 1 0 17112 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  max_cap53
timestamp 1688980957
transform 1 0 14536 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  max_cap54
timestamp 1688980957
transform -1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  max_cap55
timestamp 1688980957
transform 1 0 21804 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  max_cap56
timestamp 1688980957
transform 1 0 15916 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1688980957
transform -1 0 18032 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output13
timestamp 1688980957
transform -1 0 1932 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output14
timestamp 1688980957
transform 1 0 37444 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output15
timestamp 1688980957
transform -1 0 1932 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output16
timestamp 1688980957
transform 1 0 37628 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output17
timestamp 1688980957
transform -1 0 1932 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output18
timestamp 1688980957
transform 1 0 26956 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output19
timestamp 1688980957
transform 1 0 17480 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output20
timestamp 1688980957
transform -1 0 1932 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output21
timestamp 1688980957
transform -1 0 1932 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output22
timestamp 1688980957
transform -1 0 22540 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output23
timestamp 1688980957
transform -1 0 1932 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output24
timestamp 1688980957
transform 1 0 37444 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output25
timestamp 1688980957
transform 1 0 12972 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output26
timestamp 1688980957
transform -1 0 4508 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output27
timestamp 1688980957
transform -1 0 2576 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output28
timestamp 1688980957
transform 1 0 37628 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output29
timestamp 1688980957
transform -1 0 1932 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output30
timestamp 1688980957
transform 1 0 14904 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output31
timestamp 1688980957
transform 1 0 37444 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output32
timestamp 1688980957
transform 1 0 37444 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output33
timestamp 1688980957
transform 1 0 9108 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output34
timestamp 1688980957
transform 1 0 37444 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output35
timestamp 1688980957
transform -1 0 7084 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output36
timestamp 1688980957
transform 1 0 12972 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output37
timestamp 1688980957
transform -1 0 1932 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output38
timestamp 1688980957
transform 1 0 37628 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output39
timestamp 1688980957
transform -1 0 19964 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output40
timestamp 1688980957
transform 1 0 35512 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output41
timestamp 1688980957
transform 1 0 32936 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output42
timestamp 1688980957
transform -1 0 5152 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output43
timestamp 1688980957
transform -1 0 12052 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output44
timestamp 1688980957
transform 1 0 26956 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output45
timestamp 1688980957
transform -1 0 1932 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output46
timestamp 1688980957
transform 1 0 37444 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 38272 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 38272 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 38272 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 38272 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 38272 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 38272 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 38272 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 38272 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 38272 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 38272 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 38272 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 38272 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 38272 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 38272 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 38272 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 38272 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 38272 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 38272 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 38272 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 38272 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 38272 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 38272 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 38272 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 38272 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 38272 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 38272 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 38272 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 38272 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 38272 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 38272 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 38272 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 38272 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 38272 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 38272 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 38272 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 38272 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 38272 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 38272 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 38272 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 38272 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 38272 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 38272 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 38272 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 38272 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 38272 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 38272 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 38272 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1688980957
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1688980957
transform -1 0 38272 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1688980957
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1688980957
transform -1 0 38272 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1688980957
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1688980957
transform -1 0 38272 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1688980957
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1688980957
transform -1 0 38272 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1688980957
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1688980957
transform -1 0 38272 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1688980957
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1688980957
transform -1 0 38272 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1688980957
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1688980957
transform -1 0 38272 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1688980957
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1688980957
transform -1 0 38272 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1688980957
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1688980957
transform -1 0 38272 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1688980957
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1688980957
transform -1 0 38272 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1688980957
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1688980957
transform -1 0 38272 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1688980957
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1688980957
transform -1 0 38272 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1688980957
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1688980957
transform -1 0 38272 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1688980957
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1688980957
transform -1 0 38272 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1688980957
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1688980957
transform -1 0 38272 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1688980957
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1688980957
transform -1 0 38272 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1688980957
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1688980957
transform -1 0 38272 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1688980957
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1688980957
transform -1 0 38272 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1688980957
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1688980957
transform -1 0 38272 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1688980957
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1688980957
transform -1 0 38272 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1688980957
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1688980957
transform -1 0 38272 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1688980957
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1688980957
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1688980957
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1688980957
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1688980957
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1688980957
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1688980957
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1688980957
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1688980957
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1688980957
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1688980957
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1688980957
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1688980957
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1688980957
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1688980957
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1688980957
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1688980957
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1688980957
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1688980957
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1688980957
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1688980957
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1688980957
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1688980957
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1688980957
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1688980957
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1688980957
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1688980957
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1688980957
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1688980957
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1688980957
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1688980957
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1688980957
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1688980957
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1688980957
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1688980957
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1688980957
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1688980957
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1688980957
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1688980957
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1688980957
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1688980957
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1688980957
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1688980957
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1688980957
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1688980957
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1688980957
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1688980957
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1688980957
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1688980957
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1688980957
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1688980957
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1688980957
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1688980957
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1688980957
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1688980957
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1688980957
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1688980957
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1688980957
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1688980957
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1688980957
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1688980957
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1688980957
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1688980957
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1688980957
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1688980957
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1688980957
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1688980957
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1688980957
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1688980957
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1688980957
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1688980957
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1688980957
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1688980957
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1688980957
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1688980957
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1688980957
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1688980957
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1688980957
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1688980957
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1688980957
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1688980957
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1688980957
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1688980957
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1688980957
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1688980957
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1688980957
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1688980957
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1688980957
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1688980957
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1688980957
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1688980957
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1688980957
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1688980957
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1688980957
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1688980957
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1688980957
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1688980957
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1688980957
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1688980957
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1688980957
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1688980957
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1688980957
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1688980957
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1688980957
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1688980957
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1688980957
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1688980957
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1688980957
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1688980957
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1688980957
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1688980957
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1688980957
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1688980957
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1688980957
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1688980957
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1688980957
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1688980957
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1688980957
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1688980957
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1688980957
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1688980957
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1688980957
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1688980957
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1688980957
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1688980957
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1688980957
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1688980957
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1688980957
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1688980957
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1688980957
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1688980957
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1688980957
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1688980957
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1688980957
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1688980957
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1688980957
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1688980957
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1688980957
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1688980957
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1688980957
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1688980957
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1688980957
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1688980957
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1688980957
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1688980957
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1688980957
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1688980957
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1688980957
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1688980957
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1688980957
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1688980957
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1688980957
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1688980957
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1688980957
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1688980957
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1688980957
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1688980957
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1688980957
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1688980957
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1688980957
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1688980957
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1688980957
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1688980957
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1688980957
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1688980957
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1688980957
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1688980957
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1688980957
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1688980957
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1688980957
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1688980957
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1688980957
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1688980957
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1688980957
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1688980957
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1688980957
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1688980957
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1688980957
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1688980957
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1688980957
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1688980957
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1688980957
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1688980957
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1688980957
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1688980957
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1688980957
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1688980957
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1688980957
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1688980957
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1688980957
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1688980957
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1688980957
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1688980957
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1688980957
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1688980957
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1688980957
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1688980957
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1688980957
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1688980957
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1688980957
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1688980957
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1688980957
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1688980957
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1688980957
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1688980957
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1688980957
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1688980957
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1688980957
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1688980957
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1688980957
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1688980957
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1688980957
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1688980957
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1688980957
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1688980957
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1688980957
transform 1 0 26864 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1688980957
transform 1 0 32016 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1688980957
transform 1 0 37168 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1688980957
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1688980957
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1688980957
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1688980957
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1688980957
transform 1 0 24288 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1688980957
transform 1 0 29440 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1688980957
transform 1 0 34592 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1688980957
transform 1 0 3680 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1688980957
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1688980957
transform 1 0 8832 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1688980957
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1688980957
transform 1 0 13984 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1688980957
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1688980957
transform 1 0 19136 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1688980957
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1688980957
transform 1 0 24288 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1688980957
transform 1 0 26864 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1688980957
transform 1 0 29440 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1688980957
transform 1 0 32016 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1688980957
transform 1 0 34592 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1688980957
transform 1 0 37168 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  wire50
timestamp 1688980957
transform -1 0 17572 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  wire51
timestamp 1688980957
transform -1 0 15824 0 -1 27200
box -38 -48 406 592
<< labels >>
flabel metal4 s 4868 2128 5188 39216 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 35588 2128 35908 39216 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 6006 38320 6326 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal5 s 1056 36642 38320 36962 0 FreeSans 2560 0 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 4208 2128 4528 39216 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal4 s 34928 2128 35248 39216 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 5346 38320 5666 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal5 s 1056 35982 38320 36302 0 FreeSans 2560 0 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 27208 800 27328 0 FreeSans 480 0 0 0 clk
port 2 nsew signal input
flabel metal3 s 38618 8848 39418 8968 0 FreeSans 480 0 0 0 cs
port 3 nsew signal input
flabel metal3 s 0 11568 800 11688 0 FreeSans 480 0 0 0 gpi[0]
port 4 nsew signal input
flabel metal3 s 38618 29248 39418 29368 0 FreeSans 480 0 0 0 gpi[10]
port 5 nsew signal input
flabel metal3 s 0 31968 800 32088 0 FreeSans 480 0 0 0 gpi[11]
port 6 nsew signal input
flabel metal3 s 38618 13608 39418 13728 0 FreeSans 480 0 0 0 gpi[12]
port 7 nsew signal input
flabel metal2 s 1950 40762 2006 41562 0 FreeSans 224 90 0 0 gpi[13]
port 8 nsew signal input
flabel metal2 s 28354 0 28410 800 0 FreeSans 224 90 0 0 gpi[14]
port 9 nsew signal input
flabel metal3 s 38618 25168 39418 25288 0 FreeSans 480 0 0 0 gpi[15]
port 10 nsew signal input
flabel metal3 s 0 23128 800 23248 0 FreeSans 480 0 0 0 gpi[16]
port 11 nsew signal input
flabel metal3 s 38618 4088 39418 4208 0 FreeSans 480 0 0 0 gpi[17]
port 12 nsew signal input
flabel metal2 s 30286 0 30342 800 0 FreeSans 224 90 0 0 gpi[18]
port 13 nsew signal input
flabel metal2 s 23846 0 23902 800 0 FreeSans 224 90 0 0 gpi[19]
port 14 nsew signal input
flabel metal3 s 0 6808 800 6928 0 FreeSans 480 0 0 0 gpi[1]
port 15 nsew signal input
flabel metal2 s 39302 0 39358 800 0 FreeSans 224 90 0 0 gpi[20]
port 16 nsew signal input
flabel metal3 s 38618 6128 39418 6248 0 FreeSans 480 0 0 0 gpi[21]
port 17 nsew signal input
flabel metal2 s 34794 0 34850 800 0 FreeSans 224 90 0 0 gpi[22]
port 18 nsew signal input
flabel metal2 s 30930 40762 30986 41562 0 FreeSans 224 90 0 0 gpi[23]
port 19 nsew signal input
flabel metal2 s 28354 40762 28410 41562 0 FreeSans 224 90 0 0 gpi[24]
port 20 nsew signal input
flabel metal3 s 0 29928 800 30048 0 FreeSans 480 0 0 0 gpi[25]
port 21 nsew signal input
flabel metal3 s 38618 27208 39418 27328 0 FreeSans 480 0 0 0 gpi[26]
port 22 nsew signal input
flabel metal3 s 38618 31968 39418 32088 0 FreeSans 480 0 0 0 gpi[27]
port 23 nsew signal input
flabel metal3 s 0 34688 800 34808 0 FreeSans 480 0 0 0 gpi[28]
port 24 nsew signal input
flabel metal2 s 21914 0 21970 800 0 FreeSans 224 90 0 0 gpi[29]
port 25 nsew signal input
flabel metal2 s 10966 0 11022 800 0 FreeSans 224 90 0 0 gpi[2]
port 26 nsew signal input
flabel metal3 s 0 39448 800 39568 0 FreeSans 480 0 0 0 gpi[30]
port 27 nsew signal input
flabel metal3 s 0 2048 800 2168 0 FreeSans 480 0 0 0 gpi[31]
port 28 nsew signal input
flabel metal2 s 24490 40762 24546 41562 0 FreeSans 224 90 0 0 gpi[32]
port 29 nsew signal input
flabel metal2 s 6458 40762 6514 41562 0 FreeSans 224 90 0 0 gpi[33]
port 30 nsew signal input
flabel metal2 s 8390 0 8446 800 0 FreeSans 224 90 0 0 gpi[3]
port 31 nsew signal input
flabel metal2 s 15474 40762 15530 41562 0 FreeSans 224 90 0 0 gpi[4]
port 32 nsew signal input
flabel metal2 s 37370 40762 37426 41562 0 FreeSans 224 90 0 0 gpi[5]
port 33 nsew signal input
flabel metal2 s 37370 0 37426 800 0 FreeSans 224 90 0 0 gpi[6]
port 34 nsew signal input
flabel metal2 s 19982 40762 20038 41562 0 FreeSans 224 90 0 0 gpi[7]
port 35 nsew signal input
flabel metal2 s 39302 40762 39358 41562 0 FreeSans 224 90 0 0 gpi[8]
port 36 nsew signal input
flabel metal2 s 32862 0 32918 800 0 FreeSans 224 90 0 0 gpi[9]
port 37 nsew signal input
flabel metal2 s 17406 40762 17462 41562 0 FreeSans 224 90 0 0 gpo[0]
port 38 nsew signal tristate
flabel metal3 s 0 4088 800 4208 0 FreeSans 480 0 0 0 gpo[10]
port 39 nsew signal tristate
flabel metal3 s 38618 10888 39418 11008 0 FreeSans 480 0 0 0 gpo[11]
port 40 nsew signal tristate
flabel metal3 s 0 8848 800 8968 0 FreeSans 480 0 0 0 gpo[12]
port 41 nsew signal tristate
flabel metal3 s 38618 15648 39418 15768 0 FreeSans 480 0 0 0 gpo[13]
port 42 nsew signal tristate
flabel metal2 s 18 40762 74 41562 0 FreeSans 224 90 0 0 gpo[14]
port 43 nsew signal tristate
flabel metal2 s 26422 40762 26478 41562 0 FreeSans 224 90 0 0 gpo[15]
port 44 nsew signal tristate
flabel metal2 s 17406 0 17462 800 0 FreeSans 224 90 0 0 gpo[16]
port 45 nsew signal tristate
flabel metal2 s 18 0 74 800 0 FreeSans 224 90 0 0 gpo[17]
port 46 nsew signal tristate
flabel metal3 s 0 25168 800 25288 0 FreeSans 480 0 0 0 gpo[18]
port 47 nsew signal tristate
flabel metal2 s 21914 40762 21970 41562 0 FreeSans 224 90 0 0 gpo[19]
port 48 nsew signal tristate
flabel metal3 s 0 15648 800 15768 0 FreeSans 480 0 0 0 gpo[1]
port 49 nsew signal tristate
flabel metal3 s 38618 38768 39418 38888 0 FreeSans 480 0 0 0 gpo[20]
port 50 nsew signal tristate
flabel metal2 s 12898 40762 12954 41562 0 FreeSans 224 90 0 0 gpo[21]
port 51 nsew signal tristate
flabel metal2 s 3882 0 3938 800 0 FreeSans 224 90 0 0 gpo[22]
port 52 nsew signal tristate
flabel metal2 s 1950 0 2006 800 0 FreeSans 224 90 0 0 gpo[23]
port 53 nsew signal tristate
flabel metal3 s 38618 36728 39418 36848 0 FreeSans 480 0 0 0 gpo[24]
port 54 nsew signal tristate
flabel metal3 s 0 18368 800 18488 0 FreeSans 480 0 0 0 gpo[25]
port 55 nsew signal tristate
flabel metal2 s 14830 0 14886 800 0 FreeSans 224 90 0 0 gpo[26]
port 56 nsew signal tristate
flabel metal3 s 38618 34008 39418 34128 0 FreeSans 480 0 0 0 gpo[27]
port 57 nsew signal tristate
flabel metal3 s 38618 1368 39418 1488 0 FreeSans 480 0 0 0 gpo[28]
port 58 nsew signal tristate
flabel metal2 s 9034 40762 9090 41562 0 FreeSans 224 90 0 0 gpo[29]
port 59 nsew signal tristate
flabel metal3 s 38618 20408 39418 20528 0 FreeSans 480 0 0 0 gpo[2]
port 60 nsew signal tristate
flabel metal2 s 6458 0 6514 800 0 FreeSans 224 90 0 0 gpo[30]
port 61 nsew signal tristate
flabel metal2 s 12898 0 12954 800 0 FreeSans 224 90 0 0 gpo[31]
port 62 nsew signal tristate
flabel metal3 s 0 20408 800 20528 0 FreeSans 480 0 0 0 gpo[32]
port 63 nsew signal tristate
flabel metal3 s 38618 22448 39418 22568 0 FreeSans 480 0 0 0 gpo[33]
port 64 nsew signal tristate
flabel metal2 s 19338 0 19394 800 0 FreeSans 224 90 0 0 gpo[3]
port 65 nsew signal tristate
flabel metal2 s 35438 40762 35494 41562 0 FreeSans 224 90 0 0 gpo[4]
port 66 nsew signal tristate
flabel metal2 s 32862 40762 32918 41562 0 FreeSans 224 90 0 0 gpo[5]
port 67 nsew signal tristate
flabel metal2 s 4526 40762 4582 41562 0 FreeSans 224 90 0 0 gpo[6]
port 68 nsew signal tristate
flabel metal2 s 10966 40762 11022 41562 0 FreeSans 224 90 0 0 gpo[7]
port 69 nsew signal tristate
flabel metal2 s 26422 0 26478 800 0 FreeSans 224 90 0 0 gpo[8]
port 70 nsew signal tristate
flabel metal3 s 0 13608 800 13728 0 FreeSans 480 0 0 0 gpo[9]
port 71 nsew signal tristate
flabel metal3 s 0 36728 800 36848 0 FreeSans 480 0 0 0 nrst
port 72 nsew signal input
flabel metal3 s 38618 17688 39418 17808 0 FreeSans 480 0 0 0 store_en
port 73 nsew signal tristate
rlabel metal1 19688 39168 19688 39168 0 VGND
rlabel metal1 19688 38624 19688 38624 0 VPWR
rlabel viali 22310 25262 22310 25262 0 ALU.flags_to_alu\[0\]
rlabel metal2 18446 33150 18446 33150 0 ALU.flags_to_alu\[1\]
rlabel metal1 17434 27370 17434 27370 0 ALU.flags_to_alu\[2\]
rlabel metal1 6670 30158 6670 30158 0 ALU.flags_to_alu\[3\]
rlabel metal1 8740 28662 8740 28662 0 ALU.flags_to_alu\[4\]
rlabel metal1 11592 32402 11592 32402 0 ALU.flags_to_alu\[5\]
rlabel metal2 13018 35751 13018 35751 0 ALU.flags_to_alu\[6\]
rlabel metal1 17250 35020 17250 35020 0 ALU.flags_to_alu\[7\]
rlabel metal2 9614 12920 9614 12920 0 ALU.immediate\[0\]
rlabel metal1 6348 13362 6348 13362 0 ALU.immediate\[10\]
rlabel metal1 17894 21624 17894 21624 0 ALU.immediate\[11\]
rlabel metal2 19734 23358 19734 23358 0 ALU.immediate\[12\]
rlabel metal1 7774 17850 7774 17850 0 ALU.immediate\[13\]
rlabel metal1 8096 12954 8096 12954 0 ALU.immediate\[14\]
rlabel metal2 26082 19975 26082 19975 0 ALU.immediate\[15\]
rlabel metal1 17802 7888 17802 7888 0 ALU.immediate\[1\]
rlabel metal1 17894 9146 17894 9146 0 ALU.immediate\[2\]
rlabel metal1 16836 8602 16836 8602 0 ALU.immediate\[3\]
rlabel metal1 14030 11288 14030 11288 0 ALU.immediate\[4\]
rlabel metal2 17618 11458 17618 11458 0 ALU.immediate\[5\]
rlabel metal1 14122 15572 14122 15572 0 ALU.immediate\[6\]
rlabel metal2 12282 16031 12282 16031 0 ALU.immediate\[7\]
rlabel metal1 14122 17136 14122 17136 0 ALU.immediate\[8\]
rlabel metal1 4462 19958 4462 19958 0 ALU.immediate\[9\]
rlabel metal1 13110 7174 13110 7174 0 ByteBuffer.counter\[0\]
rlabel metal1 13202 6834 13202 6834 0 ByteBuffer.counter\[1\]
rlabel metal1 12926 12818 12926 12818 0 ByteBuffer.instr\[16\]
rlabel metal1 17388 17646 17388 17646 0 ByteBuffer.instr\[17\]
rlabel metal2 16882 12614 16882 12614 0 ByteBuffer.instr\[18\]
rlabel via1 19734 17170 19734 17170 0 ByteBuffer.instr\[19\]
rlabel metal1 20654 16524 20654 16524 0 ByteBuffer.instr\[20\]
rlabel metal2 19550 13600 19550 13600 0 ByteBuffer.instr\[21\]
rlabel metal1 16652 18258 16652 18258 0 ByteBuffer.instr\[22\]
rlabel metal2 15226 13090 15226 13090 0 ByteBuffer.instr\[23\]
rlabel metal1 11914 8466 11914 8466 0 ByteBuffer.next_counter\[0\]
rlabel metal1 9706 7480 9706 7480 0 ByteBuffer.next_counter\[1\]
rlabel metal2 8234 5372 8234 5372 0 ByteDecoder.num_bytes\[1\]
rlabel metal1 9982 5134 9982 5134 0 ByteDecoder.num_bytes\[2\]
rlabel metal1 9062 5780 9062 5780 0 ByteDecoder.num_bytes\[3\]
rlabel metal1 12742 5644 12742 5644 0 ByteDecoder.state\[0\]
rlabel metal1 12512 5746 12512 5746 0 ByteDecoder.state\[1\]
rlabel metal1 10304 5202 10304 5202 0 FSM.next_state\[0\]
rlabel metal1 11776 5270 11776 5270 0 FSM.next_state\[1\]
rlabel metal1 15364 6222 15364 6222 0 MemControl.state\[0\]
rlabel metal2 15870 4964 15870 4964 0 MemControl.state\[1\]
rlabel metal1 15042 6222 15042 6222 0 MemControl.state\[2\]
rlabel via1 8694 8262 8694 8262 0 PC.i_mem_addr\[0\]
rlabel metal2 3818 21454 3818 21454 0 PC.i_mem_addr\[10\]
rlabel metal1 3910 20876 3910 20876 0 PC.i_mem_addr\[11\]
rlabel metal1 8004 23018 8004 23018 0 PC.i_mem_addr\[12\]
rlabel metal2 4738 25296 4738 25296 0 PC.i_mem_addr\[13\]
rlabel metal2 5244 21556 5244 21556 0 PC.i_mem_addr\[14\]
rlabel metal1 5152 19822 5152 19822 0 PC.i_mem_addr\[15\]
rlabel metal1 5796 7378 5796 7378 0 PC.i_mem_addr\[1\]
rlabel metal1 4462 8466 4462 8466 0 PC.i_mem_addr\[2\]
rlabel metal1 6624 10778 6624 10778 0 PC.i_mem_addr\[3\]
rlabel metal1 4324 12138 4324 12138 0 PC.i_mem_addr\[4\]
rlabel metal1 3588 12954 3588 12954 0 PC.i_mem_addr\[5\]
rlabel metal1 3358 14994 3358 14994 0 PC.i_mem_addr\[6\]
rlabel metal1 5842 17238 5842 17238 0 PC.i_mem_addr\[7\]
rlabel metal1 17296 14042 17296 14042 0 PC.i_mem_addr\[8\]
rlabel metal1 3680 20366 3680 20366 0 PC.i_mem_addr\[9\]
rlabel metal1 18906 24140 18906 24140 0 RegFile.A\[0\]
rlabel metal1 22034 33456 22034 33456 0 RegFile.A\[1\]
rlabel metal1 19044 26894 19044 26894 0 RegFile.A\[2\]
rlabel metal1 34178 29648 34178 29648 0 RegFile.A\[3\]
rlabel metal2 13018 24463 13018 24463 0 RegFile.A\[4\]
rlabel metal1 32246 31246 32246 31246 0 RegFile.A\[5\]
rlabel metal1 13202 37774 13202 37774 0 RegFile.A\[6\]
rlabel metal1 25806 35054 25806 35054 0 RegFile.A\[7\]
rlabel metal2 28290 26367 28290 26367 0 RegFile.B\[0\]
rlabel metal1 20102 33898 20102 33898 0 RegFile.B\[1\]
rlabel metal1 15042 26418 15042 26418 0 RegFile.B\[2\]
rlabel metal2 29026 29478 29026 29478 0 RegFile.B\[3\]
rlabel metal2 30038 28832 30038 28832 0 RegFile.B\[4\]
rlabel metal2 29486 30872 29486 30872 0 RegFile.B\[5\]
rlabel metal1 17526 37876 17526 37876 0 RegFile.B\[6\]
rlabel metal2 29670 36074 29670 36074 0 RegFile.B\[7\]
rlabel metal1 12466 25262 12466 25262 0 RegFile.C\[0\]
rlabel metal2 18078 35054 18078 35054 0 RegFile.C\[1\]
rlabel metal1 16514 28458 16514 28458 0 RegFile.C\[2\]
rlabel metal1 13386 30838 13386 30838 0 RegFile.C\[3\]
rlabel metal1 20792 29138 20792 29138 0 RegFile.C\[4\]
rlabel metal2 20746 31025 20746 31025 0 RegFile.C\[5\]
rlabel metal2 16238 36992 16238 36992 0 RegFile.C\[6\]
rlabel metal2 21022 38080 21022 38080 0 RegFile.C\[7\]
rlabel metal1 22126 27030 22126 27030 0 RegFile.D\[0\]
rlabel metal1 15456 33898 15456 33898 0 RegFile.D\[1\]
rlabel metal1 33672 26350 33672 26350 0 RegFile.D\[2\]
rlabel metal2 30682 29954 30682 29954 0 RegFile.D\[3\]
rlabel metal2 22034 28900 22034 28900 0 RegFile.D\[4\]
rlabel metal1 29946 31858 29946 31858 0 RegFile.D\[5\]
rlabel metal1 15962 37910 15962 37910 0 RegFile.D\[6\]
rlabel metal2 30038 35904 30038 35904 0 RegFile.D\[7\]
rlabel metal1 13110 25296 13110 25296 0 RegFile.E\[0\]
rlabel metal1 16468 33966 16468 33966 0 RegFile.E\[1\]
rlabel metal1 14858 26350 14858 26350 0 RegFile.E\[2\]
rlabel metal1 14674 30668 14674 30668 0 RegFile.E\[3\]
rlabel metal1 7406 28186 7406 28186 0 RegFile.E\[4\]
rlabel via1 12098 32827 12098 32827 0 RegFile.E\[5\]
rlabel metal2 16882 36992 16882 36992 0 RegFile.E\[6\]
rlabel metal1 23323 33932 23323 33932 0 RegFile.E\[7\]
rlabel metal2 22586 24718 22586 24718 0 RegFile.H\[0\]
rlabel metal1 20516 33966 20516 33966 0 RegFile.H\[1\]
rlabel metal1 17158 26384 17158 26384 0 RegFile.H\[2\]
rlabel metal1 17710 31280 17710 31280 0 RegFile.H\[3\]
rlabel metal1 26082 28628 26082 28628 0 RegFile.H\[4\]
rlabel metal2 31878 32504 31878 32504 0 RegFile.H\[5\]
rlabel metal1 15410 36176 15410 36176 0 RegFile.H\[6\]
rlabel metal1 33580 36142 33580 36142 0 RegFile.H\[7\]
rlabel metal1 12466 24752 12466 24752 0 RegFile.L\[0\]
rlabel metal1 16882 34578 16882 34578 0 RegFile.L\[1\]
rlabel via1 16790 28050 16790 28050 0 RegFile.L\[2\]
rlabel metal2 9430 31008 9430 31008 0 RegFile.L\[3\]
rlabel metal1 7176 29478 7176 29478 0 RegFile.L\[4\]
rlabel metal1 6440 32946 6440 32946 0 RegFile.L\[5\]
rlabel metal2 10718 36992 10718 36992 0 RegFile.L\[6\]
rlabel metal1 22540 37298 22540 37298 0 RegFile.L\[7\]
rlabel metal1 16652 4794 16652 4794 0 _0000_
rlabel metal1 13708 5270 13708 5270 0 _0001_
rlabel metal1 14536 4250 14536 4250 0 _0066_
rlabel metal1 7728 5746 7728 5746 0 _0067_
rlabel metal1 8326 4216 8326 4216 0 _0068_
rlabel metal1 6072 5338 6072 5338 0 _0069_
rlabel metal1 6578 15130 6578 15130 0 _0070_
rlabel metal1 6164 14042 6164 14042 0 _0071_
rlabel metal1 4830 12954 4830 12954 0 _0072_
rlabel metal1 6900 21114 6900 21114 0 _0073_
rlabel metal1 8004 17850 8004 17850 0 _0074_
rlabel metal1 6486 17306 6486 17306 0 _0075_
rlabel metal1 6440 12750 6440 12750 0 _0076_
rlabel metal1 6992 19482 6992 19482 0 _0077_
rlabel metal1 11270 13192 11270 13192 0 _0078_
rlabel metal1 13202 15130 13202 15130 0 _0079_
rlabel metal1 15180 12138 15180 12138 0 _0080_
rlabel metal1 12489 11798 12489 11798 0 _0081_
rlabel metal1 10212 14450 10212 14450 0 _0082_
rlabel metal1 14168 10710 14168 10710 0 _0083_
rlabel metal1 11822 9962 11822 9962 0 _0084_
rlabel metal1 13478 12920 13478 12920 0 _0085_
rlabel metal2 8602 13022 8602 13022 0 _0086_
rlabel metal1 15676 6970 15676 6970 0 _0087_
rlabel metal2 16054 9282 16054 9282 0 _0088_
rlabel metal1 13570 8534 13570 8534 0 _0089_
rlabel metal1 10258 11186 10258 11186 0 _0090_
rlabel metal1 16054 11186 16054 11186 0 _0091_
rlabel metal2 10074 9180 10074 9180 0 _0092_
rlabel metal1 9476 16218 9476 16218 0 _0093_
rlabel metal2 11086 22882 11086 22882 0 _0094_
rlabel metal1 7498 33082 7498 33082 0 _0095_
rlabel metal1 7360 26554 7360 26554 0 _0096_
rlabel metal1 5290 30158 5290 30158 0 _0097_
rlabel metal1 6532 28594 6532 28594 0 _0098_
rlabel metal1 5934 31654 5934 31654 0 _0099_
rlabel metal2 9338 23460 9338 23460 0 _0100_
rlabel metal1 5428 26010 5428 26010 0 _0101_
rlabel metal2 7958 24548 7958 24548 0 _0102_
rlabel metal1 7452 34714 7452 34714 0 _0103_
rlabel metal2 8326 27812 8326 27812 0 _0104_
rlabel metal2 8326 31552 8326 31552 0 _0105_
rlabel metal1 4646 28730 4646 28730 0 _0106_
rlabel metal1 4876 32538 4876 32538 0 _0107_
rlabel metal1 9246 37128 9246 37128 0 _0108_
rlabel metal1 20838 36890 20838 36890 0 _0109_
rlabel metal1 25944 24242 25944 24242 0 _0110_
rlabel metal1 31004 35122 31004 35122 0 _0111_
rlabel metal1 31372 26418 31372 26418 0 _0112_
rlabel metal2 35282 31450 35282 31450 0 _0113_
rlabel metal2 34454 28322 34454 28322 0 _0114_
rlabel metal1 31510 32776 31510 32776 0 _0115_
rlabel metal2 28198 35394 28198 35394 0 _0116_
rlabel metal2 32246 36516 32246 36516 0 _0117_
rlabel metal1 9016 25466 9016 25466 0 _0118_
rlabel metal1 6440 35802 6440 35802 0 _0119_
rlabel metal1 10166 27098 10166 27098 0 _0120_
rlabel metal1 6348 30362 6348 30362 0 _0121_
rlabel metal1 4692 27642 4692 27642 0 _0122_
rlabel metal1 5336 34034 5336 34034 0 _0123_
rlabel metal2 12834 38488 12834 38488 0 _0124_
rlabel metal1 22126 38216 22126 38216 0 _0125_
rlabel metal1 26680 27098 26680 27098 0 _0126_
rlabel metal1 33166 35122 33166 35122 0 _0127_
rlabel metal1 33534 26894 33534 26894 0 _0128_
rlabel metal1 34132 30906 34132 30906 0 _0129_
rlabel metal1 32246 28594 32246 28594 0 _0130_
rlabel metal1 28566 32538 28566 32538 0 _0131_
rlabel metal1 25944 37978 25944 37978 0 _0132_
rlabel metal1 30590 37298 30590 37298 0 _0133_
rlabel metal1 10580 24922 10580 24922 0 _0134_
rlabel metal1 9568 35734 9568 35734 0 _0135_
rlabel metal1 10580 28186 10580 28186 0 _0136_
rlabel metal1 9844 31450 9844 31450 0 _0137_
rlabel metal1 8878 29682 8878 29682 0 _0138_
rlabel metal1 9246 33592 9246 33592 0 _0139_
rlabel metal1 9706 37978 9706 37978 0 _0140_
rlabel metal1 19596 38386 19596 38386 0 _0141_
rlabel metal1 27876 26894 27876 26894 0 _0142_
rlabel metal2 28106 34272 28106 34272 0 _0143_
rlabel metal1 29762 27064 29762 27064 0 _0144_
rlabel metal1 27738 29206 27738 29206 0 _0145_
rlabel metal2 29302 28798 29302 28798 0 _0146_
rlabel metal1 28060 31654 28060 31654 0 _0147_
rlabel metal1 27186 37978 27186 37978 0 _0148_
rlabel metal1 29210 37774 29210 37774 0 _0149_
rlabel metal1 29026 24718 29026 24718 0 _0150_
rlabel metal1 34914 32946 34914 32946 0 _0151_
rlabel metal1 35098 26418 35098 26418 0 _0152_
rlabel metal1 34914 29002 34914 29002 0 _0153_
rlabel metal1 34776 25194 34776 25194 0 _0154_
rlabel metal1 30038 31246 30038 31246 0 _0155_
rlabel metal1 27048 33422 27048 33422 0 _0156_
rlabel metal1 34546 34034 34546 34034 0 _0157_
rlabel metal1 7452 7514 7452 7514 0 _0158_
rlabel metal1 4646 6426 4646 6426 0 _0159_
rlabel metal1 2944 7446 2944 7446 0 _0160_
rlabel metal1 4692 10234 4692 10234 0 _0161_
rlabel metal1 1748 10778 1748 10778 0 _0162_
rlabel metal1 1840 12410 1840 12410 0 _0163_
rlabel metal1 1840 14042 1840 14042 0 _0164_
rlabel metal2 4278 17442 4278 17442 0 _0165_
rlabel metal1 2024 16422 2024 16422 0 _0166_
rlabel metal1 1748 19414 1748 19414 0 _0167_
rlabel metal1 1748 24378 1748 24378 0 _0168_
rlabel metal1 1702 21624 1702 21624 0 _0169_
rlabel metal1 5612 24242 5612 24242 0 _0170_
rlabel metal1 3772 25466 3772 25466 0 _0171_
rlabel metal2 2898 25500 2898 25500 0 _0172_
rlabel metal1 4784 18938 4784 18938 0 _0173_
rlabel metal1 27968 4250 27968 4250 0 _0174_
rlabel metal1 27968 6698 27968 6698 0 _0175_
rlabel metal1 26082 8976 26082 8976 0 _0176_
rlabel metal1 26772 8466 26772 8466 0 _0177_
rlabel metal1 27554 6834 27554 6834 0 _0178_
rlabel metal1 27554 6732 27554 6732 0 _0179_
rlabel metal1 28382 6732 28382 6732 0 _0180_
rlabel metal1 27922 7344 27922 7344 0 _0181_
rlabel metal1 28520 7378 28520 7378 0 _0182_
rlabel metal1 17664 10642 17664 10642 0 _0183_
rlabel metal1 36202 21658 36202 21658 0 _0184_
rlabel metal1 35696 20910 35696 20910 0 _0185_
rlabel metal1 35190 20876 35190 20876 0 _0186_
rlabel metal2 34454 20621 34454 20621 0 _0187_
rlabel metal2 33350 30022 33350 30022 0 _0188_
rlabel metal1 34592 29138 34592 29138 0 _0189_
rlabel metal2 23046 5644 23046 5644 0 _0190_
rlabel metal1 23368 5338 23368 5338 0 _0191_
rlabel metal1 23414 5100 23414 5100 0 _0192_
rlabel metal2 24426 4896 24426 4896 0 _0193_
rlabel metal1 20654 4794 20654 4794 0 _0194_
rlabel metal1 24886 5644 24886 5644 0 _0195_
rlabel metal1 25392 6426 25392 6426 0 _0196_
rlabel metal1 24702 7310 24702 7310 0 _0197_
rlabel metal1 25116 8806 25116 8806 0 _0198_
rlabel metal1 25392 7310 25392 7310 0 _0199_
rlabel metal1 25484 7446 25484 7446 0 _0200_
rlabel metal1 24702 5678 24702 5678 0 _0201_
rlabel metal1 24058 5134 24058 5134 0 _0202_
rlabel metal2 23690 5508 23690 5508 0 _0203_
rlabel metal1 21758 18768 21758 18768 0 _0204_
rlabel metal1 36064 19482 36064 19482 0 _0205_
rlabel metal1 35650 19686 35650 19686 0 _0206_
rlabel viali 35374 19817 35374 19817 0 _0207_
rlabel metal1 34822 19754 34822 19754 0 _0208_
rlabel via1 25346 21590 25346 21590 0 _0209_
rlabel metal1 32200 25874 32200 25874 0 _0210_
rlabel metal1 34776 26010 34776 26010 0 _0211_
rlabel metal2 22034 7854 22034 7854 0 _0212_
rlabel metal1 22356 8262 22356 8262 0 _0213_
rlabel metal1 19964 6426 19964 6426 0 _0214_
rlabel metal1 20884 6834 20884 6834 0 _0215_
rlabel metal2 22402 7650 22402 7650 0 _0216_
rlabel metal1 20102 7820 20102 7820 0 _0217_
rlabel metal1 23552 8466 23552 8466 0 _0218_
rlabel metal1 22908 8942 22908 8942 0 _0219_
rlabel metal1 23230 8500 23230 8500 0 _0220_
rlabel metal1 22402 7854 22402 7854 0 _0221_
rlabel metal1 22448 7378 22448 7378 0 _0222_
rlabel metal1 23184 7514 23184 7514 0 _0223_
rlabel via2 9062 19363 9062 19363 0 _0224_
rlabel metal1 34362 18190 34362 18190 0 _0225_
rlabel metal1 35190 18190 35190 18190 0 _0226_
rlabel metal1 34822 18326 34822 18326 0 _0227_
rlabel metal1 34040 17646 34040 17646 0 _0228_
rlabel metal2 17250 19074 17250 19074 0 _0229_
rlabel metal1 28290 19482 28290 19482 0 _0230_
rlabel metal1 34684 33490 34684 33490 0 _0231_
rlabel viali 22121 10642 22121 10642 0 _0232_
rlabel metal1 21022 10166 21022 10166 0 _0233_
rlabel metal1 21022 10098 21022 10098 0 _0234_
rlabel metal1 21528 10098 21528 10098 0 _0235_
rlabel metal1 21482 10234 21482 10234 0 _0236_
rlabel metal1 22586 10098 22586 10098 0 _0237_
rlabel metal1 22448 9690 22448 9690 0 _0238_
rlabel metal1 21896 11118 21896 11118 0 _0239_
rlabel metal1 21758 11016 21758 11016 0 _0240_
rlabel metal2 22310 10642 22310 10642 0 _0241_
rlabel metal2 22678 10438 22678 10438 0 _0242_
rlabel metal2 22034 19907 22034 19907 0 _0243_
rlabel metal1 32200 17238 32200 17238 0 _0244_
rlabel metal1 32292 17170 32292 17170 0 _0245_
rlabel metal1 32706 17102 32706 17102 0 _0246_
rlabel metal1 33074 17136 33074 17136 0 _0247_
rlabel metal2 17894 14552 17894 14552 0 _0248_
rlabel metal1 27370 24820 27370 24820 0 _0249_
rlabel metal1 28888 23834 28888 23834 0 _0250_
rlabel metal1 25530 21386 25530 21386 0 _0251_
rlabel metal1 28842 34034 28842 34034 0 _0252_
rlabel metal1 29118 36890 29118 36890 0 _0253_
rlabel metal1 27002 37434 27002 37434 0 _0254_
rlabel metal1 28198 30906 28198 30906 0 _0255_
rlabel metal1 29348 28526 29348 28526 0 _0256_
rlabel metal1 28428 29614 28428 29614 0 _0257_
rlabel metal1 30176 26554 30176 26554 0 _0258_
rlabel metal1 28198 33966 28198 33966 0 _0259_
rlabel metal1 28014 26554 28014 26554 0 _0260_
rlabel metal1 13708 17510 13708 17510 0 _0261_
rlabel metal1 13386 21454 13386 21454 0 _0262_
rlabel metal1 14490 20026 14490 20026 0 _0263_
rlabel metal1 15548 21046 15548 21046 0 _0264_
rlabel metal1 23736 23698 23736 23698 0 _0265_
rlabel metal1 22586 21658 22586 21658 0 _0266_
rlabel metal2 22954 22916 22954 22916 0 _0267_
rlabel metal1 22724 23562 22724 23562 0 _0268_
rlabel metal1 23276 23086 23276 23086 0 _0269_
rlabel metal3 19711 33116 19711 33116 0 _0270_
rlabel metal2 19458 38454 19458 38454 0 _0271_
rlabel metal1 10166 36754 10166 36754 0 _0272_
rlabel metal1 10120 37842 10120 37842 0 _0273_
rlabel metal1 9016 21658 9016 21658 0 _0274_
rlabel metal1 10028 33082 10028 33082 0 _0275_
rlabel metal1 9706 21658 9706 21658 0 _0276_
rlabel metal1 8556 29002 8556 29002 0 _0277_
rlabel metal1 10304 20026 10304 20026 0 _0278_
rlabel metal1 10120 31314 10120 31314 0 _0279_
rlabel metal1 9660 21114 9660 21114 0 _0280_
rlabel metal1 11178 28050 11178 28050 0 _0281_
rlabel metal1 8740 19482 8740 19482 0 _0282_
rlabel metal1 9660 35258 9660 35258 0 _0283_
rlabel metal1 11132 19958 11132 19958 0 _0284_
rlabel metal1 11408 24786 11408 24786 0 _0285_
rlabel metal1 24978 23290 24978 23290 0 _0286_
rlabel metal1 24702 23732 24702 23732 0 _0287_
rlabel metal2 23506 24004 23506 24004 0 _0288_
rlabel metal1 33166 34476 33166 34476 0 _0289_
rlabel metal1 31280 36890 31280 36890 0 _0290_
rlabel metal1 26266 37434 26266 37434 0 _0291_
rlabel metal1 29072 32402 29072 32402 0 _0292_
rlabel metal1 33028 28186 33028 28186 0 _0293_
rlabel metal1 33856 30702 33856 30702 0 _0294_
rlabel metal1 33212 26554 33212 26554 0 _0295_
rlabel metal1 33626 34714 33626 34714 0 _0296_
rlabel metal1 27002 26962 27002 26962 0 _0297_
rlabel metal1 13662 37944 13662 37944 0 _0298_
rlabel metal1 21666 37978 21666 37978 0 _0299_
rlabel metal1 12190 37978 12190 37978 0 _0300_
rlabel metal1 5566 33626 5566 33626 0 _0301_
rlabel metal1 5612 27438 5612 27438 0 _0302_
rlabel metal1 6946 30226 6946 30226 0 _0303_
rlabel metal1 11040 26962 11040 26962 0 _0304_
rlabel metal1 7038 35666 7038 35666 0 _0305_
rlabel metal1 9292 25262 9292 25262 0 _0306_
rlabel metal2 23966 23324 23966 23324 0 _0307_
rlabel metal2 32706 25194 32706 25194 0 _0308_
rlabel metal1 32338 36142 32338 36142 0 _0309_
rlabel metal1 28382 35020 28382 35020 0 _0310_
rlabel metal1 31096 32266 31096 32266 0 _0311_
rlabel metal1 34408 28050 34408 28050 0 _0312_
rlabel metal2 35466 31348 35466 31348 0 _0313_
rlabel metal2 32154 26486 32154 26486 0 _0314_
rlabel metal1 31326 34714 31326 34714 0 _0315_
rlabel metal1 26588 24786 26588 24786 0 _0316_
rlabel metal1 8602 34476 8602 34476 0 _0317_
rlabel metal1 21597 36754 21597 36754 0 _0318_
rlabel metal1 8832 36890 8832 36890 0 _0319_
rlabel metal1 5750 32402 5750 32402 0 _0320_
rlabel metal1 5106 28526 5106 28526 0 _0321_
rlabel metal1 8740 30906 8740 30906 0 _0322_
rlabel metal1 8510 27506 8510 27506 0 _0323_
rlabel metal1 7912 34578 7912 34578 0 _0324_
rlabel metal1 8142 24242 8142 24242 0 _0325_
rlabel metal2 6026 18785 6026 18785 0 _0326_
rlabel metal1 13018 20434 13018 20434 0 _0327_
rlabel metal1 11362 21658 11362 21658 0 _0328_
rlabel metal1 18124 18870 18124 18870 0 _0329_
rlabel metal2 18078 18122 18078 18122 0 _0330_
rlabel metal2 17710 18292 17710 18292 0 _0331_
rlabel metal1 15870 17714 15870 17714 0 _0332_
rlabel metal3 13892 20604 13892 20604 0 _0333_
rlabel metal2 13754 23545 13754 23545 0 _0334_
rlabel metal1 12190 22066 12190 22066 0 _0335_
rlabel metal1 6302 25874 6302 25874 0 _0336_
rlabel metal1 9476 23086 9476 23086 0 _0337_
rlabel metal1 24702 20366 24702 20366 0 _0338_
rlabel metal2 23966 20128 23966 20128 0 _0339_
rlabel metal2 23874 19584 23874 19584 0 _0340_
rlabel metal1 22770 19482 22770 19482 0 _0341_
rlabel metal1 23644 19754 23644 19754 0 _0342_
rlabel metal1 13294 19142 13294 19142 0 _0343_
rlabel metal1 10028 22202 10028 22202 0 _0344_
rlabel metal1 9706 22746 9706 22746 0 _0345_
rlabel metal1 35742 15436 35742 15436 0 _0346_
rlabel metal1 28566 15028 28566 15028 0 _0347_
rlabel metal1 30084 7514 30084 7514 0 _0348_
rlabel metal2 33074 7378 33074 7378 0 _0349_
rlabel metal1 23966 6358 23966 6358 0 _0350_
rlabel metal1 24613 6426 24613 6426 0 _0351_
rlabel metal1 24150 7412 24150 7412 0 _0352_
rlabel metal2 24886 7004 24886 7004 0 _0353_
rlabel metal2 32522 6664 32522 6664 0 _0354_
rlabel metal1 34040 6630 34040 6630 0 _0355_
rlabel metal2 33534 10438 33534 10438 0 _0356_
rlabel metal1 33810 10438 33810 10438 0 _0357_
rlabel metal1 33994 10540 33994 10540 0 _0358_
rlabel metal1 34546 10506 34546 10506 0 _0359_
rlabel metal1 35512 15538 35512 15538 0 _0360_
rlabel metal1 34914 16626 34914 16626 0 _0361_
rlabel metal2 34546 18700 34546 18700 0 _0362_
rlabel metal1 34270 16966 34270 16966 0 _0363_
rlabel metal1 34316 17170 34316 17170 0 _0364_
rlabel metal1 34914 16490 34914 16490 0 _0365_
rlabel metal1 35236 16762 35236 16762 0 _0366_
rlabel metal1 33994 15028 33994 15028 0 _0367_
rlabel metal2 31234 14586 31234 14586 0 _0368_
rlabel metal1 32476 14586 32476 14586 0 _0369_
rlabel metal1 33442 14892 33442 14892 0 _0370_
rlabel metal1 34592 15130 34592 15130 0 _0371_
rlabel metal1 35282 16082 35282 16082 0 _0372_
rlabel metal1 35144 15946 35144 15946 0 _0373_
rlabel metal1 34914 16694 34914 16694 0 _0374_
rlabel metal1 32430 16524 32430 16524 0 _0375_
rlabel metal1 33212 16694 33212 16694 0 _0376_
rlabel metal1 28704 17238 28704 17238 0 _0377_
rlabel metal1 28240 17306 28240 17306 0 _0378_
rlabel metal2 28382 17476 28382 17476 0 _0379_
rlabel metal1 23138 16966 23138 16966 0 _0380_
rlabel metal1 25254 17714 25254 17714 0 _0381_
rlabel metal1 25070 17714 25070 17714 0 _0382_
rlabel metal1 25944 17646 25944 17646 0 _0383_
rlabel metal1 26312 17714 26312 17714 0 _0384_
rlabel metal1 27002 17748 27002 17748 0 _0385_
rlabel metal1 27692 17850 27692 17850 0 _0386_
rlabel metal2 27922 17850 27922 17850 0 _0387_
rlabel metal3 17204 17884 17204 17884 0 _0388_
rlabel metal1 8970 21862 8970 21862 0 _0389_
rlabel metal1 8004 26350 8004 26350 0 _0390_
rlabel metal1 8280 32946 8280 32946 0 _0391_
rlabel metal1 30360 16218 30360 16218 0 _0392_
rlabel metal1 29670 16762 29670 16762 0 _0393_
rlabel metal1 29670 12614 29670 12614 0 _0394_
rlabel metal1 22954 12138 22954 12138 0 _0395_
rlabel metal1 23414 12206 23414 12206 0 _0396_
rlabel metal2 26818 12036 26818 12036 0 _0397_
rlabel metal1 29670 12410 29670 12410 0 _0398_
rlabel metal1 29026 17204 29026 17204 0 _0399_
rlabel metal1 28750 19822 28750 19822 0 _0400_
rlabel metal2 29302 19550 29302 19550 0 _0401_
rlabel metal1 29210 19380 29210 19380 0 _0402_
rlabel metal1 29624 17170 29624 17170 0 _0403_
rlabel metal1 16606 17000 16606 17000 0 _0404_
rlabel metal1 12098 22202 12098 22202 0 _0405_
rlabel metal1 11362 22610 11362 22610 0 _0406_
rlabel metal1 7222 13804 7222 13804 0 _0407_
rlabel metal2 12374 7378 12374 7378 0 _0408_
rlabel metal1 15318 9452 15318 9452 0 _0409_
rlabel metal1 14260 7378 14260 7378 0 _0410_
rlabel metal1 16008 13158 16008 13158 0 _0411_
rlabel metal1 14674 6426 14674 6426 0 _0412_
rlabel metal1 12972 21454 12972 21454 0 _0413_
rlabel metal1 9706 5576 9706 5576 0 _0414_
rlabel metal2 9430 6018 9430 6018 0 _0415_
rlabel metal1 9798 5202 9798 5202 0 _0416_
rlabel metal1 13064 19686 13064 19686 0 _0417_
rlabel metal2 13202 19992 13202 19992 0 _0418_
rlabel metal1 8280 9622 8280 9622 0 _0419_
rlabel metal1 8924 14790 8924 14790 0 _0420_
rlabel metal1 14674 11118 14674 11118 0 _0421_
rlabel metal1 11500 15062 11500 15062 0 _0422_
rlabel metal1 8602 10608 8602 10608 0 _0423_
rlabel metal1 9246 10778 9246 10778 0 _0424_
rlabel metal1 8096 9554 8096 9554 0 _0425_
rlabel metal1 7912 14790 7912 14790 0 _0426_
rlabel metal1 7682 11152 7682 11152 0 _0427_
rlabel metal1 7912 11118 7912 11118 0 _0428_
rlabel metal1 8464 13226 8464 13226 0 _0429_
rlabel metal1 7820 9554 7820 9554 0 _0430_
rlabel metal1 7728 6222 7728 6222 0 _0431_
rlabel metal1 8326 6290 8326 6290 0 _0432_
rlabel metal1 9568 10098 9568 10098 0 _0433_
rlabel metal1 7958 9894 7958 9894 0 _0434_
rlabel metal1 15686 12818 15686 12818 0 _0435_
rlabel metal1 13570 14246 13570 14246 0 _0436_
rlabel metal1 9062 10132 9062 10132 0 _0437_
rlabel metal1 9338 6766 9338 6766 0 _0438_
rlabel metal1 9200 5202 9200 5202 0 _0439_
rlabel metal1 14260 18666 14260 18666 0 _0440_
rlabel metal1 14490 18292 14490 18292 0 _0441_
rlabel via2 20194 18411 20194 18411 0 _0442_
rlabel metal1 16468 4590 16468 4590 0 _0443_
rlabel metal1 16100 4522 16100 4522 0 _0444_
rlabel metal1 2162 18156 2162 18156 0 _0445_
rlabel metal2 15180 12444 15180 12444 0 _0446_
rlabel metal1 36386 32538 36386 32538 0 _0447_
rlabel metal1 37030 18258 37030 18258 0 _0448_
rlabel metal2 8602 35564 8602 35564 0 _0449_
rlabel via3 12581 4012 12581 4012 0 _0450_
rlabel metal3 13271 4012 13271 4012 0 _0451_
rlabel metal1 1978 23800 1978 23800 0 _0452_
rlabel metal1 37352 28050 37352 28050 0 _0453_
rlabel metal1 2162 17646 2162 17646 0 _0454_
rlabel metal2 12742 8772 12742 8772 0 _0455_
rlabel metal1 14306 8908 14306 8908 0 _0456_
rlabel metal1 6532 8874 6532 8874 0 _0457_
rlabel metal1 4370 8976 4370 8976 0 _0458_
rlabel metal2 13846 10574 13846 10574 0 _0459_
rlabel metal1 3450 9588 3450 9588 0 _0460_
rlabel metal1 6670 13498 6670 13498 0 _0461_
rlabel metal2 3450 17476 3450 17476 0 _0462_
rlabel metal1 17250 16728 17250 16728 0 _0463_
rlabel metal2 17434 11084 17434 11084 0 _0464_
rlabel metal1 17250 3094 17250 3094 0 _0465_
rlabel metal1 1886 17646 1886 17646 0 _0466_
rlabel metal2 1978 4963 1978 4963 0 _0467_
rlabel metal2 2714 22916 2714 22916 0 _0468_
rlabel via2 5658 20859 5658 20859 0 _0469_
rlabel metal1 24840 21998 24840 21998 0 _0470_
rlabel metal1 7958 22644 7958 22644 0 _0471_
rlabel metal1 5934 21488 5934 21488 0 _0472_
rlabel metal1 2346 18326 2346 18326 0 _0473_
rlabel metal2 2530 17307 2530 17307 0 _0474_
rlabel metal1 27370 21318 27370 21318 0 _0475_
rlabel metal1 25760 22610 25760 22610 0 _0476_
rlabel metal1 20470 37876 20470 37876 0 _0477_
rlabel metal2 2162 16286 2162 16286 0 _0478_
rlabel metal1 34822 20910 34822 20910 0 _0479_
rlabel metal2 25622 7723 25622 7723 0 _0480_
rlabel metal1 34730 38284 34730 38284 0 _0481_
rlabel metal1 28934 37978 28934 37978 0 _0482_
rlabel metal2 5198 38369 5198 38369 0 _0483_
rlabel via2 13202 37859 13202 37859 0 _0484_
rlabel metal2 14398 4828 14398 4828 0 _0485_
rlabel metal1 7038 5202 7038 5202 0 _0486_
rlabel metal1 6992 14994 6992 14994 0 _0487_
rlabel metal1 6624 13906 6624 13906 0 _0488_
rlabel metal1 5520 12818 5520 12818 0 _0489_
rlabel metal1 13110 11118 13110 11118 0 _0490_
rlabel metal1 7176 20910 7176 20910 0 _0491_
rlabel metal1 8602 17646 8602 17646 0 _0492_
rlabel metal1 6854 17170 6854 17170 0 _0493_
rlabel metal1 6026 12852 6026 12852 0 _0494_
rlabel metal1 7222 19414 7222 19414 0 _0495_
rlabel metal1 13294 8058 13294 8058 0 _0496_
rlabel metal1 12512 9486 12512 9486 0 _0497_
rlabel metal1 10948 13226 10948 13226 0 _0498_
rlabel metal1 13800 14586 13800 14586 0 _0499_
rlabel metal2 15088 12580 15088 12580 0 _0500_
rlabel metal2 12006 11526 12006 11526 0 _0501_
rlabel metal1 11040 14994 11040 14994 0 _0502_
rlabel metal1 13938 11118 13938 11118 0 _0503_
rlabel metal1 11638 9690 11638 9690 0 _0504_
rlabel metal1 13708 13294 13708 13294 0 _0505_
rlabel metal1 8970 13294 8970 13294 0 _0506_
rlabel metal1 15456 7378 15456 7378 0 _0507_
rlabel metal2 15962 9486 15962 9486 0 _0508_
rlabel metal1 13202 8500 13202 8500 0 _0509_
rlabel metal1 9798 11220 9798 11220 0 _0510_
rlabel metal2 15594 11322 15594 11322 0 _0511_
rlabel metal1 10350 9486 10350 9486 0 _0512_
rlabel metal1 9752 16082 9752 16082 0 _0513_
rlabel metal2 30958 28747 30958 28747 0 _0514_
rlabel via2 19090 30651 19090 30651 0 _0515_
rlabel metal2 33810 30005 33810 30005 0 _0516_
rlabel metal1 21528 31790 21528 31790 0 _0517_
rlabel metal1 18354 16150 18354 16150 0 _0518_
rlabel metal1 17434 7854 17434 7854 0 _0519_
rlabel metal1 10488 13498 10488 13498 0 _0520_
rlabel metal1 10304 12818 10304 12818 0 _0521_
rlabel metal1 10120 8602 10120 8602 0 _0522_
rlabel metal1 11454 18258 11454 18258 0 _0523_
rlabel metal1 12696 17850 12696 17850 0 _0524_
rlabel metal2 11638 20196 11638 20196 0 _0525_
rlabel metal1 11270 17680 11270 17680 0 _0526_
rlabel metal1 12466 17272 12466 17272 0 _0527_
rlabel metal2 12006 17442 12006 17442 0 _0528_
rlabel metal1 11408 17850 11408 17850 0 _0529_
rlabel metal2 11914 19754 11914 19754 0 _0530_
rlabel metal1 12052 18734 12052 18734 0 _0531_
rlabel metal1 12190 19346 12190 19346 0 _0532_
rlabel metal1 12190 18326 12190 18326 0 _0533_
rlabel metal1 11040 17714 11040 17714 0 _0534_
rlabel metal1 11132 18666 11132 18666 0 _0535_
rlabel metal1 11132 18734 11132 18734 0 _0536_
rlabel metal1 10396 17646 10396 17646 0 _0537_
rlabel metal1 12650 17680 12650 17680 0 _0538_
rlabel metal1 10764 17170 10764 17170 0 _0539_
rlabel metal1 10304 17714 10304 17714 0 _0540_
rlabel metal1 9108 8330 9108 8330 0 _0541_
rlabel metal1 3036 16626 3036 16626 0 _0542_
rlabel metal1 7958 7378 7958 7378 0 _0543_
rlabel metal1 17618 7786 17618 7786 0 _0544_
rlabel metal1 6486 7956 6486 7956 0 _0545_
rlabel metal1 6486 7310 6486 7310 0 _0546_
rlabel metal1 5888 7514 5888 7514 0 _0547_
rlabel metal1 4876 6290 4876 6290 0 _0548_
rlabel metal1 13570 8364 13570 8364 0 _0549_
rlabel metal1 5888 7854 5888 7854 0 _0550_
rlabel metal1 6210 10064 6210 10064 0 _0551_
rlabel metal1 5612 8058 5612 8058 0 _0552_
rlabel metal1 4692 8602 4692 8602 0 _0553_
rlabel metal1 3634 8466 3634 8466 0 _0554_
rlabel metal2 13110 9248 13110 9248 0 _0555_
rlabel metal1 3713 12070 3713 12070 0 _0556_
rlabel metal2 6210 10438 6210 10438 0 _0557_
rlabel metal1 6486 10574 6486 10574 0 _0558_
rlabel metal1 5658 10132 5658 10132 0 _0559_
rlabel metal1 5014 10030 5014 10030 0 _0560_
rlabel metal1 8234 10506 8234 10506 0 _0561_
rlabel metal1 3726 10642 3726 10642 0 _0562_
rlabel metal1 3312 10778 3312 10778 0 _0563_
rlabel metal1 2162 10642 2162 10642 0 _0564_
rlabel metal1 18078 12308 18078 12308 0 _0565_
rlabel metal1 17020 12342 17020 12342 0 _0566_
rlabel metal1 4646 12750 4646 12750 0 _0567_
rlabel metal2 4554 12818 4554 12818 0 _0568_
rlabel metal1 4324 12886 4324 12886 0 _0569_
rlabel metal1 3358 12614 3358 12614 0 _0570_
rlabel metal1 2392 12206 2392 12206 0 _0571_
rlabel metal1 4738 15130 4738 15130 0 _0572_
rlabel metal1 4554 15572 4554 15572 0 _0573_
rlabel metal1 3864 14382 3864 14382 0 _0574_
rlabel metal2 4094 14722 4094 14722 0 _0575_
rlabel metal1 3358 15130 3358 15130 0 _0576_
rlabel metal1 2346 13906 2346 13906 0 _0577_
rlabel metal1 8740 15946 8740 15946 0 _0578_
rlabel metal1 5336 15674 5336 15674 0 _0579_
rlabel metal1 5244 16218 5244 16218 0 _0580_
rlabel metal1 4508 17170 4508 17170 0 _0581_
rlabel metal1 3588 19346 3588 19346 0 _0582_
rlabel metal1 4094 16456 4094 16456 0 _0583_
rlabel metal1 3910 15674 3910 15674 0 _0584_
rlabel metal2 9706 18598 9706 18598 0 _0585_
rlabel metal1 2806 16660 2806 16660 0 _0586_
rlabel metal1 2346 16490 2346 16490 0 _0587_
rlabel metal1 3964 21862 3964 21862 0 _0588_
rlabel metal1 4094 19788 4094 19788 0 _0589_
rlabel metal2 3910 19550 3910 19550 0 _0590_
rlabel metal1 3358 20026 3358 20026 0 _0591_
rlabel metal1 2208 19822 2208 19822 0 _0592_
rlabel metal2 4002 22848 4002 22848 0 _0593_
rlabel metal1 3312 22746 3312 22746 0 _0594_
rlabel metal1 2898 23290 2898 23290 0 _0595_
rlabel metal1 2162 24174 2162 24174 0 _0596_
rlabel metal1 4232 21998 4232 21998 0 _0597_
rlabel metal1 4370 21590 4370 21590 0 _0598_
rlabel metal1 4508 21114 4508 21114 0 _0599_
rlabel metal1 3910 21522 3910 21522 0 _0600_
rlabel metal2 1978 21828 1978 21828 0 _0601_
rlabel metal1 7084 23018 7084 23018 0 _0602_
rlabel metal1 7222 23120 7222 23120 0 _0603_
rlabel metal2 7038 23494 7038 23494 0 _0604_
rlabel metal1 6164 23834 6164 23834 0 _0605_
rlabel metal1 5980 23290 5980 23290 0 _0606_
rlabel metal2 5290 23256 5290 23256 0 _0607_
rlabel metal1 5252 23096 5252 23096 0 _0608_
rlabel metal1 4922 23290 4922 23290 0 _0609_
rlabel metal2 4370 25092 4370 25092 0 _0610_
rlabel metal1 5382 22746 5382 22746 0 _0611_
rlabel metal1 4784 22746 4784 22746 0 _0612_
rlabel metal1 4462 23290 4462 23290 0 _0613_
rlabel metal1 3450 24378 3450 24378 0 _0614_
rlabel metal2 6394 19992 6394 19992 0 _0615_
rlabel metal1 5842 19686 5842 19686 0 _0616_
rlabel metal1 5106 18734 5106 18734 0 _0617_
rlabel metal1 21114 18734 21114 18734 0 _0618_
rlabel metal1 20332 17578 20332 17578 0 _0619_
rlabel metal1 20792 17646 20792 17646 0 _0620_
rlabel metal1 21160 17850 21160 17850 0 _0621_
rlabel metal1 20378 15878 20378 15878 0 _0622_
rlabel metal1 14214 22644 14214 22644 0 _0623_
rlabel metal1 17618 12920 17618 12920 0 _0624_
rlabel metal1 15364 13498 15364 13498 0 _0625_
rlabel metal1 19412 21522 19412 21522 0 _0626_
rlabel metal1 14260 15674 14260 15674 0 _0627_
rlabel metal1 13754 17680 13754 17680 0 _0628_
rlabel metal1 18538 31246 18538 31246 0 _0629_
rlabel metal1 29026 19380 29026 19380 0 _0630_
rlabel metal1 24012 18870 24012 18870 0 _0631_
rlabel metal1 15870 15436 15870 15436 0 _0632_
rlabel metal1 16422 20842 16422 20842 0 _0633_
rlabel metal1 16054 21046 16054 21046 0 _0634_
rlabel metal1 15739 16490 15739 16490 0 _0635_
rlabel metal1 12052 19210 12052 19210 0 _0636_
rlabel metal1 15042 20570 15042 20570 0 _0637_
rlabel metal1 13800 33558 13800 33558 0 _0638_
rlabel metal1 15686 18190 15686 18190 0 _0639_
rlabel viali 15131 21522 15131 21522 0 _0640_
rlabel metal2 19458 19788 19458 19788 0 _0641_
rlabel metal1 18998 20774 18998 20774 0 _0642_
rlabel metal1 16054 19278 16054 19278 0 _0643_
rlabel metal2 16422 20638 16422 20638 0 _0644_
rlabel metal1 20102 21522 20102 21522 0 _0645_
rlabel metal1 16100 23494 16100 23494 0 _0646_
rlabel metal1 19918 17272 19918 17272 0 _0647_
rlabel metal2 17572 21658 17572 21658 0 _0648_
rlabel metal1 20792 18938 20792 18938 0 _0649_
rlabel metal1 20424 23086 20424 23086 0 _0650_
rlabel metal2 20838 23494 20838 23494 0 _0651_
rlabel metal1 20194 33014 20194 33014 0 _0652_
rlabel metal1 14168 23290 14168 23290 0 _0653_
rlabel metal1 21804 25262 21804 25262 0 _0654_
rlabel metal1 29302 17646 29302 17646 0 _0655_
rlabel metal1 17066 14416 17066 14416 0 _0656_
rlabel metal2 17066 14790 17066 14790 0 _0657_
rlabel metal1 12512 6290 12512 6290 0 _0658_
rlabel metal1 13938 7820 13938 7820 0 _0659_
rlabel metal1 16330 15504 16330 15504 0 _0660_
rlabel metal2 16698 16864 16698 16864 0 _0661_
rlabel metal1 16652 14382 16652 14382 0 _0662_
rlabel metal1 16284 14586 16284 14586 0 _0663_
rlabel metal1 19366 15504 19366 15504 0 _0664_
rlabel metal1 19918 19890 19918 19890 0 _0665_
rlabel metal1 19826 19822 19826 19822 0 _0666_
rlabel metal2 19550 17884 19550 17884 0 _0667_
rlabel metal1 18722 18734 18722 18734 0 _0668_
rlabel metal1 18630 16082 18630 16082 0 _0669_
rlabel metal1 18860 20978 18860 20978 0 _0670_
rlabel metal1 18262 16048 18262 16048 0 _0671_
rlabel metal2 18170 16252 18170 16252 0 _0672_
rlabel metal1 18722 15538 18722 15538 0 _0673_
rlabel metal2 18630 13668 18630 13668 0 _0674_
rlabel metal1 18998 15368 18998 15368 0 _0675_
rlabel metal1 30222 25228 30222 25228 0 _0676_
rlabel metal1 14904 23698 14904 23698 0 _0677_
rlabel metal1 17020 22066 17020 22066 0 _0678_
rlabel metal1 14582 23698 14582 23698 0 _0679_
rlabel viali 27648 25262 27648 25262 0 _0680_
rlabel metal1 13386 33898 13386 33898 0 _0681_
rlabel metal1 13662 35734 13662 35734 0 _0682_
rlabel metal1 12558 26894 12558 26894 0 _0683_
rlabel metal1 19780 24038 19780 24038 0 _0684_
rlabel metal2 12650 28492 12650 28492 0 _0685_
rlabel metal1 14674 24378 14674 24378 0 _0686_
rlabel via1 23692 33966 23692 33966 0 _0687_
rlabel metal1 28106 36346 28106 36346 0 _0688_
rlabel metal3 29279 33116 29279 33116 0 _0689_
rlabel metal2 30222 23324 30222 23324 0 _0690_
rlabel metal1 30498 22576 30498 22576 0 _0691_
rlabel metal1 19826 15470 19826 15470 0 _0692_
rlabel metal1 18170 16626 18170 16626 0 _0693_
rlabel metal1 17342 22576 17342 22576 0 _0694_
rlabel metal1 18814 19822 18814 19822 0 _0695_
rlabel metal1 18170 19754 18170 19754 0 _0696_
rlabel metal2 12190 20128 12190 20128 0 _0697_
rlabel metal2 17158 22848 17158 22848 0 _0698_
rlabel metal1 16054 32878 16054 32878 0 _0699_
rlabel metal1 17342 16558 17342 16558 0 _0700_
rlabel metal1 19918 21556 19918 21556 0 _0701_
rlabel metal1 19688 21454 19688 21454 0 _0702_
rlabel metal2 18906 21835 18906 21835 0 _0703_
rlabel metal2 24334 27183 24334 27183 0 _0704_
rlabel metal1 20930 25874 20930 25874 0 _0705_
rlabel metal1 16882 26894 16882 26894 0 _0706_
rlabel metal1 16974 28016 16974 28016 0 _0707_
rlabel metal1 20746 33966 20746 33966 0 _0708_
rlabel metal2 17066 36346 17066 36346 0 _0709_
rlabel metal2 26220 35666 26220 35666 0 _0710_
rlabel via1 17319 36142 17319 36142 0 _0711_
rlabel metal1 26588 35054 26588 35054 0 _0712_
rlabel metal1 26082 37808 26082 37808 0 _0713_
rlabel metal1 29670 22644 29670 22644 0 _0714_
rlabel metal1 30636 20434 30636 20434 0 _0715_
rlabel metal1 29624 22406 29624 22406 0 _0716_
rlabel metal1 30130 22746 30130 22746 0 _0717_
rlabel metal1 30222 22066 30222 22066 0 _0718_
rlabel metal1 31786 29172 31786 29172 0 _0719_
rlabel metal1 32062 29138 32062 29138 0 _0720_
rlabel metal1 33764 29002 33764 29002 0 _0721_
rlabel metal1 26726 29648 26726 29648 0 _0722_
rlabel metal1 25990 29580 25990 29580 0 _0723_
rlabel via1 25806 21999 25806 21999 0 _0724_
rlabel metal1 27554 21046 27554 21046 0 _0725_
rlabel metal1 35052 22746 35052 22746 0 _0726_
rlabel metal2 31786 26588 31786 26588 0 _0727_
rlabel metal1 32982 25908 32982 25908 0 _0728_
rlabel metal1 35190 22984 35190 22984 0 _0729_
rlabel metal1 26542 26384 26542 26384 0 _0730_
rlabel metal1 26128 25874 26128 25874 0 _0731_
rlabel metal1 26956 22066 26956 22066 0 _0732_
rlabel metal2 27554 22984 27554 22984 0 _0733_
rlabel metal1 36754 22066 36754 22066 0 _0734_
rlabel metal1 36892 21998 36892 21998 0 _0735_
rlabel metal1 36570 19890 36570 19890 0 _0736_
rlabel metal1 36294 20026 36294 20026 0 _0737_
rlabel metal1 31786 34000 31786 34000 0 _0738_
rlabel metal1 32338 32402 32338 32402 0 _0739_
rlabel metal1 33258 19822 33258 19822 0 _0740_
rlabel metal1 21528 33354 21528 33354 0 _0741_
rlabel metal1 25898 34000 25898 34000 0 _0742_
rlabel metal1 25254 33320 25254 33320 0 _0743_
rlabel metal3 25277 33252 25277 33252 0 _0744_
rlabel metal1 33626 19856 33626 19856 0 _0745_
rlabel metal1 34868 19346 34868 19346 0 _0746_
rlabel metal2 28750 25466 28750 25466 0 _0747_
rlabel metal1 30038 25296 30038 25296 0 _0748_
rlabel metal1 31050 18258 31050 18258 0 _0749_
rlabel metal1 25254 25228 25254 25228 0 _0750_
rlabel metal2 24794 25568 24794 25568 0 _0751_
rlabel metal2 25116 21284 25116 21284 0 _0752_
rlabel metal1 31004 18326 31004 18326 0 _0753_
rlabel metal1 31947 18326 31947 18326 0 _0754_
rlabel metal1 31464 18258 31464 18258 0 _0755_
rlabel metal1 32016 17646 32016 17646 0 _0756_
rlabel metal1 17204 19958 17204 19958 0 _0757_
rlabel metal1 17848 21522 17848 21522 0 _0758_
rlabel metal1 17434 23630 17434 23630 0 _0759_
rlabel metal1 13662 33830 13662 33830 0 _0760_
rlabel via2 14306 23749 14306 23749 0 _0761_
rlabel via1 13938 31654 13938 31654 0 _0762_
rlabel metal1 15640 36074 15640 36074 0 _0763_
rlabel metal2 22862 31756 22862 31756 0 _0764_
rlabel metal1 14996 36142 14996 36142 0 _0765_
rlabel metal1 17618 23494 17618 23494 0 _0766_
rlabel metal1 14996 28050 14996 28050 0 _0767_
rlabel metal1 21620 30906 21620 30906 0 _0768_
rlabel metal2 22586 31450 22586 31450 0 _0769_
rlabel metal2 15778 36346 15778 36346 0 _0770_
rlabel metal1 14996 37706 14996 37706 0 _0771_
rlabel metal1 15732 23834 15732 23834 0 _0772_
rlabel metal1 23276 31654 23276 31654 0 _0773_
rlabel metal1 14858 29614 14858 29614 0 _0774_
rlabel metal1 22356 18938 22356 18938 0 _0775_
rlabel metal1 12466 32504 12466 32504 0 _0776_
rlabel metal1 12282 32504 12282 32504 0 _0777_
rlabel metal3 16399 32164 16399 32164 0 _0778_
rlabel metal1 19044 11118 19044 11118 0 _0779_
rlabel metal2 18216 12852 18216 12852 0 _0780_
rlabel metal2 32706 12036 32706 12036 0 _0781_
rlabel via2 18722 11611 18722 11611 0 _0782_
rlabel metal1 18308 24174 18308 24174 0 _0783_
rlabel metal1 17756 36142 17756 36142 0 _0784_
rlabel metal1 17020 21114 17020 21114 0 _0785_
rlabel metal1 16284 28526 16284 28526 0 _0786_
rlabel metal1 25438 31824 25438 31824 0 _0787_
rlabel metal1 18538 37196 18538 37196 0 _0788_
rlabel metal2 20194 26792 20194 26792 0 _0789_
rlabel metal1 23920 32436 23920 32436 0 _0790_
rlabel metal1 25346 31960 25346 31960 0 _0791_
rlabel metal1 18584 26758 18584 26758 0 _0792_
rlabel metal2 18722 36448 18722 36448 0 _0793_
rlabel metal1 17802 32538 17802 32538 0 _0794_
rlabel metal2 23368 31790 23368 31790 0 _0795_
rlabel metal1 25254 31722 25254 31722 0 _0796_
rlabel metal1 25024 30906 25024 30906 0 _0797_
rlabel metal2 25622 31484 25622 31484 0 _0798_
rlabel metal1 20792 31314 20792 31314 0 _0799_
rlabel metal1 21022 31314 21022 31314 0 _0800_
rlabel metal1 21229 31110 21229 31110 0 _0801_
rlabel via3 26749 30396 26749 30396 0 _0802_
rlabel metal1 32338 10676 32338 10676 0 _0803_
rlabel metal1 32338 11152 32338 11152 0 _0804_
rlabel metal1 33442 13260 33442 13260 0 _0805_
rlabel metal1 29716 9622 29716 9622 0 _0806_
rlabel metal2 14674 27846 14674 27846 0 _0807_
rlabel metal1 14352 27914 14352 27914 0 _0808_
rlabel metal1 14352 27642 14352 27642 0 _0809_
rlabel metal2 15134 26690 15134 26690 0 _0810_
rlabel metal1 14582 26554 14582 26554 0 _0811_
rlabel metal1 14076 26554 14076 26554 0 _0812_
rlabel metal1 13248 26350 13248 26350 0 _0813_
rlabel metal2 13662 27098 13662 27098 0 _0814_
rlabel metal2 15410 9231 15410 9231 0 _0815_
rlabel metal2 21850 8160 21850 8160 0 _0816_
rlabel metal1 16974 27472 16974 27472 0 _0817_
rlabel metal2 16698 27268 16698 27268 0 _0818_
rlabel metal1 17802 26996 17802 26996 0 _0819_
rlabel metal1 16744 26282 16744 26282 0 _0820_
rlabel metal1 17572 26554 17572 26554 0 _0821_
rlabel metal1 17480 26962 17480 26962 0 _0822_
rlabel metal1 18308 27098 18308 27098 0 _0823_
rlabel metal1 18906 27098 18906 27098 0 _0824_
rlabel metal1 16376 27574 16376 27574 0 _0825_
rlabel metal1 17572 27438 17572 27438 0 _0826_
rlabel metal1 18354 27404 18354 27404 0 _0827_
rlabel metal1 17986 15674 17986 15674 0 _0828_
rlabel via2 18906 9469 18906 9469 0 _0829_
rlabel metal2 18078 10234 18078 10234 0 _0830_
rlabel metal1 19504 4658 19504 4658 0 _0831_
rlabel metal1 30268 5202 30268 5202 0 _0832_
rlabel metal1 16652 29818 16652 29818 0 _0833_
rlabel metal1 17526 30158 17526 30158 0 _0834_
rlabel metal1 17066 30906 17066 30906 0 _0835_
rlabel metal1 17802 30056 17802 30056 0 _0836_
rlabel metal1 17112 30226 17112 30226 0 _0837_
rlabel metal1 18630 29682 18630 29682 0 _0838_
rlabel metal1 18814 29274 18814 29274 0 _0839_
rlabel metal1 16698 31280 16698 31280 0 _0840_
rlabel metal2 18630 30430 18630 30430 0 _0841_
rlabel metal2 18354 29818 18354 29818 0 _0842_
rlabel metal3 17365 10948 17365 10948 0 _0843_
rlabel metal2 18722 9792 18722 9792 0 _0844_
rlabel metal1 14260 30770 14260 30770 0 _0845_
rlabel metal1 14076 30906 14076 30906 0 _0846_
rlabel metal1 14214 29614 14214 29614 0 _0847_
rlabel metal1 14398 29784 14398 29784 0 _0848_
rlabel metal1 14490 29716 14490 29716 0 _0849_
rlabel metal1 13938 29750 13938 29750 0 _0850_
rlabel metal1 13478 29648 13478 29648 0 _0851_
rlabel metal2 13570 30362 13570 30362 0 _0852_
rlabel metal2 13248 17204 13248 17204 0 _0853_
rlabel metal1 18676 9962 18676 9962 0 _0854_
rlabel metal1 26634 7412 26634 7412 0 _0855_
rlabel metal1 28750 5270 28750 5270 0 _0856_
rlabel metal1 14628 33626 14628 33626 0 _0857_
rlabel metal1 14260 34034 14260 34034 0 _0858_
rlabel metal1 18285 34034 18285 34034 0 _0859_
rlabel metal1 19688 34102 19688 34102 0 _0860_
rlabel metal1 19274 33966 19274 33966 0 _0861_
rlabel metal2 20378 33660 20378 33660 0 _0862_
rlabel metal1 20286 33524 20286 33524 0 _0863_
rlabel metal1 11592 33966 11592 33966 0 _0864_
rlabel metal1 19918 33558 19918 33558 0 _0865_
rlabel metal2 19734 33252 19734 33252 0 _0866_
rlabel via3 19067 33252 19067 33252 0 _0867_
rlabel metal1 19642 5746 19642 5746 0 _0868_
rlabel metal2 17894 7004 17894 7004 0 _0869_
rlabel metal1 18860 35734 18860 35734 0 _0870_
rlabel metal1 18998 35598 18998 35598 0 _0871_
rlabel metal1 16974 34034 16974 34034 0 _0872_
rlabel metal1 16468 34102 16468 34102 0 _0873_
rlabel metal1 16790 34170 16790 34170 0 _0874_
rlabel metal1 17112 34714 17112 34714 0 _0875_
rlabel metal1 18630 32436 18630 32436 0 _0876_
rlabel metal1 17664 33626 17664 33626 0 _0877_
rlabel metal1 18492 33082 18492 33082 0 _0878_
rlabel metal2 18860 32402 18860 32402 0 _0879_
rlabel via3 18469 32028 18469 32028 0 _0880_
rlabel metal1 18906 5678 18906 5678 0 _0881_
rlabel metal1 20102 5338 20102 5338 0 _0882_
rlabel metal1 18860 7310 18860 7310 0 _0883_
rlabel metal1 18630 7378 18630 7378 0 _0884_
rlabel metal2 20102 11628 20102 11628 0 _0885_
rlabel metal1 22356 25874 22356 25874 0 _0886_
rlabel metal1 21942 24582 21942 24582 0 _0887_
rlabel metal1 22724 25466 22724 25466 0 _0888_
rlabel metal1 20838 26282 20838 26282 0 _0889_
rlabel metal2 22678 26180 22678 26180 0 _0890_
rlabel metal1 22770 25806 22770 25806 0 _0891_
rlabel metal2 22310 24378 22310 24378 0 _0892_
rlabel metal2 21022 25500 21022 25500 0 _0893_
rlabel metal1 21022 25398 21022 25398 0 _0894_
rlabel metal1 20930 23086 20930 23086 0 _0895_
rlabel metal1 20010 11152 20010 11152 0 _0896_
rlabel metal2 19826 25942 19826 25942 0 _0897_
rlabel metal1 18998 24378 18998 24378 0 _0898_
rlabel metal2 19182 23902 19182 23902 0 _0899_
rlabel metal1 19090 23732 19090 23732 0 _0900_
rlabel metal1 19274 23562 19274 23562 0 _0901_
rlabel metal2 18722 24004 18722 24004 0 _0902_
rlabel metal1 18722 24038 18722 24038 0 _0903_
rlabel metal1 13018 24888 13018 24888 0 _0904_
rlabel metal1 12788 24786 12788 24786 0 _0905_
rlabel metal2 13110 22080 13110 22080 0 _0906_
rlabel metal2 19366 12818 19366 12818 0 _0907_
rlabel metal1 20148 9486 20148 9486 0 _0908_
rlabel metal1 19642 7854 19642 7854 0 _0909_
rlabel metal1 20608 5678 20608 5678 0 _0910_
rlabel metal1 20056 4522 20056 4522 0 _0911_
rlabel metal2 29854 4624 29854 4624 0 _0912_
rlabel metal1 30912 5202 30912 5202 0 _0913_
rlabel metal1 23092 28186 23092 28186 0 _0914_
rlabel metal1 21528 29138 21528 29138 0 _0915_
rlabel metal1 22724 29002 22724 29002 0 _0916_
rlabel metal1 22816 29138 22816 29138 0 _0917_
rlabel metal1 23046 28050 23046 28050 0 _0918_
rlabel metal1 21781 27914 21781 27914 0 _0919_
rlabel metal2 22494 28662 22494 28662 0 _0920_
rlabel metal1 14030 10540 14030 10540 0 _0921_
rlabel metal2 26542 9146 26542 9146 0 _0922_
rlabel metal1 23874 26010 23874 26010 0 _0923_
rlabel metal1 24242 27914 24242 27914 0 _0924_
rlabel metal1 24196 28050 24196 28050 0 _0925_
rlabel metal1 23276 27370 23276 27370 0 _0926_
rlabel metal1 24012 27642 24012 27642 0 _0927_
rlabel metal1 24196 26350 24196 26350 0 _0928_
rlabel metal1 23092 15470 23092 15470 0 _0929_
rlabel metal1 19918 28084 19918 28084 0 _0930_
rlabel metal2 19826 28135 19826 28135 0 _0931_
rlabel metal1 19872 27914 19872 27914 0 _0932_
rlabel metal2 21574 17068 21574 17068 0 _0933_
rlabel metal1 23736 15878 23736 15878 0 _0934_
rlabel metal2 31878 9792 31878 9792 0 _0935_
rlabel metal1 33258 8874 33258 8874 0 _0936_
rlabel metal1 28566 8908 28566 8908 0 _0937_
rlabel metal2 30314 5474 30314 5474 0 _0938_
rlabel metal1 23966 35054 23966 35054 0 _0939_
rlabel metal1 21666 35666 21666 35666 0 _0940_
rlabel metal1 23690 35156 23690 35156 0 _0941_
rlabel via1 23598 35139 23598 35139 0 _0942_
rlabel metal2 23598 34170 23598 34170 0 _0943_
rlabel metal2 23874 33660 23874 33660 0 _0944_
rlabel metal2 23782 33932 23782 33932 0 _0945_
rlabel via2 12374 16099 12374 16099 0 _0946_
rlabel metal1 25300 12274 25300 12274 0 _0947_
rlabel metal1 24196 29478 24196 29478 0 _0948_
rlabel metal1 24794 36788 24794 36788 0 _0949_
rlabel metal2 24702 36992 24702 36992 0 _0950_
rlabel metal1 24012 37910 24012 37910 0 _0951_
rlabel metal1 24656 36754 24656 36754 0 _0952_
rlabel metal1 24334 36346 24334 36346 0 _0953_
rlabel via3 24955 35972 24955 35972 0 _0954_
rlabel via1 23426 16558 23426 16558 0 _0955_
rlabel metal1 21666 34578 21666 34578 0 _0956_
rlabel metal2 22678 34170 22678 34170 0 _0957_
rlabel metal3 24725 17612 24725 17612 0 _0958_
rlabel metal1 25070 16082 25070 16082 0 _0959_
rlabel metal1 27416 15470 27416 15470 0 _0960_
rlabel metal1 14674 37842 14674 37842 0 _0961_
rlabel metal1 14122 35802 14122 35802 0 _0962_
rlabel metal2 13846 37094 13846 37094 0 _0963_
rlabel metal1 13754 37910 13754 37910 0 _0964_
rlabel metal1 13800 37774 13800 37774 0 _0965_
rlabel metal2 12466 36856 12466 36856 0 _0966_
rlabel metal1 12696 36210 12696 36210 0 _0967_
rlabel metal1 11822 36244 11822 36244 0 _0968_
rlabel metal2 11454 16541 11454 16541 0 _0969_
rlabel metal1 26910 16014 26910 16014 0 _0970_
rlabel metal2 18722 31688 18722 31688 0 _0971_
rlabel metal1 18216 37230 18216 37230 0 _0972_
rlabel metal1 17158 37434 17158 37434 0 _0973_
rlabel metal1 17250 37910 17250 37910 0 _0974_
rlabel metal1 17848 37298 17848 37298 0 _0975_
rlabel metal1 17940 36346 17940 36346 0 _0976_
rlabel metal1 18630 37094 18630 37094 0 _0977_
rlabel via3 18285 17884 18285 17884 0 _0978_
rlabel metal1 16790 36210 16790 36210 0 _0979_
rlabel metal3 17503 35972 17503 35972 0 _0980_
rlabel metal2 18630 17034 18630 17034 0 _0981_
rlabel metal2 19090 16354 19090 16354 0 _0982_
rlabel metal1 30544 12818 30544 12818 0 _0983_
rlabel metal1 30544 11730 30544 11730 0 _0984_
rlabel metal1 31050 11322 31050 11322 0 _0985_
rlabel metal1 30682 16014 30682 16014 0 _0986_
rlabel metal1 26772 16082 26772 16082 0 _0987_
rlabel metal2 30084 15878 30084 15878 0 _0988_
rlabel metal1 30130 11220 30130 11220 0 _0989_
rlabel metal1 32660 16490 32660 16490 0 _0990_
rlabel metal2 33166 18972 33166 18972 0 _0991_
rlabel metal1 31372 17850 31372 17850 0 _0992_
rlabel metal1 32430 18700 32430 18700 0 _0993_
rlabel metal1 35420 19346 35420 19346 0 _0994_
rlabel metal1 36294 22678 36294 22678 0 _0995_
rlabel metal2 35972 20434 35972 20434 0 _0996_
rlabel metal1 35696 21522 35696 21522 0 _0997_
rlabel metal1 36386 23154 36386 23154 0 _0998_
rlabel metal1 35604 22678 35604 22678 0 _0999_
rlabel metal1 34960 21998 34960 21998 0 _1000_
rlabel metal1 31786 31824 31786 31824 0 _1001_
rlabel metal2 32062 30940 32062 30940 0 _1002_
rlabel metal1 33212 24786 33212 24786 0 _1003_
rlabel metal1 26082 31654 26082 31654 0 _1004_
rlabel metal1 26910 30906 26910 30906 0 _1005_
rlabel metal3 27945 37332 27945 37332 0 _1006_
rlabel metal2 33074 23936 33074 23936 0 _1007_
rlabel metal2 33350 24378 33350 24378 0 _1008_
rlabel metal1 34178 24242 34178 24242 0 _1009_
rlabel metal1 34178 24106 34178 24106 0 _1010_
rlabel metal1 32798 24276 32798 24276 0 _1011_
rlabel metal1 31188 28526 31188 28526 0 _1012_
rlabel metal2 31142 26588 31142 26588 0 _1013_
rlabel metal1 31786 24344 31786 24344 0 _1014_
rlabel metal1 25714 28730 25714 28730 0 _1015_
rlabel metal1 26358 29172 26358 29172 0 _1016_
rlabel metal1 27324 37774 27324 37774 0 _1017_
rlabel metal1 31694 24140 31694 24140 0 _1018_
rlabel metal1 31947 23698 31947 23698 0 _1019_
rlabel metal1 32568 23834 32568 23834 0 _1020_
rlabel metal1 32890 23120 32890 23120 0 _1021_
rlabel metal1 33396 22610 33396 22610 0 _1022_
rlabel metal2 33166 24412 33166 24412 0 _1023_
rlabel metal2 32706 22039 32706 22039 0 _1024_
rlabel metal1 31372 21998 31372 21998 0 _1025_
rlabel metal1 30774 21114 30774 21114 0 _1026_
rlabel metal1 30452 35666 30452 35666 0 _1027_
rlabel metal1 30268 35462 30268 35462 0 _1028_
rlabel metal1 29072 20434 29072 20434 0 _1029_
rlabel metal1 25944 35666 25944 35666 0 _1030_
rlabel metal2 25530 35326 25530 35326 0 _1031_
rlabel metal2 25990 34816 25990 34816 0 _1032_
rlabel metal1 29026 19856 29026 19856 0 _1033_
rlabel metal1 29854 19788 29854 19788 0 _1034_
rlabel metal1 30038 19856 30038 19856 0 _1035_
rlabel metal1 29946 19346 29946 19346 0 _1036_
rlabel metal1 30360 20434 30360 20434 0 _1037_
rlabel metal1 30360 19822 30360 19822 0 _1038_
rlabel metal2 20746 16626 20746 16626 0 _1039_
rlabel metal1 21022 17068 21022 17068 0 _1040_
rlabel via1 20378 16558 20378 16558 0 _1041_
rlabel metal1 21114 16082 21114 16082 0 _1042_
rlabel metal1 33810 9996 33810 9996 0 _1043_
rlabel metal1 20562 14348 20562 14348 0 _1044_
rlabel metal1 20792 14450 20792 14450 0 _1045_
rlabel metal2 19734 13702 19734 13702 0 _1046_
rlabel metal2 21114 13668 21114 13668 0 _1047_
rlabel metal2 21942 13872 21942 13872 0 _1048_
rlabel metal2 32338 17442 32338 17442 0 _1049_
rlabel metal1 31096 20434 31096 20434 0 _1050_
rlabel metal1 30682 19924 30682 19924 0 _1051_
rlabel metal1 35236 21658 35236 21658 0 _1052_
rlabel metal1 34638 19346 34638 19346 0 _1053_
rlabel metal1 34960 18598 34960 18598 0 _1054_
rlabel metal1 32338 17850 32338 17850 0 _1055_
rlabel metal2 29026 8398 29026 8398 0 _1056_
rlabel metal1 25898 6698 25898 6698 0 _1057_
rlabel metal1 21206 6732 21206 6732 0 _1058_
rlabel metal2 21666 10693 21666 10693 0 _1059_
rlabel metal1 25990 5202 25990 5202 0 _1060_
rlabel metal1 27048 7514 27048 7514 0 _1061_
rlabel metal1 25990 5134 25990 5134 0 _1062_
rlabel metal1 28290 8466 28290 8466 0 _1063_
rlabel metal1 29532 9146 29532 9146 0 _1064_
rlabel metal1 29854 11730 29854 11730 0 _1065_
rlabel metal1 25806 14960 25806 14960 0 _1066_
rlabel metal1 25668 13294 25668 13294 0 _1067_
rlabel metal1 26358 15470 26358 15470 0 _1068_
rlabel metal1 26220 12274 26220 12274 0 _1069_
rlabel viali 27196 13294 27196 13294 0 _1070_
rlabel metal1 27416 11118 27416 11118 0 _1071_
rlabel metal1 27002 9520 27002 9520 0 _1072_
rlabel metal1 27186 11696 27186 11696 0 _1073_
rlabel metal2 26680 12852 26680 12852 0 _1074_
rlabel metal1 26542 13974 26542 13974 0 _1075_
rlabel metal1 26910 12818 26910 12818 0 _1076_
rlabel metal1 26082 12954 26082 12954 0 _1077_
rlabel metal1 27646 12682 27646 12682 0 _1078_
rlabel metal2 32614 17952 32614 17952 0 _1079_
rlabel metal1 33534 18394 33534 18394 0 _1080_
rlabel metal1 34454 19380 34454 19380 0 _1081_
rlabel metal1 35328 19142 35328 19142 0 _1082_
rlabel metal1 35926 23154 35926 23154 0 _1083_
rlabel metal1 36064 22066 36064 22066 0 _1084_
rlabel metal1 33764 21930 33764 21930 0 _1085_
rlabel metal1 33258 24140 33258 24140 0 _1086_
rlabel metal1 33442 21998 33442 21998 0 _1087_
rlabel via2 31234 22083 31234 22083 0 _1088_
rlabel metal2 29670 20842 29670 20842 0 _1089_
rlabel metal1 30636 20230 30636 20230 0 _1090_
rlabel metal1 22448 14994 22448 14994 0 _1091_
rlabel metal1 29670 7310 29670 7310 0 _1092_
rlabel metal1 30314 19754 30314 19754 0 _1093_
rlabel metal1 31970 19788 31970 19788 0 _1094_
rlabel metal1 30130 16150 30130 16150 0 _1095_
rlabel metal1 30820 16218 30820 16218 0 _1096_
rlabel metal1 31694 15504 31694 15504 0 _1097_
rlabel metal1 32798 15538 32798 15538 0 _1098_
rlabel metal1 29854 16014 29854 16014 0 _1099_
rlabel metal1 32844 13906 32844 13906 0 _1100_
rlabel metal1 32706 15470 32706 15470 0 _1101_
rlabel metal2 33258 13702 33258 13702 0 _1102_
rlabel metal1 33166 12886 33166 12886 0 _1103_
rlabel metal1 30866 5542 30866 5542 0 _1104_
rlabel metal1 32614 6256 32614 6256 0 _1105_
rlabel metal2 26358 4420 26358 4420 0 _1106_
rlabel metal1 24058 4590 24058 4590 0 _1107_
rlabel metal1 19872 6290 19872 6290 0 _1108_
rlabel metal1 20240 10030 20240 10030 0 _1109_
rlabel metal1 19688 6290 19688 6290 0 _1110_
rlabel metal1 24196 4658 24196 4658 0 _1111_
rlabel metal1 26174 4556 26174 4556 0 _1112_
rlabel metal1 27048 5134 27048 5134 0 _1113_
rlabel metal1 32338 5644 32338 5644 0 _1114_
rlabel metal2 32154 5508 32154 5508 0 _1115_
rlabel metal1 32384 6290 32384 6290 0 _1116_
rlabel metal1 32706 6358 32706 6358 0 _1117_
rlabel metal1 32752 8942 32752 8942 0 _1118_
rlabel metal1 33488 12750 33488 12750 0 _1119_
rlabel metal1 33442 15538 33442 15538 0 _1120_
rlabel metal1 33028 15402 33028 15402 0 _1121_
rlabel metal2 23230 12784 23230 12784 0 _1122_
rlabel metal1 20470 10064 20470 10064 0 _1123_
rlabel metal1 32660 15674 32660 15674 0 _1124_
rlabel metal1 32292 15674 32292 15674 0 _1125_
rlabel metal2 32614 15232 32614 15232 0 _1126_
rlabel metal1 29716 11322 29716 11322 0 _1127_
rlabel metal1 29762 13498 29762 13498 0 _1128_
rlabel metal1 29072 13498 29072 13498 0 _1129_
rlabel metal2 28566 13498 28566 13498 0 _1130_
rlabel metal1 31280 12818 31280 12818 0 _1131_
rlabel metal1 32706 10642 32706 10642 0 _1132_
rlabel metal1 30774 9350 30774 9350 0 _1133_
rlabel metal1 32522 9418 32522 9418 0 _1134_
rlabel metal1 29992 8942 29992 8942 0 _1135_
rlabel metal2 30406 8364 30406 8364 0 _1136_
rlabel metal1 23000 6290 23000 6290 0 _1137_
rlabel metal1 19780 7446 19780 7446 0 _1138_
rlabel metal1 21758 7888 21758 7888 0 _1139_
rlabel via1 21030 10710 21030 10710 0 _1140_
rlabel metal1 21574 9962 21574 9962 0 _1141_
rlabel metal2 22678 7922 22678 7922 0 _1142_
rlabel metal1 27600 6222 27600 6222 0 _1143_
rlabel metal1 26542 5270 26542 5270 0 _1144_
rlabel metal2 27646 5712 27646 5712 0 _1145_
rlabel metal1 27922 6800 27922 6800 0 _1146_
rlabel metal1 31786 12818 31786 12818 0 _1147_
rlabel metal1 29762 13328 29762 13328 0 _1148_
rlabel metal1 29394 12818 29394 12818 0 _1149_
rlabel metal2 22310 16388 22310 16388 0 _1150_
rlabel metal2 32016 18292 32016 18292 0 _1151_
rlabel metal1 28014 13498 28014 13498 0 _1152_
rlabel metal1 28566 15470 28566 15470 0 _1153_
rlabel metal1 32568 11118 32568 11118 0 _1154_
rlabel metal1 30682 14382 30682 14382 0 _1155_
rlabel metal2 30774 15198 30774 15198 0 _1156_
rlabel metal1 27876 15538 27876 15538 0 _1157_
rlabel metal1 27416 15130 27416 15130 0 _1158_
rlabel metal1 21988 12818 21988 12818 0 _1159_
rlabel metal2 24150 13600 24150 13600 0 _1160_
rlabel metal2 26680 9588 26680 9588 0 _1161_
rlabel metal1 23736 13974 23736 13974 0 _1162_
rlabel metal1 21206 13192 21206 13192 0 _1163_
rlabel metal1 23046 13430 23046 13430 0 _1164_
rlabel metal1 24518 12818 24518 12818 0 _1165_
rlabel metal2 32614 13498 32614 13498 0 _1166_
rlabel metal1 25898 13974 25898 13974 0 _1167_
rlabel via1 22218 7395 22218 7395 0 _1168_
rlabel metal1 25990 13940 25990 13940 0 _1169_
rlabel metal1 24886 13940 24886 13940 0 _1170_
rlabel metal1 21712 12954 21712 12954 0 _1171_
rlabel metal2 21942 7718 21942 7718 0 _1172_
rlabel metal1 21896 11730 21896 11730 0 _1173_
rlabel via1 26450 11662 26450 11662 0 _1174_
rlabel metal1 26220 10982 26220 10982 0 _1175_
rlabel metal2 25254 12580 25254 12580 0 _1176_
rlabel metal2 24426 12580 24426 12580 0 _1177_
rlabel metal1 24840 12614 24840 12614 0 _1178_
rlabel metal1 25668 13770 25668 13770 0 _1179_
rlabel metal1 27738 14858 27738 14858 0 _1180_
rlabel metal1 28290 14960 28290 14960 0 _1181_
rlabel metal1 18630 21012 18630 21012 0 _1182_
rlabel metal1 25300 19890 25300 19890 0 _1183_
rlabel metal1 33304 36006 33304 36006 0 _1184_
rlabel metal2 20378 20604 20378 20604 0 _1185_
rlabel viali 21116 20434 21116 20434 0 _1186_
rlabel metal2 20930 20706 20930 20706 0 _1187_
rlabel metal1 23000 21522 23000 21522 0 _1188_
rlabel metal1 19918 19482 19918 19482 0 _1189_
rlabel metal1 20516 20026 20516 20026 0 _1190_
rlabel metal2 23138 21046 23138 21046 0 _1191_
rlabel metal1 25254 23120 25254 23120 0 _1192_
rlabel metal1 22126 21998 22126 21998 0 _1193_
rlabel metal1 14904 15062 14904 15062 0 _1194_
rlabel metal1 15134 14926 15134 14926 0 _1195_
rlabel metal1 14858 14892 14858 14892 0 _1196_
rlabel metal1 16606 16626 16606 16626 0 _1197_
rlabel metal1 15962 15538 15962 15538 0 _1198_
rlabel metal1 14214 15504 14214 15504 0 _1199_
rlabel metal1 15134 15674 15134 15674 0 _1200_
rlabel metal1 22724 21454 22724 21454 0 _1201_
rlabel metal2 24058 22338 24058 22338 0 _1202_
rlabel metal1 33258 33388 33258 33388 0 _1203_
rlabel metal1 33856 33626 33856 33626 0 _1204_
rlabel metal2 32890 13124 32890 13124 0 _1205_
rlabel metal1 32798 13498 32798 13498 0 _1206_
rlabel metal1 29762 12750 29762 12750 0 _1207_
rlabel metal1 32124 12886 32124 12886 0 _1208_
rlabel metal2 31878 13328 31878 13328 0 _1209_
rlabel metal1 25300 13362 25300 13362 0 _1210_
rlabel metal1 30636 14314 30636 14314 0 _1211_
rlabel metal1 30728 14246 30728 14246 0 _1212_
rlabel metal1 23966 8466 23966 8466 0 _1213_
rlabel metal1 25162 9078 25162 9078 0 _1214_
rlabel metal1 25990 13328 25990 13328 0 _1215_
rlabel metal1 27002 13328 27002 13328 0 _1216_
rlabel metal1 26864 12410 26864 12410 0 _1217_
rlabel metal1 27646 13498 27646 13498 0 _1218_
rlabel metal1 31464 13906 31464 13906 0 _1219_
rlabel metal1 31464 14042 31464 14042 0 _1220_
rlabel metal1 9798 20910 9798 20910 0 _1221_
rlabel metal1 30498 22073 30498 22073 0 _1222_
rlabel metal1 33304 17646 33304 17646 0 _1223_
rlabel metal2 5750 21335 5750 21335 0 _1224_
rlabel metal1 27094 21114 27094 21114 0 _1225_
rlabel metal2 26634 33286 26634 33286 0 _1226_
rlabel metal1 31832 8058 31832 8058 0 _1227_
rlabel metal1 31602 9452 31602 9452 0 _1228_
rlabel metal1 32936 10438 32936 10438 0 _1229_
rlabel metal1 26910 11084 26910 11084 0 _1230_
rlabel metal1 27186 10676 27186 10676 0 _1231_
rlabel metal1 26910 10642 26910 10642 0 _1232_
rlabel metal1 30130 10064 30130 10064 0 _1233_
rlabel metal1 30958 9554 30958 9554 0 _1234_
rlabel metal1 33626 9690 33626 9690 0 _1235_
rlabel metal1 32522 6732 32522 6732 0 _1236_
rlabel metal1 32936 6834 32936 6834 0 _1237_
rlabel metal1 30774 9112 30774 9112 0 _1238_
rlabel metal2 9430 21267 9430 21267 0 _1239_
rlabel metal2 33258 23052 33258 23052 0 _1240_
rlabel metal1 32798 22644 32798 22644 0 _1241_
rlabel metal1 32384 22746 32384 22746 0 _1242_
rlabel metal1 32292 22542 32292 22542 0 _1243_
rlabel metal1 32150 21862 32150 21862 0 _1244_
rlabel metal2 32614 21828 32614 21828 0 _1245_
rlabel metal1 12742 22576 12742 22576 0 _1246_
rlabel metal2 30866 32071 30866 32071 0 _1247_
rlabel metal1 29900 30906 29900 30906 0 _1248_
rlabel metal1 31878 7412 31878 7412 0 _1249_
rlabel metal1 30314 4692 30314 4692 0 _1250_
rlabel metal2 30222 5100 30222 5100 0 _1251_
rlabel metal1 30452 6766 30452 6766 0 _1252_
rlabel metal1 23046 9146 23046 9146 0 _1253_
rlabel metal1 23345 10710 23345 10710 0 _1254_
rlabel metal2 22218 11594 22218 11594 0 _1255_
rlabel metal1 24656 8602 24656 8602 0 _1256_
rlabel metal1 27784 8874 27784 8874 0 _1257_
rlabel metal1 26818 8976 26818 8976 0 _1258_
rlabel metal1 28382 8908 28382 8908 0 _1259_
rlabel metal2 27462 9486 27462 9486 0 _1260_
rlabel metal1 28198 8976 28198 8976 0 _1261_
rlabel metal1 29394 6766 29394 6766 0 _1262_
rlabel metal1 31004 6902 31004 6902 0 _1263_
rlabel metal1 31464 6970 31464 6970 0 _1264_
rlabel metal2 20194 20757 20194 20757 0 _1265_
rlabel metal1 34362 21522 34362 21522 0 _1266_
rlabel metal2 33534 21420 33534 21420 0 _1267_
rlabel metal2 33258 20842 33258 20842 0 _1268_
rlabel metal1 33350 28050 33350 28050 0 _1269_
rlabel metal1 34316 24922 34316 24922 0 _1270_
rlabel metal1 26726 4522 26726 4522 0 _1271_
rlabel metal1 27600 4794 27600 4794 0 _1272_
rlabel metal1 28106 5066 28106 5066 0 _1273_
rlabel metal2 28014 6596 28014 6596 0 _1274_
rlabel metal1 8418 15470 8418 15470 0 clk
rlabel metal1 31280 29614 31280 29614 0 clknet_0__0514_
rlabel metal1 18998 30566 18998 30566 0 clknet_0__0515_
rlabel metal2 20010 31807 20010 31807 0 clknet_0__0516_
rlabel metal1 20148 31926 20148 31926 0 clknet_0__0517_
rlabel metal1 9522 18360 9522 18360 0 clknet_0_clk
rlabel metal1 35098 29172 35098 29172 0 clknet_1_0__leaf__0514_
rlabel metal1 6670 35088 6670 35088 0 clknet_1_0__leaf__0515_
rlabel metal1 15916 38318 15916 38318 0 clknet_1_0__leaf__0516_
rlabel metal2 12742 37094 12742 37094 0 clknet_1_0__leaf__0517_
rlabel metal1 33948 32878 33948 32878 0 clknet_1_1__leaf__0514_
rlabel metal3 20263 35972 20263 35972 0 clknet_1_1__leaf__0515_
rlabel metal1 32798 35666 32798 35666 0 clknet_1_1__leaf__0516_
rlabel metal1 29578 38420 29578 38420 0 clknet_1_1__leaf__0517_
rlabel metal1 2622 7446 2622 7446 0 clknet_2_0__leaf_clk
rlabel metal1 13202 12852 13202 12852 0 clknet_2_1__leaf_clk
rlabel metal1 1426 19414 1426 19414 0 clknet_2_2__leaf_clk
rlabel metal1 15042 25874 15042 25874 0 clknet_2_3__leaf_clk
rlabel metal1 38134 8942 38134 8942 0 cs
rlabel metal3 820 11628 820 11628 0 gpi[0]
rlabel metal3 1096 6868 1096 6868 0 gpi[1]
rlabel metal1 31096 38998 31096 38998 0 gpi[23]
rlabel metal2 10994 1554 10994 1554 0 gpi[2]
rlabel metal2 8418 1027 8418 1027 0 gpi[3]
rlabel metal1 15640 38998 15640 38998 0 gpi[4]
rlabel metal1 37444 38930 37444 38930 0 gpi[5]
rlabel metal2 37398 1027 37398 1027 0 gpi[6]
rlabel metal2 20102 39899 20102 39899 0 gpi[7]
rlabel metal1 17618 39066 17618 39066 0 gpo[0]
rlabel metal3 820 4148 820 4148 0 gpo[10]
rlabel metal2 37950 10999 37950 10999 0 gpo[11]
rlabel metal3 820 8908 820 8908 0 gpo[12]
rlabel metal2 37858 15793 37858 15793 0 gpo[13]
rlabel metal1 782 39066 782 39066 0 gpo[14]
rlabel metal1 26818 39066 26818 39066 0 gpo[15]
rlabel metal2 17434 1520 17434 1520 0 gpo[16]
rlabel metal2 46 1554 46 1554 0 gpo[17]
rlabel metal3 820 25228 820 25228 0 gpo[18]
rlabel metal2 21942 39960 21942 39960 0 gpo[19]
rlabel metal3 820 15708 820 15708 0 gpo[1]
rlabel metal1 37904 38522 37904 38522 0 gpo[20]
rlabel metal2 13202 39967 13202 39967 0 gpo[21]
rlabel metal2 3910 959 3910 959 0 gpo[22]
rlabel metal2 1978 959 1978 959 0 gpo[23]
rlabel metal2 37858 36941 37858 36941 0 gpo[24]
rlabel metal3 820 18428 820 18428 0 gpo[25]
rlabel metal2 14858 959 14858 959 0 gpo[26]
rlabel metal1 37904 34510 37904 34510 0 gpo[27]
rlabel metal3 37958 1428 37958 1428 0 gpo[28]
rlabel metal1 9200 39066 9200 39066 0 gpo[29]
rlabel metal1 38134 20774 38134 20774 0 gpo[2]
rlabel metal2 6486 959 6486 959 0 gpo[30]
rlabel metal2 12926 1520 12926 1520 0 gpo[31]
rlabel metal3 751 20468 751 20468 0 gpo[32]
rlabel via2 37858 22491 37858 22491 0 gpo[33]
rlabel metal2 19366 959 19366 959 0 gpo[3]
rlabel metal1 35604 39066 35604 39066 0 gpo[4]
rlabel metal2 33166 39423 33166 39423 0 gpo[5]
rlabel metal1 4738 39066 4738 39066 0 gpo[6]
rlabel metal1 11362 39066 11362 39066 0 gpo[7]
rlabel metal2 26450 1520 26450 1520 0 gpo[8]
rlabel metal3 1096 13668 1096 13668 0 gpo[9]
rlabel metal1 36892 18734 36892 18734 0 net1
rlabel metal2 14950 20094 14950 20094 0 net10
rlabel metal1 4922 33966 4922 33966 0 net100
rlabel metal1 13202 38318 13202 38318 0 net101
rlabel metal1 21758 38318 21758 38318 0 net102
rlabel metal1 25714 27438 25714 27438 0 net103
rlabel metal1 32752 35122 32752 35122 0 net104
rlabel metal1 33442 26996 33442 26996 0 net105
rlabel metal1 34454 31348 34454 31348 0 net106
rlabel metal1 31832 28186 31832 28186 0 net107
rlabel metal1 27692 32538 27692 32538 0 net108
rlabel metal1 25254 38318 25254 38318 0 net109
rlabel metal1 20378 37400 20378 37400 0 net11
rlabel metal1 29854 37230 29854 37230 0 net110
rlabel metal1 10258 24922 10258 24922 0 net111
rlabel metal2 9246 35802 9246 35802 0 net112
rlabel metal1 10166 28526 10166 28526 0 net113
rlabel metal1 9430 31790 9430 31790 0 net114
rlabel metal1 8832 29614 8832 29614 0 net115
rlabel metal1 8832 33490 8832 33490 0 net116
rlabel metal1 9246 38318 9246 38318 0 net117
rlabel metal1 19136 38318 19136 38318 0 net118
rlabel metal1 27554 26996 27554 26996 0 net119
rlabel metal1 18170 38522 18170 38522 0 net12
rlabel metal1 28658 34612 28658 34612 0 net120
rlabel metal1 29486 26996 29486 26996 0 net121
rlabel metal1 27278 29172 27278 29172 0 net122
rlabel metal1 29210 29172 29210 29172 0 net123
rlabel metal2 27738 31450 27738 31450 0 net124
rlabel metal1 27462 38386 27462 38386 0 net125
rlabel metal1 29118 37876 29118 37876 0 net126
rlabel metal1 28934 24820 28934 24820 0 net127
rlabel metal2 8878 5848 8878 5848 0 net128
rlabel metal1 11079 4794 11079 4794 0 net129
rlabel metal2 3910 6698 3910 6698 0 net13
rlabel metal1 9614 5270 9614 5270 0 net130
rlabel metal1 8740 6222 8740 6222 0 net131
rlabel metal1 12696 8058 12696 8058 0 net132
rlabel metal1 14076 5542 14076 5542 0 net133
rlabel metal1 16054 4624 16054 4624 0 net134
rlabel metal1 17250 5338 17250 5338 0 net135
rlabel metal1 7958 32980 7958 32980 0 net136
rlabel metal1 7498 29138 7498 29138 0 net137
rlabel metal1 8050 30260 8050 30260 0 net138
rlabel metal1 7866 31824 7866 31824 0 net139
rlabel via2 17526 10523 17526 10523 0 net14
rlabel metal1 9706 23086 9706 23086 0 net140
rlabel metal1 11270 5610 11270 5610 0 net141
rlabel metal1 2277 8942 2277 8942 0 net15
rlabel metal1 34730 16048 34730 16048 0 net16
rlabel metal2 1794 37405 1794 37405 0 net17
rlabel metal1 23092 17850 23092 17850 0 net18
rlabel metal1 17526 2414 17526 2414 0 net19
rlabel metal1 9062 19890 9062 19890 0 net2
rlabel metal2 1794 2618 1794 2618 0 net20
rlabel metal1 2024 23290 2024 23290 0 net21
rlabel metal2 22862 21267 22862 21267 0 net22
rlabel metal2 1794 15946 1794 15946 0 net23
rlabel metal1 37582 38216 37582 38216 0 net24
rlabel metal1 12788 38930 12788 38930 0 net25
rlabel metal1 4922 2414 4922 2414 0 net26
rlabel metal1 2346 2414 2346 2414 0 net27
rlabel via3 13915 21692 13915 21692 0 net28
rlabel metal1 1932 17850 1932 17850 0 net29
rlabel metal1 8602 14994 8602 14994 0 net3
rlabel metal1 14996 2414 14996 2414 0 net30
rlabel metal2 36938 34102 36938 34102 0 net31
rlabel metal1 37352 18054 37352 18054 0 net32
rlabel metal1 9016 38522 9016 38522 0 net33
rlabel metal1 37490 20842 37490 20842 0 net34
rlabel metal1 7682 2414 7682 2414 0 net35
rlabel metal1 13064 2414 13064 2414 0 net36
rlabel metal1 1840 20910 1840 20910 0 net37
rlabel metal1 37628 22610 37628 22610 0 net38
rlabel metal2 19826 2618 19826 2618 0 net39
rlabel metal2 13570 20621 13570 20621 0 net4
rlabel metal1 35282 38522 35282 38522 0 net40
rlabel metal1 32660 38522 32660 38522 0 net41
rlabel metal1 5060 38522 5060 38522 0 net42
rlabel metal2 12374 38488 12374 38488 0 net43
rlabel metal1 19366 2312 19366 2312 0 net44
rlabel metal1 1794 13872 1794 13872 0 net45
rlabel metal1 2622 23018 2622 23018 0 net46
rlabel metal1 6670 7854 6670 7854 0 net47
rlabel metal2 13938 26741 13938 26741 0 net48
rlabel metal1 33580 18190 33580 18190 0 net49
rlabel metal1 10672 2618 10672 2618 0 net5
rlabel metal1 18216 35258 18216 35258 0 net50
rlabel metal1 15318 36176 15318 36176 0 net51
rlabel metal2 19090 25381 19090 25381 0 net52
rlabel metal2 18262 27455 18262 27455 0 net53
rlabel metal2 13754 29546 13754 29546 0 net54
rlabel metal2 21942 33422 21942 33422 0 net55
rlabel metal1 20010 24276 20010 24276 0 net56
rlabel metal2 2806 13600 2806 13600 0 net57
rlabel metal1 12558 15368 12558 15368 0 net58
rlabel metal2 8326 35326 8326 35326 0 net59
rlabel metal1 8740 2618 8740 2618 0 net6
rlabel metal1 10297 37230 10297 37230 0 net60
rlabel metal1 15555 5270 15555 5270 0 net61
rlabel metal2 33718 35938 33718 35938 0 net62
rlabel metal1 21068 37774 21068 37774 0 net63
rlabel metal1 34592 32878 34592 32878 0 net64
rlabel metal1 35144 26010 35144 26010 0 net65
rlabel metal1 34914 29274 34914 29274 0 net66
rlabel metal1 34730 25330 34730 25330 0 net67
rlabel metal1 29854 31314 29854 31314 0 net68
rlabel metal1 27002 33524 27002 33524 0 net69
rlabel metal2 15594 38743 15594 38743 0 net7
rlabel metal1 34592 33966 34592 33966 0 net70
rlabel metal1 10718 23086 10718 23086 0 net71
rlabel metal1 7038 33524 7038 33524 0 net72
rlabel metal1 6670 26996 6670 26996 0 net73
rlabel metal2 4278 30362 4278 30362 0 net74
rlabel metal1 6118 28594 6118 28594 0 net75
rlabel metal1 4186 31790 4186 31790 0 net76
rlabel metal1 8694 23732 8694 23732 0 net77
rlabel metal1 4738 26350 4738 26350 0 net78
rlabel metal2 7314 24922 7314 24922 0 net79
rlabel via2 37674 38811 37674 38811 0 net8
rlabel metal1 6854 35054 6854 35054 0 net80
rlabel metal1 7682 28084 7682 28084 0 net81
rlabel metal2 7866 31450 7866 31450 0 net82
rlabel metal1 3910 29172 3910 29172 0 net83
rlabel metal1 4278 32878 4278 32878 0 net84
rlabel metal1 8832 37230 8832 37230 0 net85
rlabel metal1 20378 37230 20378 37230 0 net86
rlabel metal1 25668 24242 25668 24242 0 net87
rlabel metal1 30590 35054 30590 35054 0 net88
rlabel metal1 30958 26350 30958 26350 0 net89
rlabel metal1 17595 2482 17595 2482 0 net9
rlabel metal2 34546 31518 34546 31518 0 net90
rlabel metal1 34822 28186 34822 28186 0 net91
rlabel metal1 31326 32538 31326 32538 0 net92
rlabel metal2 27462 36074 27462 36074 0 net93
rlabel metal1 32338 36788 32338 36788 0 net94
rlabel metal2 8694 26010 8694 26010 0 net95
rlabel metal1 5934 36142 5934 36142 0 net96
rlabel metal1 9706 27438 9706 27438 0 net97
rlabel metal1 5842 30702 5842 30702 0 net98
rlabel metal1 4094 28084 4094 28084 0 net99
rlabel metal3 820 36788 820 36788 0 nrst
rlabel metal1 38134 18054 38134 18054 0 store_en
<< properties >>
string FIXED_BBOX 0 0 39418 41562
<< end >>
