* NGSPICE file created from Guitar_Villains.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_12 abstract view
.subckt sky130_fd_sc_hd__buf_12 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_4 abstract view
.subckt sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_4 abstract view
.subckt sky130_fd_sc_hd__nor2b_4 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_12 abstract view
.subckt sky130_fd_sc_hd__inv_12 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_4 abstract view
.subckt sky130_fd_sc_hd__o32a_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

.subckt Guitar_Villains VGND VPWR bottom_row[0] bottom_row[1] bottom_row[2] bottom_row[3]
+ bottom_row[4] bottom_row[5] bottom_row[6] button[0] button[1] button[2] button[3]
+ chip_select clk green_disp n_rst red_disp ss0[0] ss0[1] ss0[2] ss0[3] ss0[4] ss0[5]
+ ss0[6] ss1[0] ss1[1] ss1[2] ss1[3] ss1[4] ss1[5] ss1[6] top_row[0] top_row[1] top_row[2]
+ top_row[3] top_row[4] top_row[5] top_row[6]
XFILLER_0_94_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3155_ game.addmisses.a\[15\] game.addmisses.add4.b\[3\] VGND VGND VPWR VPWR _0518_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_27_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3086_ _0447_ _0448_ VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__nand2_2
XFILLER_0_89_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3988_ _0209_ _2658_ VGND VGND VPWR VPWR _1303_ sky130_fd_sc_hd__nand2_2
XFILLER_0_91_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2939_ _0276_ _0339_ disp_song.note2\[26\] VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_17_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5727_ clknet_leaf_4_clk _0002_ net49 VGND VGND VPWR VPWR lvls.level\[2\] sky130_fd_sc_hd__dfrtp_4
X_5658_ game.flash_counter\[15\] game.flash_counter\[14\] game.flash_counter\[13\]
+ VGND VGND VPWR VPWR _2627_ sky130_fd_sc_hd__and3_1
XFILLER_0_13_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4609_ game.scoring_button_1.flash_counter_1\[17\] game.scoring_button_1.flash_counter_1\[16\]
+ game.scoring_button_1.flash_counter_1\[19\] game.scoring_button_1.flash_counter_1\[18\]
+ VGND VGND VPWR VPWR _1797_ sky130_fd_sc_hd__and4_1
X_5589_ _2584_ game.padded_notes1\[27\] _2472_ VGND VGND VPWR VPWR _2585_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_578 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4960_ disp_song.um.drum.next_note2\[10\] disp_song.um.drum.next_note2\[11\] _1956_
+ VGND VGND VPWR VPWR _2054_ sky130_fd_sc_hd__mux2_1
X_4891_ _1956_ disp_song.um.drum.next_note2\[11\] _1985_ VGND VGND VPWR VPWR _1986_
+ sky130_fd_sc_hd__o21ai_1
X_3911_ _1237_ _1240_ VGND VGND VPWR VPWR _1241_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3842_ _0966_ disp_song.toggle_green _0262_ modetrans.mode\[3\] _1190_ VGND VGND
+ VPWR VPWR _1191_ sky130_fd_sc_hd__a221o_2
XFILLER_0_46_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5512_ disp_song.note1\[2\] game.padded_notes1\[1\] _2497_ VGND VGND VPWR VPWR _2533_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3773_ _0261_ _1122_ _1124_ _1126_ VGND VGND VPWR VPWR _1127_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2724_ _0169_ VGND VGND VPWR VPWR disp_song.um.drum.next_idx2\[2\] sky130_fd_sc_hd__inv_4
X_5443_ _2491_ net231 _2473_ VGND VGND VPWR VPWR _2492_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5374_ _0858_ highest_score.highest_score\[6\] _2434_ VGND VGND VPWR VPWR _2446_
+ sky130_fd_sc_hd__mux2_1
X_4325_ game.scoring_button_2.flash_counter_1\[3\] _1562_ VGND VGND VPWR VPWR _1565_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_10_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4256_ net201 _1514_ _1517_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_2\[4\]
+ sky130_fd_sc_hd__o21a_1
X_4187_ _1460_ _1461_ VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__nor2_1
X_3207_ game.addhits.a\[7\] game.addhits.add2.b\[3\] VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__nor2_1
X_3138_ _0495_ _0497_ _0493_ VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__or3b_1
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3069_ _0400_ _0419_ _0433_ net197 VGND VGND VPWR VPWR disp_song.um.drum.next_note1\[30\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold170 game.padded_notes1\[13\] VGND VGND VPWR VPWR net243 sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 game.padded_notes2\[4\] VGND VGND VPWR VPWR net254 sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 pulseout.fin_pulse\[5\] VGND VGND VPWR VPWR net265 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5090_ _2176_ _2178_ disp_song.um.drum.next_idx2\[4\] VGND VGND VPWR VPWR _2179_
+ sky130_fd_sc_hd__mux2_1
X_4110_ game.scoring_button_2.flash_counter_1\[8\] game.scoring_button_2.flash_counter_1\[11\]
+ game.scoring_button_2.flash_counter_1\[10\] game.scoring_button_2.flash_counter_1\[9\]
+ VGND VGND VPWR VPWR _1409_ sky130_fd_sc_hd__or4b_1
XFILLER_0_75_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4041_ game.addmisses.add2.b\[2\] game.addmisses.add2.b\[1\] _1327_ game.addmisses.add2.b\[3\]
+ VGND VGND VPWR VPWR _1349_ sky130_fd_sc_hd__a31o_1
XFILLER_0_38_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5992_ clknet_leaf_37_clk _0101_ net71 VGND VGND VPWR VPWR game.padded_notes1\[11\]
+ sky130_fd_sc_hd__dfstp_1
X_4943_ _1956_ disp_song.um.drum.next_note2\[23\] _1968_ _2036_ disp_song.um.drum.next_note2\[22\]
+ VGND VGND VPWR VPWR _2037_ sky130_fd_sc_hd__a32o_1
XFILLER_0_59_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4874_ disp_song.um.drum.next_note2\[16\] disp_song.um.drum.next_note2\[17\] _2670_
+ VGND VGND VPWR VPWR _1969_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3825_ disp_song.mi6.in\[2\] _1105_ _1104_ disp_song.mi6.in\[3\] VGND VGND VPWR VPWR
+ _1176_ sky130_fd_sc_hd__a211o_1
X_3756_ disp_song.mi6.in\[3\] _1105_ _1110_ _1081_ _0925_ VGND VGND VPWR VPWR _1111_
+ sky130_fd_sc_hd__a2111o_1
X_2707_ _2678_ VGND VGND VPWR VPWR _2679_ sky130_fd_sc_hd__clkbuf_4
X_5426_ _2480_ VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3687_ _0642_ _1040_ VGND VGND VPWR VPWR _1043_ sky130_fd_sc_hd__or2b_1
XFILLER_0_100_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5357_ _1034_ highest_score.highest_score\[0\] _2434_ VGND VGND VPWR VPWR _2435_
+ sky130_fd_sc_hd__mux2_1
X_5288_ _2185_ _2192_ _2197_ VGND VGND VPWR VPWR _2372_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_10_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4308_ game.scoring_button_2.flash_counter_2\[19\] game.scoring_button_2.flash_counter_2\[18\]
+ _1546_ game.scoring_button_2.flash_counter_2\[20\] VGND VGND VPWR VPWR _1554_ sky130_fd_sc_hd__a31o_1
X_4239_ game.counter\[15\] _0222_ _0229_ _0230_ _1505_ VGND VGND VPWR VPWR _1506_
+ sky130_fd_sc_hd__o2111a_1
XFILLER_0_97_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4590_ game.addmisses.a\[14\] _1767_ _1771_ VGND VGND VPWR VPWR _1780_ sky130_fd_sc_hd__and3_1
X_3610_ _0914_ _0969_ VGND VGND VPWR VPWR _0970_ sky130_fd_sc_hd__and2b_1
XFILLER_0_101_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3541_ _0901_ _0903_ VGND VGND VPWR VPWR _0904_ sky130_fd_sc_hd__nand2_1
XFILLER_0_52_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3472_ _0821_ _0828_ _0830_ _0834_ VGND VGND VPWR VPWR _0835_ sky130_fd_sc_hd__a2bb2o_1
X_5211_ disp_song.um.drum.next_note1\[1\] _2191_ disp_song.um.drum.next_idx1\[0\]
+ VGND VGND VPWR VPWR _2298_ sky130_fd_sc_hd__a21oi_1
X_5142_ _0198_ _2208_ VGND VGND VPWR VPWR _2230_ sky130_fd_sc_hd__and2_1
X_5073_ _2157_ _2160_ _2161_ _2162_ VGND VGND VPWR VPWR _2163_ sky130_fd_sc_hd__o22a_1
X_4024_ game.addmisses.add2.b\[1\] _1327_ VGND VGND VPWR VPWR _1334_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5975_ clknet_leaf_34_clk game.scoring_button_1.next_flash_counter_2\[20\] net72
+ VGND VGND VPWR VPWR game.scoring_button_1.flash_counter_2\[20\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4926_ _2009_ _2019_ VGND VGND VPWR VPWR _2020_ sky130_fd_sc_hd__nand2_4
X_4857_ _0162_ _1951_ VGND VGND VPWR VPWR _1952_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3808_ _0966_ _1114_ _1159_ modetrans.mode\[5\] lvls.level\[1\] VGND VGND VPWR VPWR
+ _1160_ sky130_fd_sc_hd__a32o_1
XFILLER_0_105_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4788_ game.scoring_button_1.flash_counter_1\[13\] game.scoring_button_1.flash_counter_1\[12\]
+ _1905_ game.scoring_button_1.flash_counter_1\[14\] VGND VGND VPWR VPWR _1913_ sky130_fd_sc_hd__a31o_1
XFILLER_0_43_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3739_ _1070_ _1093_ _1065_ VGND VGND VPWR VPWR _1094_ sky130_fd_sc_hd__a21o_1
X_5409_ _2468_ VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2972_ _2661_ _0352_ VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__or2_1
X_5760_ clknet_leaf_47_clk game.scoring_button_2.next_missed net56 VGND VGND VPWR
+ VPWR game.missed_2 sky130_fd_sc_hd__dfrtp_4
X_4711_ net184 _1857_ game.missed_1 VGND VGND VPWR VPWR _1860_ sky130_fd_sc_hd__a21boi_1
XTAP_1290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5691_ disp_song.next_red disp_song.next_green _2650_ VGND VGND VPWR VPWR _2651_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4642_ _1814_ VGND VGND VPWR VPWR game.scoring_button_1.next_count\[14\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4573_ game.addmisses.a\[12\] _1749_ VGND VGND VPWR VPWR _1765_ sky130_fd_sc_hd__and2_1
XFILLER_0_52_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3524_ _0608_ _0675_ _0886_ VGND VGND VPWR VPWR _0887_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3455_ _0791_ _0817_ _0793_ VGND VGND VPWR VPWR _0818_ sky130_fd_sc_hd__o21ai_1
X_3386_ _0527_ _0748_ _0524_ VGND VGND VPWR VPWR _0749_ sky130_fd_sc_hd__and3_1
X_6174_ clknet_leaf_45_clk disp_song.um.drum.next_d1\[6\] net54 VGND VGND VPWR VPWR
+ disp_song.display_note1\[6\] sky130_fd_sc_hd__dfrtp_1
X_5125_ disp_song.um.drum.next_idx1\[1\] _2210_ _2212_ _2189_ VGND VGND VPWR VPWR
+ _2213_ sky130_fd_sc_hd__o211a_1
X_5056_ disp_song.um.drum.next_idx2\[1\] _2081_ _1995_ VGND VGND VPWR VPWR _2147_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_98_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4007_ _1305_ _1317_ VGND VGND VPWR VPWR _1320_ sky130_fd_sc_hd__nor2_1
X_5958_ clknet_leaf_36_clk game.scoring_button_1.next_flash_counter_2\[3\] net72 VGND
+ VGND VPWR VPWR game.scoring_button_1.flash_counter_2\[3\] sky130_fd_sc_hd__dfrtp_1
X_4909_ disp_song.um.drum.next_note2\[4\] disp_song.um.drum.next_note2\[5\] disp_song.um.drum.next_idx2\[0\]
+ VGND VGND VPWR VPWR _2004_ sky130_fd_sc_hd__mux2_1
X_5889_ clknet_leaf_31_clk _0072_ net69 VGND VGND VPWR VPWR game.padded_notes2\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_586 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold41 modetrans.u2.Q2 VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__dlygate4sd3_1
Xhold30 game.scoring_button_2.flash_counter_1\[1\] VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 pulseout.fin_pulse\[4\] VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 game.flash_counter\[22\] VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold63 _0087_ VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__dlygate4sd3_1
Xhold85 game.scoring_button_1.flash_counter_2\[10\] VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold96 game.scoring_button_2.flash_counter_2\[19\] VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_5 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_111_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3240_ _0576_ _0577_ _0537_ VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__a21oi_1
X_3171_ _0532_ _0533_ VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__nand2_1
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5812_ clknet_leaf_47_clk game.scoring_button_2.next_flash_counter_2\[3\] net56 VGND
+ VGND VPWR VPWR game.scoring_button_2.flash_counter_2\[3\] sky130_fd_sc_hd__dfrtp_1
X_5743_ clknet_leaf_69_clk game.scoring_button_2.next_num_misses\[15\] net46 VGND
+ VGND VPWR VPWR game.addmisses.add4.b\[3\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_8_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2955_ _2661_ _0183_ _0264_ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__or3b_1
XFILLER_0_57_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_223 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2886_ _0279_ _0298_ VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__nor2_1
X_5674_ _2614_ _2637_ _2638_ VGND VGND VPWR VPWR _2639_ sky130_fd_sc_hd__and3_1
X_4625_ _1791_ _1426_ VGND VGND VPWR VPWR _1806_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4556_ game.addmisses.a\[11\] _1747_ _1748_ VGND VGND VPWR VPWR _1751_ sky130_fd_sc_hd__and3b_1
XFILLER_0_25_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3507_ game.flash_counter\[9\] game.flash_counter\[8\] _0869_ VGND VGND VPWR VPWR
+ _0870_ sky130_fd_sc_hd__and3_1
XFILLER_0_12_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4487_ _1690_ VGND VGND VPWR VPWR _1691_ sky130_fd_sc_hd__clkbuf_4
X_3438_ _0800_ _0693_ VGND VGND VPWR VPWR _0801_ sky130_fd_sc_hd__xnor2_1
X_6157_ clknet_leaf_13_clk net76 net58 VGND VGND VPWR VPWR disp_song.um.boton1e.edge_1
+ sky130_fd_sc_hd__dfrtp_2
X_3369_ game.addhits.a\[14\] game.addhits.add4.b\[2\] VGND VGND VPWR VPWR _0732_ sky130_fd_sc_hd__nor2_1
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5108_ disp_song.um.drum.next_note1\[14\] disp_song.um.drum.next_note1\[15\] disp_song.um.drum.next_idx1\[0\]
+ VGND VGND VPWR VPWR _2196_ sky130_fd_sc_hd__mux2_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6088_ clknet_leaf_23_clk disp_song.um.drum.next_note1\[0\] net64 VGND VGND VPWR
+ VPWR disp_song.note1\[0\] sky130_fd_sc_hd__dfrtp_1
X_5039_ _2109_ _2118_ _2130_ _1950_ VGND VGND VPWR VPWR _2131_ sky130_fd_sc_hd__a211o_1
XFILLER_0_95_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput20 net20 VGND VGND VPWR VPWR ss0[4] sky130_fd_sc_hd__clkbuf_4
Xoutput31 net31 VGND VGND VPWR VPWR top_row[1] sky130_fd_sc_hd__clkbuf_4
Xoutput7 net7 VGND VGND VPWR VPWR bottom_row[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2740_ _0170_ _0182_ disp_song.um.idx_note1\[4\] VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_26_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4410_ game.addhits.a\[3\] _1620_ VGND VGND VPWR VPWR _1629_ sky130_fd_sc_hd__nand2_1
X_5390_ net147 _2454_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_111_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4341_ game.scoring_button_2.flash_counter_1\[7\] game.scoring_button_2.flash_counter_1\[8\]
+ _1572_ VGND VGND VPWR VPWR _1576_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4272_ game.scoring_button_2.flash_counter_2\[9\] _1525_ VGND VGND VPWR VPWR _1529_
+ sky130_fd_sc_hd__or2_1
X_3223_ game.addhits.a\[11\] game.addhits.add3.b\[3\] VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__nor2_1
X_6011_ clknet_leaf_48_clk _0120_ net56 VGND VGND VPWR VPWR game.padded_notes1\[30\]
+ sky130_fd_sc_hd__dfstp_1
X_3154_ game.addmisses.a\[15\] game.addmisses.add4.b\[3\] VGND VGND VPWR VPWR _0517_
+ sky130_fd_sc_hd__nand2_1
X_3085_ game.addmisses.a\[4\] game.addmisses.add2.b\[0\] VGND VGND VPWR VPWR _0448_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_49_304 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3987_ _1290_ _1292_ _1296_ _1301_ VGND VGND VPWR VPWR _1302_ sky130_fd_sc_hd__o31a_1
XFILLER_0_91_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2938_ _2656_ _0335_ VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__or2_1
X_5726_ clknet_leaf_4_clk _0001_ net49 VGND VGND VPWR VPWR lvls.level\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_60_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2869_ _0290_ VGND VGND VPWR VPWR disp_song.um.drum.next_note2\[6\] sky130_fd_sc_hd__buf_1
X_5657_ net121 _2624_ VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5588_ disp_song.note1\[27\] game.padded_notes1\[26\] _0209_ VGND VGND VPWR VPWR
+ _2584_ sky130_fd_sc_hd__mux2_1
X_4608_ game.scoring_button_1.flash_counter_1\[21\] game.scoring_button_1.flash_counter_1\[20\]
+ game.scoring_button_1.flash_counter_1\[22\] VGND VGND VPWR VPWR _1796_ sky130_fd_sc_hd__or3_1
XFILLER_0_13_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4539_ _1675_ _1721_ VGND VGND VPWR VPWR _1736_ sky130_fd_sc_hd__nor2_1
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_3_6__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_6__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_68_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4890_ disp_song.um.drum.next_idx2\[0\] disp_song.um.drum.next_note2\[10\] VGND VGND
+ VPWR VPWR _1985_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3910_ _1232_ _1239_ VGND VGND VPWR VPWR _1240_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_58_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3841_ game.hit_1 game.hit_2 _0210_ VGND VGND VPWR VPWR _1190_ sky130_fd_sc_hd__o21a_1
XFILLER_0_104_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3772_ _0258_ _1125_ VGND VGND VPWR VPWR _1126_ sky130_fd_sc_hd__nand2_1
X_5511_ _2532_ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__clkbuf_1
X_2723_ _0168_ VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_42_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5442_ disp_song.note2\[14\] game.padded_notes2\[13\] _0219_ VGND VGND VPWR VPWR
+ _2491_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5373_ _2445_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__clkbuf_1
X_4324_ _1564_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_1\[2\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_22_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4255_ game.scoring_button_2.flash_counter_2\[4\] _1514_ game.missed_2 VGND VGND
+ VPWR VPWR _1517_ sky130_fd_sc_hd__a21boi_1
X_4186_ game.counter\[17\] _1457_ VGND VGND VPWR VPWR _1461_ sky130_fd_sc_hd__and2_1
X_3206_ _0563_ _0568_ VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__nor2_2
XFILLER_0_38_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3137_ _0493_ _0498_ _0499_ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3068_ _0400_ _0421_ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5709_ clknet_leaf_23_clk modetrans.pushed_4 net64 VGND VGND VPWR VPWR modetrans.u3.sync_pb
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold160 game.padded_notes2\[28\] VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 disp_song.note2\[29\] VGND VGND VPWR VPWR net244 sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 disp_song.note2\[31\] VGND VGND VPWR VPWR net255 sky130_fd_sc_hd__dlygate4sd3_1
Xhold193 disp_song.um.idx_note2\[2\] VGND VGND VPWR VPWR net266 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4040_ _1348_ VGND VGND VPWR VPWR game.scoring_button_2.next_num_misses\[6\] sky130_fd_sc_hd__clkbuf_1
X_5991_ clknet_leaf_37_clk _0100_ net71 VGND VGND VPWR VPWR game.padded_notes1\[10\]
+ sky130_fd_sc_hd__dfstp_1
X_4942_ _2035_ _2016_ VGND VGND VPWR VPWR _2036_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4873_ _1967_ VGND VGND VPWR VPWR _1968_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_74_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3824_ _1086_ _0927_ _1116_ VGND VGND VPWR VPWR _1175_ sky130_fd_sc_hd__and3b_1
XFILLER_0_104_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3755_ _1105_ _1107_ disp_song.mi6.in\[3\] VGND VGND VPWR VPWR _1110_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2706_ _2654_ _2677_ VGND VGND VPWR VPWR _2678_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3686_ _0642_ _1040_ _1041_ VGND VGND VPWR VPWR _1042_ sky130_fd_sc_hd__a21oi_1
X_5425_ _2479_ net209 _2473_ VGND VGND VPWR VPWR _2480_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5356_ _2433_ VGND VGND VPWR VPWR _2434_ sky130_fd_sc_hd__buf_2
X_5287_ _2201_ _2220_ _2365_ VGND VGND VPWR VPWR _2371_ sky130_fd_sc_hd__mux2_1
X_4307_ game.scoring_button_2.flash_counter_2\[19\] game.scoring_button_2.flash_counter_2\[20\]
+ _1549_ VGND VGND VPWR VPWR _1553_ sky130_fd_sc_hd__and3_1
X_4238_ _0249_ _0223_ VGND VGND VPWR VPWR _1505_ sky130_fd_sc_hd__and2b_1
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4169_ _1405_ _0013_ VGND VGND VPWR VPWR _1448_ sky130_fd_sc_hd__and2_1
XFILLER_0_92_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3540_ highest_score.highest_score\[6\] highest_score.highest_score\[5\] highest_score.highest_score\[4\]
+ _0899_ VGND VGND VPWR VPWR _0903_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_101_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3471_ _0833_ VGND VGND VPWR VPWR _0834_ sky130_fd_sc_hd__buf_2
XFILLER_0_51_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5210_ _2295_ _2296_ _2254_ VGND VGND VPWR VPWR _2297_ sky130_fd_sc_hd__mux2_1
X_5141_ _2227_ _2228_ disp_song.um.drum.next_idx1\[1\] VGND VGND VPWR VPWR _2229_
+ sky130_fd_sc_hd__mux2_1
X_5072_ _2034_ _2021_ _2157_ VGND VGND VPWR VPWR _2162_ sky130_fd_sc_hd__o21ai_1
X_4023_ _1326_ _1328_ _1333_ _1289_ VGND VGND VPWR VPWR game.scoring_button_2.next_num_misses\[4\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5974_ clknet_leaf_32_clk game.scoring_button_1.next_flash_counter_2\[19\] net71
+ VGND VGND VPWR VPWR game.scoring_button_1.flash_counter_2\[19\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4925_ _2667_ _2670_ VGND VGND VPWR VPWR _2019_ sky130_fd_sc_hd__nand2_2
X_4856_ disp_song.um.drum.next_idx2\[3\] _1948_ VGND VGND VPWR VPWR _1951_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3807_ _0925_ _1084_ _1158_ VGND VGND VPWR VPWR _1159_ sky130_fd_sc_hd__o21ai_1
X_4787_ game.scoring_button_1.flash_counter_1\[13\] game.scoring_button_1.flash_counter_1\[14\]
+ _1908_ VGND VGND VPWR VPWR _1912_ sky130_fd_sc_hd__and3_1
XFILLER_0_55_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3738_ _0629_ _1092_ VGND VGND VPWR VPWR _1093_ sky130_fd_sc_hd__nand2_1
X_3669_ _1021_ _1022_ _1024_ VGND VGND VPWR VPWR _1025_ sky130_fd_sc_hd__and3_1
X_5408_ _2467_ game.padded_notes2\[3\] _2462_ VGND VGND VPWR VPWR _2468_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5339_ highest_score.highest_score\[1\] _1028_ _1029_ _1030_ VGND VGND VPWR VPWR
+ _2417_ sky130_fd_sc_hd__or4_1
XFILLER_0_108_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_58_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_58_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_88_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2971_ _0194_ _0363_ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__nand2_2
XFILLER_0_29_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4710_ _1859_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_2\[12\]
+ sky130_fd_sc_hd__clkbuf_1
X_5690_ disp_song.um.boton2e.edge_2 disp_song.um.boton2e.edge_1 VGND VGND VPWR VPWR
+ _2650_ sky130_fd_sc_hd__and2b_1
XTAP_1291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4641_ _1791_ _1452_ VGND VGND VPWR VPWR _1814_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4572_ _1764_ VGND VGND VPWR VPWR game.scoring_button_1.next_num_misses\[11\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3523_ _0686_ _0885_ VGND VGND VPWR VPWR _0886_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_52_493 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3454_ _0692_ _0683_ _0816_ _0680_ VGND VGND VPWR VPWR _0817_ sky130_fd_sc_hd__a22oi_2
XFILLER_0_110_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3385_ _0730_ _0747_ VGND VGND VPWR VPWR _0748_ sky130_fd_sc_hd__xor2_1
X_6173_ clknet_leaf_45_clk disp_song.um.drum.next_d1\[5\] net54 VGND VGND VPWR VPWR
+ disp_song.display_note1\[5\] sky130_fd_sc_hd__dfrtp_1
X_5124_ _2185_ _2211_ VGND VGND VPWR VPWR _2212_ sky130_fd_sc_hd__or2_1
X_5055_ _1983_ _2142_ _2143_ _2145_ VGND VGND VPWR VPWR _2146_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_49_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_49_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_27_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4006_ game.addmisses.add1.b\[3\] _1315_ VGND VGND VPWR VPWR _1319_ sky130_fd_sc_hd__and2_2
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5957_ clknet_leaf_34_clk game.scoring_button_1.next_flash_counter_2\[2\] net72 VGND
+ VGND VPWR VPWR game.scoring_button_1.flash_counter_2\[2\] sky130_fd_sc_hd__dfrtp_1
X_4908_ disp_song.um.drum.next_note2\[6\] disp_song.um.drum.next_note2\[7\] disp_song.um.drum.next_idx2\[0\]
+ VGND VGND VPWR VPWR _2003_ sky130_fd_sc_hd__mux2_1
X_5888_ clknet_leaf_30_clk _0071_ net69 VGND VGND VPWR VPWR game.padded_notes2\[21\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_7_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4839_ _0032_ _1471_ VGND VGND VPWR VPWR _1942_ sky130_fd_sc_hd__and2b_1
XFILLER_0_31_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold31 game.scoring_button_2.next_flash_counter_1\[1\] VGND VGND VPWR VPWR net104
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold20 game.out\[6\] VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 game.out\[4\] VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 game.flash_counter\[17\] VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 game.flash_counter\[11\] VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 disp_song.um.boton1e.edge_2 VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__buf_1
Xhold97 game.scoring_button_1.hit VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 game.scoring_button_2.flash_counter_2\[13\] VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_6 net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3170_ game.addhits.a\[9\] game.addhits.add3.b\[1\] VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__or2_1
XFILLER_0_88_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5811_ clknet_leaf_47_clk game.scoring_button_2.next_flash_counter_2\[2\] net56 VGND
+ VGND VPWR VPWR game.scoring_button_2.flash_counter_2\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5742_ clknet_leaf_69_clk game.scoring_button_2.next_num_misses\[14\] net46 VGND
+ VGND VPWR VPWR game.addmisses.add4.b\[2\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_84_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2954_ _2661_ _0183_ _0265_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__or3_1
XFILLER_0_8_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2885_ _0302_ VGND VGND VPWR VPWR disp_song.um.drum.next_note2\[10\] sky130_fd_sc_hd__buf_1
XFILLER_0_72_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5673_ game.flash_counter\[19\] _2636_ VGND VGND VPWR VPWR _2638_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4624_ _1805_ VGND VGND VPWR VPWR game.scoring_button_1.next_count\[5\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_600 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4555_ _1747_ _1748_ _1749_ VGND VGND VPWR VPWR _1750_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_52_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3506_ game.flash_counter\[1\] game.flash_counter\[0\] game.flash_counter\[5\] VGND
+ VGND VPWR VPWR _0869_ sky130_fd_sc_hd__and3_1
XFILLER_0_40_441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4486_ _1688_ _1689_ VGND VGND VPWR VPWR _1690_ sky130_fd_sc_hd__or2_1
XFILLER_0_40_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3437_ _0694_ _0799_ VGND VGND VPWR VPWR _0800_ sky130_fd_sc_hd__and2_1
X_6156_ clknet_3_5__leaf_clk disp_song.um.boton1e.edge_1 net63 VGND VGND VPWR VPWR
+ disp_song.um.boton1e.edge_2 sky130_fd_sc_hd__dfrtp_1
X_3368_ _0728_ _0729_ _0726_ VGND VGND VPWR VPWR _0731_ sky130_fd_sc_hd__o21a_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5107_ _0185_ _2194_ VGND VGND VPWR VPWR _2195_ sky130_fd_sc_hd__nand2_4
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6087_ clknet_leaf_43_clk disp_song.um.next_position\[4\] net65 VGND VGND VPWR VPWR
+ disp_song.mi6.in\[4\] sky130_fd_sc_hd__dfstp_1
X_3299_ _0646_ _0655_ VGND VGND VPWR VPWR _0662_ sky130_fd_sc_hd__xnor2_1
X_5038_ _2020_ _2123_ _2128_ _2129_ VGND VGND VPWR VPWR _2130_ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput10 net10 VGND VGND VPWR VPWR bottom_row[3] sky130_fd_sc_hd__clkbuf_4
Xoutput32 net32 VGND VGND VPWR VPWR top_row[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput21 net21 VGND VGND VPWR VPWR ss0[5] sky130_fd_sc_hd__clkbuf_4
Xoutput8 net8 VGND VGND VPWR VPWR bottom_row[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4340_ net192 _1572_ _1575_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_1\[7\]
+ sky130_fd_sc_hd__o21a_1
X_4271_ game.scoring_button_2.flash_counter_2\[9\] _1525_ VGND VGND VPWR VPWR _1528_
+ sky130_fd_sc_hd__and2_1
X_3222_ _0579_ _0584_ VGND VGND VPWR VPWR _0585_ sky130_fd_sc_hd__nor2_1
X_6010_ clknet_leaf_48_clk _0119_ net56 VGND VGND VPWR VPWR game.padded_notes1\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_3153_ _0508_ _0510_ _0509_ VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_89_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3084_ game.addmisses.a\[4\] game.addmisses.add2.b\[0\] VGND VGND VPWR VPWR _0447_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_76_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3986_ game.scoring_button_2.counts\[22\] _1300_ VGND VGND VPWR VPWR _1301_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2937_ _0269_ _0271_ _0334_ _0338_ VGND VGND VPWR VPWR disp_song.um.drum.next_note2\[25\]
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5725_ clknet_leaf_4_clk _0000_ net49 VGND VGND VPWR VPWR lvls.level\[0\] sky130_fd_sc_hd__dfstp_2
XFILLER_0_94_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5656_ _2626_ VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__clkbuf_1
X_2868_ _0269_ disp_song.note2\[6\] _0289_ VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4607_ game.scoring_button_1.flash_counter_1\[8\] game.scoring_button_1.flash_counter_1\[11\]
+ game.scoring_button_1.flash_counter_1\[10\] game.scoring_button_1.flash_counter_1\[9\]
+ VGND VGND VPWR VPWR _1795_ sky130_fd_sc_hd__or4b_1
X_2799_ game.counter\[10\] _0227_ VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__xor2_1
X_5587_ _2583_ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__clkbuf_1
X_4538_ game.addmisses.a\[6\] game.addmisses.a\[5\] _1713_ game.addmisses.a\[7\] VGND
+ VGND VPWR VPWR _1735_ sky130_fd_sc_hd__a31o_1
X_4469_ game.scoring_button_1.check_hit.edge_1 game.scoring_button_1.check_hit.edge_2
+ VGND VGND VPWR VPWR _1673_ sky130_fd_sc_hd__or2b_2
XFILLER_0_68_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6139_ clknet_leaf_28_clk disp_song.um.drum.next_note2\[19\] net68 VGND VGND VPWR
+ VPWR disp_song.note2\[19\] sky130_fd_sc_hd__dfstp_1
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3840_ _1076_ _1185_ _1188_ _1189_ _0935_ VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__o41a_2
XFILLER_0_104_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3771_ _1047_ _1096_ VGND VGND VPWR VPWR _1125_ sky130_fd_sc_hd__and2b_1
X_5510_ _2531_ net232 _2515_ VGND VGND VPWR VPWR _2532_ sky130_fd_sc_hd__mux2_1
X_2722_ _2662_ _0166_ _0167_ _2654_ VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__o211a_1
XFILLER_0_6_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5441_ _2490_ VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_81_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5372_ _2444_ highest_score.highest_score\[5\] _2434_ VGND VGND VPWR VPWR _2445_
+ sky130_fd_sc_hd__mux2_1
X_4323_ _1562_ game.hit_2 _1563_ VGND VGND VPWR VPWR _1564_ sky130_fd_sc_hd__and3b_1
X_4254_ _1516_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_2\[3\]
+ sky130_fd_sc_hd__clkbuf_1
X_4185_ game.counter\[17\] _1457_ VGND VGND VPWR VPWR _1460_ sky130_fd_sc_hd__nor2_1
X_3205_ _0566_ _0567_ VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__xor2_1
X_3136_ _0494_ _0497_ _0495_ VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__o21ai_1
X_3067_ _0398_ _0419_ _0432_ net165 VGND VGND VPWR VPWR disp_song.um.drum.next_note1\[29\]
+ sky130_fd_sc_hd__a22o_1
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5708_ clknet_leaf_43_clk net80 net65 VGND VGND VPWR VPWR modetrans.u3.Q2 sky130_fd_sc_hd__dfrtp_1
X_3969_ game.addhits.add4.b\[3\] _1278_ _1282_ VGND VGND VPWR VPWR _1285_ sky130_fd_sc_hd__a21oi_1
X_5639_ net129 game.flash_counter\[8\] _2612_ _2613_ net37 VGND VGND VPWR VPWR _0138_
+ sky130_fd_sc_hd__a311oi_1
XFILLER_0_103_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold161 game.padded_notes2\[30\] VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__dlygate4sd3_1
Xhold150 game.padded_notes1\[29\] VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 game.padded_notes1\[5\] VGND VGND VPWR VPWR net256 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 disp_song.note1\[21\] VGND VGND VPWR VPWR net245 sky130_fd_sc_hd__dlygate4sd3_1
Xhold194 game.addhits.a\[4\] VGND VGND VPWR VPWR net267 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5990_ clknet_leaf_33_clk _0099_ net71 VGND VGND VPWR VPWR game.padded_notes1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_4941_ _2666_ _2669_ VGND VGND VPWR VPWR _2035_ sky130_fd_sc_hd__nor2_2
X_4872_ disp_song.um.drum.next_idx2\[2\] _1949_ VGND VGND VPWR VPWR _1967_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3823_ disp_song.mi6.in\[3\] _1116_ _1080_ _1114_ _0925_ VGND VGND VPWR VPWR _1174_
+ sky130_fd_sc_hd__o221a_1
X_3754_ _1106_ _1108_ _0925_ VGND VGND VPWR VPWR _1109_ sky130_fd_sc_hd__a21bo_1
X_2705_ _2671_ _2675_ _2676_ VGND VGND VPWR VPWR _2677_ sky130_fd_sc_hd__mux2_2
X_3685_ _0625_ _0880_ net44 VGND VGND VPWR VPWR _1041_ sky130_fd_sc_hd__o21ai_1
X_5424_ disp_song.note2\[8\] game.padded_notes2\[7\] _0219_ VGND VGND VPWR VPWR _2479_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5355_ net42 _2428_ _2432_ VGND VGND VPWR VPWR _2433_ sky130_fd_sc_hd__or3b_1
X_5286_ _2368_ _2369_ _2365_ VGND VGND VPWR VPWR _2370_ sky130_fd_sc_hd__mux2_1
X_4306_ net169 _1549_ _1552_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_2\[19\]
+ sky130_fd_sc_hd__o21a_1
X_4237_ game.counter\[9\] _0245_ _1503_ _0236_ VGND VGND VPWR VPWR _1504_ sky130_fd_sc_hd__a211oi_1
X_4168_ _1443_ _1446_ _1447_ VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__o21a_1
XFILLER_0_65_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4099_ _1396_ _1399_ net45 VGND VGND VPWR VPWR _1400_ sky130_fd_sc_hd__mux2_1
X_3119_ _0480_ _0481_ VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_28 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3470_ _0775_ _0831_ _0832_ VGND VGND VPWR VPWR _0833_ sky130_fd_sc_hd__or3_1
XFILLER_0_86_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5140_ disp_song.um.drum.next_note1\[16\] disp_song.um.drum.next_note1\[17\] disp_song.um.drum.next_idx1\[0\]
+ VGND VGND VPWR VPWR _2228_ sky130_fd_sc_hd__mux2_1
X_5071_ _2026_ _2111_ _2031_ _2034_ VGND VGND VPWR VPWR _2161_ sky130_fd_sc_hd__o211a_1
X_4022_ game.addmisses.add2.b\[0\] _1331_ _1332_ VGND VGND VPWR VPWR _1333_ sky130_fd_sc_hd__a21bo_1
X_5973_ clknet_leaf_31_clk game.scoring_button_1.next_flash_counter_2\[18\] net70
+ VGND VGND VPWR VPWR game.scoring_button_1.flash_counter_2\[18\] sky130_fd_sc_hd__dfrtp_1
X_4924_ _2017_ VGND VGND VPWR VPWR _2018_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4855_ _1948_ _1949_ VGND VGND VPWR VPWR _1950_ sky130_fd_sc_hd__nor2_2
XFILLER_0_74_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3806_ _0926_ _1082_ _0925_ VGND VGND VPWR VPWR _1158_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_34_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4786_ net155 _1908_ _1911_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_1\[13\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_27_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3737_ _0912_ _0636_ VGND VGND VPWR VPWR _1092_ sky130_fd_sc_hd__and2b_1
XFILLER_0_42_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3668_ _0830_ _0834_ _1019_ _1023_ VGND VGND VPWR VPWR _1024_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_30_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5407_ disp_song.note2\[3\] game.padded_notes2\[2\] _0219_ VGND VGND VPWR VPWR _2467_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3599_ _0255_ _0958_ _0959_ _0258_ VGND VGND VPWR VPWR _0960_ sky130_fd_sc_hd__a22o_1
X_5338_ _1012_ _1028_ _1057_ VGND VGND VPWR VPWR _2416_ sky130_fd_sc_hd__o21ai_1
X_5269_ _2268_ _2272_ _2271_ _2254_ VGND VGND VPWR VPWR _2354_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_19_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2970_ _0362_ VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4640_ _1813_ VGND VGND VPWR VPWR game.scoring_button_1.next_count\[13\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4571_ _1755_ _1760_ _1762_ _1763_ _1675_ game.addmisses.a\[11\] VGND VGND VPWR VPWR
+ _1764_ sky130_fd_sc_hd__mux4_1
XFILLER_0_24_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3522_ _0754_ _0884_ _0766_ VGND VGND VPWR VPWR _0885_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_4_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3453_ _0682_ _0815_ VGND VGND VPWR VPWR _0816_ sky130_fd_sc_hd__nand2_1
X_6172_ clknet_leaf_43_clk disp_song.um.drum.next_d1\[4\] net65 VGND VGND VPWR VPWR
+ disp_song.display_note1\[4\] sky130_fd_sc_hd__dfrtp_1
X_5123_ disp_song.um.drum.next_note1\[0\] disp_song.um.drum.next_note1\[1\] _0176_
+ VGND VGND VPWR VPWR _2211_ sky130_fd_sc_hd__mux2_1
X_3384_ _0735_ _0746_ VGND VGND VPWR VPWR _0747_ sky130_fd_sc_hd__and2_1
X_5054_ _2666_ _2076_ _2141_ _2144_ VGND VGND VPWR VPWR _2145_ sky130_fd_sc_hd__a211o_1
XFILLER_0_79_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4005_ _1312_ _1317_ VGND VGND VPWR VPWR _1318_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5956_ clknet_leaf_34_clk net106 net71 VGND VGND VPWR VPWR game.scoring_button_1.flash_counter_2\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5887_ clknet_leaf_30_clk _0070_ net69 VGND VGND VPWR VPWR game.padded_notes2\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_4907_ _1992_ _2000_ _2001_ _2666_ VGND VGND VPWR VPWR _2002_ sky130_fd_sc_hd__a2bb2o_1
X_4838_ _1941_ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_620 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4769_ _1898_ game.hit_1 _1899_ VGND VGND VPWR VPWR _1900_ sky130_fd_sc_hd__and3b_1
XFILLER_0_101_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold32 game.scoring_button_1.flash_counter_2\[1\] VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 disp_song.um.boton0e.edge_1 VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 _0128_ VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 game.out\[0\] VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 _0126_ VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 game.out\[5\] VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__buf_1
Xhold76 disp_song.um.drum.next_note2\[26\] VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__dlygate4sd3_1
Xhold87 disp_song.note1\[31\] VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 game.scoring_button_2.flash_counter_1\[19\] VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5810_ clknet_leaf_47_clk net108 net55 VGND VGND VPWR VPWR game.scoring_button_2.flash_counter_2\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_2953_ _0291_ _0345_ _0348_ net255 VGND VGND VPWR VPWR disp_song.um.drum.next_note2\[31\]
+ sky130_fd_sc_hd__a22o_1
X_5741_ clknet_leaf_69_clk game.scoring_button_2.next_num_misses\[13\] net46 VGND
+ VGND VPWR VPWR game.addmisses.add4.b\[1\] sky130_fd_sc_hd__dfrtp_2
X_2884_ disp_song.note2\[10\] _0269_ _0301_ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__mux2_1
X_5672_ game.flash_counter\[19\] _2636_ VGND VGND VPWR VPWR _2637_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4623_ _1791_ _0027_ VGND VGND VPWR VPWR _1805_ sky130_fd_sc_hd__and2_1
XFILLER_0_72_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4554_ game.addmisses.a\[10\] _1748_ game.addmisses.a\[11\] VGND VGND VPWR VPWR _1749_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_25_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3505_ game.flash_counter\[3\] game.flash_counter\[2\] game.flash_counter\[4\] VGND
+ VGND VPWR VPWR _0868_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4485_ _0209_ _2656_ VGND VGND VPWR VPWR _1689_ sky130_fd_sc_hd__nand2_2
XFILLER_0_0_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3436_ _0597_ _0601_ _0605_ VGND VGND VPWR VPWR _0799_ sky130_fd_sc_hd__o21ai_1
X_6155_ clknet_leaf_13_clk net2 net58 VGND VGND VPWR VPWR disp_song.um.boton1e.sync_b
+ sky130_fd_sc_hd__dfrtp_1
X_3367_ _0728_ _0729_ VGND VGND VPWR VPWR _0730_ sky130_fd_sc_hd__xnor2_2
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5106_ _0197_ _2187_ VGND VGND VPWR VPWR _2194_ sky130_fd_sc_hd__and2_1
X_6086_ clknet_leaf_23_clk disp_song.um.next_position\[3\] net65 VGND VGND VPWR VPWR
+ disp_song.mi6.in\[3\] sky130_fd_sc_hd__dfstp_4
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5037_ _2107_ _2117_ VGND VGND VPWR VPWR _2129_ sky130_fd_sc_hd__nor2_1
X_3298_ _0640_ _0645_ VGND VGND VPWR VPWR _0661_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_79_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5939_ clknet_leaf_52_clk game.scoring_button_1.next_flash_counter_1\[7\] net55 VGND
+ VGND VPWR VPWR game.scoring_button_1.flash_counter_1\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput22 net22 VGND VGND VPWR VPWR ss0[6] sky130_fd_sc_hd__clkbuf_4
Xoutput9 net9 VGND VGND VPWR VPWR bottom_row[2] sky130_fd_sc_hd__clkbuf_4
Xoutput33 net33 VGND VGND VPWR VPWR top_row[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput11 net11 VGND VGND VPWR VPWR bottom_row[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_109_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4270_ _1527_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_2\[8\]
+ sky130_fd_sc_hd__clkbuf_1
X_3221_ _0580_ _0583_ VGND VGND VPWR VPWR _0584_ sky130_fd_sc_hd__xnor2_1
X_3152_ _0514_ _0512_ VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__nor2_1
X_3083_ _0444_ _0445_ VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__nand2_2
XFILLER_0_77_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3985_ game.scoring_button_2.counts\[20\] game.scoring_button_2.counts\[19\] _1299_
+ game.scoring_button_2.counts\[21\] VGND VGND VPWR VPWR _1300_ sky130_fd_sc_hd__a31o_1
XFILLER_0_9_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2936_ _0270_ _0337_ disp_song.note2\[25\] VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__o21a_1
X_5724_ clknet_leaf_6_clk _0048_ net59 VGND VGND VPWR VPWR pulseout.fin_pulse\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2867_ _0273_ _0288_ VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__nand2_1
X_5655_ _2624_ _2625_ VGND VGND VPWR VPWR _2626_ sky130_fd_sc_hd__and2_1
XFILLER_0_87_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4606_ game.scoring_button_1.flash_counter_1\[13\] game.scoring_button_1.flash_counter_1\[12\]
+ game.scoring_button_1.flash_counter_1\[15\] game.scoring_button_1.flash_counter_1\[14\]
+ VGND VGND VPWR VPWR _1794_ sky130_fd_sc_hd__or4b_1
XFILLER_0_103_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2798_ game.counter\[8\] _0227_ VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__xor2_1
X_5586_ _2582_ game.padded_notes1\[26\] _2472_ VGND VGND VPWR VPWR _2583_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4537_ _1734_ VGND VGND VPWR VPWR game.scoring_button_1.next_num_misses\[6\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4468_ game.addhits.a\[15\] _1613_ _1672_ _1612_ VGND VGND VPWR VPWR game.scoring_button_1.next_num_hits\[15\]
+ sky130_fd_sc_hd__a22o_1
X_3419_ _0673_ _0665_ _0672_ VGND VGND VPWR VPWR _0782_ sky130_fd_sc_hd__and3_1
X_6138_ clknet_leaf_29_clk disp_song.um.drum.next_note2\[18\] net69 VGND VGND VPWR
+ VPWR disp_song.note2\[18\] sky130_fd_sc_hd__dfrtp_1
X_4399_ game.addhits.a\[0\] _1616_ _1617_ VGND VGND VPWR VPWR _1618_ sky130_fd_sc_hd__a21boi_1
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6069_ clknet_leaf_62_clk highest_score.nxt_mode\[0\] net54 VGND VGND VPWR VPWR highest_score.score_mode\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_67_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_480 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3770_ _0895_ _1123_ _0255_ VGND VGND VPWR VPWR _1124_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_109_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2721_ disp_song.um.idx_note2\[2\] _2662_ VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__nand2_1
X_5440_ _2489_ game.padded_notes2\[13\] _2473_ VGND VGND VPWR VPWR _2490_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5371_ _2443_ VGND VGND VPWR VPWR _2444_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4322_ game.scoring_button_2.flash_counter_1\[1\] game.scoring_button_2.flash_counter_1\[0\]
+ game.scoring_button_2.flash_counter_1\[2\] VGND VGND VPWR VPWR _1563_ sky130_fd_sc_hd__a21o_1
XFILLER_0_22_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4253_ _1514_ game.missed_2 _1515_ VGND VGND VPWR VPWR _1516_ sky130_fd_sc_hd__and3b_1
X_3204_ _0540_ _0562_ _0538_ VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__o21a_1
X_4184_ _1459_ VGND VGND VPWR VPWR game.scoring_button_2.next_count\[16\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3135_ _0496_ _0497_ VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__xor2_2
X_3066_ _0398_ _0421_ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_72 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3968_ _1226_ _1283_ _1284_ _1227_ net213 VGND VGND VPWR VPWR game.scoring_button_2.next_num_hits\[14\]
+ sky130_fd_sc_hd__a32o_1
X_2919_ _0325_ VGND VGND VPWR VPWR disp_song.next_red sky130_fd_sc_hd__inv_2
X_5707_ clknet_leaf_23_clk net77 net65 VGND VGND VPWR VPWR modetrans.u3.Q1 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3899_ game.addhits.add1.b\[2\] game.scoring_button_2.acc\[2\] VGND VGND VPWR VPWR
+ _1229_ sky130_fd_sc_hd__nor2_1
X_5638_ game.flash_counter\[8\] _2612_ game.flash_counter\[9\] VGND VGND VPWR VPWR
+ _2613_ sky130_fd_sc_hd__a21oi_1
X_5569_ _2571_ VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__clkbuf_1
Xhold162 game.padded_notes2\[12\] VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 game.padded_notes1\[8\] VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__dlygate4sd3_1
Xhold140 game.addhits.add4.b\[2\] VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 disp_song.note1\[13\] VGND VGND VPWR VPWR net246 sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 disp_song.note1\[7\] VGND VGND VPWR VPWR net268 sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 game.addhits.a\[6\] VGND VGND VPWR VPWR net257 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4940_ _2010_ _2012_ VGND VGND VPWR VPWR _2034_ sky130_fd_sc_hd__nor2_2
XFILLER_0_59_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4871_ disp_song.um.drum.next_note2\[18\] disp_song.um.drum.next_note2\[19\] disp_song.um.drum.next_idx2\[0\]
+ VGND VGND VPWR VPWR _1966_ sky130_fd_sc_hd__mux2_2
XFILLER_0_24_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3822_ _1161_ _1037_ _1162_ _1172_ net38 VGND VGND VPWR VPWR _1173_ sky130_fd_sc_hd__o311a_1
XFILLER_0_74_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3753_ disp_song.mi6.in\[3\] disp_song.mi6.in\[2\] _1107_ VGND VGND VPWR VPWR _1108_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_40_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2704_ _2657_ _2660_ _2661_ VGND VGND VPWR VPWR _2676_ sky130_fd_sc_hd__o21a_1
XFILLER_0_70_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3684_ _0625_ _0649_ net44 VGND VGND VPWR VPWR _1040_ sky130_fd_sc_hd__and3_1
XFILLER_0_54_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5423_ _2478_ VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5354_ _2429_ _2430_ _2431_ _0921_ _2423_ VGND VGND VPWR VPWR _2432_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_10_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4305_ net169 _1549_ _1486_ VGND VGND VPWR VPWR _1552_ sky130_fd_sc_hd__a21boi_1
X_5285_ _0191_ _2316_ _2237_ VGND VGND VPWR VPWR _2369_ sky130_fd_sc_hd__o21ba_1
X_4236_ game.counter\[21\] _0241_ _0243_ game.counter\[14\] VGND VGND VPWR VPWR _1503_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4167_ game.counter\[11\] game.counter\[12\] _1439_ game.counter\[13\] VGND VGND
+ VPWR VPWR _1447_ sky130_fd_sc_hd__a31o_1
XFILLER_0_4_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3118_ _0472_ _0473_ _0474_ VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__o21a_1
X_4098_ game.addmisses.add4.b\[3\] _1397_ _1398_ VGND VGND VPWR VPWR _1399_ sky130_fd_sc_hd__mux2_1
X_3049_ _0381_ _0421_ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5070_ _2041_ _2159_ _2034_ VGND VGND VPWR VPWR _2160_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4021_ game.addmisses.add2.b\[0\] _1305_ _1319_ VGND VGND VPWR VPWR _1332_ sky130_fd_sc_hd__or3b_1
X_5972_ clknet_leaf_31_clk game.scoring_button_1.next_flash_counter_2\[17\] net72
+ VGND VGND VPWR VPWR game.scoring_button_1.flash_counter_2\[17\] sky130_fd_sc_hd__dfrtp_1
X_4923_ _1956_ disp_song.um.drum.next_note2\[31\] _1965_ _2016_ disp_song.um.drum.next_note2\[30\]
+ VGND VGND VPWR VPWR _2017_ sky130_fd_sc_hd__a32o_1
X_4854_ _2677_ _0162_ VGND VGND VPWR VPWR _1949_ sky130_fd_sc_hd__nand2_4
XFILLER_0_62_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4785_ net155 _1908_ game.hit_1 VGND VGND VPWR VPWR _1911_ sky130_fd_sc_hd__a21boi_1
X_3805_ _0259_ _1154_ VGND VGND VPWR VPWR _1157_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3736_ _0806_ _1025_ _1035_ VGND VGND VPWR VPWR _1091_ sky130_fd_sc_hd__and3_1
X_3667_ _0762_ _0824_ _0825_ _0826_ _0786_ VGND VGND VPWR VPWR _1023_ sky130_fd_sc_hd__o311a_1
XFILLER_0_30_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5406_ _2466_ VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__clkbuf_1
X_3598_ _0939_ _0675_ _0889_ VGND VGND VPWR VPWR _0959_ sky130_fd_sc_hd__and3b_1
XFILLER_0_11_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5337_ _1028_ _1029_ _1030_ highest_score.highest_score\[1\] VGND VGND VPWR VPWR
+ _2415_ sky130_fd_sc_hd__o31a_1
X_5268_ _2267_ _2269_ _2256_ VGND VGND VPWR VPWR _2353_ sky130_fd_sc_hd__mux2_1
X_4219_ _1405_ _1303_ _1486_ VGND VGND VPWR VPWR game.scoring_button_2.next_missed
+ sky130_fd_sc_hd__o21bai_1
X_5199_ _2283_ _2285_ _2254_ VGND VGND VPWR VPWR _2286_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4570_ _1744_ _1760_ VGND VGND VPWR VPWR _1763_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3521_ _0748_ _0594_ _0704_ _0883_ VGND VGND VPWR VPWR _0884_ sky130_fd_sc_hd__or4_1
XFILLER_0_24_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3452_ _0693_ VGND VGND VPWR VPWR _0815_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6171_ clknet_leaf_43_clk disp_song.um.drum.next_d1\[3\] net65 VGND VGND VPWR VPWR
+ disp_song.display_note1\[3\] sky130_fd_sc_hd__dfrtp_1
X_3383_ _0739_ _0745_ _0743_ VGND VGND VPWR VPWR _0746_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_110_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5122_ disp_song.note1\[2\] _2209_ disp_song.um.drum.next_idx1\[0\] VGND VGND VPWR
+ VPWR _2210_ sky130_fd_sc_hd__mux2_1
X_5053_ _2666_ _1973_ VGND VGND VPWR VPWR _2144_ sky130_fd_sc_hd__nor2_1
X_4004_ _1315_ _1316_ VGND VGND VPWR VPWR _1317_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5955_ clknet_leaf_33_clk game.scoring_button_1.next_flash_counter_2\[0\] net71 VGND
+ VGND VPWR VPWR game.scoring_button_1.flash_counter_2\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_87_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5886_ clknet_leaf_30_clk _0069_ net69 VGND VGND VPWR VPWR game.padded_notes2\[19\]
+ sky130_fd_sc_hd__dfstp_1
X_4906_ disp_song.um.drum.next_note2\[2\] disp_song.um.drum.next_note2\[3\] _2670_
+ VGND VGND VPWR VPWR _2001_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4837_ _0032_ _1467_ VGND VGND VPWR VPWR _1941_ sky130_fd_sc_hd__and2b_1
XFILLER_0_16_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4768_ game.scoring_button_1.flash_counter_1\[7\] game.scoring_button_1.flash_counter_1\[6\]
+ _1891_ game.scoring_button_1.flash_counter_1\[8\] VGND VGND VPWR VPWR _1899_ sky130_fd_sc_hd__a31o_1
X_4699_ _1850_ _1830_ _1851_ VGND VGND VPWR VPWR _1852_ sky130_fd_sc_hd__and3b_1
X_3719_ _1032_ _1037_ _1039_ _1074_ net38 VGND VGND VPWR VPWR _1075_ sky130_fd_sc_hd__o311a_1
XFILLER_0_101_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold22 game.scoring_button_1.check_hit.in VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 game.scoring_button_2.check_hit.edge_1 VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 game.scoring_button_1.next_flash_counter_2\[1\] VGND VGND VPWR VPWR net106
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 pulseout.fin_pulse\[2\] VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 game.out\[11\] VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 game.scoring_button_1.flash_counter_2\[7\] VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 disp_song.note1\[25\] VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 _0122_ VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__dlygate4sd3_1
Xhold99 game.scoring_button_1.flash_counter_1\[19\] VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2952_ _0313_ _0337_ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5740_ clknet_leaf_70_clk game.scoring_button_2.next_num_misses\[12\] net46 VGND
+ VGND VPWR VPWR game.addmisses.add4.b\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_84_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2883_ _0276_ _0298_ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__nor2_1
X_5671_ net264 _2636_ VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__nor2_1
X_4622_ _1804_ VGND VGND VPWR VPWR game.scoring_button_1.next_count\[4\] sky130_fd_sc_hd__clkbuf_1
X_4553_ game.addmisses.a\[9\] _1741_ VGND VGND VPWR VPWR _1748_ sky130_fd_sc_hd__or2_1
XFILLER_0_40_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4484_ _1676_ _1678_ _1682_ _1687_ VGND VGND VPWR VPWR _1688_ sky130_fd_sc_hd__o31a_1
X_3504_ game.flash_counter\[20\] _0866_ game.flash_counter\[22\] VGND VGND VPWR VPWR
+ _0867_ sky130_fd_sc_hd__o21a_1
XFILLER_0_4_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3435_ _0797_ _0723_ VGND VGND VPWR VPWR _0798_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6154_ clknet_leaf_31_clk net79 net70 VGND VGND VPWR VPWR disp_song.um.boton0e.edge_1
+ sky130_fd_sc_hd__dfrtp_1
X_3366_ _0531_ _0593_ _0529_ VGND VGND VPWR VPWR _0729_ sky130_fd_sc_hd__a21oi_2
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6085_ clknet_leaf_43_clk disp_song.um.next_position\[2\] net65 VGND VGND VPWR VPWR
+ disp_song.mi6.in\[2\] sky130_fd_sc_hd__dfstp_2
X_5105_ _2191_ _2192_ disp_song.um.drum.next_idx1\[2\] VGND VGND VPWR VPWR _2193_
+ sky130_fd_sc_hd__a21oi_1
X_3297_ _0632_ _0657_ VGND VGND VPWR VPWR _0660_ sky130_fd_sc_hd__xnor2_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5036_ _2100_ _2124_ _2125_ _2127_ _2026_ VGND VGND VPWR VPWR _2128_ sky130_fd_sc_hd__a221o_1
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5938_ clknet_leaf_56_clk game.scoring_button_1.next_flash_counter_1\[6\] net73 VGND
+ VGND VPWR VPWR game.scoring_button_1.flash_counter_1\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5869_ clknet_leaf_22_clk _0052_ net59 VGND VGND VPWR VPWR game.padded_notes2\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput12 net12 VGND VGND VPWR VPWR bottom_row[5] sky130_fd_sc_hd__clkbuf_4
Xoutput23 net23 VGND VGND VPWR VPWR ss1[0] sky130_fd_sc_hd__buf_2
XFILLER_0_31_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput34 net34 VGND VGND VPWR VPWR top_row[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_598 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3220_ _0581_ _0582_ VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__and2b_1
X_3151_ _0505_ _0513_ VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__xnor2_2
X_3082_ game.addmisses.a\[5\] game.addmisses.add2.b\[1\] VGND VGND VPWR VPWR _0445_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_77_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_74 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3984_ game.scoring_button_2.counts\[17\] game.scoring_button_2.counts\[16\] game.scoring_button_2.counts\[15\]
+ _1298_ game.scoring_button_2.counts\[18\] VGND VGND VPWR VPWR _1299_ sky130_fd_sc_hd__a41o_1
X_2935_ _2658_ _0336_ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__or2_2
X_5723_ clknet_leaf_6_clk _0047_ net59 VGND VGND VPWR VPWR pulseout.fin_pulse\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_524 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2866_ disp_song.um.idx_note2\[0\] disp_song.um.idx_note2\[2\] disp_song.um.idx_note2\[1\]
+ VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__and3b_1
X_5654_ game.flash_counter\[13\] _2623_ VGND VGND VPWR VPWR _2625_ sky130_fd_sc_hd__or2_1
X_4605_ game.scoring_button_1.flash_counter_1\[1\] game.scoring_button_1.flash_counter_1\[0\]
+ game.scoring_button_1.flash_counter_1\[3\] game.scoring_button_1.flash_counter_1\[2\]
+ VGND VGND VPWR VPWR _1793_ sky130_fd_sc_hd__or4_1
XFILLER_0_103_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2797_ game.counter\[11\] _0227_ VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__xor2_1
X_5585_ disp_song.note1\[26\] game.padded_notes1\[25\] _0209_ VGND VGND VPWR VPWR
+ _2582_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4536_ _1729_ _1733_ _1675_ VGND VGND VPWR VPWR _1734_ sky130_fd_sc_hd__mux2_1
XFILLER_0_40_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4467_ _1669_ _1671_ VGND VGND VPWR VPWR _1672_ sky130_fd_sc_hd__nor2_1
X_3418_ _0683_ _0780_ _0691_ VGND VGND VPWR VPWR _0781_ sky130_fd_sc_hd__mux2_2
X_4398_ game.addhits.a\[1\] game.scoring_button_1.acc\[1\] VGND VGND VPWR VPWR _1617_
+ sky130_fd_sc_hd__nand2_1
X_6137_ clknet_leaf_28_clk disp_song.um.drum.next_note2\[17\] net68 VGND VGND VPWR
+ VPWR disp_song.note2\[17\] sky130_fd_sc_hd__dfstp_1
X_3349_ _0708_ VGND VGND VPWR VPWR _0712_ sky130_fd_sc_hd__inv_2
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6068_ clknet_leaf_25_clk _0153_ net64 VGND VGND VPWR VPWR disp_song.toggle_state
+ sky130_fd_sc_hd__dfrtp_1
X_5019_ _1968_ _2035_ _2023_ _2024_ VGND VGND VPWR VPWR _2111_ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2720_ _0164_ _0165_ VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__or2_2
XFILLER_0_89_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_77 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5370_ _0830_ _0791_ _0857_ _2442_ VGND VGND VPWR VPWR _2443_ sky130_fd_sc_hd__a211o_1
X_4321_ game.scoring_button_2.flash_counter_1\[1\] game.scoring_button_2.flash_counter_1\[0\]
+ game.scoring_button_2.flash_counter_1\[2\] VGND VGND VPWR VPWR _1562_ sky130_fd_sc_hd__and3_1
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4252_ game.scoring_button_2.flash_counter_2\[3\] _1511_ VGND VGND VPWR VPWR _1515_
+ sky130_fd_sc_hd__or2_1
X_3203_ _0564_ _0565_ VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__or2b_1
XFILLER_0_38_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4183_ _1405_ _1458_ VGND VGND VPWR VPWR _1459_ sky130_fd_sc_hd__and2_1
X_3134_ _0488_ _0489_ _0490_ VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__o21a_1
X_3065_ _0374_ _0425_ _0431_ VGND VGND VPWR VPWR disp_song.um.drum.next_note1\[28\]
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_77_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3967_ _1279_ _1282_ VGND VGND VPWR VPWR _1284_ sky130_fd_sc_hd__or2_1
X_2918_ _0160_ _0325_ VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__nor2_1
XFILLER_0_57_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5706_ clknet_leaf_60_clk _0042_ net51 VGND VGND VPWR VPWR highest_score.highest_score\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_30_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_30_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_60_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3898_ _1228_ VGND VGND VPWR VPWR game.scoring_button_2.next_num_hits\[0\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_415 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2849_ _0275_ VGND VGND VPWR VPWR disp_song.um.drum.next_note2\[1\] sky130_fd_sc_hd__buf_1
XFILLER_0_60_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5637_ net187 _2612_ VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__xor2_1
X_5568_ _2570_ net222 _2472_ VGND VGND VPWR VPWR _2571_ sky130_fd_sc_hd__mux2_1
Xhold141 game.padded_notes1\[9\] VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__dlygate4sd3_1
Xhold152 game.padded_notes1\[21\] VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__dlygate4sd3_1
X_4519_ game.addmisses.a\[4\] _1717_ _1718_ VGND VGND VPWR VPWR _1719_ sky130_fd_sc_hd__a21bo_1
Xhold130 game.scoring_button_1.acc\[1\] VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 disp_song.note2\[23\] VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 disp_song.note1\[8\] VGND VGND VPWR VPWR net247 sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 game.addhits.add3.b\[1\] VGND VGND VPWR VPWR net258 sky130_fd_sc_hd__dlygate4sd3_1
X_5499_ net133 _2460_ _2462_ net143 VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__a22o_1
Xhold196 game.out\[12\] VGND VGND VPWR VPWR net269 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_21_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_21_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_63_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4870_ _1964_ VGND VGND VPWR VPWR _1965_ sky130_fd_sc_hd__buf_4
X_3821_ _0879_ _1171_ VGND VGND VPWR VPWR _1172_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_12_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_12_clk sky130_fd_sc_hd__clkbuf_16
X_3752_ _1077_ _0926_ VGND VGND VPWR VPWR _1107_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2703_ _2673_ _2674_ VGND VGND VPWR VPWR _2675_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3683_ _1035_ _1033_ _1038_ VGND VGND VPWR VPWR _1039_ sky130_fd_sc_hd__a21o_1
X_5422_ _2477_ game.padded_notes2\[7\] _2473_ VGND VGND VPWR VPWR _2478_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5353_ _2423_ highest_score.highest_score\[6\] _0835_ _2424_ VGND VGND VPWR VPWR
+ _2431_ sky130_fd_sc_hd__and4b_1
X_4304_ _1551_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_2\[18\]
+ sky130_fd_sc_hd__clkbuf_1
X_5284_ _0191_ _2203_ _2206_ VGND VGND VPWR VPWR _2368_ sky130_fd_sc_hd__o21a_1
XFILLER_0_10_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4235_ game.counter\[17\] game.counter\[18\] game.counter\[20\] _0240_ _1501_ VGND
+ VGND VPWR VPWR _1502_ sky130_fd_sc_hd__o221a_1
X_4166_ game.counter\[13\] game.counter\[12\] VGND VGND VPWR VPWR _1446_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3117_ _0478_ _0479_ VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__or2b_1
X_4097_ game.addmisses.add4.b\[2\] _1385_ VGND VGND VPWR VPWR _1398_ sky130_fd_sc_hd__nand2_1
X_3048_ _0420_ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_77_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4999_ _2090_ _2091_ _0169_ VGND VGND VPWR VPWR _2092_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4020_ _1305_ _1329_ _1330_ VGND VGND VPWR VPWR _1331_ sky130_fd_sc_hd__o21a_1
Xclkbuf_leaf_1_clk clknet_3_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_1_clk sky130_fd_sc_hd__clkbuf_16
X_5971_ clknet_leaf_31_clk net195 net70 VGND VGND VPWR VPWR game.scoring_button_1.flash_counter_2\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4922_ _2669_ _1992_ VGND VGND VPWR VPWR _2016_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4853_ _2666_ _0169_ VGND VGND VPWR VPWR _1948_ sky130_fd_sc_hd__nor2_2
XFILLER_0_74_279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4784_ _1910_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_1\[12\]
+ sky130_fd_sc_hd__clkbuf_1
X_3804_ _1037_ _1120_ _1130_ _1155_ net38 VGND VGND VPWR VPWR _1156_ sky130_fd_sc_hd__o311a_1
XFILLER_0_51_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3735_ net38 VGND VGND VPWR VPWR _1090_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5405_ _2465_ net242 _2462_ VGND VGND VPWR VPWR _2466_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3666_ _0834_ _1015_ _0830_ VGND VGND VPWR VPWR _1022_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_530 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3597_ highest_score.highest_score\[4\] _0906_ _0895_ VGND VGND VPWR VPWR _0958_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5336_ _1021_ _1022_ VGND VGND VPWR VPWR _2414_ sky130_fd_sc_hd__nand2_1
X_5267_ _2348_ _2351_ _2339_ VGND VGND VPWR VPWR _2352_ sky130_fd_sc_hd__mux2_1
X_4218_ _1479_ _1480_ _1485_ game.missed_2 VGND VGND VPWR VPWR _1486_ sky130_fd_sc_hd__o31a_2
X_5198_ _2232_ disp_song.um.drum.next_note1\[14\] _2195_ _2284_ VGND VGND VPWR VPWR
+ _2285_ sky130_fd_sc_hd__o211a_1
X_4149_ game.counter\[8\] _1429_ game.counter\[9\] VGND VGND VPWR VPWR _1434_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_97_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_235 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3520_ _0697_ _0604_ _0882_ _0716_ VGND VGND VPWR VPWR _0883_ sky130_fd_sc_hd__or4b_1
XFILLER_0_21_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3451_ _0781_ _0791_ _0813_ VGND VGND VPWR VPWR _0814_ sky130_fd_sc_hd__or3_2
X_6170_ clknet_leaf_44_clk disp_song.um.drum.next_d1\[2\] net65 VGND VGND VPWR VPWR
+ disp_song.display_note1\[2\] sky130_fd_sc_hd__dfrtp_1
X_3382_ _0734_ _0744_ VGND VGND VPWR VPWR _0745_ sky130_fd_sc_hd__xnor2_1
X_5121_ _0373_ _2208_ VGND VGND VPWR VPWR _2209_ sky130_fd_sc_hd__nor2_1
X_5052_ _1980_ _2141_ _1983_ VGND VGND VPWR VPWR _2143_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4003_ game.addmisses.add1.b\[1\] game.addmisses.add1.b\[0\] game.addmisses.add1.b\[2\]
+ VGND VGND VPWR VPWR _1316_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5954_ clknet_leaf_61_clk game.scoring_button_1.next_flash_counter_1\[22\] net53
+ VGND VGND VPWR VPWR game.scoring_button_1.flash_counter_1\[22\] sky130_fd_sc_hd__dfrtp_1
X_5885_ clknet_leaf_29_clk _0068_ net69 VGND VGND VPWR VPWR game.padded_notes2\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4905_ disp_song.um.drum.next_idx2\[1\] _1999_ VGND VGND VPWR VPWR _2000_ sky130_fd_sc_hd__nand2_1
X_4836_ _1940_ VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4767_ game.scoring_button_1.flash_counter_1\[7\] game.scoring_button_1.flash_counter_1\[8\]
+ _1894_ VGND VGND VPWR VPWR _1898_ sky130_fd_sc_hd__and3_1
XFILLER_0_43_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4698_ game.scoring_button_1.flash_counter_2\[9\] _1847_ VGND VGND VPWR VPWR _1851_
+ sky130_fd_sc_hd__or2_1
X_3718_ _0879_ _1073_ VGND VGND VPWR VPWR _1074_ sky130_fd_sc_hd__nand2_1
XFILLER_0_70_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3649_ _0906_ _0996_ _0258_ VGND VGND VPWR VPWR _1006_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5319_ _0179_ _2232_ disp_song.um.drum.next_note1\[2\] _2208_ _2400_ VGND VGND VPWR
+ VPWR _2401_ sky130_fd_sc_hd__a41o_1
XFILLER_0_11_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold23 game.flash_counter\[4\] VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__dlygate4sd3_1
Xhold12 game.scoring_button_1.flash_counter_1\[22\] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 game.flash_counter\[9\] VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 game.scoring_button_2.flash_counter_2\[1\] VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 _0086_ VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 game.scoring_button_1.flash_counter_1\[7\] VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__dlygate4sd3_1
Xhold78 game.scoring_button_2.flash_counter_2\[7\] VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__dlygate4sd3_1
Xhold67 game.out\[9\] VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2951_ _0288_ _0345_ _0347_ net200 VGND VGND VPWR VPWR disp_song.um.drum.next_note2\[30\]
+ sky130_fd_sc_hd__a22o_1
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_588 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5670_ game.flash_counter\[18\] game.flash_counter\[17\] game.flash_counter\[16\]
+ _2629_ VGND VGND VPWR VPWR _2636_ sky130_fd_sc_hd__and4_1
XFILLER_0_29_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2882_ _0300_ VGND VGND VPWR VPWR disp_song.um.drum.next_note2\[9\] sky130_fd_sc_hd__buf_1
X_4621_ _1791_ _0026_ VGND VGND VPWR VPWR _1804_ sky130_fd_sc_hd__and2_1
XFILLER_0_84_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4552_ game.addmisses.a\[9\] _1741_ VGND VGND VPWR VPWR _1747_ sky130_fd_sc_hd__nand2_1
X_4483_ game.scoring_button_1.counts\[22\] _1686_ VGND VGND VPWR VPWR _1687_ sky130_fd_sc_hd__nand2_1
X_3503_ game.flash_counter\[19\] game.flash_counter\[18\] _0865_ game.flash_counter\[21\]
+ VGND VGND VPWR VPWR _0866_ sky130_fd_sc_hd__a31o_1
XFILLER_0_40_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3434_ _0724_ _0595_ VGND VGND VPWR VPWR _0797_ sky130_fd_sc_hd__or2_1
X_6153_ clknet_leaf_26_clk net83 net70 VGND VGND VPWR VPWR disp_song.um.boton0e.edge_2
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3365_ _0726_ _0727_ VGND VGND VPWR VPWR _0728_ sky130_fd_sc_hd__nand2_1
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6084_ clknet_leaf_23_clk disp_song.um.next_position\[1\] net65 VGND VGND VPWR VPWR
+ disp_song.mi6.in\[1\] sky130_fd_sc_hd__dfstp_1
X_5104_ disp_song.um.drum.next_note1\[12\] disp_song.um.drum.next_note1\[13\] _0176_
+ VGND VGND VPWR VPWR _2192_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3296_ _0625_ _0631_ _0658_ VGND VGND VPWR VPWR _0659_ sky130_fd_sc_hd__o21ai_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5035_ _2126_ _2110_ _2100_ VGND VGND VPWR VPWR _2127_ sky130_fd_sc_hd__a21oi_1
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5937_ clknet_leaf_61_clk game.scoring_button_1.next_flash_counter_1\[5\] net53 VGND
+ VGND VPWR VPWR game.scoring_button_1.flash_counter_1\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5868_ clknet_leaf_22_clk _0051_ net65 VGND VGND VPWR VPWR game.padded_notes2\[1\]
+ sky130_fd_sc_hd__dfstp_1
X_4819_ _1933_ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5799_ clknet_leaf_56_clk game.scoring_button_2.next_flash_counter_1\[13\] net52
+ VGND VGND VPWR VPWR game.scoring_button_2.flash_counter_1\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_422 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput24 net24 VGND VGND VPWR VPWR ss1[1] sky130_fd_sc_hd__clkbuf_4
Xoutput13 net13 VGND VGND VPWR VPWR bottom_row[6] sky130_fd_sc_hd__clkbuf_4
Xoutput35 net35 VGND VGND VPWR VPWR top_row[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_3_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_41_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3150_ _0507_ _0506_ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__or2b_1
X_3081_ game.addmisses.a\[5\] game.addmisses.add2.b\[1\] VGND VGND VPWR VPWR _0444_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_9_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3983_ game.scoring_button_2.counts\[11\] game.scoring_button_2.counts\[10\] _1297_
+ _1290_ VGND VGND VPWR VPWR _1298_ sky130_fd_sc_hd__a31o_1
X_5722_ clknet_leaf_6_clk _0046_ net59 VGND VGND VPWR VPWR pulseout.fin_pulse\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2934_ _2659_ _0335_ VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_536 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2865_ _0287_ VGND VGND VPWR VPWR disp_song.um.drum.next_note2\[5\] sky130_fd_sc_hd__buf_1
XFILLER_0_17_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5653_ game.flash_counter\[13\] _2623_ VGND VGND VPWR VPWR _2624_ sky130_fd_sc_hd__nand2_1
X_5584_ _2581_ VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4604_ game.scoring_button_1.flash_counter_1\[5\] game.scoring_button_1.flash_counter_1\[4\]
+ game.scoring_button_1.flash_counter_1\[7\] game.scoring_button_1.flash_counter_1\[6\]
+ VGND VGND VPWR VPWR _1792_ sky130_fd_sc_hd__or4b_1
X_2796_ _0226_ VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4535_ game.addmisses.a\[6\] _1693_ _1732_ VGND VGND VPWR VPWR _1733_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_111_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4466_ game.addhits.a\[15\] _1664_ _1668_ VGND VGND VPWR VPWR _1671_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3417_ _0692_ _0779_ VGND VGND VPWR VPWR _0780_ sky130_fd_sc_hd__and2_1
X_4397_ game.addhits.a\[1\] game.scoring_button_1.acc\[1\] VGND VGND VPWR VPWR _1616_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_110_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6136_ clknet_leaf_25_clk disp_song.um.drum.next_note2\[16\] net64 VGND VGND VPWR
+ VPWR disp_song.note2\[16\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3348_ _0702_ _0710_ VGND VGND VPWR VPWR _0711_ sky130_fd_sc_hd__or2_2
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6067_ clknet_leaf_7_clk _0032_ net59 VGND VGND VPWR VPWR game.beat_clk sky130_fd_sc_hd__dfrtp_2
X_3279_ _0546_ _0560_ VGND VGND VPWR VPWR _0642_ sky130_fd_sc_hd__xor2_4
X_5018_ _0162_ _2107_ VGND VGND VPWR VPWR _2110_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4320_ net103 game.scoring_button_2.flash_counter_1\[0\] _1561_ VGND VGND VPWR VPWR
+ game.scoring_button_2.next_flash_counter_1\[1\] sky130_fd_sc_hd__a21oi_1
XFILLER_0_10_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4251_ game.scoring_button_2.flash_counter_2\[3\] _1511_ VGND VGND VPWR VPWR _1514_
+ sky130_fd_sc_hd__and2_1
X_3202_ game.addhits.a\[6\] game.addhits.add2.b\[2\] VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__nand2_1
X_4182_ _1456_ _1457_ VGND VGND VPWR VPWR _1458_ sky130_fd_sc_hd__nor2_1
X_3133_ _0494_ _0495_ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__or2b_1
X_3064_ _0374_ _0426_ net122 VGND VGND VPWR VPWR _0431_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_54_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3966_ _0742_ _1282_ _1277_ VGND VGND VPWR VPWR _1283_ sky130_fd_sc_hd__a21oi_1
X_2917_ _2661_ modetrans.mode\[2\] VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__nand2_2
XFILLER_0_73_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5705_ clknet_leaf_60_clk _0041_ net50 VGND VGND VPWR VPWR highest_score.highest_score\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_92_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5636_ _2603_ net37 _2612_ VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__nor3_1
XFILLER_0_33_528 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3897_ _1226_ _1227_ game.addhits.add1.b\[0\] VGND VGND VPWR VPWR _1228_ sky130_fd_sc_hd__mux2_1
X_2848_ _0269_ disp_song.note2\[1\] _0274_ VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5567_ disp_song.note1\[20\] game.padded_notes1\[19\] _2541_ VGND VGND VPWR VPWR
+ _2570_ sky130_fd_sc_hd__mux2_1
X_2779_ modetrans.u2.Q2 modetrans.u2.Q1 VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__and2b_1
Xhold153 game.padded_notes1\[16\] VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__dlygate4sd3_1
Xhold131 disp_song.note1\[23\] VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 game.addhits.a\[13\] VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__dlygate4sd3_1
Xhold120 game.scoring_button_2.next_flash_counter_1\[7\] VGND VGND VPWR VPWR net193
+ sky130_fd_sc_hd__dlygate4sd3_1
X_4518_ game.addmisses.a\[4\] _1691_ _1705_ VGND VGND VPWR VPWR _1718_ sky130_fd_sc_hd__or3b_1
X_5498_ game.padded_notes2\[31\] _2460_ _2462_ net133 VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__a22o_1
Xhold164 disp_song.note1\[15\] VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 disp_song.note1\[24\] VGND VGND VPWR VPWR net259 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4449_ _1655_ game.addhits.a\[11\] _1658_ VGND VGND VPWR VPWR _1659_ sky130_fd_sc_hd__mux2_1
Xhold175 game.addmisses.a\[12\] VGND VGND VPWR VPWR net248 sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 modetrans.mode\[4\] VGND VGND VPWR VPWR net270 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6119_ clknet_leaf_48_clk disp_song.um.drum.next_note1\[31\] net56 VGND VGND VPWR
+ VPWR disp_song.note1\[31\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_95_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_303 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3820_ _1165_ _1168_ _1170_ _0921_ VGND VGND VPWR VPWR _1171_ sky130_fd_sc_hd__a31o_1
XFILLER_0_6_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3751_ _1104_ _1082_ _1105_ VGND VGND VPWR VPWR _1106_ sky130_fd_sc_hd__or3b_1
X_2702_ disp_song.um.idx_note2\[3\] _2672_ VGND VGND VPWR VPWR _2674_ sky130_fd_sc_hd__and2_1
XFILLER_0_70_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3682_ _1025_ _1031_ _1034_ VGND VGND VPWR VPWR _1038_ sky130_fd_sc_hd__and3_1
X_5421_ disp_song.note2\[7\] game.padded_notes2\[6\] _0219_ VGND VGND VPWR VPWR _2477_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5352_ _2426_ _2421_ VGND VGND VPWR VPWR _2430_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4303_ _1549_ _1486_ _1550_ VGND VGND VPWR VPWR _1551_ sky130_fd_sc_hd__and3b_1
X_5283_ _2212_ _2361_ _2363_ _2366_ VGND VGND VPWR VPWR _2367_ sky130_fd_sc_hd__a31o_1
X_4234_ game.counter\[4\] game.counter\[22\] game.counter\[19\] game.counter\[5\]
+ VGND VGND VPWR VPWR _1501_ sky130_fd_sc_hd__and4bb_1
X_4165_ _1445_ VGND VGND VPWR VPWR game.scoring_button_2.next_count\[12\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3116_ game.addmisses.a\[7\] game.addmisses.add2.b\[3\] VGND VGND VPWR VPWR _0479_
+ sky130_fd_sc_hd__nand2_1
X_4096_ game.addmisses.add4.b\[2\] _1385_ _1388_ VGND VGND VPWR VPWR _1397_ sky130_fd_sc_hd__o21a_1
XFILLER_0_77_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3047_ _2654_ _2660_ _0409_ VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__and3_1
XFILLER_0_37_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4998_ _1978_ _1979_ _2666_ VGND VGND VPWR VPWR _2091_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3949_ net258 _1227_ _1270_ _1226_ VGND VGND VPWR VPWR game.scoring_button_2.next_num_hits\[9\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5619_ _2599_ VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout70 net73 VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_24_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5970_ clknet_leaf_31_clk game.scoring_button_1.next_flash_counter_2\[15\] net70
+ VGND VGND VPWR VPWR game.scoring_button_1.flash_counter_2\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4921_ _1968_ _2014_ VGND VGND VPWR VPWR _2015_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_564 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4852_ _1947_ VGND VGND VPWR VPWR disp_song.um.next_position\[4\] sky130_fd_sc_hd__clkbuf_1
X_3803_ _0879_ _1154_ VGND VGND VPWR VPWR _1155_ sky130_fd_sc_hd__nand2_1
X_4783_ _1908_ game.hit_1 _1909_ VGND VGND VPWR VPWR _1910_ sky130_fd_sc_hd__and3b_1
XFILLER_0_15_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3734_ _1075_ _1076_ _1089_ _0935_ VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__o31a_2
XFILLER_0_15_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3665_ _0786_ _1011_ _1019_ _1020_ _0830_ VGND VGND VPWR VPWR _1021_ sky130_fd_sc_hd__a41o_1
XFILLER_0_70_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5404_ disp_song.note2\[2\] game.padded_notes2\[1\] _0219_ VGND VGND VPWR VPWR _2465_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3596_ _0955_ _0956_ VGND VGND VPWR VPWR _0957_ sky130_fd_sc_hd__or2_1
X_5335_ _2413_ VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5266_ _2254_ _2336_ _2349_ _2350_ VGND VGND VPWR VPWR _2351_ sky130_fd_sc_hd__a31o_1
XFILLER_0_55_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4217_ _1481_ _1482_ _1483_ _1484_ VGND VGND VPWR VPWR _1485_ sky130_fd_sc_hd__or4b_1
X_5197_ _0176_ disp_song.um.drum.next_note1\[15\] VGND VGND VPWR VPWR _2284_ sky130_fd_sc_hd__or2_1
X_4148_ _1433_ VGND VGND VPWR VPWR game.scoring_button_2.next_count\[8\] sky130_fd_sc_hd__clkbuf_1
X_4079_ game.addmisses.add4.b\[0\] _1381_ VGND VGND VPWR VPWR _1382_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3450_ _0808_ _0812_ VGND VGND VPWR VPWR _0813_ sky130_fd_sc_hd__or2_1
X_3381_ _0740_ _0743_ VGND VGND VPWR VPWR _0744_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5120_ _2207_ VGND VGND VPWR VPWR _2208_ sky130_fd_sc_hd__clkbuf_2
X_5051_ _1959_ _2140_ _2141_ VGND VGND VPWR VPWR _2142_ sky130_fd_sc_hd__mux2_1
X_4002_ game.addmisses.add1.b\[2\] game.addmisses.add1.b\[1\] game.addmisses.add1.b\[0\]
+ VGND VGND VPWR VPWR _1315_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_79_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5953_ clknet_leaf_45_clk game.scoring_button_1.next_flash_counter_1\[21\] net53
+ VGND VGND VPWR VPWR game.scoring_button_1.flash_counter_1\[21\] sky130_fd_sc_hd__dfrtp_1
X_5884_ clknet_leaf_29_clk _0067_ net69 VGND VGND VPWR VPWR game.padded_notes2\[17\]
+ sky130_fd_sc_hd__dfstp_1
X_4904_ disp_song.um.drum.next_note2\[0\] disp_song.um.drum.next_note2\[1\] _2670_
+ VGND VGND VPWR VPWR _1999_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4835_ _0032_ _1463_ VGND VGND VPWR VPWR _1940_ sky130_fd_sc_hd__and2b_1
XFILLER_0_28_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4766_ net162 _1894_ _1897_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_1\[7\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_7_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3717_ _1051_ _1063_ _1072_ _0921_ VGND VGND VPWR VPWR _1073_ sky130_fd_sc_hd__a31o_1
X_4697_ game.scoring_button_1.flash_counter_2\[9\] _1847_ VGND VGND VPWR VPWR _1850_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_31_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_637 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3648_ _0918_ _0992_ _0261_ VGND VGND VPWR VPWR _1005_ sky130_fd_sc_hd__o21ai_1
X_3579_ _0255_ _0895_ VGND VGND VPWR VPWR _0941_ sky130_fd_sc_hd__nor2_2
X_5318_ disp_song.um.drum.next_note1\[3\] _2208_ _2252_ _2314_ disp_song.um.drum.next_note1\[4\]
+ VGND VGND VPWR VPWR _2400_ sky130_fd_sc_hd__a32o_1
XFILLER_0_11_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold13 game.scoring_button_1.flash_counter_2\[22\] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 disp_song.note1\[0\] VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 game.out\[1\] VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 game.scoring_button_2.next_flash_counter_2\[1\] VGND VGND VPWR VPWR net108
+ sky130_fd_sc_hd__dlygate4sd3_1
X_5249_ _2283_ _2285_ _2256_ VGND VGND VPWR VPWR _2334_ sky130_fd_sc_hd__mux2_1
Xhold57 _0138_ VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 highest_score.highest_score\[7\] VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__dlygate4sd3_1
Xhold68 _0084_ VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2950_ _0310_ _0337_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2881_ disp_song.note2\[9\] _0269_ _0299_ VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__mux2_1
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4620_ _1803_ VGND VGND VPWR VPWR game.scoring_button_1.next_count\[3\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4551_ _1699_ _1740_ _1742_ _1746_ VGND VGND VPWR VPWR game.scoring_button_1.next_num_misses\[8\]
+ sky130_fd_sc_hd__a31o_1
X_4482_ game.scoring_button_1.counts\[19\] game.scoring_button_1.counts\[20\] _1685_
+ game.scoring_button_1.counts\[21\] VGND VGND VPWR VPWR _1686_ sky130_fd_sc_hd__a31o_1
XFILLER_0_12_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3502_ game.flash_counter\[17\] game.flash_counter\[16\] game.flash_counter\[15\]
+ _0864_ VGND VGND VPWR VPWR _0865_ sky130_fd_sc_hd__or4_1
XFILLER_0_0_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3433_ _0702_ _0723_ _0795_ VGND VGND VPWR VPWR _0796_ sky130_fd_sc_hd__o21bai_1
X_6152_ clknet_leaf_31_clk net1 net70 VGND VGND VPWR VPWR disp_song.um.boton0e.sync_b
+ sky130_fd_sc_hd__dfrtp_1
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3364_ game.addhits.a\[13\] game.addhits.add4.b\[1\] VGND VGND VPWR VPWR _0727_ sky130_fd_sc_hd__or2_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5103_ _2190_ VGND VGND VPWR VPWR _2191_ sky130_fd_sc_hd__clkbuf_4
X_6083_ clknet_leaf_23_clk disp_song.um.next_position\[0\] net64 VGND VGND VPWR VPWR
+ disp_song.mi6.in\[0\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_57_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3295_ _0632_ _0657_ VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__nand2_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5034_ _2043_ _2063_ VGND VGND VPWR VPWR _2126_ sky130_fd_sc_hd__nand2_1
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5936_ clknet_leaf_56_clk game.scoring_button_1.next_flash_counter_1\[4\] net51 VGND
+ VGND VPWR VPWR game.scoring_button_1.flash_counter_1\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5867_ clknet_leaf_23_clk net92 net64 VGND VGND VPWR VPWR game.padded_notes2\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4818_ _0248_ _1415_ VGND VGND VPWR VPWR _1933_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5798_ clknet_leaf_53_clk game.scoring_button_2.next_flash_counter_1\[12\] net52
+ VGND VGND VPWR VPWR game.scoring_button_2.flash_counter_1\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4749_ _1884_ game.hit_1 _1885_ VGND VGND VPWR VPWR _1886_ sky130_fd_sc_hd__and3b_1
XFILLER_0_31_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput14 net14 VGND VGND VPWR VPWR green_disp sky130_fd_sc_hd__clkbuf_4
Xoutput25 net25 VGND VGND VPWR VPWR ss1[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput36 net36 VGND VGND VPWR VPWR top_row[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3080_ _0441_ _0442_ VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__nand2_2
XFILLER_0_27_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3982_ game.scoring_button_2.counts\[8\] game.scoring_button_2.counts\[7\] _1294_
+ game.scoring_button_2.counts\[9\] VGND VGND VPWR VPWR _1297_ sky130_fd_sc_hd__a31o_1
XFILLER_0_9_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2933_ _0297_ _0326_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__nand2_1
X_5721_ clknet_leaf_7_clk _0045_ net59 VGND VGND VPWR VPWR pulseout.fin_pulse\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_2864_ _0269_ disp_song.note2\[5\] _0286_ VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__mux2_1
X_5652_ _2610_ _2619_ _2623_ VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__nor3_1
XFILLER_0_45_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4603_ game.scoring_button_1.check_hit.in VGND VGND VPWR VPWR _1791_ sky130_fd_sc_hd__buf_6
X_2795_ lvls.level\[0\] lvls.level\[1\] lvls.level\[2\] VGND VGND VPWR VPWR _0226_
+ sky130_fd_sc_hd__or3b_1
X_5583_ _2580_ net217 _2472_ VGND VGND VPWR VPWR _2581_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4534_ _1691_ _1730_ _1731_ VGND VGND VPWR VPWR _1732_ sky130_fd_sc_hd__or3b_1
XFILLER_0_40_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4465_ _1612_ _1669_ _1670_ _1613_ net206 VGND VGND VPWR VPWR game.scoring_button_1.next_num_hits\[14\]
+ sky130_fd_sc_hd__a32o_1
X_4396_ game.addhits.a\[2\] game.scoring_button_1.acc\[2\] VGND VGND VPWR VPWR _1615_
+ sky130_fd_sc_hd__nor2_1
X_3416_ _0683_ VGND VGND VPWR VPWR _0779_ sky130_fd_sc_hd__inv_2
X_6135_ clknet_leaf_29_clk disp_song.um.drum.next_note2\[15\] net69 VGND VGND VPWR
+ VPWR disp_song.note2\[15\] sky130_fd_sc_hd__dfstp_1
X_3347_ _0708_ _0709_ VGND VGND VPWR VPWR _0710_ sky130_fd_sc_hd__xnor2_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6066_ clknet_leaf_12_clk _0023_ net57 VGND VGND VPWR VPWR game.counter\[22\] sky130_fd_sc_hd__dfrtp_2
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5017_ _2100_ _2101_ _2106_ _2108_ VGND VGND VPWR VPWR _2109_ sky130_fd_sc_hd__a211o_1
X_3278_ _0454_ _0468_ VGND VGND VPWR VPWR _0641_ sky130_fd_sc_hd__xor2_2
XFILLER_0_95_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5919_ clknet_leaf_21_clk game.scoring_button_1.next_count\[10\] net60 VGND VGND
+ VPWR VPWR game.scoring_button_1.counts\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4250_ _1513_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_2\[2\]
+ sky130_fd_sc_hd__clkbuf_1
X_4181_ game.counter\[15\] game.counter\[16\] _1451_ VGND VGND VPWR VPWR _1457_ sky130_fd_sc_hd__and3_1
X_3201_ game.addhits.a\[6\] game.addhits.add2.b\[2\] VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__nor2_1
X_3132_ game.addmisses.a\[11\] game.addmisses.add3.b\[3\] VGND VGND VPWR VPWR _0495_
+ sky130_fd_sc_hd__nand2_1
X_3063_ _0430_ VGND VGND VPWR VPWR disp_song.um.drum.next_note1\[27\] sky130_fd_sc_hd__inv_2
XFILLER_0_54_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3965_ game.addhits.add4.b\[1\] game.addhits.add4.b\[2\] _1275_ VGND VGND VPWR VPWR
+ _1282_ sky130_fd_sc_hd__and3_1
X_2916_ _0324_ VGND VGND VPWR VPWR disp_song.um.drum.next_note2\[19\] sky130_fd_sc_hd__buf_1
XFILLER_0_72_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5704_ clknet_leaf_60_clk _0040_ net50 VGND VGND VPWR VPWR highest_score.highest_score\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_3896_ _0208_ _1226_ VGND VGND VPWR VPWR _1227_ sky130_fd_sc_hd__nor2_8
X_2847_ _0271_ _0273_ VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__nand2_1
X_5635_ _2611_ VGND VGND VPWR VPWR _2612_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_85_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold110 disp_song.note1\[12\] VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__dlygate4sd3_1
X_5566_ _2569_ VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__clkbuf_1
X_2778_ _0214_ _0213_ VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__nand2_1
Xhold121 game.scoring_button_1.flash_counter_2\[16\] VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__dlygate4sd3_1
X_5497_ _2528_ VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold132 disp_song.note1\[22\] VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__dlygate4sd3_1
Xhold143 game.addhits.a\[8\] VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__dlygate4sd3_1
X_4517_ _1691_ _1715_ _1716_ VGND VGND VPWR VPWR _1717_ sky130_fd_sc_hd__o21a_1
XFILLER_0_41_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold154 game.padded_notes2\[6\] VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 game.padded_notes1\[17\] VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4448_ game.addhits.a\[10\] _1653_ VGND VGND VPWR VPWR _1658_ sky130_fd_sc_hd__and2_1
Xhold176 game.addhits.add3.b\[0\] VGND VGND VPWR VPWR net249 sky130_fd_sc_hd__dlygate4sd3_1
Xhold187 game.addhits.a\[9\] VGND VGND VPWR VPWR net260 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_95_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4379_ net171 _1600_ _1413_ VGND VGND VPWR VPWR _1603_ sky130_fd_sc_hd__a21boi_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6118_ clknet_leaf_48_clk disp_song.um.drum.next_note1\[30\] net56 VGND VGND VPWR
+ VPWR disp_song.note1\[30\] sky130_fd_sc_hd__dfstp_1
X_6049_ clknet_leaf_15_clk _0027_ net62 VGND VGND VPWR VPWR game.counter\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3750_ _1077_ _0926_ VGND VGND VPWR VPWR _1105_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2701_ disp_song.um.idx_note2\[3\] _2672_ VGND VGND VPWR VPWR _2673_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_55 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3681_ _1031_ _1033_ _1034_ _1036_ _1032_ VGND VGND VPWR VPWR _1037_ sky130_fd_sc_hd__a311oi_4
X_5420_ _2476_ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5351_ _2423_ _2424_ _2425_ VGND VGND VPWR VPWR _2429_ sky130_fd_sc_hd__and3b_1
X_5282_ _2185_ _2228_ _2364_ _0191_ _2365_ VGND VGND VPWR VPWR _2366_ sky130_fd_sc_hd__o221a_1
XFILLER_0_2_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4302_ game.scoring_button_2.flash_counter_2\[18\] _1546_ VGND VGND VPWR VPWR _1550_
+ sky130_fd_sc_hd__or2_1
X_4233_ _0241_ _1446_ _1497_ _1499_ VGND VGND VPWR VPWR _1500_ sky130_fd_sc_hd__a211oi_1
X_4164_ _1405_ _0012_ VGND VGND VPWR VPWR _1445_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4095_ game.addmisses.add4.b\[2\] _1393_ _1395_ VGND VGND VPWR VPWR _1396_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3115_ game.addmisses.a\[7\] game.addmisses.add2.b\[3\] VGND VGND VPWR VPWR _0478_
+ sky130_fd_sc_hd__nor2_1
X_3046_ _0418_ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_77_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4997_ disp_song.um.drum.next_idx2\[1\] _1965_ _1966_ _2089_ VGND VGND VPWR VPWR
+ _2090_ sky130_fd_sc_hd__a31o_1
X_3948_ game.addhits.add3.b\[3\] _1266_ _1267_ _1269_ VGND VGND VPWR VPWR _1270_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_60_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3879_ _0933_ _1215_ VGND VGND VPWR VPWR _1216_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5618_ _2597_ _2598_ VGND VGND VPWR VPWR _2599_ sky130_fd_sc_hd__and2b_1
XFILLER_0_103_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5549_ disp_song.note1\[14\] game.padded_notes1\[13\] _2541_ VGND VGND VPWR VPWR
+ _2558_ sky130_fd_sc_hd__mux2_1
XTAP_1433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout71 net73 VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__buf_6
Xfanout60 net61 VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__buf_8
XFILLER_0_36_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4920_ disp_song.um.drum.next_note2\[28\] disp_song.um.drum.next_note2\[29\] _1956_
+ VGND VGND VPWR VPWR _2014_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4851_ _0405_ _0352_ _0316_ VGND VGND VPWR VPWR _1947_ sky130_fd_sc_hd__or3b_1
XFILLER_0_28_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3802_ _1151_ _1152_ _1153_ _0921_ VGND VGND VPWR VPWR _1154_ sky130_fd_sc_hd__a31o_1
X_4782_ game.scoring_button_1.flash_counter_1\[12\] _1905_ VGND VGND VPWR VPWR _1909_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_55_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3733_ _0259_ _1073_ _1088_ VGND VGND VPWR VPWR _1089_ sky130_fd_sc_hd__o21ai_1
X_3664_ _0806_ _1015_ _1016_ VGND VGND VPWR VPWR _1020_ sky130_fd_sc_hd__or3b_1
X_5403_ _2464_ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3595_ _0909_ _0913_ _0936_ VGND VGND VPWR VPWR _0956_ sky130_fd_sc_hd__and3_1
XFILLER_0_100_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5334_ game.scoring_button_2.acc\[2\] _2410_ VGND VGND VPWR VPWR _2413_ sky130_fd_sc_hd__and2_1
X_5265_ _2254_ _2260_ VGND VGND VPWR VPWR _2350_ sky130_fd_sc_hd__nor2_1
X_5196_ disp_song.um.drum.next_idx1\[0\] disp_song.um.drum.next_note1\[13\] _2191_
+ _2282_ VGND VGND VPWR VPWR _2283_ sky130_fd_sc_hd__o211a_1
X_4216_ game.scoring_button_2.flash_counter_2\[17\] game.scoring_button_2.flash_counter_2\[16\]
+ game.scoring_button_2.flash_counter_2\[19\] game.scoring_button_2.flash_counter_2\[18\]
+ VGND VGND VPWR VPWR _1484_ sky130_fd_sc_hd__and4_1
XFILLER_0_48_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4147_ _1405_ _1432_ VGND VGND VPWR VPWR _1433_ sky130_fd_sc_hd__and2_1
X_4078_ game.addmisses.add3.b\[3\] _1357_ _1369_ VGND VGND VPWR VPWR _1381_ sky130_fd_sc_hd__and3_1
XFILLER_0_92_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3029_ _0357_ _0355_ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3380_ _0741_ _0742_ VGND VGND VPWR VPWR _0743_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5050_ _2666_ _2085_ _1982_ _2679_ VGND VGND VPWR VPWR _2141_ sky130_fd_sc_hd__o2bb2a_2
X_4001_ _1289_ _1310_ _1312_ _1314_ VGND VGND VPWR VPWR game.scoring_button_2.next_num_misses\[1\]
+ sky130_fd_sc_hd__o2bb2a_1
X_5952_ clknet_leaf_45_clk game.scoring_button_1.next_flash_counter_1\[20\] net53
+ VGND VGND VPWR VPWR game.scoring_button_1.flash_counter_1\[20\] sky130_fd_sc_hd__dfrtp_1
X_4903_ _1990_ _1997_ _1983_ VGND VGND VPWR VPWR _1998_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5883_ clknet_leaf_30_clk _0066_ net69 VGND VGND VPWR VPWR game.padded_notes2\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4834_ _1939_ VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4765_ net162 _1894_ game.hit_1 VGND VGND VPWR VPWR _1897_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_16_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3716_ _1069_ _1071_ _0261_ VGND VGND VPWR VPWR _1072_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4696_ _1849_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_2\[8\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3647_ _0892_ _0994_ _0941_ VGND VGND VPWR VPWR _1004_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_31_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3578_ _0671_ _0939_ _0675_ VGND VGND VPWR VPWR _0940_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5317_ _2379_ _2388_ _2393_ _2399_ _0214_ VGND VGND VPWR VPWR disp_song.um.drum.next_d1\[5\]
+ sky130_fd_sc_hd__o221a_1
Xhold14 game.scoring_button_2.flash_counter_2\[22\] VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 game.counter\[0\] VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 _0090_ VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 _0123_ VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__dlygate4sd3_1
X_5248_ _2252_ _2323_ disp_song.um.drum.next_idx1\[4\] VGND VGND VPWR VPWR _2333_
+ sky130_fd_sc_hd__o21ai_1
X_5179_ _0175_ disp_song.um.drum.next_note1\[21\] VGND VGND VPWR VPWR _2266_ sky130_fd_sc_hd__nand2_1
Xhold69 game.flash_counter\[6\] VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 game.scoring_button_2.hit VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_159 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2880_ _0270_ _0298_ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4550_ game.addmisses.a\[8\] _1743_ _1745_ _1675_ VGND VGND VPWR VPWR _1746_ sky130_fd_sc_hd__o211a_1
XFILLER_0_40_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4481_ game.scoring_button_1.counts\[15\] game.scoring_button_1.counts\[17\] game.scoring_button_1.counts\[16\]
+ _1684_ game.scoring_button_1.counts\[18\] VGND VGND VPWR VPWR _1685_ sky130_fd_sc_hd__a41o_1
X_3501_ game.flash_counter\[12\] game.flash_counter\[13\] _0863_ game.flash_counter\[14\]
+ VGND VGND VPWR VPWR _0864_ sky130_fd_sc_hd__o31a_1
X_3432_ _0702_ _0723_ _0781_ _0794_ _0710_ VGND VGND VPWR VPWR _0795_ sky130_fd_sc_hd__a221o_1
X_6151_ clknet_leaf_29_clk disp_song.um.drum.next_note2\[31\] net69 VGND VGND VPWR
+ VPWR disp_song.note2\[31\] sky130_fd_sc_hd__dfstp_1
X_3363_ game.addhits.a\[13\] game.addhits.add4.b\[1\] VGND VGND VPWR VPWR _0726_ sky130_fd_sc_hd__nand2_1
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5102_ disp_song.um.drum.next_idx1\[4\] disp_song.um.drum.next_idx1\[2\] disp_song.um.drum.next_idx1\[3\]
+ VGND VGND VPWR VPWR _2190_ sky130_fd_sc_hd__or3_1
X_6082_ clknet_leaf_42_clk disp_song.um.drum.next_idx1\[4\] net64 VGND VGND VPWR VPWR
+ disp_song.um.idx_note1\[4\] sky130_fd_sc_hd__dfstp_1
X_3294_ _0646_ _0655_ _0656_ VGND VGND VPWR VPWR _0657_ sky130_fd_sc_hd__a21o_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5033_ _2045_ _2110_ VGND VGND VPWR VPWR _2125_ sky130_fd_sc_hd__or2_1
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5935_ clknet_leaf_60_clk game.scoring_button_1.next_flash_counter_1\[3\] net51 VGND
+ VGND VPWR VPWR game.scoring_button_1.flash_counter_1\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5866_ clknet_leaf_64_clk game.scoring_button_1.next_num_hits\[15\] net50 VGND VGND
+ VPWR VPWR game.addhits.a\[15\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_48_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4817_ net109 _0032_ VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__nor2_1
XFILLER_0_63_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_60_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_60_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_28_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5797_ clknet_leaf_53_clk game.scoring_button_2.next_flash_counter_1\[11\] net52
+ VGND VGND VPWR VPWR game.scoring_button_2.flash_counter_1\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4748_ game.scoring_button_1.flash_counter_1\[1\] game.scoring_button_1.flash_counter_1\[0\]
+ game.scoring_button_1.flash_counter_1\[2\] VGND VGND VPWR VPWR _1885_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4679_ _1836_ game.missed_1 _1837_ VGND VGND VPWR VPWR _1838_ sky130_fd_sc_hd__and3b_1
XFILLER_0_31_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput15 net15 VGND VGND VPWR VPWR red_disp sky130_fd_sc_hd__clkbuf_4
XFILLER_0_31_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput26 net26 VGND VGND VPWR VPWR ss1[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_51_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_51_clk sky130_fd_sc_hd__clkbuf_16
XPHY_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3981_ game.scoring_button_2.counts\[21\] game.scoring_button_2.counts\[22\] _1294_
+ _1295_ VGND VGND VPWR VPWR _1296_ sky130_fd_sc_hd__or4_1
XFILLER_0_57_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2932_ disp_song.um.idx_note2\[3\] disp_song.um.idx_note2\[4\] disp_song.next_red
+ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__and3_1
X_5720_ clknet_leaf_6_clk _0044_ net59 VGND VGND VPWR VPWR pulseout.fin_pulse\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_42_clk clknet_3_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_42_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_45_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2863_ _0273_ _0285_ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5651_ _0842_ _2622_ VGND VGND VPWR VPWR _2623_ sky130_fd_sc_hd__and2_1
X_2794_ game.counter\[14\] _0223_ _0224_ VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__o21a_1
X_5582_ disp_song.note1\[25\] game.padded_notes1\[24\] _2541_ VGND VGND VPWR VPWR
+ _2580_ sky130_fd_sc_hd__mux2_1
X_4602_ _1675_ _1788_ _1790_ VGND VGND VPWR VPWR game.scoring_button_1.next_num_misses\[15\]
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_13_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4533_ game.addmisses.a\[5\] game.addmisses.a\[4\] _1705_ game.addmisses.a\[6\] VGND
+ VGND VPWR VPWR _1731_ sky130_fd_sc_hd__a31o_1
XFILLER_0_53_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4464_ _1665_ _1668_ VGND VGND VPWR VPWR _1670_ sky130_fd_sc_hd__or2_1
XFILLER_0_110_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3415_ _0763_ _0772_ _0771_ VGND VGND VPWR VPWR _0778_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_7_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4395_ _1614_ VGND VGND VPWR VPWR game.scoring_button_1.next_num_hits\[0\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6134_ clknet_leaf_20_clk disp_song.um.drum.next_note2\[14\] net63 VGND VGND VPWR
+ VPWR disp_song.note2\[14\] sky130_fd_sc_hd__dfrtp_1
X_3346_ _0695_ _0701_ _0699_ VGND VGND VPWR VPWR _0709_ sky130_fd_sc_hd__a21o_1
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6065_ clknet_leaf_12_clk _0022_ net57 VGND VGND VPWR VPWR game.counter\[21\] sky130_fd_sc_hd__dfrtp_4
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5016_ _0162_ _2107_ VGND VGND VPWR VPWR _2108_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3277_ _0634_ _0636_ _0639_ VGND VGND VPWR VPWR _0640_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_95_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5918_ clknet_leaf_15_clk game.scoring_button_1.next_count\[9\] net62 VGND VGND VPWR
+ VPWR game.scoring_button_1.counts\[9\] sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_33_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_33_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_75_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5849_ clknet_leaf_69_clk game.scoring_button_1.next_num_misses\[14\] net46 VGND
+ VGND VPWR VPWR game.addmisses.a\[14\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_86_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_24_clk clknet_3_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_24_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_27_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4180_ game.counter\[15\] _1451_ game.counter\[16\] VGND VGND VPWR VPWR _1456_ sky130_fd_sc_hd__a21oi_1
X_3200_ _0540_ _0562_ VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__xor2_4
X_3131_ game.addmisses.a\[11\] game.addmisses.add3.b\[3\] VGND VGND VPWR VPWR _0494_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3062_ _0370_ _0425_ _0429_ VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__o21a_1
XFILLER_0_89_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_118 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_15_clk clknet_3_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_15_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_70_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3964_ net190 _1227_ _1281_ _1226_ VGND VGND VPWR VPWR game.scoring_button_2.next_num_hits\[13\]
+ sky130_fd_sc_hd__a22o_1
X_2915_ _0269_ disp_song.note2\[19\] _0323_ VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5703_ clknet_leaf_60_clk _0039_ net50 VGND VGND VPWR VPWR highest_score.highest_score\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_3895_ _1225_ VGND VGND VPWR VPWR _1226_ sky130_fd_sc_hd__buf_6
X_2846_ _0272_ VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_72_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5634_ game.flash_counter\[6\] game.flash_counter\[7\] game.flash_counter\[5\] _2601_
+ VGND VGND VPWR VPWR _2611_ sky130_fd_sc_hd__and4_1
X_5565_ _2568_ game.padded_notes1\[19\] _2472_ VGND VGND VPWR VPWR _2569_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold100 game.scoring_button_2.flash_counter_1\[13\] VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__dlygate4sd3_1
X_2777_ _2654_ VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__buf_6
Xhold111 game.scoring_button_1.flash_counter_2\[13\] VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__dlygate4sd3_1
Xhold122 game.scoring_button_1.next_flash_counter_2\[16\] VGND VGND VPWR VPWR net195
+ sky130_fd_sc_hd__dlygate4sd3_1
X_5496_ _2527_ game.padded_notes2\[31\] _2515_ VGND VGND VPWR VPWR _2528_ sky130_fd_sc_hd__mux2_1
Xhold144 game.padded_notes1\[25\] VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 game.addhits.a\[14\] VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__dlygate4sd3_1
X_4516_ modetrans.mode\[0\] _1691_ VGND VGND VPWR VPWR _1716_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold166 game.padded_notes2\[26\] VGND VGND VPWR VPWR net239 sky130_fd_sc_hd__dlygate4sd3_1
Xhold177 disp_song.note1\[14\] VGND VGND VPWR VPWR net250 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4447_ game.addhits.a\[10\] _1653_ VGND VGND VPWR VPWR _1657_ sky130_fd_sc_hd__or2_1
Xhold155 game.addhits.a\[11\] VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 game.padded_notes2\[16\] VGND VGND VPWR VPWR net261 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4378_ _1602_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_1\[18\]
+ sky130_fd_sc_hd__clkbuf_1
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6117_ clknet_leaf_40_clk disp_song.um.drum.next_note1\[29\] net66 VGND VGND VPWR
+ VPWR disp_song.note1\[29\] sky130_fd_sc_hd__dfrtp_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3329_ _0684_ _0689_ _0688_ VGND VGND VPWR VPWR _0692_ sky130_fd_sc_hd__a21o_1
X_6048_ clknet_leaf_15_clk _0026_ net62 VGND VGND VPWR VPWR game.counter\[4\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_48_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2700_ disp_song.um.idx_note2\[1\] disp_song.um.idx_note2\[0\] disp_song.um.idx_note2\[2\]
+ VGND VGND VPWR VPWR _2672_ sky130_fd_sc_hd__or3_2
XFILLER_0_54_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3680_ _1025_ _1033_ _1035_ VGND VGND VPWR VPWR _1036_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5350_ _2418_ _2419_ _2420_ _2422_ _2427_ VGND VGND VPWR VPWR _2428_ sky130_fd_sc_hd__o2111a_1
X_5281_ _2361_ VGND VGND VPWR VPWR _2365_ sky130_fd_sc_hd__inv_2
X_4301_ game.scoring_button_2.flash_counter_2\[18\] _1546_ VGND VGND VPWR VPWR _1549_
+ sky130_fd_sc_hd__and2_1
X_4232_ game.counter\[13\] game.counter\[12\] _1498_ _0227_ VGND VGND VPWR VPWR _1499_
+ sky130_fd_sc_hd__o31a_1
Xclkbuf_leaf_4_clk clknet_3_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_4_clk sky130_fd_sc_hd__clkbuf_16
X_4163_ net144 _1443_ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4094_ _1358_ _1394_ VGND VGND VPWR VPWR _1395_ sky130_fd_sc_hd__or2_1
X_3114_ _0471_ _0476_ VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__and2_1
X_3045_ _0264_ _0409_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__and2_1
X_4996_ _2088_ VGND VGND VPWR VPWR _2089_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3947_ _1266_ _1267_ _1268_ VGND VGND VPWR VPWR _1269_ sky130_fd_sc_hd__o21ai_1
X_3878_ _0966_ disp_song.display_note2\[3\] _0211_ game.out\[3\] _0208_ VGND VGND
+ VPWR VPWR _1215_ sky130_fd_sc_hd__a221o_2
XFILLER_0_61_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5617_ game.flash_counter\[2\] _2595_ game.flash_counter\[3\] VGND VGND VPWR VPWR
+ _2598_ sky130_fd_sc_hd__a21o_1
X_2829_ highest_score.score_mode\[1\] VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_103_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5548_ _2557_ VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5479_ _2516_ VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__clkbuf_1
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout72 net73 VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__buf_4
Xfanout61 net73 VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__clkbuf_8
Xfanout50 net52 VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__buf_8
XFILLER_0_107_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_3_7__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_7__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_99_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4850_ _1946_ VGND VGND VPWR VPWR disp_song.um.next_position\[3\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3801_ _1122_ _1133_ _0955_ VGND VGND VPWR VPWR _1153_ sky130_fd_sc_hd__a21o_1
X_4781_ game.scoring_button_1.flash_counter_1\[12\] _1905_ VGND VGND VPWR VPWR _1908_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3732_ _0352_ _1085_ _1087_ VGND VGND VPWR VPWR _1088_ sky130_fd_sc_hd__or3b_1
XFILLER_0_82_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3663_ _0775_ _1018_ _0776_ net43 VGND VGND VPWR VPWR _1019_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_43_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5402_ _2463_ game.padded_notes2\[1\] _2462_ VGND VGND VPWR VPWR _2464_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3594_ _0255_ _0258_ VGND VGND VPWR VPWR _0955_ sky130_fd_sc_hd__nand2_2
X_5333_ _2412_ VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__clkbuf_1
X_5264_ disp_song.note1\[24\] disp_song.um.drum.next_note1\[25\] _0175_ VGND VGND
+ VPWR VPWR _2349_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5195_ _0175_ disp_song.um.drum.next_note1\[12\] VGND VGND VPWR VPWR _2282_ sky130_fd_sc_hd__or2_1
X_4215_ game.scoring_button_2.flash_counter_2\[21\] game.scoring_button_2.flash_counter_2\[20\]
+ game.scoring_button_2.flash_counter_2\[22\] VGND VGND VPWR VPWR _1483_ sky130_fd_sc_hd__or3_1
X_4146_ game.counter\[8\] _1429_ VGND VGND VPWR VPWR _1432_ sky130_fd_sc_hd__xor2_1
XFILLER_0_97_308 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4077_ game.addmisses.add4.b\[0\] _1363_ VGND VGND VPWR VPWR _1380_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_544 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3028_ _0177_ _0181_ _0264_ _0405_ _0406_ VGND VGND VPWR VPWR disp_song.um.drum.next_note1\[16\]
+ sky130_fd_sc_hd__a41o_1
XFILLER_0_108_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4979_ _2011_ _2072_ VGND VGND VPWR VPWR _2073_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4000_ game.addmisses.add1.b\[3\] _1309_ _1313_ VGND VGND VPWR VPWR _1314_ sky130_fd_sc_hd__o21ai_1
X_5951_ clknet_leaf_61_clk game.scoring_button_1.next_flash_counter_1\[19\] net53
+ VGND VGND VPWR VPWR game.scoring_button_1.flash_counter_1\[19\] sky130_fd_sc_hd__dfrtp_1
X_4902_ _2666_ _1965_ _1991_ _1996_ VGND VGND VPWR VPWR _1997_ sky130_fd_sc_hd__a31o_1
XFILLER_0_75_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5882_ clknet_leaf_30_clk _0065_ net69 VGND VGND VPWR VPWR game.padded_notes2\[15\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_62_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4833_ _0032_ _1458_ VGND VGND VPWR VPWR _1939_ sky130_fd_sc_hd__and2b_1
XFILLER_0_47_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4764_ _1896_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_1\[6\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3715_ _1067_ _1070_ _1066_ _1068_ VGND VGND VPWR VPWR _1071_ sky130_fd_sc_hd__o211a_1
XFILLER_0_55_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4695_ _1847_ game.missed_1 _1848_ VGND VGND VPWR VPWR _1849_ sky130_fd_sc_hd__and3b_1
XFILLER_0_31_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3646_ _0840_ _0859_ VGND VGND VPWR VPWR _1003_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3577_ _0671_ net44 VGND VGND VPWR VPWR _0939_ sky130_fd_sc_hd__nand2_1
XFILLER_0_87_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5316_ _2387_ _2398_ _2379_ VGND VGND VPWR VPWR _2399_ sky130_fd_sc_hd__o21ai_1
X_5247_ disp_song.um.drum.next_note1\[0\] _2208_ _2252_ _2312_ disp_song.um.drum.next_note1\[2\]
+ VGND VGND VPWR VPWR _2332_ sky130_fd_sc_hd__a32o_1
Xhold26 game.flash_counter\[1\] VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 game.scoring_button_2.next_flash_counter_2\[22\] VGND VGND VPWR VPWR net88
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 game.out\[13\] VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 game.flash_counter\[14\] VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__dlygate4sd3_1
X_5178_ _2247_ _2255_ _2264_ VGND VGND VPWR VPWR _2265_ sky130_fd_sc_hd__o21ba_1
Xhold59 _0049_ VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4129_ _1421_ VGND VGND VPWR VPWR game.scoring_button_2.next_count\[3\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_107_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3500_ game.flash_counter\[10\] _0862_ game.flash_counter\[11\] VGND VGND VPWR VPWR
+ _0863_ sky130_fd_sc_hd__o21a_1
XFILLER_0_25_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4480_ game.scoring_button_1.counts\[11\] game.scoring_button_1.counts\[10\] _1683_
+ _1676_ VGND VGND VPWR VPWR _1684_ sky130_fd_sc_hd__a31o_1
XFILLER_0_40_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3431_ _0784_ _0790_ _0793_ VGND VGND VPWR VPWR _0794_ sky130_fd_sc_hd__a21o_1
X_6150_ clknet_leaf_32_clk disp_song.um.drum.next_note2\[30\] net70 VGND VGND VPWR
+ VPWR disp_song.note2\[30\] sky130_fd_sc_hd__dfrtp_1
X_3362_ _0595_ _0723_ _0724_ VGND VGND VPWR VPWR _0725_ sky130_fd_sc_hd__o21bai_4
XFILLER_0_0_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5101_ _2188_ VGND VGND VPWR VPWR _2189_ sky130_fd_sc_hd__inv_2
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6081_ clknet_leaf_43_clk disp_song.um.drum.next_idx1\[3\] net65 VGND VGND VPWR VPWR
+ disp_song.um.idx_note1\[3\] sky130_fd_sc_hd__dfstp_2
X_3293_ _0649_ _0654_ VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__and2_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5032_ _2040_ _2069_ _2110_ VGND VGND VPWR VPWR _2124_ sky130_fd_sc_hd__mux2_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_75 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5934_ clknet_leaf_60_clk game.scoring_button_1.next_flash_counter_1\[2\] net51 VGND
+ VGND VPWR VPWR game.scoring_button_1.flash_counter_1\[2\] sky130_fd_sc_hd__dfrtp_1
X_5865_ clknet_leaf_64_clk game.scoring_button_1.next_num_hits\[14\] net47 VGND VGND
+ VPWR VPWR game.addhits.a\[14\] sky130_fd_sc_hd__dfrtp_2
X_4816_ net85 _1929_ _1932_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_1\[22\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5796_ clknet_leaf_53_clk game.scoring_button_2.next_flash_counter_1\[10\] net52
+ VGND VGND VPWR VPWR game.scoring_button_2.flash_counter_1\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4747_ game.scoring_button_1.flash_counter_1\[1\] game.scoring_button_1.flash_counter_1\[0\]
+ game.scoring_button_1.flash_counter_1\[2\] VGND VGND VPWR VPWR _1884_ sky130_fd_sc_hd__and3_1
XFILLER_0_43_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4678_ game.scoring_button_1.flash_counter_2\[3\] _1833_ VGND VGND VPWR VPWR _1837_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_71_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3629_ _0928_ _0965_ VGND VGND VPWR VPWR _0988_ sky130_fd_sc_hd__or2b_1
XFILLER_0_101_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput16 net16 VGND VGND VPWR VPWR ss0[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput27 net27 VGND VGND VPWR VPWR ss1[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3980_ game.scoring_button_2.counts\[20\] game.scoring_button_2.counts\[19\] game.scoring_button_2.counts\[18\]
+ game.scoring_button_2.counts\[17\] VGND VGND VPWR VPWR _1295_ sky130_fd_sc_hd__or4_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2931_ _0294_ _0330_ _0333_ disp_song.note2\[24\] VGND VGND VPWR VPWR disp_song.um.drum.next_note2\[24\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5650_ _0868_ _0870_ _2621_ VGND VGND VPWR VPWR _2622_ sky130_fd_sc_hd__and3_1
XFILLER_0_45_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
X_2862_ disp_song.um.idx_note2\[1\] disp_song.um.idx_note2\[0\] disp_song.um.idx_note2\[2\]
+ VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__and3b_1
X_4601_ game.addmisses.a\[15\] _1781_ _1789_ _1699_ VGND VGND VPWR VPWR _1790_ sky130_fd_sc_hd__a211o_1
XFILLER_0_38_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2793_ game.counter\[20\] _0222_ VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__or2_1
X_5581_ _2579_ VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_25_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4532_ game.addmisses.a\[6\] game.addmisses.a\[5\] game.addmisses.a\[4\] _1705_ VGND
+ VGND VPWR VPWR _1730_ sky130_fd_sc_hd__and4_1
XFILLER_0_13_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4463_ _0741_ _1668_ _1663_ VGND VGND VPWR VPWR _1669_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_111_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3414_ _0763_ _0771_ VGND VGND VPWR VPWR _0777_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4394_ _1612_ _1613_ game.addhits.a\[0\] VGND VGND VPWR VPWR _1614_ sky130_fd_sc_hd__mux2_1
X_6133_ clknet_leaf_19_clk disp_song.um.drum.next_note2\[13\] net63 VGND VGND VPWR
+ VPWR disp_song.note2\[13\] sky130_fd_sc_hd__dfstp_1
X_3345_ _0704_ _0707_ VGND VGND VPWR VPWR _0708_ sky130_fd_sc_hd__xnor2_2
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6064_ clknet_leaf_12_clk _0021_ net57 VGND VGND VPWR VPWR game.counter\[20\] sky130_fd_sc_hd__dfrtp_2
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3276_ _0638_ VGND VGND VPWR VPWR _0639_ sky130_fd_sc_hd__inv_2
X_5015_ _2019_ _2085_ VGND VGND VPWR VPWR _2107_ sky130_fd_sc_hd__and2_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5917_ clknet_leaf_15_clk game.scoring_button_1.next_count\[8\] net58 VGND VGND VPWR
+ VPWR game.scoring_button_1.counts\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5848_ clknet_leaf_69_clk game.scoring_button_1.next_num_misses\[13\] net46 VGND
+ VGND VPWR VPWR game.addmisses.a\[13\] sky130_fd_sc_hd__dfrtp_2
X_5779_ clknet_leaf_11_clk game.scoring_button_2.next_count\[16\] net57 VGND VGND
+ VPWR VPWR game.scoring_button_2.counts\[16\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3130_ _0487_ _0492_ VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3061_ _0370_ _0426_ disp_song.note1\[27\] VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3963_ _1277_ _1279_ _1280_ VGND VGND VPWR VPWR _1281_ sky130_fd_sc_hd__o21ai_1
X_2914_ disp_song.um.idx_note2\[3\] _0318_ _0160_ _0279_ VGND VGND VPWR VPWR _0323_
+ sky130_fd_sc_hd__or4_1
XFILLER_0_70_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5702_ clknet_leaf_61_clk _0038_ net53 VGND VGND VPWR VPWR highest_score.highest_score\[3\]
+ sky130_fd_sc_hd__dfrtp_2
X_3894_ game.scoring_button_2.check_hit.edge_1 game.scoring_button_2.check_hit.edge_2
+ game.scoring_button_2.hit VGND VGND VPWR VPWR _1225_ sky130_fd_sc_hd__and3b_1
X_2845_ _2654_ _0156_ _2676_ _2675_ VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__and4_1
XFILLER_0_72_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5633_ _2602_ _2604_ _2605_ _2609_ VGND VGND VPWR VPWR _2610_ sky130_fd_sc_hd__nor4_1
X_5564_ disp_song.note1\[19\] game.padded_notes1\[18\] _2541_ VGND VGND VPWR VPWR
+ _2568_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2776_ modetrans.mode\[3\] _0207_ _0212_ _0213_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__o31a_1
Xhold101 game.scoring_button_2.flash_counter_1\[16\] VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__dlygate4sd3_1
X_4515_ game.addmisses.a\[4\] _1705_ VGND VGND VPWR VPWR _1715_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5495_ disp_song.note2\[31\] game.padded_notes2\[30\] _2497_ VGND VGND VPWR VPWR
+ _2527_ sky130_fd_sc_hd__mux2_1
Xhold123 game.addhits.a\[10\] VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__dlygate4sd3_1
Xhold134 game.scoring_button_1.flash_counter_1\[4\] VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__dlygate4sd3_1
Xhold112 game.scoring_button_2.flash_counter_2\[16\] VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold156 game.padded_notes2\[10\] VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 game.padded_notes1\[4\] VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 disp_song.note1\[18\] VGND VGND VPWR VPWR net240 sky130_fd_sc_hd__dlygate4sd3_1
X_4446_ net260 _1613_ _1656_ _1612_ VGND VGND VPWR VPWR game.scoring_button_1.next_num_hits\[9\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold178 game.padded_notes2\[20\] VGND VGND VPWR VPWR net251 sky130_fd_sc_hd__dlygate4sd3_1
Xhold189 disp_song.note1\[6\] VGND VGND VPWR VPWR net262 sky130_fd_sc_hd__dlygate4sd3_1
X_4377_ _1600_ _1413_ _1601_ VGND VGND VPWR VPWR _1602_ sky130_fd_sc_hd__and3b_1
XFILLER_0_95_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3328_ _0684_ _0690_ VGND VGND VPWR VPWR _0691_ sky130_fd_sc_hd__xnor2_1
X_6116_ clknet_leaf_48_clk disp_song.um.drum.next_note1\[28\] net56 VGND VGND VPWR
+ VPWR disp_song.note1\[28\] sky130_fd_sc_hd__dfrtp_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6047_ clknet_leaf_16_clk _0025_ net62 VGND VGND VPWR VPWR game.counter\[3\] sky130_fd_sc_hd__dfrtp_1
X_3259_ _0620_ _0621_ VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5280_ disp_song.note1\[18\] disp_song.um.drum.next_note1\[19\] disp_song.um.drum.next_idx1\[0\]
+ VGND VGND VPWR VPWR _2364_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4300_ _1548_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_2\[17\]
+ sky130_fd_sc_hd__clkbuf_1
X_4231_ game.counter\[21\] VGND VGND VPWR VPWR _1498_ sky130_fd_sc_hd__inv_2
X_4162_ _1444_ VGND VGND VPWR VPWR game.scoring_button_2.next_count\[11\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4093_ game.addmisses.add4.b\[2\] _1381_ _1385_ VGND VGND VPWR VPWR _1394_ sky130_fd_sc_hd__and3_1
X_3113_ _0472_ _0475_ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__xnor2_2
X_3044_ _0377_ _0410_ _0417_ VGND VGND VPWR VPWR disp_song.um.drum.next_note1\[21\]
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_81_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4995_ _2666_ _1969_ VGND VGND VPWR VPWR _2088_ sky130_fd_sc_hd__nand2_1
XFILLER_0_105_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3946_ game.addhits.add3.b\[2\] game.addhits.add3.b\[1\] _1264_ game.addhits.add3.b\[3\]
+ VGND VGND VPWR VPWR _1268_ sky130_fd_sc_hd__o31a_1
XFILLER_0_45_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3877_ _1214_ VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_475 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5616_ game.flash_counter\[3\] game.flash_counter\[2\] _2595_ VGND VGND VPWR VPWR
+ _2597_ sky130_fd_sc_hd__and3_1
X_2828_ _0256_ _0257_ VGND VGND VPWR VPWR highest_score.nxt_mode\[0\] sky130_fd_sc_hd__nand2_1
XFILLER_0_45_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5547_ _2556_ net243 _2515_ VGND VGND VPWR VPWR _2557_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2759_ _0199_ VGND VGND VPWR VPWR disp_song.um.drum.next_idx1\[1\] sky130_fd_sc_hd__inv_6
X_5478_ _2514_ game.padded_notes2\[25\] _2515_ VGND VGND VPWR VPWR _2516_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4429_ game.addhits.a\[5\] VGND VGND VPWR VPWR _1643_ sky130_fd_sc_hd__inv_2
XFILLER_0_111_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout62 net63 VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__buf_6
Xfanout73 net6 VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__buf_12
Xfanout51 net52 VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_8
XFILLER_0_107_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4780_ _1907_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_1\[11\]
+ sky130_fd_sc_hd__clkbuf_1
X_3800_ _1060_ _1123_ _1135_ _0258_ VGND VGND VPWR VPWR _1152_ sky130_fd_sc_hd__a31o_1
XFILLER_0_7_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3731_ _1077_ _1084_ _1086_ _0925_ _1080_ VGND VGND VPWR VPWR _1087_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_43_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3662_ _1012_ _0807_ _1015_ _1017_ VGND VGND VPWR VPWR _1018_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5401_ disp_song.note2\[1\] game.padded_notes2\[0\] _0219_ VGND VGND VPWR VPWR _2463_
+ sky130_fd_sc_hd__mux2_1
X_3593_ _0951_ _0954_ _0935_ VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__o21a_1
X_5332_ net252 _2411_ VGND VGND VPWR VPWR _2412_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5263_ _2249_ _2251_ _2256_ VGND VGND VPWR VPWR _2348_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4214_ game.scoring_button_2.flash_counter_2\[8\] game.scoring_button_2.flash_counter_2\[11\]
+ game.scoring_button_2.flash_counter_2\[10\] game.scoring_button_2.flash_counter_2\[9\]
+ VGND VGND VPWR VPWR _1482_ sky130_fd_sc_hd__or4b_1
X_5194_ _2265_ _2279_ _2280_ VGND VGND VPWR VPWR _2281_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4145_ _1431_ VGND VGND VPWR VPWR game.scoring_button_2.next_count\[7\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_92_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4076_ game.addmisses.add4.b\[0\] _1363_ VGND VGND VPWR VPWR _1379_ sky130_fd_sc_hd__and2_1
X_3027_ _2661_ _0404_ _0182_ _0265_ disp_song.note1\[16\] VGND VGND VPWR VPWR _0406_
+ sky130_fd_sc_hd__o41a_1
XFILLER_0_78_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4978_ _2062_ _2071_ _2032_ VGND VGND VPWR VPWR _2072_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3929_ _1253_ _1254_ VGND VGND VPWR VPWR _1255_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5950_ clknet_leaf_61_clk game.scoring_button_1.next_flash_counter_1\[18\] net53
+ VGND VGND VPWR VPWR game.scoring_button_1.flash_counter_1\[18\] sky130_fd_sc_hd__dfrtp_1
X_4901_ _1992_ _1995_ VGND VGND VPWR VPWR _1996_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5881_ clknet_leaf_20_clk _0064_ net69 VGND VGND VPWR VPWR game.padded_notes2\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_4832_ _1938_ VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4763_ _1894_ _1799_ _1895_ VGND VGND VPWR VPWR _1896_ sky130_fd_sc_hd__and3b_1
XFILLER_0_43_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4694_ game.scoring_button_1.flash_counter_2\[7\] game.scoring_button_1.flash_counter_2\[6\]
+ _1840_ game.scoring_button_1.flash_counter_2\[8\] VGND VGND VPWR VPWR _1848_ sky130_fd_sc_hd__a31o_1
XFILLER_0_15_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3714_ _0629_ _0636_ VGND VGND VPWR VPWR _1070_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3645_ _1001_ _1002_ _0935_ VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__o21a_1
XFILLER_0_43_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3576_ _0614_ _0914_ _0937_ _0261_ VGND VGND VPWR VPWR _0938_ sky130_fd_sc_hd__o31a_1
XFILLER_0_11_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5315_ _2397_ VGND VGND VPWR VPWR _2398_ sky130_fd_sc_hd__inv_2
X_5246_ disp_song.um.drum.next_note1\[1\] _2314_ VGND VGND VPWR VPWR _2331_ sky130_fd_sc_hd__and2_1
XFILLER_0_53_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold27 _2596_ VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 game.scoring_button_2.flash_counter_1\[22\] VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 game.scoring_button_1.flash_counter_1\[1\] VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 disp_song.note1\[28\] VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__dlygate4sd3_1
X_5177_ _2256_ _2260_ _2262_ _2263_ _2247_ VGND VGND VPWR VPWR _2264_ sky130_fd_sc_hd__o221a_1
X_4128_ _1405_ _0025_ VGND VGND VPWR VPWR _1421_ sky130_fd_sc_hd__and2_1
X_4059_ game.addmisses.add3.b\[3\] _1361_ _1362_ VGND VGND VPWR VPWR _1365_ sky130_fd_sc_hd__and3b_1
XFILLER_0_109_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3430_ _0680_ _0792_ VGND VGND VPWR VPWR _0793_ sky130_fd_sc_hd__or2_1
X_3361_ _0594_ _0504_ _0528_ VGND VGND VPWR VPWR _0724_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6080_ clknet_leaf_43_clk disp_song.um.drum.next_idx1\[2\] net64 VGND VGND VPWR VPWR
+ disp_song.um.idx_note1\[2\] sky130_fd_sc_hd__dfstp_4
XFILLER_0_0_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5100_ _2185_ _2186_ _2187_ _0197_ VGND VGND VPWR VPWR _2188_ sky130_fd_sc_hd__a2bb2o_1
X_5031_ _2120_ _2122_ _2108_ VGND VGND VPWR VPWR _2123_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3292_ _0649_ _0654_ VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__xor2_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5933_ clknet_leaf_60_clk net112 net51 VGND VGND VPWR VPWR game.scoring_button_1.flash_counter_1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5864_ clknet_leaf_59_clk game.scoring_button_1.next_num_hits\[13\] net47 VGND VGND
+ VPWR VPWR game.addhits.a\[13\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_75_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4815_ net85 _1929_ game.hit_1 VGND VGND VPWR VPWR _1932_ sky130_fd_sc_hd__o21ai_1
X_5795_ clknet_leaf_53_clk game.scoring_button_2.next_flash_counter_1\[9\] net52 VGND
+ VGND VPWR VPWR game.scoring_button_2.flash_counter_1\[9\] sky130_fd_sc_hd__dfrtp_1
X_4746_ net111 game.scoring_button_1.flash_counter_1\[0\] _1883_ VGND VGND VPWR VPWR
+ game.scoring_button_1.next_flash_counter_1\[1\] sky130_fd_sc_hd__a21oi_1
X_4677_ game.scoring_button_1.flash_counter_2\[3\] _1833_ VGND VGND VPWR VPWR _1836_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_43_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3628_ _0981_ _0985_ _0986_ _0949_ modetrans.mode\[3\] VGND VGND VPWR VPWR _0987_
+ sky130_fd_sc_hd__o221a_1
Xoutput17 net17 VGND VGND VPWR VPWR ss0[1] sky130_fd_sc_hd__clkbuf_4
Xoutput28 net28 VGND VGND VPWR VPWR ss1[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3559_ _0897_ _0908_ _0920_ _0921_ VGND VGND VPWR VPWR _0922_ sky130_fd_sc_hd__a31o_1
X_5229_ disp_song.um.drum.next_note1\[1\] _2312_ _2314_ disp_song.um.drum.next_note1\[0\]
+ VGND VGND VPWR VPWR _2315_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_570 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2930_ _2672_ _0158_ _0327_ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__or3_1
XFILLER_0_85_643 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2861_ _0264_ _0283_ _0284_ disp_song.note2\[4\] VGND VGND VPWR VPWR disp_song.um.drum.next_note2\[4\]
+ sky130_fd_sc_hd__a22o_1
X_4600_ game.addmisses.a\[15\] _1780_ VGND VGND VPWR VPWR _1789_ sky130_fd_sc_hd__nor2_1
X_2792_ game.counter\[20\] _0222_ VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__nand2_1
X_5580_ _2578_ net210 _2472_ VGND VGND VPWR VPWR _2579_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4531_ game.addmisses.a\[6\] _1728_ VGND VGND VPWR VPWR _1729_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_111_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4462_ game.addhits.a\[13\] game.addhits.a\[14\] _1661_ VGND VGND VPWR VPWR _1668_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_68_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3413_ _0763_ _0771_ _0772_ _0752_ VGND VGND VPWR VPWR _0776_ sky130_fd_sc_hd__a211o_1
XFILLER_0_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4393_ _0208_ _1612_ VGND VGND VPWR VPWR _1613_ sky130_fd_sc_hd__nor2_8
XFILLER_0_110_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6132_ clknet_leaf_20_clk disp_song.um.drum.next_note2\[12\] net63 VGND VGND VPWR
+ VPWR disp_song.note2\[12\] sky130_fd_sc_hd__dfrtp_1
X_3344_ _0600_ _0706_ VGND VGND VPWR VPWR _0707_ sky130_fd_sc_hd__nor2_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6063_ clknet_leaf_12_clk _0019_ net58 VGND VGND VPWR VPWR game.counter\[19\] sky130_fd_sc_hd__dfrtp_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3275_ _0544_ _0637_ VGND VGND VPWR VPWR _0638_ sky130_fd_sc_hd__nand2_2
X_5014_ _2042_ _2103_ _2104_ _2020_ _2105_ VGND VGND VPWR VPWR _2106_ sky130_fd_sc_hd__o221a_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5916_ clknet_leaf_14_clk game.scoring_button_1.next_count\[7\] net58 VGND VGND VPWR
+ VPWR game.scoring_button_1.counts\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5847_ clknet_3_0__leaf_clk game.scoring_button_1.next_num_misses\[12\] net46 VGND
+ VGND VPWR VPWR game.addmisses.a\[12\] sky130_fd_sc_hd__dfrtp_2
X_5778_ clknet_leaf_11_clk game.scoring_button_2.next_count\[15\] net57 VGND VGND
+ VPWR VPWR game.scoring_button_2.counts\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4729_ _1871_ _1830_ _1872_ VGND VGND VPWR VPWR _1873_ sky130_fd_sc_hd__and3b_1
XFILLER_0_16_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_495 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3060_ _0362_ _0425_ _0428_ VGND VGND VPWR VPWR disp_song.um.drum.next_note1\[26\]
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3962_ game.addhits.add4.b\[3\] _1278_ VGND VGND VPWR VPWR _1280_ sky130_fd_sc_hd__or2_1
X_5701_ clknet_leaf_62_clk _0037_ net53 VGND VGND VPWR VPWR highest_score.highest_score\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_2913_ _0322_ VGND VGND VPWR VPWR disp_song.um.drum.next_note2\[18\] sky130_fd_sc_hd__buf_1
X_3893_ _1224_ VGND VGND VPWR VPWR modetrans.pushed_3 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2844_ _0270_ VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__inv_2
X_5632_ _2606_ _2607_ _2608_ VGND VGND VPWR VPWR _2609_ sky130_fd_sc_hd__or3_1
X_5563_ _2567_ VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2775_ net114 modetrans.u2.Q1 VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__or2b_1
XFILLER_0_5_467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4514_ _1675_ _1713_ VGND VGND VPWR VPWR _1714_ sky130_fd_sc_hd__nor2_1
X_5494_ _2526_ VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__clkbuf_1
Xhold124 disp_song.note1\[30\] VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__dlygate4sd3_1
Xhold102 game.flash_counter\[21\] VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold113 game.scoring_button_2.next_flash_counter_2\[16\] VGND VGND VPWR VPWR net186
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 game.addhits.a\[2\] VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold157 game.padded_notes2\[18\] VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__dlygate4sd3_1
Xhold168 game.padded_notes1\[12\] VGND VGND VPWR VPWR net241 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold146 game.addhits.add3.b\[3\] VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__dlygate4sd3_1
X_4445_ game.addhits.a\[11\] _1652_ _1653_ _1655_ VGND VGND VPWR VPWR _1656_ sky130_fd_sc_hd__o31ai_1
X_4376_ game.scoring_button_2.flash_counter_1\[18\] _1597_ VGND VGND VPWR VPWR _1601_
+ sky130_fd_sc_hd__or2_1
Xhold179 game.scoring_button_2.acc\[1\] VGND VGND VPWR VPWR net252 sky130_fd_sc_hd__dlygate4sd3_1
X_6115_ clknet_leaf_40_clk disp_song.um.drum.next_note1\[27\] net66 VGND VGND VPWR
+ VPWR disp_song.note1\[27\] sky130_fd_sc_hd__dfstp_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3327_ _0688_ _0689_ VGND VGND VPWR VPWR _0690_ sky130_fd_sc_hd__and2b_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6046_ clknet_leaf_16_clk _0024_ net62 VGND VGND VPWR VPWR game.counter\[2\] sky130_fd_sc_hd__dfrtp_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3258_ _0608_ _0619_ VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__or2_1
X_3189_ _0548_ _0551_ VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_76_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_587 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4230_ game.counter\[16\] game.counter\[17\] game.counter\[18\] _0245_ VGND VGND
+ VPWR VPWR _1497_ sky130_fd_sc_hd__o22a_1
X_4161_ game.scoring_button_2.check_hit.in _1442_ _1443_ VGND VGND VPWR VPWR _1444_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_65_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4092_ _1381_ _1385_ VGND VGND VPWR VPWR _1393_ sky130_fd_sc_hd__and2_1
X_3112_ _0473_ _0474_ VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__or2b_1
X_3043_ _0377_ _0412_ net245 VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_81_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4994_ _2079_ _2084_ _2086_ VGND VGND VPWR VPWR _2087_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3945_ game.addhits.add3.b\[1\] game.addhits.add3.b\[0\] _1253_ VGND VGND VPWR VPWR
+ _1267_ sky130_fd_sc_hd__and3_1
XFILLER_0_18_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3876_ _0933_ _1213_ VGND VGND VPWR VPWR _1214_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5615_ net113 _2595_ VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__xor2_1
XFILLER_0_45_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2827_ _0255_ _2659_ VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5546_ disp_song.note1\[13\] game.padded_notes1\[12\] _2541_ VGND VGND VPWR VPWR
+ _2556_ sky130_fd_sc_hd__mux2_1
X_2758_ _2654_ _0198_ VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__and2_2
X_5477_ _2472_ VGND VGND VPWR VPWR _2515_ sky130_fd_sc_hd__buf_8
XFILLER_0_14_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2689_ disp_song.um.idx_note2\[0\] _2662_ VGND VGND VPWR VPWR _2663_ sky130_fd_sc_hd__or2_1
X_4428_ game.addhits.a\[6\] VGND VGND VPWR VPWR _1642_ sky130_fd_sc_hd__inv_2
X_4359_ net173 _1586_ game.hit_2 VGND VGND VPWR VPWR _1589_ sky130_fd_sc_hd__a21boi_1
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6029_ clknet_leaf_59_clk net130 net51 VGND VGND VPWR VPWR game.flash_counter\[9\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_1414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout63 net73 VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__buf_8
XFILLER_0_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout52 net73 VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__buf_8
XFILLER_0_52_616 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3730_ disp_song.mi6.in\[2\] _1077_ VGND VGND VPWR VPWR _1086_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3661_ _0786_ _0806_ _1016_ VGND VGND VPWR VPWR _1017_ sky130_fd_sc_hd__and3_1
X_5400_ disp_song.note2\[0\] _2458_ _2462_ net91 VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__a22o_1
X_3592_ _0211_ net39 _0948_ _0953_ _0214_ VGND VGND VPWR VPWR _0954_ sky130_fd_sc_hd__a311o_1
X_5331_ _2410_ VGND VGND VPWR VPWR _2411_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5262_ _2340_ _2344_ _2346_ VGND VGND VPWR VPWR _2347_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4213_ game.scoring_button_2.flash_counter_2\[13\] game.scoring_button_2.flash_counter_2\[12\]
+ game.scoring_button_2.flash_counter_2\[15\] game.scoring_button_2.flash_counter_2\[14\]
+ VGND VGND VPWR VPWR _1481_ sky130_fd_sc_hd__or4b_1
X_5193_ _2186_ _2244_ _2257_ VGND VGND VPWR VPWR _2280_ sky130_fd_sc_hd__o21a_1
X_4144_ _1405_ _1430_ VGND VGND VPWR VPWR _1431_ sky130_fd_sc_hd__and2_1
XFILLER_0_92_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4075_ _1378_ VGND VGND VPWR VPWR game.scoring_button_2.next_num_misses\[11\] sky130_fd_sc_hd__clkbuf_1
X_3026_ _2661_ _0404_ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4977_ _2066_ _2070_ _2034_ VGND VGND VPWR VPWR _2071_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3928_ game.addhits.add2.b\[1\] _1251_ VGND VGND VPWR VPWR _1254_ sky130_fd_sc_hd__xnor2_1
X_3859_ _1202_ VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5529_ _2544_ game.padded_notes1\[7\] _2515_ VGND VGND VPWR VPWR _2545_ sky130_fd_sc_hd__mux2_1
XTAP_1222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5880_ clknet_leaf_20_clk _0063_ net63 VGND VGND VPWR VPWR game.padded_notes2\[13\]
+ sky130_fd_sc_hd__dfstp_1
X_4900_ _2666_ _1994_ VGND VGND VPWR VPWR _1995_ sky130_fd_sc_hd__or2_1
XFILLER_0_75_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4831_ _0032_ _1454_ VGND VGND VPWR VPWR _1938_ sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_72_clk clknet_3_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_72_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4762_ game.scoring_button_1.flash_counter_1\[6\] _1891_ VGND VGND VPWR VPWR _1895_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_55_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4693_ game.scoring_button_1.flash_counter_2\[7\] game.scoring_button_1.flash_counter_2\[8\]
+ _1843_ VGND VGND VPWR VPWR _1847_ sky130_fd_sc_hd__and3_1
X_3713_ _0636_ _1066_ _1068_ VGND VGND VPWR VPWR _1069_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3644_ _0214_ _0928_ _1000_ _0949_ VGND VGND VPWR VPWR _1002_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3575_ _0909_ _0936_ _0917_ VGND VGND VPWR VPWR _0937_ sky130_fd_sc_hd__a21oi_1
X_5314_ _2297_ _2396_ _2274_ VGND VGND VPWR VPWR _2397_ sky130_fd_sc_hd__mux2_1
X_5245_ _2195_ _2315_ _2330_ _0214_ VGND VGND VPWR VPWR disp_song.um.drum.next_d1\[2\]
+ sky130_fd_sc_hd__o211a_1
Xhold28 game.out\[2\] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__dlygate4sd3_1
Xhold17 game.scoring_button_2.check_hit.in VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold39 game.scoring_button_1.next_flash_counter_1\[1\] VGND VGND VPWR VPWR net112
+ sky130_fd_sc_hd__dlygate4sd3_1
X_5176_ disp_song.note1\[24\] _2232_ _2256_ VGND VGND VPWR VPWR _2263_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_98_608 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4127_ _1420_ VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__buf_1
XFILLER_0_78_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4058_ _1361_ _1362_ _1363_ VGND VGND VPWR VPWR _1364_ sky130_fd_sc_hd__a21boi_1
X_3009_ _2654_ _0389_ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_54_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_54_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_96_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3360_ _0711_ _0721_ _0722_ VGND VGND VPWR VPWR _0723_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_0_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5030_ _2037_ _2121_ disp_song.um.drum.next_idx2\[2\] VGND VGND VPWR VPWR _2122_
+ sky130_fd_sc_hd__mux2_1
X_3291_ _0628_ _0650_ _0653_ VGND VGND VPWR VPWR _0654_ sky130_fd_sc_hd__and3_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5932_ clknet_leaf_61_clk game.scoring_button_1.next_flash_counter_1\[0\] net53 VGND
+ VGND VPWR VPWR game.scoring_button_1.flash_counter_1\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_73_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_45_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_45_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_48_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5863_ clknet_leaf_65_clk game.scoring_button_1.next_num_hits\[12\] net47 VGND VGND
+ VPWR VPWR game.addhits.a\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5794_ clknet_leaf_53_clk game.scoring_button_2.next_flash_counter_1\[8\] net52 VGND
+ VGND VPWR VPWR game.scoring_button_2.flash_counter_1\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4814_ _1931_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_1\[21\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4745_ net111 game.scoring_button_1.flash_counter_1\[0\] game.hit_1 VGND VGND VPWR
+ VPWR _1883_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4676_ _1835_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_2\[2\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3627_ _0849_ _0850_ _0855_ net39 VGND VGND VPWR VPWR _0986_ sky130_fd_sc_hd__o211a_1
XFILLER_0_31_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput29 net29 VGND VGND VPWR VPWR ss1[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput18 net18 VGND VGND VPWR VPWR ss0[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3558_ modetrans.mode\[3\] VGND VGND VPWR VPWR _0921_ sky130_fd_sc_hd__inv_2
XFILLER_0_101_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3489_ _0813_ _0851_ _0775_ _0831_ _0844_ VGND VGND VPWR VPWR _0852_ sky130_fd_sc_hd__a2111oi_1
X_5228_ _2313_ VGND VGND VPWR VPWR _2314_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5159_ _0175_ _0191_ _0198_ VGND VGND VPWR VPWR _2246_ sky130_fd_sc_hd__and3_2
Xclkbuf_leaf_36_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_36_clk sky130_fd_sc_hd__clkbuf_16
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_27_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_27_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_84_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2860_ _0163_ _0265_ _0282_ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__or3_1
XFILLER_0_57_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2791_ lvls.level\[0\] lvls.level\[1\] VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__nor2b_2
XFILLER_0_104_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_649 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4530_ game.addmisses.a\[7\] _1720_ _1727_ _1722_ VGND VGND VPWR VPWR _1728_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4461_ net215 _1613_ _1667_ _1612_ VGND VGND VPWR VPWR game.scoring_button_1.next_num_hits\[13\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3412_ _0752_ _0773_ _0774_ VGND VGND VPWR VPWR _0775_ sky130_fd_sc_hd__a21o_1
X_6131_ clknet_leaf_19_clk disp_song.um.drum.next_note2\[11\] net63 VGND VGND VPWR
+ VPWR disp_song.note2\[11\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4392_ _1611_ VGND VGND VPWR VPWR _1612_ sky130_fd_sc_hd__buf_6
XFILLER_0_110_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3343_ _0492_ _0705_ VGND VGND VPWR VPWR _0706_ sky130_fd_sc_hd__xnor2_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6062_ clknet_leaf_12_clk _0018_ net58 VGND VGND VPWR VPWR game.counter\[18\] sky130_fd_sc_hd__dfrtp_4
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3274_ game.addhits.add1.b\[0\] game.addhits.a\[0\] VGND VGND VPWR VPWR _0637_ sky130_fd_sc_hd__or2_1
X_5013_ _2100_ VGND VGND VPWR VPWR _2105_ sky130_fd_sc_hd__inv_2
XFILLER_0_84_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5915_ clknet_leaf_17_clk game.scoring_button_1.next_count\[6\] net62 VGND VGND VPWR
+ VPWR game.scoring_button_1.counts\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5846_ clknet_leaf_71_clk game.scoring_button_1.next_num_misses\[11\] net46 VGND
+ VGND VPWR VPWR game.addmisses.a\[11\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_91_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2989_ _0367_ _0377_ _0378_ disp_song.note1\[5\] VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__a2bb2o_1
X_5777_ clknet_leaf_7_clk game.scoring_button_2.next_count\[14\] net59 VGND VGND VPWR
+ VPWR game.scoring_button_2.counts\[14\] sky130_fd_sc_hd__dfrtp_1
X_4728_ game.scoring_button_1.flash_counter_2\[18\] _1868_ VGND VGND VPWR VPWR _1872_
+ sky130_fd_sc_hd__or2_1
X_4659_ game.scoring_button_1.flash_counter_2\[5\] game.scoring_button_1.flash_counter_2\[4\]
+ game.scoring_button_1.flash_counter_2\[7\] game.scoring_button_1.flash_counter_2\[6\]
+ VGND VGND VPWR VPWR _1823_ sky130_fd_sc_hd__or4b_1
XFILLER_0_71_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3961_ game.addhits.add4.b\[3\] _1278_ VGND VGND VPWR VPWR _1279_ sky130_fd_sc_hd__nand2_1
X_2912_ _0269_ disp_song.note2\[18\] _0321_ VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5700_ clknet_leaf_62_clk _0036_ net53 VGND VGND VPWR VPWR highest_score.highest_score\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_3892_ _0933_ net3 VGND VGND VPWR VPWR _1224_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2843_ disp_song.um.idx_note2\[1\] disp_song.um.idx_note2\[2\] disp_song.um.idx_note2\[0\]
+ VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__or3b_2
X_5631_ game.flash_counter\[18\] game.flash_counter\[14\] game.flash_counter\[15\]
+ game.flash_counter\[19\] VGND VGND VPWR VPWR _2608_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_26_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5562_ _2566_ game.padded_notes1\[18\] _2472_ VGND VGND VPWR VPWR _2567_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2774_ modetrans.mode\[5\] _0208_ _0211_ _0203_ VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__o31a_1
XFILLER_0_5_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4513_ game.addmisses.a\[4\] _1697_ VGND VGND VPWR VPWR _1713_ sky130_fd_sc_hd__and2_1
XFILLER_0_41_522 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5493_ _2525_ net234 _2515_ VGND VGND VPWR VPWR _2526_ sky130_fd_sc_hd__mux2_1
Xhold125 game.addhits.add3.b\[2\] VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__dlygate4sd3_1
Xhold103 game.scoring_button_2.flash_counter_1\[4\] VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__dlygate4sd3_1
Xhold114 game.flash_counter\[8\] VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__dlygate4sd3_1
Xhold158 game.padded_notes2\[14\] VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 game.padded_notes2\[8\] VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_7_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_7_clk sky130_fd_sc_hd__clkbuf_16
X_4444_ _1652_ _1653_ _1654_ VGND VGND VPWR VPWR _1655_ sky130_fd_sc_hd__o21ai_1
Xhold147 game.addhits.a\[7\] VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__dlygate4sd3_1
Xhold169 game.padded_notes2\[2\] VGND VGND VPWR VPWR net242 sky130_fd_sc_hd__dlygate4sd3_1
X_4375_ game.scoring_button_2.flash_counter_1\[18\] _1597_ VGND VGND VPWR VPWR _1600_
+ sky130_fd_sc_hd__and2_1
X_6114_ clknet_leaf_39_clk disp_song.um.drum.next_note1\[26\] net66 VGND VGND VPWR
+ VPWR disp_song.note1\[26\] sky130_fd_sc_hd__dfstp_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3326_ _0686_ _0687_ VGND VGND VPWR VPWR _0689_ sky130_fd_sc_hd__or2_1
X_6045_ clknet_leaf_16_clk _0020_ net62 VGND VGND VPWR VPWR game.counter\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3257_ _0608_ _0619_ VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__nand2_1
X_3188_ _0549_ _0550_ VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__and2b_1
XFILLER_0_49_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5829_ clknet_leaf_52_clk game.scoring_button_2.next_flash_counter_2\[20\] net55
+ VGND VGND VPWR VPWR game.scoring_button_2.flash_counter_2\[20\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_522 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_216 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4160_ game.counter\[11\] _1439_ VGND VGND VPWR VPWR _1443_ sky130_fd_sc_hd__nand2_2
XFILLER_0_4_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3111_ game.addmisses.a\[6\] game.addmisses.add2.b\[2\] VGND VGND VPWR VPWR _0474_
+ sky130_fd_sc_hd__nand2_1
X_4091_ _1289_ _1390_ _1391_ _1392_ VGND VGND VPWR VPWR game.scoring_button_2.next_num_misses\[13\]
+ sky130_fd_sc_hd__o22a_1
X_3042_ _0375_ _0410_ _0416_ VGND VGND VPWR VPWR disp_song.um.drum.next_note1\[20\]
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_65_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4993_ _0162_ _2085_ VGND VGND VPWR VPWR _2086_ sky130_fd_sc_hd__or2_1
XFILLER_0_81_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3944_ game.addhits.add3.b\[1\] _1264_ VGND VGND VPWR VPWR _1266_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3875_ _0966_ disp_song.display_note2\[2\] _0211_ game.out\[2\] _0208_ VGND VGND
+ VPWR VPWR _1213_ sky130_fd_sc_hd__a221o_1
XFILLER_0_18_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5614_ _2595_ net100 VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__nor2_1
X_2826_ _0255_ _2659_ VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5545_ _2555_ VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__clkbuf_1
X_2757_ _0179_ _0171_ VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_30_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5476_ disp_song.note2\[25\] game.padded_notes2\[24\] _2497_ VGND VGND VPWR VPWR
+ _2514_ sky130_fd_sc_hd__mux2_1
X_2688_ _2657_ _2660_ _2661_ VGND VGND VPWR VPWR _2662_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_76_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4427_ game.addhits.a\[5\] _1613_ _1641_ _1612_ VGND VGND VPWR VPWR game.scoring_button_1.next_num_hits\[5\]
+ sky130_fd_sc_hd__a22o_1
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4358_ _1588_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_1\[12\]
+ sky130_fd_sc_hd__clkbuf_1
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3309_ _0667_ _0668_ _0671_ VGND VGND VPWR VPWR _0672_ sky130_fd_sc_hd__o21ai_1
X_4289_ _1539_ _1486_ _1540_ VGND VGND VPWR VPWR _1541_ sky130_fd_sc_hd__and3b_1
X_6028_ clknet_leaf_59_clk _0137_ net51 VGND VGND VPWR VPWR game.flash_counter\[8\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_1415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout64 net65 VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__buf_6
XFILLER_0_36_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout53 net73 VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__buf_8
XFILLER_0_52_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_536 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3660_ _0787_ _1013_ VGND VGND VPWR VPWR _1016_ sky130_fd_sc_hd__or2_1
X_3591_ lvls.level\[1\] _0952_ modetrans.mode\[5\] VGND VGND VPWR VPWR _0953_ sky130_fd_sc_hd__o21a_2
X_5330_ _0209_ _2658_ _1302_ VGND VGND VPWR VPWR _2410_ sky130_fd_sc_hd__nand3_1
X_5261_ _2252_ _2323_ _2345_ _0197_ VGND VGND VPWR VPWR _2346_ sky130_fd_sc_hd__o22a_1
X_4212_ game.scoring_button_2.flash_counter_2\[1\] game.scoring_button_2.flash_counter_2\[0\]
+ game.scoring_button_2.flash_counter_2\[3\] game.scoring_button_2.flash_counter_2\[2\]
+ VGND VGND VPWR VPWR _1480_ sky130_fd_sc_hd__or4_1
X_5192_ _2247_ _2270_ _2275_ _2278_ VGND VGND VPWR VPWR _2279_ sky130_fd_sc_hd__o22a_1
X_4143_ _1428_ _1429_ VGND VGND VPWR VPWR _1430_ sky130_fd_sc_hd__nor2_1
X_4074_ _1369_ _1374_ _1376_ _1377_ _1289_ game.addmisses.add3.b\[3\] VGND VGND VPWR
+ VPWR _1378_ sky130_fd_sc_hd__mux4_1
X_3025_ disp_song.um.idx_note1\[4\] VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4976_ _2067_ _2069_ _2026_ VGND VGND VPWR VPWR _2070_ sky130_fd_sc_hd__mux2_1
X_3927_ game.addhits.add2.b\[2\] game.addhits.add2.b\[1\] _1251_ game.addhits.add2.b\[3\]
+ VGND VGND VPWR VPWR _1253_ sky130_fd_sc_hd__o31a_2
XFILLER_0_34_606 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3858_ _0933_ _1201_ VGND VGND VPWR VPWR _1202_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2809_ game.counter\[15\] VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3789_ _1037_ _1039_ _1130_ _1141_ net38 VGND VGND VPWR VPWR _1142_ sky130_fd_sc_hd__o311a_1
X_5528_ disp_song.note1\[7\] game.padded_notes1\[6\] _2541_ VGND VGND VPWR VPWR _2544_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5459_ _2502_ game.padded_notes2\[19\] _2473_ VGND VGND VPWR VPWR _2503_ sky130_fd_sc_hd__mux2_1
XTAP_1223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4830_ _1937_ VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4761_ game.scoring_button_1.flash_counter_1\[6\] _1891_ VGND VGND VPWR VPWR _1894_
+ sky130_fd_sc_hd__and2_1
X_4692_ net161 _1843_ _1846_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_2\[7\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_83_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3712_ _0641_ _1067_ VGND VGND VPWR VPWR _1068_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3643_ _0856_ _0991_ _1000_ _0211_ net39 VGND VGND VPWR VPWR _1001_ sky130_fd_sc_hd__o221a_1
XFILLER_0_102_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3574_ _0667_ _0912_ VGND VGND VPWR VPWR _0936_ sky130_fd_sc_hd__nor2_1
X_5313_ _2310_ _2394_ _2395_ _2254_ VGND VGND VPWR VPWR _2396_ sky130_fd_sc_hd__o22a_1
X_5244_ _2234_ _2322_ _2329_ VGND VGND VPWR VPWR _2330_ sky130_fd_sc_hd__or3_1
Xhold18 game.padded_notes2\[0\] VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 _0125_ VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__dlygate4sd3_1
X_5175_ disp_song.um.drum.next_note1\[25\] _2261_ _2185_ VGND VGND VPWR VPWR _2262_
+ sky130_fd_sc_hd__a21oi_1
X_4126_ _1418_ _1419_ VGND VGND VPWR VPWR _1420_ sky130_fd_sc_hd__and2b_1
X_4057_ game.addmisses.add3.b\[2\] _1362_ game.addmisses.add3.b\[3\] VGND VGND VPWR
+ VPWR _1363_ sky130_fd_sc_hd__o21a_1
X_3008_ _0363_ _0392_ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__nand2_1
XFILLER_0_66_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4959_ disp_song.note2\[8\] _1956_ VGND VGND VPWR VPWR _2053_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3290_ _0651_ _0652_ _0641_ VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__a21o_1
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_620 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5931_ clknet_leaf_13_clk game.scoring_button_1.next_count\[22\] net58 VGND VGND
+ VPWR VPWR game.scoring_button_1.counts\[22\] sky130_fd_sc_hd__dfrtp_1
X_5862_ clknet_leaf_65_clk game.scoring_button_1.next_num_hits\[11\] net47 VGND VGND
+ VPWR VPWR game.addhits.a\[11\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_75_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5793_ clknet_leaf_53_clk net193 net52 VGND VGND VPWR VPWR game.scoring_button_2.flash_counter_1\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_4813_ _1929_ game.hit_1 _1930_ VGND VGND VPWR VPWR _1931_ sky130_fd_sc_hd__and3b_1
X_4744_ _1882_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_1\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_83_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4675_ _1833_ game.missed_1 _1834_ VGND VGND VPWR VPWR _1835_ sky130_fd_sc_hd__and3b_1
XFILLER_0_98_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3626_ _0258_ _0982_ _0984_ _0941_ VGND VGND VPWR VPWR _0985_ sky130_fd_sc_hd__a2bb2o_1
Xoutput19 net19 VGND VGND VPWR VPWR ss0[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3557_ _0916_ _0919_ _0261_ VGND VGND VPWR VPWR _0920_ sky130_fd_sc_hd__o21ai_1
X_3488_ _0808_ _0812_ VGND VGND VPWR VPWR _0851_ sky130_fd_sc_hd__nand2_1
X_5227_ disp_song.um.drum.next_idx1\[4\] _0191_ disp_song.um.drum.next_idx1\[3\] _2244_
+ VGND VGND VPWR VPWR _2313_ sky130_fd_sc_hd__or4b_1
X_5158_ _0191_ _2244_ VGND VGND VPWR VPWR _2245_ sky130_fd_sc_hd__nor2_1
X_5089_ _2091_ _2177_ _0169_ VGND VGND VPWR VPWR _2178_ sky130_fd_sc_hd__mux2_1
X_4109_ game.scoring_button_2.flash_counter_1\[13\] game.scoring_button_2.flash_counter_1\[12\]
+ game.scoring_button_2.flash_counter_1\[15\] game.scoring_button_2.flash_counter_1\[14\]
+ VGND VGND VPWR VPWR _1408_ sky130_fd_sc_hd__or4b_1
XFILLER_0_94_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_104_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2790_ _0221_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4460_ _1663_ _1665_ _1666_ VGND VGND VPWR VPWR _1667_ sky130_fd_sc_hd__o21ai_1
X_3411_ _0762_ VGND VGND VPWR VPWR _0774_ sky130_fd_sc_hd__inv_2
XFILLER_0_40_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4391_ game.scoring_button_1.check_hit.edge_1 game.scoring_button_1.check_hit.edge_2
+ game.scoring_button_1.hit VGND VGND VPWR VPWR _1611_ sky130_fd_sc_hd__and3b_1
X_6130_ clknet_leaf_19_clk disp_song.um.drum.next_note2\[10\] net63 VGND VGND VPWR
+ VPWR disp_song.note2\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3342_ _0487_ _0500_ VGND VGND VPWR VPWR _0705_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6061_ clknet_leaf_12_clk _0017_ net58 VGND VGND VPWR VPWR game.counter\[17\] sky130_fd_sc_hd__dfrtp_2
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3273_ _0450_ _0635_ VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__nand2_2
X_5012_ disp_song.um.drum.next_idx2\[0\] _1965_ _2054_ _2043_ VGND VGND VPWR VPWR
+ _2104_ sky130_fd_sc_hd__o211a_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5914_ clknet_leaf_15_clk game.scoring_button_1.next_count\[5\] net62 VGND VGND VPWR
+ VPWR game.scoring_button_1.counts\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5845_ clknet_leaf_71_clk game.scoring_button_1.next_num_misses\[10\] net46 VGND
+ VGND VPWR VPWR game.addmisses.a\[10\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_63_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2988_ _0368_ _0377_ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__or2_1
X_5776_ clknet_leaf_7_clk game.scoring_button_2.next_count\[13\] net59 VGND VGND VPWR
+ VPWR game.scoring_button_2.counts\[13\] sky130_fd_sc_hd__dfrtp_1
X_4727_ game.scoring_button_1.flash_counter_2\[18\] _1868_ VGND VGND VPWR VPWR _1871_
+ sky130_fd_sc_hd__and2_1
X_4658_ _1822_ VGND VGND VPWR VPWR game.scoring_button_1.next_count\[22\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3609_ _0617_ _0609_ _0614_ VGND VGND VPWR VPWR _0969_ sky130_fd_sc_hd__or3_1
XFILLER_0_31_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4589_ _1767_ _1771_ VGND VGND VPWR VPWR _1779_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_98_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3960_ game.addhits.add4.b\[1\] _1275_ VGND VGND VPWR VPWR _1278_ sky130_fd_sc_hd__xnor2_1
X_2911_ disp_song.um.idx_note2\[3\] _0318_ _0160_ _0276_ VGND VGND VPWR VPWR _0321_
+ sky130_fd_sc_hd__or4_1
XFILLER_0_70_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3891_ _1223_ VGND VGND VPWR VPWR modetrans.pushed_4 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2842_ _2657_ VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__clkbuf_8
X_5630_ game.flash_counter\[13\] game.flash_counter\[11\] game.flash_counter\[10\]
+ game.flash_counter\[12\] VGND VGND VPWR VPWR _2607_ sky130_fd_sc_hd__or4bb_1
X_5561_ disp_song.note1\[18\] game.padded_notes1\[17\] _2541_ VGND VGND VPWR VPWR
+ _2566_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2773_ _0210_ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__buf_8
X_5492_ disp_song.note2\[30\] game.padded_notes2\[29\] _2497_ VGND VGND VPWR VPWR
+ _2525_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4512_ game.addmisses.a\[4\] _1697_ VGND VGND VPWR VPWR _1712_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold104 game.scoring_button_1.flash_counter_2\[4\] VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__dlygate4sd3_1
Xhold126 game.counter\[2\] VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_77 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold115 game.addhits.add2.b\[0\] VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold148 game.padded_notes2\[24\] VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__dlygate4sd3_1
Xhold159 game.padded_notes1\[1\] VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__dlygate4sd3_1
Xhold137 game.padded_notes1\[24\] VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__dlygate4sd3_1
X_4443_ game.addhits.a\[10\] game.addhits.a\[9\] _1650_ game.addhits.a\[11\] VGND
+ VGND VPWR VPWR _1654_ sky130_fd_sc_hd__o31a_1
XFILLER_0_111_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4374_ _1599_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_1\[17\]
+ sky130_fd_sc_hd__clkbuf_1
X_6113_ clknet_leaf_40_clk disp_song.um.drum.next_note1\[25\] net66 VGND VGND VPWR
+ VPWR disp_song.note1\[25\] sky130_fd_sc_hd__dfrtp_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3325_ _0686_ _0687_ VGND VGND VPWR VPWR _0688_ sky130_fd_sc_hd__and2_1
X_6044_ clknet_leaf_13_clk _0009_ net58 VGND VGND VPWR VPWR game.counter\[0\] sky130_fd_sc_hd__dfrtp_2
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3256_ _0609_ _0614_ _0615_ _0618_ VGND VGND VPWR VPWR _0619_ sky130_fd_sc_hd__o211a_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3187_ game.addhits.a\[2\] game.addhits.add1.b\[2\] VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5828_ clknet_leaf_50_clk game.scoring_button_2.next_flash_counter_2\[19\] net56
+ VGND VGND VPWR VPWR game.scoring_button_2.flash_counter_2\[19\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5759_ clknet_leaf_64_clk game.scoring_button_2.next_num_hits\[15\] net47 VGND VGND
+ VPWR VPWR game.addhits.add4.b\[3\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_32_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3110_ game.addmisses.a\[6\] game.addmisses.add2.b\[2\] VGND VGND VPWR VPWR _0473_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4090_ game.addmisses.add4.b\[1\] _1383_ _1289_ VGND VGND VPWR VPWR _1392_ sky130_fd_sc_hd__o21ai_1
X_3041_ _0375_ _0412_ net163 VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__o21ai_1
X_4992_ _2677_ _0169_ VGND VGND VPWR VPWR _2085_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3943_ _1264_ _1265_ net249 _1227_ VGND VGND VPWR VPWR game.scoring_button_2.next_num_hits\[8\]
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_46_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_626 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3874_ _1212_ VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5613_ game.flash_counter\[0\] _0842_ net99 VGND VGND VPWR VPWR _2596_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_3_2__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_2825_ highest_score.score_mode\[0\] VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__clkbuf_8
X_5544_ _2554_ net241 _2515_ VGND VGND VPWR VPWR _2555_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2756_ _0197_ VGND VGND VPWR VPWR disp_song.um.drum.next_idx1\[3\] sky130_fd_sc_hd__inv_2
X_5475_ _2513_ VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__clkbuf_1
X_2687_ disp_song.toggle_state VGND VGND VPWR VPWR _2661_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4426_ _1639_ _1640_ VGND VGND VPWR VPWR _1641_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4357_ _1586_ game.hit_2 _1587_ VGND VGND VPWR VPWR _1588_ sky130_fd_sc_hd__and3b_1
XFILLER_0_39_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4288_ game.scoring_button_2.flash_counter_2\[13\] game.scoring_button_2.flash_counter_2\[12\]
+ _1532_ game.scoring_button_2.flash_counter_2\[14\] VGND VGND VPWR VPWR _1540_ sky130_fd_sc_hd__a31o_1
X_3308_ _0669_ _0670_ VGND VGND VPWR VPWR _0671_ sky130_fd_sc_hd__or2_2
X_6027_ clknet_leaf_59_clk _0136_ net50 VGND VGND VPWR VPWR game.flash_counter\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3239_ _0537_ _0576_ _0577_ VGND VGND VPWR VPWR _0602_ sky130_fd_sc_hd__and3_1
XTAP_1405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout65 net73 VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__buf_6
XFILLER_0_9_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout54 net73 VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__buf_4
XFILLER_0_51_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3590_ lvls.level\[2\] lvls.level\[0\] VGND VGND VPWR VPWR _0952_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5260_ disp_song.um.drum.next_idx1\[2\] _2252_ VGND VGND VPWR VPWR _2345_ sky130_fd_sc_hd__nor2_1
X_4211_ game.scoring_button_2.flash_counter_2\[5\] game.scoring_button_2.flash_counter_2\[4\]
+ game.scoring_button_2.flash_counter_2\[7\] game.scoring_button_2.flash_counter_2\[6\]
+ VGND VGND VPWR VPWR _1479_ sky130_fd_sc_hd__or4b_1
X_5191_ _2256_ _2277_ VGND VGND VPWR VPWR _2278_ sky130_fd_sc_hd__nor2_1
X_4142_ game.counter\[6\] game.counter\[7\] _1423_ VGND VGND VPWR VPWR _1429_ sky130_fd_sc_hd__and3_1
X_4073_ _1358_ _1374_ VGND VGND VPWR VPWR _1377_ sky130_fd_sc_hd__nor2_1
X_3024_ _0380_ _0402_ _0403_ net237 VGND VGND VPWR VPWR disp_song.um.drum.next_note1\[15\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4975_ _2038_ _2068_ disp_song.note2\[4\] disp_song.um.drum.next_idx2\[0\] VGND VGND
+ VPWR VPWR _2069_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_19_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3926_ _1226_ _1250_ _1252_ _1227_ net188 VGND VGND VPWR VPWR game.scoring_button_2.next_num_hits\[4\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_34_618 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3857_ _0966_ disp_song.display_note1\[3\] _0211_ game.out\[10\] _0208_ VGND VGND
+ VPWR VPWR _1201_ sky130_fd_sc_hd__a221o_2
XFILLER_0_46_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2808_ game.counter\[9\] _0237_ game.counter\[15\] _0227_ _0238_ VGND VGND VPWR VPWR
+ _0239_ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3788_ _0210_ _1140_ VGND VGND VPWR VPWR _1141_ sky130_fd_sc_hd__or2_1
X_5527_ _2543_ VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__clkbuf_1
X_2739_ disp_song.um.idx_note1\[4\] _0182_ VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__or2_1
X_5458_ disp_song.note2\[19\] game.padded_notes2\[18\] _2497_ VGND VGND VPWR VPWR
+ _2502_ sky130_fd_sc_hd__mux2_1
X_5389_ _2455_ VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__clkbuf_1
X_4409_ _1627_ VGND VGND VPWR VPWR _1628_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_14 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4760_ _1893_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_1\[5\]
+ sky130_fd_sc_hd__clkbuf_1
X_4691_ net161 _1843_ game.missed_1 VGND VGND VPWR VPWR _1846_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_15_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3711_ _0633_ _1064_ _0912_ VGND VGND VPWR VPWR _1067_ sky130_fd_sc_hd__or3_1
XFILLER_0_55_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3642_ _0999_ VGND VGND VPWR VPWR _1000_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5312_ disp_song.note1\[1\] _2185_ disp_song.um.drum.next_note1\[0\] _2232_ VGND
+ VGND VPWR VPWR _2395_ sky130_fd_sc_hd__o22a_1
XFILLER_0_11_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3573_ _0924_ _0931_ _0932_ _0935_ VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__o31a_1
XFILLER_0_51_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5243_ disp_song.um.drum.next_idx1\[4\] _2323_ _2328_ VGND VGND VPWR VPWR _2329_
+ sky130_fd_sc_hd__a21boi_1
Xhold19 _0050_ VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__dlygate4sd3_1
X_5174_ _2258_ VGND VGND VPWR VPWR _2261_ sky130_fd_sc_hd__inv_2
X_4125_ game.counter\[1\] game.counter\[0\] game.counter\[2\] game.counter\[3\] VGND
+ VGND VPWR VPWR _1419_ sky130_fd_sc_hd__a31o_1
XFILLER_0_78_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4056_ game.addmisses.add3.b\[1\] _1355_ VGND VGND VPWR VPWR _1362_ sky130_fd_sc_hd__or2_1
X_3007_ _2661_ _0352_ _0194_ _0359_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__nor4_1
XFILLER_0_66_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4958_ disp_song.um.drum.next_note2\[9\] _2029_ _2666_ VGND VGND VPWR VPWR _2052_
+ sky130_fd_sc_hd__a21oi_1
X_4889_ _1972_ _1981_ _1983_ VGND VGND VPWR VPWR _1984_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3909_ _1233_ _1238_ VGND VGND VPWR VPWR _1239_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_632 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5930_ clknet_leaf_13_clk game.scoring_button_1.next_count\[21\] net58 VGND VGND
+ VPWR VPWR game.scoring_button_1.counts\[21\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5861_ clknet_leaf_65_clk game.scoring_button_1.next_num_hits\[10\] net47 VGND VGND
+ VPWR VPWR game.addhits.a\[10\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_8_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5792_ clknet_leaf_55_clk game.scoring_button_2.next_flash_counter_1\[6\] net52 VGND
+ VGND VPWR VPWR game.scoring_button_2.flash_counter_1\[6\] sky130_fd_sc_hd__dfrtp_1
X_4812_ game.scoring_button_1.flash_counter_1\[21\] _1926_ VGND VGND VPWR VPWR _1930_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_7_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4743_ game.scoring_button_1.flash_counter_1\[0\] _1799_ VGND VGND VPWR VPWR _1882_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_71_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4674_ game.scoring_button_1.flash_counter_2\[1\] game.scoring_button_1.flash_counter_2\[0\]
+ game.scoring_button_1.flash_counter_2\[2\] VGND VGND VPWR VPWR _1834_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3625_ _0893_ _0959_ _0983_ VGND VGND VPWR VPWR _0984_ sky130_fd_sc_hd__or3_1
XFILLER_0_11_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3556_ _0913_ _0917_ _0918_ VGND VGND VPWR VPWR _0919_ sky130_fd_sc_hd__a21oi_1
X_5226_ _2311_ VGND VGND VPWR VPWR _2312_ sky130_fd_sc_hd__inv_2
X_3487_ _0841_ _0847_ _0835_ VGND VGND VPWR VPWR _0850_ sky130_fd_sc_hd__and3_1
XFILLER_0_51_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5157_ _2243_ VGND VGND VPWR VPWR _2244_ sky130_fd_sc_hd__buf_2
X_5088_ disp_song.um.drum.next_idx2\[1\] _1966_ _2089_ VGND VGND VPWR VPWR _2177_
+ sky130_fd_sc_hd__a21o_1
X_4108_ game.scoring_button_2.flash_counter_1\[1\] game.scoring_button_2.flash_counter_1\[0\]
+ game.scoring_button_2.flash_counter_1\[3\] game.scoring_button_2.flash_counter_1\[2\]
+ VGND VGND VPWR VPWR _1407_ sky130_fd_sc_hd__or4_1
X_4039_ _1343_ _1347_ _1289_ VGND VGND VPWR VPWR _1348_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3410_ _0763_ _0771_ _0772_ VGND VGND VPWR VPWR _0773_ sky130_fd_sc_hd__a21o_1
X_4390_ net89 _1607_ _1610_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_1\[22\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3341_ _0585_ _0592_ _0703_ _0584_ VGND VGND VPWR VPWR _0704_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6060_ clknet_leaf_12_clk _0016_ net58 VGND VGND VPWR VPWR game.counter\[16\] sky130_fd_sc_hd__dfrtp_4
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3272_ game.addmisses.add1.b\[0\] game.addmisses.a\[0\] VGND VGND VPWR VPWR _0635_
+ sky130_fd_sc_hd__or2_1
X_5011_ _2053_ _2102_ VGND VGND VPWR VPWR _2103_ sky130_fd_sc_hd__nor2_1
XFILLER_0_84_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5913_ clknet_leaf_15_clk game.scoring_button_1.next_count\[4\] net62 VGND VGND VPWR
+ VPWR game.scoring_button_1.counts\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5844_ clknet_leaf_70_clk game.scoring_button_1.next_num_misses\[9\] net46 VGND VGND
+ VPWR VPWR game.addmisses.a\[9\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_29_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2987_ disp_song.um.idx_note1\[3\] _0179_ disp_song.um.idx_note1\[0\] disp_song.um.idx_note1\[2\]
+ VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__or4bb_2
X_5775_ clknet_leaf_7_clk game.scoring_button_2.next_count\[12\] net59 VGND VGND VPWR
+ VPWR game.scoring_button_2.counts\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4726_ _1870_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_2\[17\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4657_ game.scoring_button_1.check_hit.in _1477_ VGND VGND VPWR VPWR _1822_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3608_ _0849_ _0855_ _0856_ _0861_ VGND VGND VPWR VPWR _0968_ sky130_fd_sc_hd__a211o_1
XFILLER_0_101_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4588_ _1675_ _1776_ _1777_ _1778_ VGND VGND VPWR VPWR game.scoring_button_1.next_num_misses\[13\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_101_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3539_ _0898_ _0900_ _0901_ VGND VGND VPWR VPWR _0902_ sky130_fd_sc_hd__o21a_1
X_5209_ _2232_ disp_song.um.drum.next_note1\[7\] _2191_ _2268_ disp_song.um.drum.next_note1\[6\]
+ VGND VGND VPWR VPWR _2296_ sky130_fd_sc_hd__a32o_1
XFILLER_0_79_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_565 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2910_ _0320_ VGND VGND VPWR VPWR disp_song.um.drum.next_note2\[17\] sky130_fd_sc_hd__clkbuf_1
X_3890_ _0933_ net4 VGND VGND VPWR VPWR _1223_ sky130_fd_sc_hd__and2_1
XFILLER_0_70_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2841_ _0268_ VGND VGND VPWR VPWR disp_song.um.drum.next_note2\[0\] sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_73_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5560_ _2565_ VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__clkbuf_1
X_2772_ _0209_ modetrans.mode\[4\] VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__or2_4
X_5491_ _2524_ VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4511_ _1709_ _1710_ _1711_ _1675_ VGND VGND VPWR VPWR game.scoring_button_1.next_num_misses\[3\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4442_ game.addhits.a\[9\] game.addhits.a\[8\] _1639_ VGND VGND VPWR VPWR _1653_
+ sky130_fd_sc_hd__and3_1
Xhold116 game.addhits.a\[12\] VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__dlygate4sd3_1
Xhold105 game.addhits.add1.b\[3\] VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold138 game.padded_notes2\[22\] VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__dlygate4sd3_1
Xhold127 disp_song.note2\[30\] VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_79_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold149 game.padded_notes1\[20\] VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4373_ _1597_ _1413_ _1598_ VGND VGND VPWR VPWR _1599_ sky130_fd_sc_hd__and3b_1
XFILLER_0_21_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6112_ clknet_leaf_41_clk disp_song.um.drum.next_note1\[24\] net67 VGND VGND VPWR
+ VPWR disp_song.note1\[24\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3324_ _0617_ _0615_ VGND VGND VPWR VPWR _0687_ sky130_fd_sc_hd__nor2_1
X_6043_ clknet_leaf_58_clk _0152_ net50 VGND VGND VPWR VPWR game.flash_counter\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3255_ _0617_ VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__inv_2
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3186_ game.addhits.a\[2\] game.addhits.add1.b\[2\] VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_123 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5827_ clknet_leaf_50_clk game.scoring_button_2.next_flash_counter_2\[18\] net56
+ VGND VGND VPWR VPWR game.scoring_button_2.flash_counter_2\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5758_ clknet_leaf_65_clk game.scoring_button_2.next_num_hits\[14\] net47 VGND VGND
+ VPWR VPWR game.addhits.add4.b\[2\] sky130_fd_sc_hd__dfrtp_2
X_4709_ _1857_ game.missed_1 _1858_ VGND VGND VPWR VPWR _1859_ sky130_fd_sc_hd__and3b_1
X_5689_ _2649_ VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3040_ _0415_ VGND VGND VPWR VPWR disp_song.um.drum.next_note1\[19\] sky130_fd_sc_hd__inv_2
X_4991_ _0169_ _2080_ _2083_ VGND VGND VPWR VPWR _2084_ sky130_fd_sc_hd__o21ai_1
X_3942_ game.addhits.add3.b\[0\] _1253_ _1226_ VGND VGND VPWR VPWR _1265_ sky130_fd_sc_hd__o21ai_1
X_3873_ _0933_ _1211_ VGND VGND VPWR VPWR _1212_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2824_ _0232_ _0254_ VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__nor2_4
X_5612_ _2594_ VGND VGND VPWR VPWR _2595_ sky130_fd_sc_hd__clkbuf_2
X_5543_ disp_song.note1\[12\] game.padded_notes1\[11\] _2541_ VGND VGND VPWR VPWR
+ _2554_ sky130_fd_sc_hd__mux2_1
X_2755_ _0196_ VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__buf_4
XFILLER_0_5_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5474_ _2512_ net221 _2473_ VGND VGND VPWR VPWR _2513_ sky130_fd_sc_hd__mux2_1
X_2686_ _2658_ _2659_ VGND VGND VPWR VPWR _2660_ sky130_fd_sc_hd__nor2_4
XFILLER_0_41_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4425_ game.addhits.a\[5\] _1637_ VGND VGND VPWR VPWR _1640_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4356_ game.scoring_button_2.flash_counter_1\[12\] _1583_ VGND VGND VPWR VPWR _1587_
+ sky130_fd_sc_hd__or2_1
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3307_ _0560_ _0561_ _0543_ VGND VGND VPWR VPWR _0670_ sky130_fd_sc_hd__a21oi_1
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4287_ game.scoring_button_2.flash_counter_2\[13\] game.scoring_button_2.flash_counter_2\[14\]
+ _1535_ VGND VGND VPWR VPWR _1539_ sky130_fd_sc_hd__and3_1
X_6026_ clknet_leaf_58_clk _0135_ net50 VGND VGND VPWR VPWR game.flash_counter\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3238_ _0492_ _0598_ _0600_ VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__a21boi_1
X_3169_ game.addhits.a\[9\] game.addhits.add3.b\[1\] VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__nand2_1
XTAP_1406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout55 net56 VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__buf_6
XFILLER_0_91_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout66 net73 VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__buf_6
XFILLER_0_9_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4210_ _1478_ VGND VGND VPWR VPWR game.scoring_button_2.next_count\[22\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5190_ disp_song.note1\[18\] _2232_ _2276_ VGND VGND VPWR VPWR _2277_ sky130_fd_sc_hd__o21ai_1
X_4141_ game.counter\[6\] _1423_ game.counter\[7\] VGND VGND VPWR VPWR _1428_ sky130_fd_sc_hd__a21oi_1
X_4072_ game.addmisses.add3.b\[2\] _1362_ VGND VGND VPWR VPWR _1376_ sky130_fd_sc_hd__nor2_1
X_3023_ _0382_ _0402_ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__nand2_1
X_4974_ _1956_ disp_song.um.drum.next_note2\[5\] VGND VGND VPWR VPWR _2068_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3925_ _1251_ VGND VGND VPWR VPWR _1252_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3856_ _1200_ VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2807_ game.counter\[5\] game.counter\[13\] game.counter\[12\] _0209_ VGND VGND VPWR
+ VPWR _0238_ sky130_fd_sc_hd__or4b_1
XFILLER_0_6_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3787_ _0921_ _1139_ VGND VGND VPWR VPWR _1140_ sky130_fd_sc_hd__nor2_1
X_5526_ _2542_ game.padded_notes1\[6\] _2515_ VGND VGND VPWR VPWR _2543_ sky130_fd_sc_hd__mux2_1
X_2738_ _0177_ _0181_ VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5457_ _2501_ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__clkbuf_1
X_4408_ _1623_ _1626_ VGND VGND VPWR VPWR _1627_ sky130_fd_sc_hd__nand2_1
X_5388_ _0206_ _2452_ _2454_ VGND VGND VPWR VPWR _2455_ sky130_fd_sc_hd__and3_1
XFILLER_0_10_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4339_ game.scoring_button_2.flash_counter_1\[7\] _1572_ game.hit_2 VGND VGND VPWR
+ VPWR _1575_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_5_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6009_ clknet_leaf_49_clk _0118_ net56 VGND VGND VPWR VPWR game.padded_notes1\[28\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_66_clk clknet_3_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_66_clk sky130_fd_sc_hd__clkbuf_16
XTAP_1214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_57_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_57_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_87_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_608 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3710_ _0629_ _1065_ VGND VGND VPWR VPWR _1066_ sky130_fd_sc_hd__or2_1
X_4690_ _1845_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_2\[6\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_43_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3641_ modetrans.mode\[3\] _0998_ VGND VGND VPWR VPWR _0999_ sky130_fd_sc_hd__nand2_1
XFILLER_0_102_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3572_ _0934_ VGND VGND VPWR VPWR _0935_ sky130_fd_sc_hd__buf_4
X_5311_ disp_song.note1\[2\] _2232_ disp_song.um.drum.next_idx1\[1\] _2209_ VGND VGND
+ VPWR VPWR _2394_ sky130_fd_sc_hd__o22a_1
XFILLER_0_11_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5242_ _2324_ _2325_ _2326_ _2327_ disp_song.um.drum.next_idx1\[2\] _0197_ VGND VGND
+ VPWR VPWR _2328_ sky130_fd_sc_hd__mux4_1
X_5173_ disp_song.note1\[26\] _2232_ _2259_ VGND VGND VPWR VPWR _2260_ sky130_fd_sc_hd__o21ai_1
X_4124_ game.counter\[1\] game.counter\[0\] game.counter\[3\] game.counter\[2\] VGND
+ VGND VPWR VPWR _1418_ sky130_fd_sc_hd__and4_1
Xinput1 button[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__clkbuf_1
X_4055_ game.addmisses.add3.b\[1\] _1355_ VGND VGND VPWR VPWR _1361_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_48_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_48_clk sky130_fd_sc_hd__clkbuf_16
X_3006_ _0391_ VGND VGND VPWR VPWR disp_song.um.drum.next_note1\[9\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_108_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4957_ _2022_ _2033_ _2050_ _2032_ VGND VGND VPWR VPWR _2051_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_74_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4888_ _1948_ _1982_ VGND VGND VPWR VPWR _1983_ sky130_fd_sc_hd__nor2_4
XFILLER_0_34_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3908_ game.addhits.add1.b\[2\] game.scoring_button_2.acc\[2\] VGND VGND VPWR VPWR
+ _1238_ sky130_fd_sc_hd__or2_1
X_3839_ _0259_ _1183_ VGND VGND VPWR VPWR _1189_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5509_ disp_song.note1\[1\] game.padded_notes1\[0\] _2497_ VGND VGND VPWR VPWR _2531_
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_39_clk clknet_3_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_39_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_96_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_530 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5860_ clknet_leaf_65_clk game.scoring_button_1.next_num_hits\[9\] net47 VGND VGND
+ VPWR VPWR game.addhits.a\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4811_ game.scoring_button_1.flash_counter_1\[21\] _1926_ VGND VGND VPWR VPWR _1929_
+ sky130_fd_sc_hd__and2_1
X_5791_ clknet_leaf_54_clk game.scoring_button_2.next_flash_counter_1\[5\] net52 VGND
+ VGND VPWR VPWR game.scoring_button_2.flash_counter_1\[5\] sky130_fd_sc_hd__dfrtp_1
X_4742_ net86 _1878_ _1881_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_2\[22\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4673_ game.scoring_button_1.flash_counter_2\[1\] game.scoring_button_1.flash_counter_2\[0\]
+ game.scoring_button_1.flash_counter_2\[2\] VGND VGND VPWR VPWR _1833_ sky130_fd_sc_hd__and3_1
XFILLER_0_83_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3624_ _0887_ _0939_ VGND VGND VPWR VPWR _0983_ sky130_fd_sc_hd__nor2_1
XFILLER_0_98_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3555_ _0909_ _0913_ _0915_ VGND VGND VPWR VPWR _0918_ sky130_fd_sc_hd__a21o_1
X_3486_ _0835_ _0840_ _0848_ VGND VGND VPWR VPWR _0849_ sky130_fd_sc_hd__o21ai_1
X_5225_ disp_song.um.drum.next_idx1\[4\] _0191_ disp_song.um.drum.next_idx1\[3\] _2310_
+ VGND VGND VPWR VPWR _2311_ sky130_fd_sc_hd__or4b_1
XFILLER_0_44_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5156_ _2654_ _0173_ _0198_ VGND VGND VPWR VPWR _2243_ sky130_fd_sc_hd__and3_1
X_5087_ _2093_ _2094_ disp_song.um.drum.next_idx2\[2\] VGND VGND VPWR VPWR _2176_
+ sky130_fd_sc_hd__mux2_1
X_4107_ game.scoring_button_2.flash_counter_1\[5\] game.scoring_button_2.flash_counter_1\[4\]
+ game.scoring_button_2.flash_counter_1\[7\] game.scoring_button_2.flash_counter_1\[6\]
+ VGND VGND VPWR VPWR _1406_ sky130_fd_sc_hd__or4b_1
X_4038_ game.addmisses.add2.b\[2\] _1307_ _1346_ VGND VGND VPWR VPWR _1347_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5989_ clknet_leaf_33_clk _0098_ net71 VGND VGND VPWR VPWR game.padded_notes1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3340_ _0579_ _0696_ VGND VGND VPWR VPWR _0703_ sky130_fd_sc_hd__or2_1
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5010_ disp_song.um.drum.next_note2\[9\] _1968_ disp_song.um.drum.next_idx2\[1\]
+ VGND VGND VPWR VPWR _2102_ sky130_fd_sc_hd__a21oi_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3271_ _0460_ _0629_ _0633_ VGND VGND VPWR VPWR _0634_ sky130_fd_sc_hd__o21ai_4
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5912_ clknet_leaf_16_clk game.scoring_button_1.next_count\[3\] net62 VGND VGND VPWR
+ VPWR game.scoring_button_1.counts\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5843_ clknet_leaf_72_clk game.scoring_button_1.next_num_misses\[8\] net48 VGND VGND
+ VPWR VPWR game.addmisses.a\[8\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_33_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2986_ _0367_ _0375_ _0376_ VGND VGND VPWR VPWR disp_song.um.drum.next_note1\[4\]
+ sky130_fd_sc_hd__o21ai_2
X_5774_ clknet_leaf_7_clk game.scoring_button_2.next_count\[11\] net57 VGND VGND VPWR
+ VPWR game.scoring_button_2.counts\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4725_ _1868_ _1830_ _1869_ VGND VGND VPWR VPWR _1870_ sky130_fd_sc_hd__and3b_1
X_4656_ _1821_ VGND VGND VPWR VPWR game.scoring_button_1.next_count\[21\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4587_ game.addmisses.a\[13\] _1769_ _1675_ VGND VGND VPWR VPWR _1778_ sky130_fd_sc_hd__o21ai_1
X_3607_ _0963_ _0967_ _0935_ VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__o21a_1
XFILLER_0_101_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3538_ _0899_ highest_score.highest_score\[6\] highest_score.highest_score\[5\] VGND
+ VGND VPWR VPWR _0901_ sky130_fd_sc_hd__or3_1
X_3469_ _0796_ _0801_ _0803_ _0798_ VGND VGND VPWR VPWR _0832_ sky130_fd_sc_hd__or4b_1
X_5208_ _2230_ _2294_ disp_song.note1\[4\] disp_song.um.drum.next_idx1\[0\] VGND VGND
+ VPWR VPWR _2295_ sky130_fd_sc_hd__a2bb2o_1
X_5139_ disp_song.note1\[18\] _2226_ disp_song.um.drum.next_idx1\[0\] VGND VGND VPWR
+ VPWR _2227_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2840_ _2661_ _0158_ _0264_ _0267_ VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__a31o_1
XFILLER_0_45_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2771_ modetrans.mode\[1\] VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__buf_8
XFILLER_0_5_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5490_ _2523_ game.padded_notes2\[29\] _2515_ VGND VGND VPWR VPWR _2524_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4510_ game.addmisses.a\[3\] _1693_ _1709_ _1692_ VGND VGND VPWR VPWR _1711_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold106 pulseout.fin_pulse\[0\] VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xhold117 game.addhits.add4.b\[1\] VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__dlygate4sd3_1
X_4441_ game.addhits.a\[9\] _1650_ VGND VGND VPWR VPWR _1652_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold128 game.scoring_button_2.flash_counter_2\[4\] VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 game.padded_notes1\[28\] VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__dlygate4sd3_1
X_6111_ clknet_leaf_40_clk disp_song.um.drum.next_note1\[23\] net66 VGND VGND VPWR
+ VPWR disp_song.note1\[23\] sky130_fd_sc_hd__dfstp_1
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4372_ game.scoring_button_2.flash_counter_1\[15\] game.scoring_button_2.flash_counter_1\[16\]
+ _1590_ game.scoring_button_2.flash_counter_1\[17\] VGND VGND VPWR VPWR _1598_ sky130_fd_sc_hd__a31o_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3323_ _0569_ _0685_ _0574_ VGND VGND VPWR VPWR _0686_ sky130_fd_sc_hd__mux2_1
X_6042_ clknet_leaf_58_clk _0151_ net50 VGND VGND VPWR VPWR game.flash_counter\[22\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3254_ _0477_ _0616_ _0482_ VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__mux2_2
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3185_ game.addhits.add1.b\[0\] game.addhits.a\[0\] _0545_ _0547_ VGND VGND VPWR
+ VPWR _0548_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_95_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_603 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5826_ clknet_leaf_52_clk game.scoring_button_2.next_flash_counter_2\[17\] net55
+ VGND VGND VPWR VPWR game.scoring_button_2.flash_counter_2\[17\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2969_ disp_song.um.idx_note1\[0\] disp_song.um.idx_note1\[2\] _0179_ VGND VGND VPWR
+ VPWR _0362_ sky130_fd_sc_hd__or3b_2
X_5757_ clknet_leaf_64_clk game.scoring_button_2.next_num_hits\[13\] net47 VGND VGND
+ VPWR VPWR game.addhits.add4.b\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_29_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4708_ game.scoring_button_1.flash_counter_2\[12\] _1854_ VGND VGND VPWR VPWR _1858_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_17_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5688_ _2614_ _2647_ _2648_ VGND VGND VPWR VPWR _2649_ sky130_fd_sc_hd__and3_1
X_4639_ _1791_ _0013_ VGND VGND VPWR VPWR _1813_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4990_ disp_song.um.drum.next_idx2\[2\] _1962_ _2082_ VGND VGND VPWR VPWR _2083_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3941_ game.addhits.add3.b\[0\] _1253_ VGND VGND VPWR VPWR _1264_ sky130_fd_sc_hd__and2_1
X_3872_ _0966_ disp_song.display_note2\[1\] _0211_ game.out\[1\] _0208_ VGND VGND
+ VPWR VPWR _1211_ sky130_fd_sc_hd__a221o_1
X_2823_ _0253_ VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_73_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5611_ game.flash_counter\[1\] game.flash_counter\[0\] _0842_ VGND VGND VPWR VPWR
+ _2594_ sky130_fd_sc_hd__and3_1
X_5542_ _2553_ VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__clkbuf_1
X_2754_ modetrans.mode\[2\] _0195_ VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5473_ disp_song.note2\[24\] game.padded_notes2\[23\] _2497_ VGND VGND VPWR VPWR
+ _2512_ sky130_fd_sc_hd__mux2_1
X_2685_ disp_song.um.boton0e.edge_2 disp_song.um.boton0e.edge_1 VGND VGND VPWR VPWR
+ _2659_ sky130_fd_sc_hd__or2b_4
X_4424_ game.addhits.a\[6\] game.addhits.a\[5\] _1637_ game.addhits.a\[7\] VGND VGND
+ VPWR VPWR _1639_ sky130_fd_sc_hd__o31a_2
XFILLER_0_111_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4355_ game.scoring_button_2.flash_counter_1\[12\] _1583_ VGND VGND VPWR VPWR _1586_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_111_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3306_ _0543_ _0560_ _0561_ VGND VGND VPWR VPWR _0669_ sky130_fd_sc_hd__and3_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4286_ net159 _1535_ _1538_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_2\[13\]
+ sky130_fd_sc_hd__o21a_1
X_6025_ clknet_leaf_58_clk _0134_ net50 VGND VGND VPWR VPWR game.flash_counter\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3237_ _0493_ _0498_ _0599_ VGND VGND VPWR VPWR _0600_ sky130_fd_sc_hd__a21oi_2
X_3168_ _0529_ _0530_ VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__nor2_1
XTAP_1429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3099_ game.addmisses.a\[3\] game.addmisses.add1.b\[3\] VGND VGND VPWR VPWR _0462_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout56 net73 VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__buf_6
XFILLER_0_107_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout67 net73 VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__buf_4
XFILLER_0_9_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5809_ clknet_leaf_47_clk game.scoring_button_2.next_flash_counter_2\[0\] net56 VGND
+ VGND VPWR VPWR game.scoring_button_2.flash_counter_2\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_45_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_102_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_388 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4140_ _1427_ VGND VGND VPWR VPWR game.scoring_button_2.next_count\[6\] sky130_fd_sc_hd__clkbuf_1
X_4071_ net45 _1372_ _1373_ _1375_ VGND VGND VPWR VPWR game.scoring_button_2.next_num_misses\[10\]
+ sky130_fd_sc_hd__a22o_1
X_3022_ disp_song.um.idx_note1\[0\] disp_song.um.idx_note1\[2\] disp_song.um.idx_note1\[3\]
+ _0179_ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__and4_1
X_4973_ _1956_ disp_song.um.drum.next_note2\[7\] _1968_ _2036_ disp_song.um.drum.next_note2\[6\]
+ VGND VGND VPWR VPWR _2067_ sky130_fd_sc_hd__a32o_1
XFILLER_0_25_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3924_ game.addhits.add2.b\[0\] _1244_ VGND VGND VPWR VPWR _1251_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3855_ _0933_ _1199_ VGND VGND VPWR VPWR _1200_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2806_ game.counter\[14\] VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__inv_2
X_3786_ _0955_ _1134_ _1136_ _1138_ VGND VGND VPWR VPWR _1139_ sky130_fd_sc_hd__o211a_1
X_5525_ disp_song.note1\[6\] game.padded_notes1\[5\] _2541_ VGND VGND VPWR VPWR _2542_
+ sky130_fd_sc_hd__mux2_1
X_2737_ _0178_ _0180_ VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__and2_1
X_5456_ _2500_ net230 _2473_ VGND VGND VPWR VPWR _2501_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4407_ _1618_ _1625_ VGND VGND VPWR VPWR _1626_ sky130_fd_sc_hd__xnor2_1
X_5387_ _2447_ _2453_ VGND VGND VPWR VPWR _2454_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4338_ _1574_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_1\[6\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4269_ _1525_ game.missed_2 _1526_ VGND VGND VPWR VPWR _1527_ sky130_fd_sc_hd__and3b_1
X_6008_ clknet_leaf_49_clk _0117_ net56 VGND VGND VPWR VPWR game.padded_notes1\[27\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_96_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3640_ _0261_ _0993_ _0995_ _0997_ VGND VGND VPWR VPWR _0998_ sky130_fd_sc_hd__a211o_1
XFILLER_0_102_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3571_ _2654_ modetrans.mode\[5\] modetrans.mode\[3\] _0210_ _0933_ VGND VGND VPWR
+ VPWR _0934_ sky130_fd_sc_hd__o41a_1
XFILLER_0_23_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5310_ _2274_ _2286_ _2387_ _2392_ VGND VGND VPWR VPWR _2393_ sky130_fd_sc_hd__o211a_1
X_5241_ _2210_ _2211_ _2185_ VGND VGND VPWR VPWR _2327_ sky130_fd_sc_hd__mux2_1
X_5172_ _0430_ _2258_ _0175_ VGND VGND VPWR VPWR _2259_ sky130_fd_sc_hd__o21ai_1
X_4123_ _1417_ VGND VGND VPWR VPWR game.scoring_button_2.next_count\[2\] sky130_fd_sc_hd__clkbuf_1
Xinput2 button[1] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
X_4054_ net45 _1354_ _1356_ _1360_ VGND VGND VPWR VPWR game.scoring_button_2.next_num_misses\[8\]
+ sky130_fd_sc_hd__a31o_1
X_3005_ _2654_ _0388_ _0389_ _0390_ disp_song.note1\[9\] VGND VGND VPWR VPWR _0391_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4956_ _2034_ _2041_ _2049_ VGND VGND VPWR VPWR _2050_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_52_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4887_ _2664_ _0169_ VGND VGND VPWR VPWR _1982_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3907_ game.addhits.add1.b\[0\] _1236_ VGND VGND VPWR VPWR _1237_ sky130_fd_sc_hd__xor2_1
XFILLER_0_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3838_ _0925_ _1186_ _1187_ _0966_ VGND VGND VPWR VPWR _1188_ sky130_fd_sc_hd__o211a_1
XFILLER_0_61_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5508_ net97 _2458_ _2462_ game.padded_notes1\[0\] VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3769_ highest_score.highest_score\[0\] _1061_ VGND VGND VPWR VPWR _1123_ sky130_fd_sc_hd__or2_1
X_5439_ disp_song.note2\[13\] game.padded_notes2\[12\] _0219_ VGND VGND VPWR VPWR
+ _2489_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4810_ _1928_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_1\[20\]
+ sky130_fd_sc_hd__clkbuf_1
X_5790_ clknet_leaf_54_clk game.scoring_button_2.next_flash_counter_1\[4\] net52 VGND
+ VGND VPWR VPWR game.scoring_button_2.flash_counter_1\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4741_ net86 _1878_ game.missed_1 VGND VGND VPWR VPWR _1881_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_90_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4672_ net105 game.scoring_button_1.flash_counter_2\[0\] _1832_ VGND VGND VPWR VPWR
+ game.scoring_button_1.next_flash_counter_2\[1\] sky130_fd_sc_hd__a21oi_1
X_3623_ highest_score.highest_score\[4\] _0906_ _0975_ _0255_ _0904_ VGND VGND VPWR
+ VPWR _0982_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_12_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3554_ _0609_ _0667_ VGND VGND VPWR VPWR _0917_ sky130_fd_sc_hd__and2_1
X_3485_ _0841_ _0847_ VGND VGND VPWR VPWR _0848_ sky130_fd_sc_hd__and2_1
X_5224_ _0173_ disp_song.um.drum.next_idx1\[1\] VGND VGND VPWR VPWR _2310_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5155_ _2242_ VGND VGND VPWR VPWR disp_song.um.drum.next_d1\[0\] sky130_fd_sc_hd__clkbuf_1
X_5086_ disp_song.um.drum.next_note2\[0\] _2038_ _2174_ _1965_ VGND VGND VPWR VPWR
+ _2175_ sky130_fd_sc_hd__a211o_1
X_4106_ game.scoring_button_2.check_hit.in VGND VGND VPWR VPWR _1405_ sky130_fd_sc_hd__clkbuf_8
X_4037_ _1305_ _1344_ _1345_ VGND VGND VPWR VPWR _1346_ sky130_fd_sc_hd__or3b_1
XFILLER_0_94_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5988_ clknet_leaf_33_clk _0097_ net71 VGND VGND VPWR VPWR game.padded_notes1\[7\]
+ sky130_fd_sc_hd__dfstp_1
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4939_ _2013_ _2027_ _2031_ _2032_ VGND VGND VPWR VPWR _2033_ sky130_fd_sc_hd__a31o_1
XFILLER_0_19_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap42 _0842_ VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__buf_2
XFILLER_0_84_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_331 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3270_ _0466_ _0626_ _0627_ VGND VGND VPWR VPWR _0633_ sky130_fd_sc_hd__a21oi_4
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5911_ clknet_leaf_16_clk game.scoring_button_1.next_count\[2\] net62 VGND VGND VPWR
+ VPWR game.scoring_button_1.counts\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5842_ clknet_leaf_72_clk game.scoring_button_1.next_num_misses\[7\] net48 VGND VGND
+ VPWR VPWR game.addmisses.a\[7\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_48_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5773_ clknet_leaf_10_clk game.scoring_button_2.next_count\[10\] net57 VGND VGND
+ VPWR VPWR game.scoring_button_2.counts\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4724_ game.scoring_button_1.flash_counter_2\[15\] game.scoring_button_1.flash_counter_2\[16\]
+ _1861_ game.scoring_button_1.flash_counter_2\[17\] VGND VGND VPWR VPWR _1869_ sky130_fd_sc_hd__a31o_1
XFILLER_0_90_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2985_ _0368_ _0375_ disp_song.note1\[4\] VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__o21ai_1
X_4655_ game.scoring_button_1.check_hit.in _1475_ VGND VGND VPWR VPWR _1821_ sky130_fd_sc_hd__and2_1
X_4586_ game.addmisses.a\[13\] _1716_ _1769_ VGND VGND VPWR VPWR _1777_ sky130_fd_sc_hd__and3_1
XFILLER_0_24_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3606_ _0949_ _0961_ _0965_ _0966_ _0953_ VGND VGND VPWR VPWR _0967_ sky130_fd_sc_hd__a221o_1
XFILLER_0_101_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3537_ _0899_ highest_score.highest_score\[6\] VGND VGND VPWR VPWR _0900_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3468_ _0752_ _0773_ VGND VGND VPWR VPWR _0831_ sky130_fd_sc_hd__nor2_1
X_5207_ _0175_ disp_song.um.drum.next_note1\[5\] VGND VGND VPWR VPWR _2294_ sky130_fd_sc_hd__nand2_1
X_3399_ _0760_ _0761_ VGND VGND VPWR VPWR _0762_ sky130_fd_sc_hd__xnor2_4
X_5138_ _0415_ _2208_ VGND VGND VPWR VPWR _2226_ sky130_fd_sc_hd__nor2_1
X_5069_ _2121_ _2158_ _2026_ VGND VGND VPWR VPWR _2159_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2770_ modetrans.mode\[0\] VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_53_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4440_ _1650_ _1651_ net216 _1613_ VGND VGND VPWR VPWR game.scoring_button_1.next_num_hits\[8\]
+ sky130_fd_sc_hd__a2bb2o_1
Xhold107 game.scoring_button_1.flash_counter_1\[16\] VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold118 disp_song.note2\[22\] VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold129 game.addhits.a\[3\] VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__dlygate4sd3_1
X_6110_ clknet_leaf_38_clk disp_song.um.drum.next_note1\[22\] net66 VGND VGND VPWR
+ VPWR disp_song.note1\[22\] sky130_fd_sc_hd__dfstp_1
X_4371_ game.scoring_button_2.flash_counter_1\[17\] game.scoring_button_2.flash_counter_1\[16\]
+ _1593_ VGND VGND VPWR VPWR _1597_ sky130_fd_sc_hd__and3_1
XFILLER_0_95_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3322_ _0569_ _0575_ VGND VGND VPWR VPWR _0685_ sky130_fd_sc_hd__and2b_1
X_6041_ clknet_leaf_57_clk _0150_ net50 VGND VGND VPWR VPWR game.flash_counter\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3253_ _0610_ _0483_ VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__and2_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3184_ game.addhits.a\[1\] game.addhits.add1.b\[1\] VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5825_ clknet_leaf_52_clk net186 net55 VGND VGND VPWR VPWR game.scoring_button_2.flash_counter_2\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2968_ _0361_ VGND VGND VPWR VPWR disp_song.um.drum.next_note1\[1\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_63_139 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5756_ clknet_leaf_65_clk game.scoring_button_2.next_num_hits\[12\] net47 VGND VGND
+ VPWR VPWR game.addhits.add4.b\[0\] sky130_fd_sc_hd__dfrtp_1
X_4707_ game.scoring_button_1.flash_counter_2\[12\] _1854_ VGND VGND VPWR VPWR _1857_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_72_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5687_ game.flash_counter\[22\] _2629_ _2645_ game.flash_counter\[23\] VGND VGND
+ VPWR VPWR _2648_ sky130_fd_sc_hd__a31o_1
X_2899_ _0312_ VGND VGND VPWR VPWR disp_song.um.drum.next_note2\[14\] sky130_fd_sc_hd__buf_1
X_4638_ _1812_ VGND VGND VPWR VPWR game.scoring_button_1.next_count\[12\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4569_ game.addmisses.a\[10\] _1748_ VGND VGND VPWR VPWR _1762_ sky130_fd_sc_hd__nor2_1
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3940_ _1226_ _1259_ _1263_ net153 VGND VGND VPWR VPWR game.scoring_button_2.next_num_hits\[7\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3871_ _1210_ VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2822_ _0236_ _0239_ _0244_ _0252_ VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__or4_1
X_5610_ net124 _0830_ VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__xnor2_1
X_5541_ _2552_ game.padded_notes1\[11\] _2515_ VGND VGND VPWR VPWR _2553_ sky130_fd_sc_hd__mux2_1
X_2753_ _0194_ _0177_ _0170_ VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5472_ _2511_ VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__clkbuf_1
X_2684_ net148 disp_song.um.boton1e.edge_1 VGND VGND VPWR VPWR _2658_ sky130_fd_sc_hd__nor2b_4
XFILLER_0_30_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4423_ _1612_ _1636_ _1638_ _1613_ net267 VGND VGND VPWR VPWR game.scoring_button_1.next_num_hits\[4\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_41_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4354_ _1585_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_1\[11\]
+ sky130_fd_sc_hd__clkbuf_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3305_ _0476_ _0609_ _0617_ VGND VGND VPWR VPWR _0668_ sky130_fd_sc_hd__a21boi_1
X_6024_ clknet_leaf_58_clk _0133_ net50 VGND VGND VPWR VPWR game.flash_counter\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4285_ net159 _1535_ game.missed_2 VGND VGND VPWR VPWR _1538_ sky130_fd_sc_hd__a21boi_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3236_ _0493_ _0499_ _0498_ VGND VGND VPWR VPWR _0599_ sky130_fd_sc_hd__a21oi_1
X_3167_ game.addhits.a\[12\] game.addhits.add4.b\[0\] VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__nor2_1
X_3098_ _0454_ _0460_ VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__nor2_1
XTAP_1419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout46 net73 VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__buf_8
XFILLER_0_37_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout68 net70 VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__buf_6
Xfanout57 net61 VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__buf_6
X_5808_ clknet_leaf_55_clk game.scoring_button_2.next_flash_counter_1\[22\] net73
+ VGND VGND VPWR VPWR game.scoring_button_2.flash_counter_1\[22\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5739_ clknet_leaf_70_clk game.scoring_button_2.next_num_misses\[11\] net46 VGND
+ VGND VPWR VPWR game.addmisses.add3.b\[3\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_91_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4070_ net45 _1374_ VGND VGND VPWR VPWR _1375_ sky130_fd_sc_hd__nor2_1
X_3021_ _0380_ _0400_ _0401_ net250 VGND VGND VPWR VPWR disp_song.um.drum.next_note1\[14\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4972_ _2026_ _2043_ _2063_ _2065_ VGND VGND VPWR VPWR _2066_ sky130_fd_sc_hd__a31o_1
XFILLER_0_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3923_ game.addhits.add2.b\[0\] _1244_ VGND VGND VPWR VPWR _1250_ sky130_fd_sc_hd__or2_1
XFILLER_0_73_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3854_ _0966_ disp_song.display_note1\[2\] _0211_ game.out\[9\] _0208_ VGND VGND
+ VPWR VPWR _1199_ sky130_fd_sc_hd__a221o_2
X_2805_ _0233_ _0234_ _0235_ VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__or3_1
XFILLER_0_6_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3785_ _1050_ _1137_ _0896_ VGND VGND VPWR VPWR _1138_ sky130_fd_sc_hd__a21o_1
X_2736_ disp_song.um.idx_note1\[0\] _0179_ VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__nor2_2
X_5524_ _0209_ VGND VGND VPWR VPWR _2541_ sky130_fd_sc_hd__buf_6
XFILLER_0_6_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5455_ disp_song.note2\[18\] game.padded_notes2\[17\] _2497_ VGND VGND VPWR VPWR
+ _2500_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4406_ _1619_ _1624_ VGND VGND VPWR VPWR _1625_ sky130_fd_sc_hd__nand2_1
X_5386_ pulseout.fin_pulse\[0\] pulseout.fin_pulse\[1\] pulseout.fin_pulse\[2\] pulseout.fin_pulse\[3\]
+ VGND VGND VPWR VPWR _2453_ sky130_fd_sc_hd__and4_1
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4337_ _1572_ _1413_ _1573_ VGND VGND VPWR VPWR _1574_ sky130_fd_sc_hd__and3b_1
X_4268_ game.scoring_button_2.flash_counter_2\[7\] game.scoring_button_2.flash_counter_2\[6\]
+ _1518_ game.scoring_button_2.flash_counter_2\[8\] VGND VGND VPWR VPWR _1526_ sky130_fd_sc_hd__a31o_1
X_3219_ game.addhits.a\[10\] game.addhits.add3.b\[2\] VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__nand2_1
X_6007_ clknet_leaf_49_clk _0116_ net66 VGND VGND VPWR VPWR game.padded_notes1\[26\]
+ sky130_fd_sc_hd__dfstp_1
X_4199_ game.counter\[20\] _1466_ VGND VGND VPWR VPWR _1470_ sky130_fd_sc_hd__and2_1
XTAP_1205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_350 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3570_ net5 VGND VGND VPWR VPWR _0933_ sky130_fd_sc_hd__inv_12
XFILLER_0_24_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5240_ _2192_ _2196_ disp_song.um.drum.next_idx1\[1\] VGND VGND VPWR VPWR _2326_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5171_ disp_song.um.drum.next_idx1\[4\] _2257_ VGND VGND VPWR VPWR _2258_ sky130_fd_sc_hd__nor2_2
X_4122_ _1405_ _0024_ VGND VGND VPWR VPWR _1417_ sky130_fd_sc_hd__and2_1
X_4053_ game.addmisses.add3.b\[0\] _1357_ _1359_ _1289_ VGND VGND VPWR VPWR _1360_
+ sky130_fd_sc_hd__o211a_1
X_3004_ _2661_ _0194_ _0359_ _0354_ VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__or4_1
Xinput3 button[2] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
X_4955_ _2020_ _2045_ _2048_ _2013_ VGND VGND VPWR VPWR _2049_ sky130_fd_sc_hd__o211a_1
XFILLER_0_19_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3906_ _1231_ _1230_ VGND VGND VPWR VPWR _1236_ sky130_fd_sc_hd__nand2_1
X_4886_ _1961_ _1974_ _1977_ _1980_ _2679_ VGND VGND VPWR VPWR _1981_ sky130_fd_sc_hd__o32a_1
XFILLER_0_74_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3837_ _1080_ _1086_ _0925_ VGND VGND VPWR VPWR _1187_ sky130_fd_sc_hd__or3b_1
XFILLER_0_6_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3768_ _1067_ _1093_ VGND VGND VPWR VPWR _1122_ sky130_fd_sc_hd__or2_1
X_2719_ disp_song.um.idx_note2\[1\] disp_song.um.idx_note2\[0\] disp_song.um.idx_note2\[2\]
+ VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__o21ba_1
X_5507_ net170 _2530_ _1673_ VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__o21a_1
XFILLER_0_100_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3699_ highest_score.highest_score\[2\] highest_score.highest_score\[1\] highest_score.highest_score\[3\]
+ VGND VGND VPWR VPWR _1055_ sky130_fd_sc_hd__or3b_1
X_5438_ _2488_ VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5369_ _0830_ _0838_ VGND VGND VPWR VPWR _2442_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4740_ _1880_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_2\[21\]
+ sky130_fd_sc_hd__clkbuf_1
X_4671_ net105 game.scoring_button_1.flash_counter_2\[0\] game.missed_1 VGND VGND
+ VPWR VPWR _1832_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_83_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3622_ _0956_ _0971_ _0261_ VGND VGND VPWR VPWR _0981_ sky130_fd_sc_hd__o21a_1
XFILLER_0_71_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3553_ _0909_ _0913_ _0915_ _0667_ VGND VGND VPWR VPWR _0916_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3484_ net42 _0845_ _0846_ VGND VGND VPWR VPWR _0847_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_11_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5223_ _2309_ VGND VGND VPWR VPWR disp_song.um.drum.next_d1\[1\] sky130_fd_sc_hd__clkbuf_1
X_5154_ _0214_ _2241_ VGND VGND VPWR VPWR _2242_ sky130_fd_sc_hd__and2_1
X_4105_ _1289_ _1402_ _1404_ VGND VGND VPWR VPWR game.scoring_button_2.next_num_misses\[15\]
+ sky130_fd_sc_hd__o21ai_1
X_5085_ _2664_ _1956_ disp_song.um.drum.next_note2\[2\] _1992_ VGND VGND VPWR VPWR
+ _2174_ sky130_fd_sc_hd__and4b_1
XFILLER_0_2_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4036_ game.addmisses.add2.b\[1\] game.addmisses.add2.b\[0\] _1319_ game.addmisses.add2.b\[2\]
+ VGND VGND VPWR VPWR _1345_ sky130_fd_sc_hd__a31o_1
XFILLER_0_63_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5987_ clknet_leaf_37_clk _0096_ net71 VGND VGND VPWR VPWR game.padded_notes1\[6\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_93_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4938_ _2679_ _2010_ VGND VGND VPWR VPWR _2032_ sky130_fd_sc_hd__xnor2_1
X_4869_ _1948_ _1949_ VGND VGND VPWR VPWR _1964_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap43 _0811_ VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5910_ clknet_leaf_16_clk game.scoring_button_1.next_count\[1\] net62 VGND VGND VPWR
+ VPWR game.scoring_button_1.counts\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5841_ clknet_leaf_73_clk game.scoring_button_1.next_num_misses\[6\] net48 VGND VGND
+ VPWR VPWR game.addmisses.a\[6\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_48_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2984_ disp_song.um.idx_note1\[3\] _0374_ VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__or2_2
X_5772_ clknet_leaf_10_clk game.scoring_button_2.next_count\[9\] net57 VGND VGND VPWR
+ VPWR game.scoring_button_2.counts\[9\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_63 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4723_ game.scoring_button_1.flash_counter_2\[17\] game.scoring_button_1.flash_counter_2\[16\]
+ _1864_ VGND VGND VPWR VPWR _1868_ sky130_fd_sc_hd__and3_1
XFILLER_0_83_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4654_ _1820_ VGND VGND VPWR VPWR game.scoring_button_1.next_count\[20\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_618 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4585_ game.addmisses.a\[15\] _1773_ _1775_ VGND VGND VPWR VPWR _1776_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3605_ _2654_ VGND VGND VPWR VPWR _0966_ sky130_fd_sc_hd__buf_6
XFILLER_0_12_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3536_ net152 VGND VGND VPWR VPWR _0899_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3467_ _0829_ VGND VGND VPWR VPWR _0830_ sky130_fd_sc_hd__clkbuf_4
X_5206_ _2247_ _2286_ _2292_ VGND VGND VPWR VPWR _2293_ sky130_fd_sc_hd__o21ba_1
X_3398_ _0725_ _0750_ _0749_ VGND VGND VPWR VPWR _0761_ sky130_fd_sc_hd__a21oi_4
X_5137_ _2222_ _2224_ VGND VGND VPWR VPWR _2225_ sky130_fd_sc_hd__nor2_1
X_5068_ disp_song.note2\[16\] disp_song.um.drum.next_idx2\[1\] _2044_ VGND VGND VPWR
+ VPWR _2158_ sky130_fd_sc_hd__o21a_1
XFILLER_0_74_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4019_ modetrans.mode\[0\] _1305_ VGND VGND VPWR VPWR _1330_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_434 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold108 game.scoring_button_1.flash_counter_2\[19\] VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__dlygate4sd3_1
X_4370_ net174 _1593_ _1596_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_1\[16\]
+ sky130_fd_sc_hd__o21a_1
Xhold119 game.scoring_button_2.flash_counter_1\[7\] VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__dlygate4sd3_1
X_3321_ _0622_ _0679_ _0620_ VGND VGND VPWR VPWR _0684_ sky130_fd_sc_hd__o21ai_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_95_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6040_ clknet_leaf_57_clk _0149_ net50 VGND VGND VPWR VPWR game.flash_counter\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3252_ _0476_ _0609_ VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__nand2_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3183_ _0544_ _0545_ VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5824_ clknet_leaf_51_clk game.scoring_button_2.next_flash_counter_2\[15\] net55
+ VGND VGND VPWR VPWR game.scoring_button_2.flash_counter_2\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2967_ _0355_ _0358_ _0360_ disp_song.note1\[1\] VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_72_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5755_ clknet_leaf_68_clk game.scoring_button_2.next_num_hits\[11\] net46 VGND VGND
+ VPWR VPWR game.addhits.add3.b\[3\] sky130_fd_sc_hd__dfrtp_2
X_4706_ _1856_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_2\[11\]
+ sky130_fd_sc_hd__clkbuf_1
X_2898_ disp_song.note2\[14\] _0269_ _0311_ VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5686_ game.flash_counter\[22\] game.flash_counter\[23\] _2629_ _2645_ VGND VGND
+ VPWR VPWR _2647_ sky130_fd_sc_hd__nand4_1
XFILLER_0_32_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4637_ _1791_ _0012_ VGND VGND VPWR VPWR _1812_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4568_ _1699_ _1758_ _1759_ _1761_ VGND VGND VPWR VPWR game.scoring_button_1.next_num_misses\[10\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3519_ _0608_ _0675_ _0881_ _0686_ VGND VGND VPWR VPWR _0882_ sky130_fd_sc_hd__o31a_1
X_4499_ game.addmisses.a\[2\] game.addmisses.a\[1\] game.addmisses.a\[0\] VGND VGND
+ VPWR VPWR _1701_ sky130_fd_sc_hd__and3_1
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6169_ clknet_leaf_45_clk disp_song.um.drum.next_d1\[1\] net54 VGND VGND VPWR VPWR
+ disp_song.display_note1\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_20_clk clknet_3_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_20_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_90_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3870_ _0933_ _1209_ VGND VGND VPWR VPWR _1210_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2821_ _0246_ _0247_ _0249_ _0251_ VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__or4b_1
XFILLER_0_26_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5540_ disp_song.note1\[11\] game.padded_notes1\[10\] _2541_ VGND VGND VPWR VPWR
+ _2552_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2752_ _0193_ VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_11_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_11_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_26_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5471_ _2510_ game.padded_notes2\[23\] _2473_ VGND VGND VPWR VPWR _2511_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_302 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2683_ _2655_ _2656_ VGND VGND VPWR VPWR _2657_ sky130_fd_sc_hd__nor2_4
X_4422_ _1637_ VGND VGND VPWR VPWR _1638_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4353_ _1583_ game.hit_2 _1584_ VGND VGND VPWR VPWR _1585_ sky130_fd_sc_hd__and3b_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4284_ _1537_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_2\[12\]
+ sky130_fd_sc_hd__clkbuf_1
X_3304_ _0449_ _0666_ VGND VGND VPWR VPWR _0667_ sky130_fd_sc_hd__xnor2_4
X_6023_ clknet_leaf_64_clk _0132_ net50 VGND VGND VPWR VPWR game.flash_counter\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3235_ _0487_ _0500_ VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__xor2_1
XFILLER_0_39_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3166_ game.addhits.a\[12\] game.addhits.add4.b\[0\] VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__and2_1
XFILLER_0_96_519 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3097_ _0456_ _0459_ VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_55_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout47 net73 VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__buf_4
XFILLER_0_36_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout69 net70 VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__buf_8
XFILLER_0_91_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout58 net61 VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__buf_6
X_5807_ clknet_leaf_55_clk game.scoring_button_2.next_flash_counter_1\[21\] net52
+ VGND VGND VPWR VPWR game.scoring_button_2.flash_counter_1\[21\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3999_ game.scoring_button_2.check_hit.edge_1 _1287_ game.scoring_button_2.hit VGND
+ VGND VPWR VPWR _1313_ sky130_fd_sc_hd__nor3_1
XFILLER_0_91_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5738_ clknet_leaf_70_clk game.scoring_button_2.next_num_misses\[10\] net46 VGND
+ VGND VPWR VPWR game.addmisses.add3.b\[2\] sky130_fd_sc_hd__dfrtp_4
X_5669_ game.flash_counter\[17\] game.flash_counter\[16\] _2629_ net263 VGND VGND
+ VPWR VPWR _2635_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_32_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_69_clk clknet_3_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_69_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_55_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_154 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3020_ _0382_ _0400_ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_0_clk clknet_3_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_0_clk sky130_fd_sc_hd__clkbuf_16
X_4971_ disp_song.um.drum.next_idx2\[0\] disp_song.um.drum.next_note2\[3\] _1965_
+ _2020_ _2064_ VGND VGND VPWR VPWR _2065_ sky130_fd_sc_hd__o2111a_1
X_3922_ _1226_ _1246_ _1249_ _1227_ net178 VGND VGND VPWR VPWR game.scoring_button_2.next_num_hits\[3\]
+ sky130_fd_sc_hd__a32o_1
X_3853_ _1198_ VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
X_2804_ game.counter\[7\] _0227_ VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3784_ _0639_ _1042_ net44 VGND VGND VPWR VPWR _1137_ sky130_fd_sc_hd__or3b_1
X_5523_ _2540_ VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__clkbuf_1
X_2735_ disp_song.um.idx_note1\[1\] VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_14_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5454_ _2499_ VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5385_ pulseout.fin_pulse\[0\] pulseout.fin_pulse\[1\] pulseout.fin_pulse\[2\] game.beat_clk
+ pulseout.fin_pulse\[3\] VGND VGND VPWR VPWR _2452_ sky130_fd_sc_hd__a41o_1
X_4405_ game.addhits.a\[2\] game.scoring_button_1.acc\[2\] VGND VGND VPWR VPWR _1624_
+ sky130_fd_sc_hd__or2_1
X_4336_ game.scoring_button_2.flash_counter_1\[6\] _1569_ VGND VGND VPWR VPWR _1573_
+ sky130_fd_sc_hd__or2_1
X_4267_ game.scoring_button_2.flash_counter_2\[7\] game.scoring_button_2.flash_counter_2\[8\]
+ _1521_ VGND VGND VPWR VPWR _1525_ sky130_fd_sc_hd__and3_1
X_4198_ game.counter\[20\] _1466_ VGND VGND VPWR VPWR _1469_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6006_ clknet_leaf_39_clk _0115_ net66 VGND VGND VPWR VPWR game.padded_notes1\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_3218_ game.addhits.a\[10\] game.addhits.add3.b\[2\] VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__nor2_1
X_3149_ _0508_ _0511_ VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__xnor2_2
XTAP_1239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_530 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5170_ disp_song.um.drum.next_idx1\[3\] _2245_ VGND VGND VPWR VPWR _2257_ sky130_fd_sc_hd__or2_1
X_4121_ net199 _1415_ VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__xnor2_1
X_4052_ _1358_ _1357_ game.addmisses.add3.b\[0\] VGND VGND VPWR VPWR _1359_ sky130_fd_sc_hd__o21ai_1
Xinput4 button[3] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
X_3003_ _2661_ _0194_ _0358_ VGND VGND VPWR VPWR _0389_ sky130_fd_sc_hd__nor3_1
XFILLER_0_36_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4954_ _1965_ _2046_ _2047_ _2026_ VGND VGND VPWR VPWR _2048_ sky130_fd_sc_hd__a31o_1
XFILLER_0_74_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3905_ game.addhits.add1.b\[3\] _1234_ VGND VGND VPWR VPWR _1235_ sky130_fd_sc_hd__nor2_1
X_4885_ _1978_ _1979_ disp_song.um.drum.next_idx2\[1\] VGND VGND VPWR VPWR _1980_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3836_ _1077_ _1117_ _1080_ disp_song.mi6.in\[2\] VGND VGND VPWR VPWR _1186_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_6_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3767_ _1090_ _1120_ VGND VGND VPWR VPWR _1121_ sky130_fd_sc_hd__nor2_1
X_2718_ _0163_ VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__inv_2
X_5506_ _2529_ VGND VGND VPWR VPWR _2530_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3698_ highest_score.highest_score\[3\] _1053_ VGND VGND VPWR VPWR _1054_ sky130_fd_sc_hd__or2_1
X_5437_ _2487_ net235 _2473_ VGND VGND VPWR VPWR _2488_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5368_ _2441_ VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__clkbuf_1
X_4319_ net103 game.scoring_button_2.flash_counter_1\[0\] game.hit_2 VGND VGND VPWR
+ VPWR _1561_ sky130_fd_sc_hd__o21ai_1
X_5299_ _2310_ _2380_ _2381_ _2254_ VGND VGND VPWR VPWR _2382_ sky130_fd_sc_hd__o22a_1
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4670_ _1831_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_2\[0\]
+ sky130_fd_sc_hd__clkbuf_1
X_3621_ _0931_ _0953_ _0980_ _0935_ VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__o31a_1
XFILLER_0_71_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3552_ _0909_ _0614_ _0914_ VGND VGND VPWR VPWR _0915_ sky130_fd_sc_hd__nor3_1
XFILLER_0_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3483_ _0762_ _0824_ _0825_ _0826_ _0781_ VGND VGND VPWR VPWR _0846_ sky130_fd_sc_hd__o311a_1
X_5222_ _0214_ _2308_ VGND VGND VPWR VPWR _2309_ sky130_fd_sc_hd__and2_1
X_5153_ _2217_ _2239_ _2240_ VGND VGND VPWR VPWR _2241_ sky130_fd_sc_hd__mux2_1
X_4104_ game.addmisses.add4.b\[3\] _1395_ _1403_ net45 VGND VGND VPWR VPWR _1404_
+ sky130_fd_sc_hd__a211o_1
X_5084_ disp_song.um.drum.next_note2\[5\] _2134_ _2135_ disp_song.um.drum.next_note2\[4\]
+ _2172_ VGND VGND VPWR VPWR _2173_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4035_ game.addmisses.add2.b\[2\] game.addmisses.add2.b\[1\] game.addmisses.add2.b\[0\]
+ _1319_ VGND VGND VPWR VPWR _1344_ sky130_fd_sc_hd__and4_1
XFILLER_0_2_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5986_ clknet_leaf_33_clk _0095_ net71 VGND VGND VPWR VPWR game.padded_notes1\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4937_ _2028_ _2030_ _2020_ VGND VGND VPWR VPWR _2031_ sky130_fd_sc_hd__a21o_1
XFILLER_0_59_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4868_ _1961_ _1962_ VGND VGND VPWR VPWR _1963_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_503 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3819_ _1059_ _1098_ _1169_ _0258_ VGND VGND VPWR VPWR _1170_ sky130_fd_sc_hd__a31o_1
XFILLER_0_62_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4799_ _1919_ _1799_ _1920_ VGND VGND VPWR VPWR _1921_ sky130_fd_sc_hd__and3b_1
XFILLER_0_15_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xmax_cap44 _0885_ VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_85_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5840_ clknet_leaf_71_clk game.scoring_button_1.next_num_misses\[5\] net48 VGND VGND
+ VPWR VPWR game.addmisses.a\[5\] sky130_fd_sc_hd__dfrtp_4
X_2983_ disp_song.um.idx_note1\[2\] _0180_ VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__nand2_2
X_5771_ clknet_leaf_10_clk game.scoring_button_2.next_count\[8\] net57 VGND VGND VPWR
+ VPWR game.scoring_button_2.counts\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4722_ net194 _1864_ _1867_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_2\[16\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_8_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4653_ game.scoring_button_1.check_hit.in _1471_ VGND VGND VPWR VPWR _1820_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4584_ game.addmisses.a\[14\] _1771_ _1774_ VGND VGND VPWR VPWR _1775_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_24_271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3604_ disp_song.mi6.in\[3\] _0964_ _0929_ VGND VGND VPWR VPWR _0965_ sky130_fd_sc_hd__a21o_1
X_3535_ highest_score.highest_score\[5\] VGND VGND VPWR VPWR _0898_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3466_ _0762_ _0824_ _0825_ _0826_ VGND VGND VPWR VPWR _0829_ sky130_fd_sc_hd__o31a_1
X_5205_ _2256_ _2288_ _2289_ _2291_ _2247_ VGND VGND VPWR VPWR _2292_ sky130_fd_sc_hd__o221a_1
X_3397_ _0758_ _0759_ VGND VGND VPWR VPWR _0760_ sky130_fd_sc_hd__or2b_2
XFILLER_0_42_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5136_ _2195_ _2223_ disp_song.um.drum.next_idx1\[1\] VGND VGND VPWR VPWR _2224_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5067_ _2679_ _2012_ VGND VGND VPWR VPWR _2157_ sky130_fd_sc_hd__xnor2_2
X_4018_ game.addmisses.add2.b\[0\] _1319_ VGND VGND VPWR VPWR _1329_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5969_ clknet_leaf_31_clk game.scoring_button_1.next_flash_counter_2\[14\] net69
+ VGND VGND VPWR VPWR game.scoring_button_1.flash_counter_2\[14\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_111_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold109 game.addhits.add4.b\[0\] VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3320_ _0680_ _0682_ VGND VGND VPWR VPWR _0683_ sky130_fd_sc_hd__and2b_1
XFILLER_0_95_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3251_ _0610_ _0611_ _0613_ _0476_ VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__o22a_1
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3182_ game.addhits.a\[1\] game.addhits.add1.b\[1\] VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__xor2_4
XFILLER_0_76_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5823_ clknet_leaf_51_clk game.scoring_button_2.next_flash_counter_2\[14\] net55
+ VGND VGND VPWR VPWR game.scoring_button_2.flash_counter_2\[14\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_650 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2966_ _0359_ _0355_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__or2_1
X_5754_ clknet_leaf_68_clk game.scoring_button_2.next_num_hits\[10\] net46 VGND VGND
+ VPWR VPWR game.addhits.add3.b\[2\] sky130_fd_sc_hd__dfrtp_1
X_4705_ _1854_ game.missed_1 _1855_ VGND VGND VPWR VPWR _1856_ sky130_fd_sc_hd__and3b_1
X_2897_ _0310_ _0298_ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__nor2_1
X_5685_ net125 _2646_ VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_44_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4636_ _1811_ VGND VGND VPWR VPWR game.scoring_button_1.next_count\[11\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4567_ _1699_ _1760_ VGND VGND VPWR VPWR _1761_ sky130_fd_sc_hd__nor2_1
X_3518_ _0671_ _0624_ _0880_ VGND VGND VPWR VPWR _0881_ sky130_fd_sc_hd__and3b_1
X_4498_ _1675_ _1696_ _1698_ _1700_ VGND VGND VPWR VPWR game.scoring_button_1.next_num_misses\[1\]
+ sky130_fd_sc_hd__o2bb2a_1
X_3449_ _0781_ _0793_ _0784_ VGND VGND VPWR VPWR _0812_ sky130_fd_sc_hd__a21o_1
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6168_ clknet_leaf_44_clk disp_song.um.drum.next_d1\[0\] net54 VGND VGND VPWR VPWR
+ disp_song.display_note1\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5119_ _0185_ _0191_ _0197_ VGND VGND VPWR VPWR _2207_ sky130_fd_sc_hd__and3_1
X_6099_ clknet_leaf_37_clk disp_song.um.drum.next_note1\[11\] net67 VGND VGND VPWR
+ VPWR disp_song.note1\[11\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_79_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2820_ game.counter\[9\] _0222_ _0250_ game.counter\[19\] game.counter\[18\] VGND
+ VGND VPWR VPWR _0251_ sky130_fd_sc_hd__o2111a_1
X_2751_ _0182_ _0192_ VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5470_ disp_song.note2\[23\] game.padded_notes2\[22\] _2497_ VGND VGND VPWR VPWR
+ _2510_ sky130_fd_sc_hd__mux2_1
X_2682_ disp_song.um.boton0e.edge_2 disp_song.um.boton0e.edge_1 VGND VGND VPWR VPWR
+ _2656_ sky130_fd_sc_hd__nor2b_4
XFILLER_0_81_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4421_ game.addhits.a\[4\] _1630_ VGND VGND VPWR VPWR _1637_ sky130_fd_sc_hd__and2_1
XFILLER_0_1_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_572 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4352_ game.scoring_button_2.flash_counter_1\[9\] game.scoring_button_2.flash_counter_1\[10\]
+ _1576_ game.scoring_button_2.flash_counter_1\[11\] VGND VGND VPWR VPWR _1584_ sky130_fd_sc_hd__a31o_1
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4283_ _1535_ game.missed_2 _1536_ VGND VGND VPWR VPWR _1537_ sky130_fd_sc_hd__and3b_1
X_3303_ _0468_ _0469_ VGND VGND VPWR VPWR _0666_ sky130_fd_sc_hd__nor2_2
X_6022_ clknet_leaf_59_clk _0131_ net50 VGND VGND VPWR VPWR game.flash_counter\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3234_ _0443_ _0596_ VGND VGND VPWR VPWR _0597_ sky130_fd_sc_hd__xnor2_2
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3165_ _0512_ _0524_ _0527_ VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_55_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3096_ _0457_ _0458_ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__and2b_1
XFILLER_0_89_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xfanout59 net60 VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_6
X_5806_ clknet_leaf_55_clk game.scoring_button_2.next_flash_counter_1\[20\] net52
+ VGND VGND VPWR VPWR game.scoring_button_2.flash_counter_1\[20\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3998_ _1309_ _1311_ VGND VGND VPWR VPWR _1312_ sky130_fd_sc_hd__and2_1
Xfanout48 net49 VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__buf_8
X_2949_ _0285_ _0345_ _0346_ net244 VGND VGND VPWR VPWR disp_song.um.drum.next_note2\[29\]
+ sky130_fd_sc_hd__a22o_1
X_5737_ clknet_leaf_70_clk game.scoring_button_2.next_num_misses\[9\] net46 VGND VGND
+ VPWR VPWR game.addmisses.add3.b\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_44_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5668_ net137 _2633_ VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__xnor2_1
X_4619_ _1791_ _0025_ VGND VGND VPWR VPWR _1803_ sky130_fd_sc_hd__and2_1
X_5599_ _2591_ VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_99_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_531 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4970_ _2669_ disp_song.um.drum.next_note2\[2\] VGND VGND VPWR VPWR _2064_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3921_ _1235_ _1241_ _1243_ VGND VGND VPWR VPWR _1249_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_46_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3852_ _0933_ _1197_ VGND VGND VPWR VPWR _1198_ sky130_fd_sc_hd__and2_1
X_2803_ game.counter\[6\] _0222_ VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__and2_1
XFILLER_0_27_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5522_ _2539_ net256 _2515_ VGND VGND VPWR VPWR _2540_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3783_ _1062_ _1135_ _0258_ VGND VGND VPWR VPWR _1136_ sky130_fd_sc_hd__a21o_1
XFILLER_0_54_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2734_ disp_song.um.idx_note1\[2\] VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_347 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5453_ _2498_ game.padded_notes2\[17\] _2473_ VGND VGND VPWR VPWR _2499_ sky130_fd_sc_hd__mux2_1
X_5384_ net128 _2449_ VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_188 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4404_ game.addhits.a\[0\] _1622_ VGND VGND VPWR VPWR _1623_ sky130_fd_sc_hd__xor2_1
X_4335_ game.scoring_button_2.flash_counter_1\[6\] _1569_ VGND VGND VPWR VPWR _1572_
+ sky130_fd_sc_hd__and2_1
X_4266_ net151 _1521_ _1524_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_2\[7\]
+ sky130_fd_sc_hd__o21a_1
X_6005_ clknet_leaf_39_clk _0114_ net66 VGND VGND VPWR VPWR game.padded_notes1\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_4197_ _1468_ VGND VGND VPWR VPWR game.scoring_button_2.next_count\[19\] sky130_fd_sc_hd__clkbuf_1
X_3217_ _0533_ _0578_ _0532_ VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__a21boi_1
X_3148_ _0509_ _0510_ VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3079_ game.addmisses.a\[8\] game.addmisses.add3.b\[0\] VGND VGND VPWR VPWR _0442_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_77_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4120_ _1416_ VGND VGND VPWR VPWR game.scoring_button_2.next_count\[1\] sky130_fd_sc_hd__clkbuf_1
X_4051_ modetrans.mode\[0\] _1305_ VGND VGND VPWR VPWR _1358_ sky130_fd_sc_hd__and2_1
Xinput5 chip_select VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__buf_2
X_3002_ _0179_ disp_song.um.idx_note1\[0\] _0178_ VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__and3b_1
XFILLER_0_36_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4953_ _2669_ disp_song.um.drum.next_note2\[18\] VGND VGND VPWR VPWR _2047_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_575 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3904_ _1229_ _1232_ _1233_ VGND VGND VPWR VPWR _1234_ sky130_fd_sc_hd__o21ai_1
X_4884_ disp_song.um.drum.next_note2\[20\] disp_song.um.drum.next_note2\[21\] disp_song.um.drum.next_idx2\[0\]
+ VGND VGND VPWR VPWR _1979_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3835_ _1036_ _1162_ _1184_ net38 VGND VGND VPWR VPWR _1185_ sky130_fd_sc_hd__o211a_1
XFILLER_0_27_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3766_ _0806_ _1035_ _1033_ VGND VGND VPWR VPWR _1120_ sky130_fd_sc_hd__and3_1
X_2717_ disp_song.um.idx_note2\[1\] disp_song.um.idx_note2\[0\] disp_song.um.idx_note2\[2\]
+ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__or3b_4
X_5505_ _0209_ _2656_ _1688_ VGND VGND VPWR VPWR _2529_ sky130_fd_sc_hd__nand3_1
X_5436_ disp_song.note2\[12\] game.padded_notes2\[11\] _0219_ VGND VGND VPWR VPWR
+ _2487_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3697_ highest_score.highest_score\[2\] VGND VGND VPWR VPWR _1053_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5367_ _0946_ highest_score.highest_score\[4\] _2434_ VGND VGND VPWR VPWR _2441_
+ sky130_fd_sc_hd__mux2_1
X_4318_ _1560_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_1\[0\]
+ sky130_fd_sc_hd__clkbuf_1
X_5298_ disp_song.note1\[17\] _2185_ _2271_ VGND VGND VPWR VPWR _2381_ sky130_fd_sc_hd__o21a_1
X_4249_ _1511_ game.missed_2 _1512_ VGND VGND VPWR VPWR _1513_ sky130_fd_sc_hd__and3b_1
XFILLER_0_97_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3620_ net39 _0968_ _0978_ _0979_ VGND VGND VPWR VPWR _0980_ sky130_fd_sc_hd__a31o_1
XFILLER_0_43_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3551_ _0617_ _0912_ VGND VGND VPWR VPWR _0914_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3482_ _0809_ _0843_ _0844_ _0775_ _0831_ VGND VGND VPWR VPWR _0845_ sky130_fd_sc_hd__a2111o_1
X_5221_ _2281_ _2306_ _2307_ VGND VGND VPWR VPWR _2308_ sky130_fd_sc_hd__mux2_1
X_5152_ _0185_ _2194_ VGND VGND VPWR VPWR _2240_ sky130_fd_sc_hd__nor2_1
X_4103_ game.addmisses.add4.b\[3\] _1394_ VGND VGND VPWR VPWR _1403_ sky130_fd_sc_hd__nor2_1
X_5083_ disp_song.um.drum.next_note2\[3\] _1992_ _2035_ _2171_ disp_song.um.drum.next_note2\[1\]
+ VGND VGND VPWR VPWR _2172_ sky130_fd_sc_hd__a32o_1
XFILLER_0_79_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4034_ game.addmisses.add2.b\[2\] _1342_ VGND VGND VPWR VPWR _1343_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5985_ clknet_leaf_32_clk _0094_ net71 VGND VGND VPWR VPWR game.padded_notes1\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4936_ disp_song.um.drum.next_note2\[25\] _2029_ _2666_ VGND VGND VPWR VPWR _2030_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4867_ disp_song.um.drum.next_idx2\[1\] _1949_ VGND VGND VPWR VPWR _1962_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3818_ _0255_ _1055_ VGND VGND VPWR VPWR _1169_ sky130_fd_sc_hd__and2_1
X_4798_ game.scoring_button_1.flash_counter_1\[15\] game.scoring_button_1.flash_counter_1\[16\]
+ _1912_ game.scoring_button_1.flash_counter_1\[17\] VGND VGND VPWR VPWR _1920_ sky130_fd_sc_hd__a31o_1
X_3749_ _1077_ _0926_ VGND VGND VPWR VPWR _1104_ sky130_fd_sc_hd__nor2_1
X_5419_ _2475_ net227 _2473_ VGND VGND VPWR VPWR _2476_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap45 _1313_ VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__buf_2
XFILLER_0_69_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_68_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2982_ _0373_ VGND VGND VPWR VPWR disp_song.um.drum.next_note1\[3\] sky130_fd_sc_hd__inv_2
XFILLER_0_68_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5770_ clknet_leaf_11_clk game.scoring_button_2.next_count\[7\] net57 VGND VGND VPWR
+ VPWR game.scoring_button_2.counts\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4721_ game.scoring_button_1.flash_counter_2\[16\] _1864_ _1830_ VGND VGND VPWR VPWR
+ _1867_ sky130_fd_sc_hd__a21boi_1
XTAP_1390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4652_ _1819_ VGND VGND VPWR VPWR game.scoring_button_1.next_count\[19\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3603_ disp_song.mi6.in\[2\] _0926_ VGND VGND VPWR VPWR _0964_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4583_ game.addmisses.a\[15\] _1773_ VGND VGND VPWR VPWR _1774_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3534_ _0887_ _0894_ _0896_ VGND VGND VPWR VPWR _0897_ sky130_fd_sc_hd__a21o_1
X_3465_ _0762_ _0824_ _0825_ _0826_ _0827_ VGND VGND VPWR VPWR _0828_ sky130_fd_sc_hd__o311a_1
XFILLER_0_58_62 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5204_ _2256_ _2290_ VGND VGND VPWR VPWR _2291_ sky130_fd_sc_hd__nand2_1
X_3396_ _0754_ _0757_ VGND VGND VPWR VPWR _0759_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5135_ disp_song.um.drum.next_note1\[30\] disp_song.um.drum.next_note1\[31\] disp_song.um.drum.next_idx1\[0\]
+ VGND VGND VPWR VPWR _2223_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5066_ _2155_ VGND VGND VPWR VPWR _2156_ sky130_fd_sc_hd__inv_2
X_4017_ _1289_ _1327_ VGND VGND VPWR VPWR _1328_ sky130_fd_sc_hd__nor2_1
X_5968_ clknet_leaf_31_clk game.scoring_button_1.next_flash_counter_2\[13\] net69
+ VGND VGND VPWR VPWR game.scoring_button_1.flash_counter_2\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4919_ _2010_ _2012_ VGND VGND VPWR VPWR _2013_ sky130_fd_sc_hd__or2_2
XFILLER_0_75_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5899_ clknet_leaf_44_clk net134 net53 VGND VGND VPWR VPWR game.out\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_110_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3250_ _0612_ _0484_ VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__nor2_1
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3181_ game.addhits.add1.b\[0\] game.addhits.a\[0\] VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__nand2_2
XFILLER_0_88_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5822_ clknet_leaf_51_clk game.scoring_button_2.next_flash_counter_2\[13\] net55
+ VGND VGND VPWR VPWR game.scoring_button_2.flash_counter_2\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5753_ clknet_leaf_66_clk game.scoring_button_2.next_num_hits\[9\] net47 VGND VGND
+ VPWR VPWR game.addhits.add3.b\[1\] sky130_fd_sc_hd__dfrtp_1
X_4704_ game.scoring_button_1.flash_counter_2\[9\] game.scoring_button_1.flash_counter_2\[10\]
+ _1847_ game.scoring_button_1.flash_counter_2\[11\] VGND VGND VPWR VPWR _1855_ sky130_fd_sc_hd__a31o_1
X_2965_ _2660_ _0357_ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__nand2_2
XFILLER_0_17_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2896_ disp_song.um.idx_note2\[0\] _0166_ disp_song.um.idx_note2\[1\] VGND VGND VPWR
+ VPWR _0310_ sky130_fd_sc_hd__or3b_1
XFILLER_0_72_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5684_ _2629_ _2645_ VGND VGND VPWR VPWR _2646_ sky130_fd_sc_hd__nand2_1
X_4635_ game.scoring_button_1.check_hit.in _1442_ _1443_ VGND VGND VPWR VPWR _1811_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_4_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_581 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4566_ game.addmisses.a\[10\] game.addmisses.a\[9\] game.addmisses.a\[8\] _1743_
+ VGND VGND VPWR VPWR _1760_ sky130_fd_sc_hd__and4_1
XFILLER_0_69_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3517_ _0552_ _0642_ VGND VGND VPWR VPWR _0880_ sky130_fd_sc_hd__or2_1
X_4497_ game.addmisses.a\[3\] _1695_ _1699_ VGND VGND VPWR VPWR _1700_ sky130_fd_sc_hd__o21ai_1
X_3448_ _0777_ _0778_ _0796_ _0810_ VGND VGND VPWR VPWR _0811_ sky130_fd_sc_hd__nor4b_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6167_ clknet_leaf_5_clk disp_song.um.drum.next_d2\[6\] net60 VGND VGND VPWR VPWR
+ disp_song.display_note2\[6\] sky130_fd_sc_hd__dfrtp_1
X_3379_ game.addhits.add4.b\[3\] VGND VGND VPWR VPWR _0742_ sky130_fd_sc_hd__inv_2
X_5118_ _2185_ _2205_ VGND VGND VPWR VPWR _2206_ sky130_fd_sc_hd__or2_1
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6098_ clknet_leaf_37_clk disp_song.um.drum.next_note1\[10\] net71 VGND VGND VPWR
+ VPWR disp_song.note1\[10\] sky130_fd_sc_hd__dfstp_1
X_5049_ disp_song.um.drum.next_idx2\[1\] _1969_ _2139_ VGND VGND VPWR VPWR _2140_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2750_ disp_song.um.idx_note1\[3\] _0186_ VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2681_ net148 disp_song.um.boton1e.edge_1 VGND VGND VPWR VPWR _2655_ sky130_fd_sc_hd__nand2b_4
XFILLER_0_26_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4420_ game.addhits.a\[4\] _1630_ VGND VGND VPWR VPWR _1636_ sky130_fd_sc_hd__or2_1
XFILLER_0_111_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4351_ game.scoring_button_2.flash_counter_1\[11\] game.scoring_button_2.flash_counter_1\[10\]
+ _1579_ VGND VGND VPWR VPWR _1583_ sky130_fd_sc_hd__and3_1
X_4282_ game.scoring_button_2.flash_counter_2\[12\] _1532_ VGND VGND VPWR VPWR _1536_
+ sky130_fd_sc_hd__or2_1
X_3302_ _0659_ _0664_ VGND VGND VPWR VPWR _0665_ sky130_fd_sc_hd__or2_2
X_6021_ clknet_leaf_59_clk _0130_ net50 VGND VGND VPWR VPWR game.flash_counter\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3233_ _0484_ _0485_ VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__nor2_1
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3164_ _0525_ _0526_ _0520_ VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__mux2_2
X_3095_ game.addmisses.a\[2\] game.addmisses.add1.b\[2\] VGND VGND VPWR VPWR _0458_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5805_ clknet_leaf_57_clk game.scoring_button_2.next_flash_counter_1\[19\] net50
+ VGND VGND VPWR VPWR game.scoring_button_2.flash_counter_1\[19\] sky130_fd_sc_hd__dfrtp_1
X_3997_ game.addmisses.add1.b\[2\] game.addmisses.add1.b\[1\] game.addmisses.add1.b\[0\]
+ game.addmisses.add1.b\[3\] VGND VGND VPWR VPWR _1311_ sky130_fd_sc_hd__o31a_1
Xfanout49 net73 VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__buf_8
X_2948_ _0307_ _0337_ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__or2_1
X_5736_ clknet_leaf_70_clk game.scoring_button_2.next_num_misses\[8\] net46 VGND VGND
+ VPWR VPWR game.addmisses.add3.b\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_44_120 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5667_ _2634_ VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4618_ _1802_ VGND VGND VPWR VPWR game.scoring_button_1.next_count\[2\] sky130_fd_sc_hd__clkbuf_1
X_2879_ _0297_ _0161_ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__nand2_2
XFILLER_0_72_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5598_ _2590_ game.padded_notes1\[30\] _2472_ VGND VGND VPWR VPWR _2591_ sky130_fd_sc_hd__mux2_1
X_4549_ _1744_ _1743_ game.addmisses.a\[8\] VGND VGND VPWR VPWR _1745_ sky130_fd_sc_hd__o21ai_1
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3920_ net167 _1227_ _1248_ _1226_ VGND VGND VPWR VPWR game.scoring_button_2.next_num_hits\[2\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_598 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3851_ _0966_ disp_song.display_note1\[1\] _0211_ game.out\[8\] _0208_ VGND VGND
+ VPWR VPWR _1197_ sky130_fd_sc_hd__a221o_2
XFILLER_0_46_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2802_ game.counter\[6\] _0222_ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3782_ highest_score.highest_score\[0\] _1056_ VGND VGND VPWR VPWR _1135_ sky130_fd_sc_hd__or2_1
XFILLER_0_109_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5521_ disp_song.note1\[5\] game.padded_notes1\[4\] _2497_ VGND VGND VPWR VPWR _2539_
+ sky130_fd_sc_hd__mux2_1
X_2733_ disp_song.um.idx_note1\[3\] VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__inv_2
XFILLER_0_81_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5452_ disp_song.note2\[17\] game.padded_notes2\[16\] _2497_ VGND VGND VPWR VPWR
+ _2498_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5383_ _2451_ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__clkbuf_1
X_4403_ _1617_ _1616_ VGND VGND VPWR VPWR _1622_ sky130_fd_sc_hd__nand2_1
X_4334_ _1571_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_1\[5\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6004_ clknet_leaf_39_clk _0113_ net66 VGND VGND VPWR VPWR game.padded_notes1\[23\]
+ sky130_fd_sc_hd__dfstp_1
X_4265_ net151 _1521_ game.missed_2 VGND VGND VPWR VPWR _1524_ sky130_fd_sc_hd__a21boi_1
X_4196_ _1405_ _1467_ VGND VGND VPWR VPWR _1468_ sky130_fd_sc_hd__and2_1
X_3216_ _0534_ _0578_ VGND VGND VPWR VPWR _0579_ sky130_fd_sc_hd__xnor2_1
X_3147_ game.addmisses.a\[14\] game.addmisses.add4.b\[2\] VGND VGND VPWR VPWR _0510_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3078_ game.addmisses.a\[8\] game.addmisses.add3.b\[0\] VGND VGND VPWR VPWR _0441_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5719_ clknet_leaf_7_clk _0043_ net59 VGND VGND VPWR VPWR pulseout.fin_pulse\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4050_ _1305_ _1351_ VGND VGND VPWR VPWR _1357_ sky130_fd_sc_hd__nor2_2
X_3001_ _0367_ _0386_ _0387_ VGND VGND VPWR VPWR disp_song.um.drum.next_note1\[8\]
+ sky130_fd_sc_hd__o21ai_1
Xinput6 n_rst VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__buf_1
XFILLER_0_78_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4952_ disp_song.um.drum.next_idx2\[0\] disp_song.um.drum.next_note2\[19\] VGND VGND
+ VPWR VPWR _2046_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4883_ disp_song.um.drum.next_note2\[22\] disp_song.um.drum.next_note2\[23\] disp_song.um.drum.next_idx2\[0\]
+ VGND VGND VPWR VPWR _1978_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_502 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_587 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3903_ game.addhits.add1.b\[2\] game.scoring_button_2.acc\[2\] VGND VGND VPWR VPWR
+ _1233_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3834_ _0879_ _1183_ VGND VGND VPWR VPWR _1184_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3765_ _1114_ _1118_ _0352_ VGND VGND VPWR VPWR _1119_ sky130_fd_sc_hd__a21oi_1
X_2716_ _0162_ VGND VGND VPWR VPWR disp_song.um.drum.next_idx2\[4\] sky130_fd_sc_hd__inv_2
X_3696_ highest_score.highest_score\[1\] VGND VGND VPWR VPWR _1052_ sky130_fd_sc_hd__inv_2
X_5504_ net269 _2460_ _2462_ net110 VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5435_ _2486_ VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5366_ _2440_ VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__clkbuf_1
X_5297_ disp_song.note1\[18\] _2232_ disp_song.um.drum.next_idx1\[1\] _2226_ VGND
+ VGND VPWR VPWR _2380_ sky130_fd_sc_hd__o22a_1
X_4317_ game.scoring_button_2.flash_counter_1\[0\] _1413_ VGND VGND VPWR VPWR _1560_
+ sky130_fd_sc_hd__and2b_1
X_4248_ game.scoring_button_2.flash_counter_2\[1\] game.scoring_button_2.flash_counter_2\[0\]
+ game.scoring_button_2.flash_counter_2\[2\] VGND VGND VPWR VPWR _1512_ sky130_fd_sc_hd__a21o_1
X_4179_ _1455_ VGND VGND VPWR VPWR game.scoring_button_2.next_count\[15\] sky130_fd_sc_hd__clkbuf_1
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_3__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_37_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3550_ _0912_ _0618_ _0614_ VGND VGND VPWR VPWR _0913_ sky130_fd_sc_hd__and3b_1
XFILLER_0_3_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3481_ _0777_ _0778_ _0796_ _0810_ VGND VGND VPWR VPWR _0844_ sky130_fd_sc_hd__or4b_2
X_5220_ disp_song.um.drum.next_idx1\[4\] _2257_ VGND VGND VPWR VPWR _2307_ sky130_fd_sc_hd__nand2_1
X_5151_ _2220_ _2225_ _2229_ _2238_ _2188_ _2216_ VGND VGND VPWR VPWR _2239_ sky130_fd_sc_hd__mux4_1
XFILLER_0_47_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5082_ _2043_ VGND VGND VPWR VPWR _2171_ sky130_fd_sc_hd__inv_2
X_4102_ _1398_ _1401_ game.addmisses.add4.b\[3\] VGND VGND VPWR VPWR _1402_ sky130_fd_sc_hd__mux2_1
X_4033_ game.addmisses.add2.b\[3\] _1334_ _1341_ _1336_ VGND VGND VPWR VPWR _1342_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_649 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5984_ clknet_leaf_33_clk _0093_ net68 VGND VGND VPWR VPWR game.padded_notes1\[3\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_47_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4935_ _1949_ _2010_ VGND VGND VPWR VPWR _2029_ sky130_fd_sc_hd__or2_1
X_4866_ disp_song.um.drum.next_idx2\[1\] _1960_ _1951_ VGND VGND VPWR VPWR _1961_
+ sky130_fd_sc_hd__a21oi_2
XFILLER_0_74_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_229 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4797_ game.scoring_button_1.flash_counter_1\[17\] game.scoring_button_1.flash_counter_1\[16\]
+ _1915_ VGND VGND VPWR VPWR _1919_ sky130_fd_sc_hd__and3_1
X_3817_ _1043_ _1049_ _1167_ _0896_ VGND VGND VPWR VPWR _1168_ sky130_fd_sc_hd__a31o_1
XFILLER_0_105_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3748_ _1090_ _1038_ _1091_ _1102_ VGND VGND VPWR VPWR _1103_ sky130_fd_sc_hd__nor4_1
XFILLER_0_104_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3679_ _1028_ _1029_ _1030_ VGND VGND VPWR VPWR _1035_ sky130_fd_sc_hd__nor3_2
X_5418_ disp_song.note2\[6\] game.padded_notes2\[5\] _0219_ VGND VGND VPWR VPWR _2475_
+ sky130_fd_sc_hd__mux2_1
X_5349_ _2423_ _2424_ _2425_ _2426_ VGND VGND VPWR VPWR _2427_ sky130_fd_sc_hd__and4b_1
XFILLER_0_97_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_50_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_50_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_53_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_78 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2981_ _0367_ _0371_ _0372_ VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__o21a_1
XFILLER_0_56_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4720_ _1866_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_2\[15\]
+ sky130_fd_sc_hd__clkbuf_1
XTAP_1380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_41_clk clknet_3_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_41_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_8_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4651_ _1791_ _1467_ VGND VGND VPWR VPWR _1819_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3602_ _0211_ _0961_ _0962_ net39 VGND VGND VPWR VPWR _0963_ sky130_fd_sc_hd__o211a_1
X_4582_ _1771_ _1772_ VGND VGND VPWR VPWR _1773_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3533_ _0255_ _0895_ VGND VGND VPWR VPWR _0896_ sky130_fd_sc_hd__or2_2
XFILLER_0_52_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3464_ _0817_ VGND VGND VPWR VPWR _0827_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5203_ disp_song.note1\[8\] _0175_ VGND VGND VPWR VPWR _2290_ sky130_fd_sc_hd__or2_1
X_5134_ _2191_ _2221_ disp_song.um.drum.next_idx1\[2\] VGND VGND VPWR VPWR _2222_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_58_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3395_ _0754_ _0757_ VGND VGND VPWR VPWR _0758_ sky130_fd_sc_hd__nor2_1
X_5065_ _2679_ _2012_ _0162_ VGND VGND VPWR VPWR _2155_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4016_ game.addmisses.add2.b\[0\] _1311_ VGND VGND VPWR VPWR _1327_ sky130_fd_sc_hd__and2_1
X_5967_ clknet_leaf_35_clk game.scoring_button_1.next_flash_counter_2\[12\] net72
+ VGND VGND VPWR VPWR game.scoring_button_1.flash_counter_2\[12\] sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_32_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_32_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_90_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4918_ disp_song.um.drum.next_idx2\[2\] _2009_ VGND VGND VPWR VPWR _2012_ sky130_fd_sc_hd__nor2_2
X_5898_ clknet_leaf_26_clk _0081_ net68 VGND VGND VPWR VPWR game.padded_notes2\[31\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_74_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4849_ _0352_ _1945_ VGND VGND VPWR VPWR _1946_ sky130_fd_sc_hd__or2_1
XFILLER_0_99_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_23_clk clknet_3_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_23_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_38_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_571 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3180_ _0541_ _0542_ VGND VGND VPWR VPWR _0543_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5821_ clknet_leaf_51_clk game.scoring_button_2.next_flash_counter_2\[12\] net55
+ VGND VGND VPWR VPWR game.scoring_button_2.flash_counter_2\[12\] sky130_fd_sc_hd__dfrtp_1
X_2964_ _2657_ _0357_ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__nand2_1
X_5752_ clknet_leaf_66_clk game.scoring_button_2.next_num_hits\[8\] net46 VGND VGND
+ VPWR VPWR game.addhits.add3.b\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4703_ game.scoring_button_1.flash_counter_2\[11\] game.scoring_button_1.flash_counter_2\[10\]
+ _1850_ VGND VGND VPWR VPWR _1854_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_14_clk clknet_3_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_14_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_72_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2895_ _0309_ VGND VGND VPWR VPWR disp_song.um.drum.next_note2\[13\] sky130_fd_sc_hd__buf_1
X_5683_ game.flash_counter\[20\] game.flash_counter\[21\] _2644_ VGND VGND VPWR VPWR
+ _2645_ sky130_fd_sc_hd__and3_1
X_4634_ _1810_ VGND VGND VPWR VPWR game.scoring_button_1.next_count\[10\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_102_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_593 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4565_ game.addmisses.a\[9\] game.addmisses.a\[8\] _1743_ _1716_ game.addmisses.a\[10\]
+ VGND VGND VPWR VPWR _1759_ sky130_fd_sc_hd__a32o_1
XFILLER_0_40_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3516_ _0209_ modetrans.mode\[4\] VGND VGND VPWR VPWR _0879_ sky130_fd_sc_hd__nor2_2
XFILLER_0_40_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4496_ game.scoring_button_1.hit _1673_ VGND VGND VPWR VPWR _1699_ sky130_fd_sc_hd__nor2_4
XFILLER_0_0_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3447_ _0798_ _0801_ _0803_ _0809_ VGND VGND VPWR VPWR _0810_ sky130_fd_sc_hd__and4b_1
X_6166_ clknet_leaf_22_clk disp_song.um.drum.next_d2\[5\] net61 VGND VGND VPWR VPWR
+ disp_song.display_note2\[5\] sky130_fd_sc_hd__dfrtp_1
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3378_ game.addhits.a\[15\] VGND VGND VPWR VPWR _0741_ sky130_fd_sc_hd__inv_2
X_6097_ clknet_leaf_37_clk disp_song.um.drum.next_note1\[9\] net67 VGND VGND VPWR
+ VPWR disp_song.note1\[9\] sky130_fd_sc_hd__dfrtp_1
X_5117_ disp_song.um.drum.next_note1\[8\] disp_song.um.drum.next_note1\[9\] _0176_
+ VGND VGND VPWR VPWR _2205_ sky130_fd_sc_hd__mux2_1
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5048_ _2666_ _1968_ _1966_ VGND VGND VPWR VPWR _2139_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_630 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_105_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2680_ modetrans.mode\[2\] VGND VGND VPWR VPWR _2654_ sky130_fd_sc_hd__buf_6
XFILLER_0_26_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_552 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4350_ net156 _1579_ _1582_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_1\[10\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_111_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3301_ _0660_ _0663_ VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__and2b_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4281_ game.scoring_button_2.flash_counter_2\[12\] _1532_ VGND VGND VPWR VPWR _1535_
+ sky130_fd_sc_hd__and2_1
X_3232_ _0504_ _0528_ _0594_ VGND VGND VPWR VPWR _0595_ sky130_fd_sc_hd__a21oi_2
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6020_ clknet_leaf_59_clk _0129_ net51 VGND VGND VPWR VPWR game.flash_counter\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_3_clk clknet_3_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_3_clk sky130_fd_sc_hd__clkbuf_16
X_3163_ _0525_ _0522_ VGND VGND VPWR VPWR _0526_ sky130_fd_sc_hd__nand2_1
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3094_ game.addmisses.a\[2\] game.addmisses.add1.b\[2\] VGND VGND VPWR VPWR _0457_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5804_ clknet_leaf_56_clk game.scoring_button_2.next_flash_counter_1\[18\] net51
+ VGND VGND VPWR VPWR game.scoring_button_2.flash_counter_1\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3996_ game.addmisses.add1.b\[1\] _1307_ _1309_ _1305_ VGND VGND VPWR VPWR _1310_
+ sky130_fd_sc_hd__o2bb2a_1
X_2947_ _2655_ _0339_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5735_ clknet_leaf_72_clk game.scoring_button_2.next_num_misses\[7\] net48 VGND VGND
+ VPWR VPWR game.addmisses.add2.b\[3\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_44_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5666_ _2632_ _2633_ VGND VGND VPWR VPWR _2634_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4617_ _1791_ _0024_ VGND VGND VPWR VPWR _1802_ sky130_fd_sc_hd__and2_1
X_2878_ _2673_ _2674_ VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5597_ disp_song.note1\[30\] game.padded_notes1\[29\] _0209_ VGND VGND VPWR VPWR
+ _2590_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4548_ modetrans.mode\[0\] _1691_ VGND VGND VPWR VPWR _1744_ sky130_fd_sc_hd__and2_1
X_4479_ game.scoring_button_1.counts\[7\] game.scoring_button_1.counts\[8\] _1680_
+ game.scoring_button_1.counts\[9\] VGND VGND VPWR VPWR _1683_ sky130_fd_sc_hd__a31o_1
XFILLER_0_99_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6149_ clknet_leaf_28_clk disp_song.um.drum.next_note2\[29\] net68 VGND VGND VPWR
+ VPWR disp_song.note2\[29\] sky130_fd_sc_hd__dfstp_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3850_ _1196_ VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
X_2801_ _0231_ VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_73_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3781_ _1069_ _1133_ VGND VGND VPWR VPWR _1134_ sky130_fd_sc_hd__and2b_1
X_5520_ _2538_ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__clkbuf_1
X_2732_ _0176_ VGND VGND VPWR VPWR disp_song.um.drum.next_idx1\[0\] sky130_fd_sc_hd__clkbuf_8
XFILLER_0_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5451_ _0209_ VGND VGND VPWR VPWR _2497_ sky130_fd_sc_hd__buf_8
X_5382_ _0206_ _2449_ _2450_ VGND VGND VPWR VPWR _2451_ sky130_fd_sc_hd__and3_1
X_4402_ game.addhits.a\[3\] _1620_ VGND VGND VPWR VPWR _1621_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4333_ _1569_ game.hit_2 _1570_ VGND VGND VPWR VPWR _1571_ sky130_fd_sc_hd__and3b_1
X_4264_ _1523_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_2\[6\]
+ sky130_fd_sc_hd__clkbuf_1
X_6003_ clknet_leaf_38_clk _0112_ net66 VGND VGND VPWR VPWR game.padded_notes1\[22\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3215_ _0537_ _0576_ _0577_ _0535_ VGND VGND VPWR VPWR _0578_ sky130_fd_sc_hd__a31o_1
X_4195_ _1465_ _1466_ VGND VGND VPWR VPWR _1467_ sky130_fd_sc_hd__nor2_1
X_3146_ game.addmisses.a\[14\] game.addmisses.add4.b\[2\] VGND VGND VPWR VPWR _0509_
+ sky130_fd_sc_hd__and2_1
X_3077_ _0438_ _0439_ VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_10_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3979_ game.scoring_button_2.counts\[2\] game.scoring_button_2.counts\[1\] game.scoring_button_2.counts\[0\]
+ _1293_ VGND VGND VPWR VPWR _1294_ sky130_fd_sc_hd__or4_2
X_5718_ clknet_leaf_22_clk _0008_ net59 VGND VGND VPWR VPWR modetrans.mode\[5\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_103_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5649_ game.flash_counter\[12\] game.flash_counter\[11\] _2620_ VGND VGND VPWR VPWR
+ _2621_ sky130_fd_sc_hd__and3_1
XFILLER_0_103_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3000_ _0368_ _0386_ net247 VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_36_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_522 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4951_ _1956_ disp_song.um.drum.next_note2\[16\] _2043_ _2044_ VGND VGND VPWR VPWR
+ _2045_ sky130_fd_sc_hd__o211a_1
X_4882_ _1976_ _2666_ _1965_ VGND VGND VPWR VPWR _1977_ sky130_fd_sc_hd__and3b_1
XFILLER_0_86_385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3902_ game.addhits.add1.b\[0\] _1230_ _1231_ VGND VGND VPWR VPWR _1232_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_6_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3833_ _1180_ _1181_ _1182_ _0921_ VGND VGND VPWR VPWR _1183_ sky130_fd_sc_hd__a31o_1
XFILLER_0_27_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3764_ _1079_ _1082_ _1115_ _1117_ _0925_ VGND VGND VPWR VPWR _1118_ sky130_fd_sc_hd__a32o_1
XFILLER_0_14_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2715_ _2654_ _0156_ _2662_ _0161_ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__a31o_4
XFILLER_0_14_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3695_ _1042_ _1050_ _0896_ VGND VGND VPWR VPWR _1051_ sky130_fd_sc_hd__a21o_1
X_5503_ net117 _2460_ _2462_ game.out\[12\] VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__a22o_1
X_5434_ _2485_ game.padded_notes2\[11\] _2473_ VGND VGND VPWR VPWR _2486_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5365_ _2439_ highest_score.highest_score\[3\] _2434_ VGND VGND VPWR VPWR _2440_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4316_ net87 _1556_ _1559_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_2\[22\]
+ sky130_fd_sc_hd__a21oi_1
X_5296_ _0191_ _0197_ _2244_ _0185_ VGND VGND VPWR VPWR _2379_ sky130_fd_sc_hd__a31o_1
X_4247_ game.scoring_button_2.flash_counter_2\[1\] game.scoring_button_2.flash_counter_2\[0\]
+ game.scoring_button_2.flash_counter_2\[2\] VGND VGND VPWR VPWR _1511_ sky130_fd_sc_hd__and3_1
X_4178_ _1405_ _1454_ VGND VGND VPWR VPWR _1455_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3129_ _0488_ _0491_ VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__xnor2_2
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3480_ _0781_ _0814_ _0818_ _0804_ VGND VGND VPWR VPWR _0843_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_51_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5150_ _2235_ _2237_ VGND VGND VPWR VPWR _2238_ sky130_fd_sc_hd__nor2_1
X_5081_ _2156_ _2163_ _2170_ _0214_ VGND VGND VPWR VPWR disp_song.um.drum.next_d2\[5\]
+ sky130_fd_sc_hd__o211a_1
X_4101_ game.addmisses.add4.b\[2\] game.addmisses.add4.b\[1\] _1379_ VGND VGND VPWR
+ VPWR _1401_ sky130_fd_sc_hd__or3_1
X_4032_ _1335_ VGND VGND VPWR VPWR _1341_ sky130_fd_sc_hd__inv_2
X_5983_ clknet_leaf_26_clk _0092_ net68 VGND VGND VPWR VPWR game.padded_notes1\[2\]
+ sky130_fd_sc_hd__dfstp_1
X_4934_ disp_song.note2\[24\] _1956_ VGND VGND VPWR VPWR _2028_ sky130_fd_sc_hd__or2_1
XFILLER_0_87_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4865_ _2679_ _0169_ VGND VGND VPWR VPWR _1960_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3816_ _1166_ VGND VGND VPWR VPWR _1167_ sky130_fd_sc_hd__inv_2
X_4796_ net180 _1915_ _1918_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_1\[16\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_103_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3747_ modetrans.mode\[3\] _1101_ _0211_ VGND VGND VPWR VPWR _1102_ sky130_fd_sc_hd__a21oi_1
X_3678_ _1012_ _1028_ VGND VGND VPWR VPWR _1034_ sky130_fd_sc_hd__or2_2
XFILLER_0_42_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5417_ _2474_ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5348_ highest_score.highest_score\[5\] _0840_ VGND VGND VPWR VPWR _2426_ sky130_fd_sc_hd__or2_1
X_5279_ disp_song.note1\[2\] _2232_ _0191_ _2362_ VGND VGND VPWR VPWR _2363_ sky130_fd_sc_hd__a211o_1
XFILLER_0_65_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2980_ _0368_ _0371_ disp_song.note1\[3\] VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__o21ai_1
XTAP_1381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4650_ _1818_ VGND VGND VPWR VPWR game.scoring_button_1.next_count\[18\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3601_ _0840_ _0859_ _0946_ VGND VGND VPWR VPWR _0962_ sky130_fd_sc_hd__or3_1
XFILLER_0_71_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4581_ game.addmisses.a\[13\] _1765_ VGND VGND VPWR VPWR _1772_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3532_ _0258_ VGND VGND VPWR VPWR _0895_ sky130_fd_sc_hd__inv_2
X_3463_ _0774_ _0822_ _0823_ _0778_ _0777_ VGND VGND VPWR VPWR _0826_ sky130_fd_sc_hd__o32a_4
X_5202_ disp_song.um.drum.next_note1\[9\] _2261_ _2185_ VGND VGND VPWR VPWR _2289_
+ sky130_fd_sc_hd__a21oi_1
X_5133_ disp_song.um.drum.next_note1\[28\] disp_song.um.drum.next_note1\[29\] disp_song.um.drum.next_idx1\[0\]
+ VGND VGND VPWR VPWR _2221_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3394_ _0527_ _0756_ VGND VGND VPWR VPWR _0757_ sky130_fd_sc_hd__and2_1
X_5064_ _0352_ _2154_ VGND VGND VPWR VPWR disp_song.um.drum.next_d2\[4\] sky130_fd_sc_hd__nor2_1
X_4015_ game.addmisses.add2.b\[0\] _1311_ VGND VGND VPWR VPWR _1326_ sky130_fd_sc_hd__or2_1
X_5966_ clknet_leaf_35_clk game.scoring_button_1.next_flash_counter_2\[11\] net72
+ VGND VGND VPWR VPWR game.scoring_button_1.flash_counter_2\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5897_ clknet_leaf_31_clk _0080_ net69 VGND VGND VPWR VPWR game.padded_notes2\[30\]
+ sky130_fd_sc_hd__dfrtp_1
X_4917_ disp_song.um.drum.next_idx2\[3\] _2010_ disp_song.um.drum.next_idx2\[4\] VGND
+ VGND VPWR VPWR _2011_ sky130_fd_sc_hd__o21a_1
XFILLER_0_90_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4848_ disp_song.um.idx_note1\[3\] disp_song.um.idx_note2\[3\] _2661_ VGND VGND VPWR
+ VPWR _1945_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4779_ _1905_ game.hit_1 _1906_ VGND VGND VPWR VPWR _1907_ sky130_fd_sc_hd__and3b_1
XFILLER_0_99_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_601 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_583 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_104_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5820_ clknet_leaf_50_clk game.scoring_button_2.next_flash_counter_2\[11\] net55
+ VGND VGND VPWR VPWR game.scoring_button_2.flash_counter_2\[11\] sky130_fd_sc_hd__dfrtp_1
X_2963_ _0183_ _0356_ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__and2_2
XFILLER_0_29_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5751_ clknet_leaf_3_clk game.scoring_button_2.next_num_hits\[7\] net49 VGND VGND
+ VPWR VPWR game.addhits.add2.b\[3\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_56_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4702_ net158 _1850_ _1853_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_2\[10\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_72_612 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2894_ disp_song.note2\[13\] _0269_ _0308_ VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5682_ game.flash_counter\[19\] game.flash_counter\[18\] game.flash_counter\[17\]
+ game.flash_counter\[16\] VGND VGND VPWR VPWR _2644_ sky130_fd_sc_hd__and4_1
X_4633_ _1791_ _1440_ VGND VGND VPWR VPWR _1810_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4564_ _1750_ _1757_ _1755_ game.addmisses.a\[11\] VGND VGND VPWR VPWR _1758_ sky130_fd_sc_hd__a2bb2o_1
X_3515_ game.flash_counter\[23\] _0867_ _0877_ _0842_ VGND VGND VPWR VPWR _0878_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_4_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4495_ _1695_ _1697_ VGND VGND VPWR VPWR _1698_ sky130_fd_sc_hd__and2_1
X_3446_ _0784_ _0804_ _0808_ VGND VGND VPWR VPWR _0809_ sky130_fd_sc_hd__or3_1
X_6165_ clknet_leaf_8_clk disp_song.um.drum.next_d2\[4\] net61 VGND VGND VPWR VPWR
+ disp_song.display_note2\[4\] sky130_fd_sc_hd__dfrtp_1
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3377_ game.addhits.a\[15\] game.addhits.add4.b\[3\] VGND VGND VPWR VPWR _0740_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6096_ clknet_leaf_41_clk disp_song.um.drum.next_note1\[8\] net67 VGND VGND VPWR
+ VPWR disp_song.note1\[8\] sky130_fd_sc_hd__dfrtp_1
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5116_ _2191_ _2203_ disp_song.um.drum.next_idx1\[1\] VGND VGND VPWR VPWR _2204_
+ sky130_fd_sc_hd__a21o_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5047_ _2138_ VGND VGND VPWR VPWR disp_song.um.drum.next_d2\[3\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5949_ clknet_leaf_45_clk game.scoring_button_1.next_flash_counter_1\[17\] net53
+ VGND VGND VPWR VPWR game.scoring_button_1.flash_counter_1\[17\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_35 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3300_ _0661_ _0662_ VGND VGND VPWR VPWR _0663_ sky130_fd_sc_hd__nand2_1
X_4280_ _1534_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_2\[11\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_44 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3231_ _0531_ _0593_ VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__xor2_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3162_ _0514_ _0512_ VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__or2_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3093_ _0450_ _0455_ _0451_ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__o21a_2
XFILLER_0_71_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5803_ clknet_leaf_56_clk game.scoring_button_2.next_flash_counter_1\[17\] net51
+ VGND VGND VPWR VPWR game.scoring_button_2.flash_counter_1\[17\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3995_ game.addmisses.add1.b\[1\] game.addmisses.add1.b\[0\] VGND VGND VPWR VPWR
+ _1309_ sky130_fd_sc_hd__xnor2_1
X_2946_ _0269_ _0164_ _0334_ _0344_ VGND VGND VPWR VPWR disp_song.um.drum.next_note2\[28\]
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_29_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5734_ clknet_leaf_73_clk game.scoring_button_2.next_num_misses\[6\] net48 VGND VGND
+ VPWR VPWR game.addmisses.add2.b\[2\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_44_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2877_ _0296_ VGND VGND VPWR VPWR disp_song.um.drum.next_note2\[8\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5665_ game.flash_counter\[16\] _2629_ VGND VGND VPWR VPWR _2633_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4616_ _1801_ VGND VGND VPWR VPWR game.scoring_button_1.next_count\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5596_ _2589_ VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__clkbuf_1
X_4547_ _1691_ _1737_ VGND VGND VPWR VPWR _1743_ sky130_fd_sc_hd__nor2_2
X_4478_ game.scoring_button_1.counts\[7\] game.scoring_button_1.counts\[11\] _1680_
+ _1681_ VGND VGND VPWR VPWR _1682_ sky130_fd_sc_hd__or4_1
XFILLER_0_96_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3429_ _0791_ VGND VGND VPWR VPWR _0792_ sky130_fd_sc_hd__inv_2
X_6148_ clknet_leaf_27_clk disp_song.um.drum.next_note2\[28\] net68 VGND VGND VPWR
+ VPWR disp_song.note2\[28\] sky130_fd_sc_hd__dfrtp_1
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6079_ clknet_leaf_40_clk disp_song.um.drum.next_idx1\[1\] net66 VGND VGND VPWR VPWR
+ disp_song.um.idx_note1\[1\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2800_ _0225_ _0228_ _0229_ _0230_ VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__or4b_1
X_3780_ _1092_ _1132_ _1071_ VGND VGND VPWR VPWR _1133_ sky130_fd_sc_hd__o21ai_1
X_2731_ _0175_ VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__inv_2
X_5450_ _2496_ VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4401_ _1615_ _1618_ _1619_ VGND VGND VPWR VPWR _1620_ sky130_fd_sc_hd__o21ai_1
X_5381_ pulseout.fin_pulse\[0\] game.beat_clk pulseout.fin_pulse\[1\] VGND VGND VPWR
+ VPWR _2450_ sky130_fd_sc_hd__a21o_1
XFILLER_0_1_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4332_ game.scoring_button_2.flash_counter_1\[3\] game.scoring_button_2.flash_counter_1\[4\]
+ _1562_ game.scoring_button_2.flash_counter_1\[5\] VGND VGND VPWR VPWR _1570_ sky130_fd_sc_hd__a31o_1
X_4263_ _1521_ _1486_ _1522_ VGND VGND VPWR VPWR _1523_ sky130_fd_sc_hd__and3b_1
X_6002_ clknet_leaf_39_clk _0111_ net67 VGND VGND VPWR VPWR game.padded_notes1\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3214_ _0569_ _0571_ _0573_ VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__or3_1
X_4194_ game.counter\[19\] game.counter\[18\] _1461_ VGND VGND VPWR VPWR _1466_ sky130_fd_sc_hd__and3_1
X_3145_ _0505_ _0506_ _0507_ VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__a21oi_2
X_3076_ game.addmisses.a\[9\] game.addmisses.add3.b\[1\] VGND VGND VPWR VPWR _0439_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_82_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_217 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3978_ game.scoring_button_2.counts\[6\] game.scoring_button_2.counts\[5\] game.scoring_button_2.counts\[3\]
+ game.scoring_button_2.counts\[4\] VGND VGND VPWR VPWR _1293_ sky130_fd_sc_hd__or4_1
XFILLER_0_9_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2929_ _0291_ _0330_ _0332_ net236 VGND VGND VPWR VPWR disp_song.um.drum.next_note2\[23\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5717_ clknet_leaf_5_clk _0007_ net59 VGND VGND VPWR VPWR modetrans.mode\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5648_ game.flash_counter\[10\] game.flash_counter\[6\] game.flash_counter\[7\] VGND
+ VGND VPWR VPWR _2620_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5579_ disp_song.note1\[24\] game.padded_notes1\[23\] _2541_ VGND VGND VPWR VPWR
+ _2578_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_106_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4950_ disp_song.note2\[17\] _2670_ VGND VGND VPWR VPWR _2044_ sky130_fd_sc_hd__or2_1
XFILLER_0_59_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4881_ _2669_ disp_song.um.drum.next_note2\[31\] _1975_ VGND VGND VPWR VPWR _1976_
+ sky130_fd_sc_hd__o21ai_1
X_3901_ game.addhits.add1.b\[1\] game.scoring_button_2.acc\[1\] VGND VGND VPWR VPWR
+ _1231_ sky130_fd_sc_hd__nand2_1
XFILLER_0_86_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3832_ _1061_ _1098_ _1169_ _0258_ VGND VGND VPWR VPWR _1182_ sky130_fd_sc_hd__a31o_1
X_3763_ disp_song.mi6.in\[3\] _1116_ VGND VGND VPWR VPWR _1117_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5502_ game.out\[10\] _2460_ _2462_ net117 VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__a22o_1
X_2714_ _2654_ _2676_ _0160_ VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__and3_1
X_3694_ _0638_ _1043_ _1045_ _1049_ VGND VGND VPWR VPWR _1050_ sky130_fd_sc_hd__o211a_1
X_5433_ disp_song.note2\[11\] game.padded_notes2\[10\] _0219_ VGND VGND VPWR VPWR
+ _2485_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_607 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5364_ _1024_ VGND VGND VPWR VPWR _2439_ sky130_fd_sc_hd__inv_2
X_4315_ net87 _1556_ game.missed_2 VGND VGND VPWR VPWR _1559_ sky130_fd_sc_hd__o21ai_1
X_5295_ _2378_ VGND VGND VPWR VPWR disp_song.um.drum.next_d1\[4\] sky130_fd_sc_hd__clkbuf_1
X_4246_ net107 game.scoring_button_2.flash_counter_2\[0\] _1510_ VGND VGND VPWR VPWR
+ game.scoring_button_2.next_flash_counter_2\[1\] sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4177_ _0240_ _1451_ VGND VGND VPWR VPWR _1454_ sky130_fd_sc_hd__xnor2_1
X_3128_ _0489_ _0490_ VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__or2b_1
XFILLER_0_97_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3059_ _0362_ _0426_ net154 VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_77_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_65_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_83_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_559 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5080_ _2157_ _2164_ _2167_ _2169_ VGND VGND VPWR VPWR _2170_ sky130_fd_sc_hd__o31ai_1
X_4100_ _1400_ VGND VGND VPWR VPWR game.scoring_button_2.next_num_misses\[14\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4031_ net45 _1338_ _1340_ VGND VGND VPWR VPWR game.scoring_button_2.next_num_misses\[5\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5982_ clknet_leaf_26_clk _0091_ net68 VGND VGND VPWR VPWR game.padded_notes1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4933_ _1965_ _2023_ _2024_ _2026_ VGND VGND VPWR VPWR _2027_ sky130_fd_sc_hd__a31o_1
X_4864_ _1955_ _1958_ disp_song.um.drum.next_idx2\[1\] VGND VGND VPWR VPWR _1959_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3815_ _0642_ _0638_ _1040_ _1041_ VGND VGND VPWR VPWR _1166_ sky130_fd_sc_hd__a31o_1
X_4795_ net180 _1915_ _1799_ VGND VGND VPWR VPWR _1918_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_103_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3746_ _0261_ _1094_ _1097_ _0941_ _1100_ VGND VGND VPWR VPWR _1101_ sky130_fd_sc_hd__a221o_1
X_5416_ _2471_ game.padded_notes2\[5\] _2473_ VGND VGND VPWR VPWR _2474_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3677_ _1021_ _1022_ _1024_ VGND VGND VPWR VPWR _1033_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_10_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5347_ highest_score.highest_score\[6\] _0858_ VGND VGND VPWR VPWR _2425_ sky130_fd_sc_hd__xnor2_1
X_5278_ _2232_ _0373_ VGND VGND VPWR VPWR _2362_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4229_ game.counter\[9\] _0243_ game.counter\[14\] VGND VGND VPWR VPWR _1496_ sky130_fd_sc_hd__a21o_1
Xmax_cap37 _2610_ VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__buf_1
XFILLER_0_69_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4580_ game.addmisses.a\[12\] game.addmisses.a\[13\] _1749_ VGND VGND VPWR VPWR _1771_
+ sky130_fd_sc_hd__and3_1
X_3600_ _0957_ _0960_ _0921_ VGND VGND VPWR VPWR _0961_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_109_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3531_ _0888_ _0892_ _0893_ VGND VGND VPWR VPWR _0894_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3462_ _0776_ _0798_ VGND VGND VPWR VPWR _0825_ sky130_fd_sc_hd__and2_2
XFILLER_0_110_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5201_ disp_song.note1\[10\] _2232_ _2287_ VGND VGND VPWR VPWR _2288_ sky130_fd_sc_hd__o21ai_1
X_3393_ _0512_ _0755_ VGND VGND VPWR VPWR _0756_ sky130_fd_sc_hd__xnor2_1
X_5132_ _2218_ _2219_ disp_song.um.drum.next_idx1\[1\] VGND VGND VPWR VPWR _2220_
+ sky130_fd_sc_hd__mux2_1
X_5063_ _2146_ _2152_ _2153_ VGND VGND VPWR VPWR _2154_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_404 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4014_ _1323_ _1324_ _1325_ _1289_ VGND VGND VPWR VPWR game.scoring_button_2.next_num_misses\[3\]
+ sky130_fd_sc_hd__a22o_1
X_5965_ clknet_leaf_35_clk game.scoring_button_1.next_flash_counter_2\[10\] net72
+ VGND VGND VPWR VPWR game.scoring_button_1.flash_counter_2\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5896_ clknet_leaf_32_clk _0079_ net68 VGND VGND VPWR VPWR game.padded_notes2\[29\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_90_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4916_ disp_song.um.drum.next_idx2\[2\] _2009_ VGND VGND VPWR VPWR _2010_ sky130_fd_sc_hd__and2_2
XFILLER_0_90_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4847_ net266 _0325_ _0366_ disp_song.um.idx_note1\[2\] VGND VGND VPWR VPWR disp_song.um.next_position\[2\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_47_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4778_ game.scoring_button_1.flash_counter_1\[9\] game.scoring_button_1.flash_counter_1\[10\]
+ _1898_ game.scoring_button_1.flash_counter_1\[11\] VGND VGND VPWR VPWR _1906_ sky130_fd_sc_hd__a31o_1
XFILLER_0_43_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3729_ _1077_ _1080_ _1083_ _1084_ _0925_ VGND VGND VPWR VPWR _1085_ sky130_fd_sc_hd__o221a_1
XFILLER_0_100_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2962_ disp_song.um.idx_note1\[4\] _0182_ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__nand2_1
X_5750_ clknet_leaf_2_clk game.scoring_button_2.next_num_hits\[6\] net48 VGND VGND
+ VPWR VPWR game.addhits.add2.b\[2\] sky130_fd_sc_hd__dfrtp_2
X_4701_ net158 _1850_ game.missed_1 VGND VGND VPWR VPWR _1853_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_84_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5681_ _2604_ _2638_ _2642_ net175 VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_17_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2893_ _0307_ _0298_ VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__nor2_1
X_4632_ _1809_ VGND VGND VPWR VPWR game.scoring_button_1.next_count\[9\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4563_ _1755_ _1756_ VGND VGND VPWR VPWR _1757_ sky130_fd_sc_hd__or2_1
XFILLER_0_40_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3514_ _0868_ _0870_ _0876_ VGND VGND VPWR VPWR _0877_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4494_ game.addmisses.a\[2\] game.addmisses.a\[1\] game.addmisses.a\[0\] game.addmisses.a\[3\]
+ VGND VGND VPWR VPWR _1697_ sky130_fd_sc_hd__o31a_1
XFILLER_0_100_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3445_ _0806_ _0807_ VGND VGND VPWR VPWR _0808_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6164_ clknet_leaf_22_clk disp_song.um.drum.next_d2\[3\] net61 VGND VGND VPWR VPWR
+ disp_song.display_note2\[3\] sky130_fd_sc_hd__dfrtp_1
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3376_ _0738_ _0730_ VGND VGND VPWR VPWR _0739_ sky130_fd_sc_hd__nand2_1
X_6095_ clknet_leaf_37_clk disp_song.um.drum.next_note1\[7\] net71 VGND VGND VPWR
+ VPWR disp_song.note1\[7\] sky130_fd_sc_hd__dfstp_1
X_5115_ disp_song.um.drum.next_note1\[10\] disp_song.um.drum.next_note1\[11\] disp_song.um.drum.next_idx1\[0\]
+ VGND VGND VPWR VPWR _2203_ sky130_fd_sc_hd__mux2_1
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5046_ _0214_ _2131_ _2137_ VGND VGND VPWR VPWR _2138_ sky130_fd_sc_hd__and3_1
XFILLER_0_33_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5948_ clknet_leaf_45_clk game.scoring_button_1.next_flash_counter_1\[16\] net54
+ VGND VGND VPWR VPWR game.scoring_button_1.flash_counter_1\[16\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5879_ clknet_leaf_19_clk _0062_ net63 VGND VGND VPWR VPWR game.padded_notes2\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_542 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3230_ _0591_ _0592_ VGND VGND VPWR VPWR _0593_ sky130_fd_sc_hd__xor2_2
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3161_ _0514_ _0523_ VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__xnor2_2
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3092_ game.addmisses.a\[1\] game.addmisses.add1.b\[1\] VGND VGND VPWR VPWR _0455_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5802_ clknet_leaf_56_clk game.scoring_button_2.next_flash_counter_1\[16\] net51
+ VGND VGND VPWR VPWR game.scoring_button_2.flash_counter_1\[16\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3994_ game.addmisses.add1.b\[0\] _1289_ _1307_ _1308_ VGND VGND VPWR VPWR game.scoring_button_2.next_num_misses\[0\]
+ sky130_fd_sc_hd__a31o_1
X_2945_ _0163_ _0337_ disp_song.note2\[28\] VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__o21a_1
XFILLER_0_91_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5733_ clknet_leaf_72_clk game.scoring_button_2.next_num_misses\[5\] net48 VGND VGND
+ VPWR VPWR game.addmisses.add2.b\[1\] sky130_fd_sc_hd__dfrtp_4
X_2876_ _0269_ disp_song.note2\[8\] _0295_ VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__mux2_1
X_5664_ game.flash_counter\[16\] _2629_ VGND VGND VPWR VPWR _2632_ sky130_fd_sc_hd__or2_1
X_4615_ game.scoring_button_1.check_hit.in _0248_ _1415_ VGND VGND VPWR VPWR _1801_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_60_638 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5595_ _2588_ net223 _2472_ VGND VGND VPWR VPWR _2589_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4546_ _1741_ VGND VGND VPWR VPWR _1742_ sky130_fd_sc_hd__inv_2
XFILLER_0_110_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4477_ game.scoring_button_1.counts\[10\] game.scoring_button_1.counts\[9\] game.scoring_button_1.counts\[8\]
+ game.scoring_button_1.counts\[15\] VGND VGND VPWR VPWR _1681_ sky130_fd_sc_hd__or4_1
X_3428_ _0682_ _0693_ VGND VGND VPWR VPWR _0791_ sky130_fd_sc_hd__xnor2_2
X_6147_ clknet_leaf_26_clk disp_song.um.drum.next_note2\[27\] net68 VGND VGND VPWR
+ VPWR disp_song.note2\[27\] sky130_fd_sc_hd__dfstp_1
X_3359_ _0714_ _0720_ _0718_ VGND VGND VPWR VPWR _0722_ sky130_fd_sc_hd__a21o_1
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6078_ clknet_leaf_40_clk disp_song.um.drum.next_idx1\[0\] net66 VGND VGND VPWR VPWR
+ disp_song.um.idx_note1\[0\] sky130_fd_sc_hd__dfstp_4
X_5029_ disp_song.note2\[19\] disp_song.um.drum.next_idx2\[0\] _2047_ _2043_ VGND
+ VGND VPWR VPWR _2121_ sky130_fd_sc_hd__o211a_1
XFILLER_0_75_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2730_ _0174_ VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__buf_4
XFILLER_0_14_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4400_ game.addhits.a\[2\] game.scoring_button_1.acc\[2\] VGND VGND VPWR VPWR _1619_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5380_ pulseout.fin_pulse\[0\] pulseout.fin_pulse\[1\] game.beat_clk VGND VGND VPWR
+ VPWR _2449_ sky130_fd_sc_hd__nand3_1
XFILLER_0_1_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4331_ game.scoring_button_2.flash_counter_1\[5\] game.scoring_button_2.flash_counter_1\[4\]
+ _1565_ VGND VGND VPWR VPWR _1569_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4262_ game.scoring_button_2.flash_counter_2\[6\] _1518_ VGND VGND VPWR VPWR _1522_
+ sky130_fd_sc_hd__or2_1
X_6001_ clknet_leaf_38_clk _0110_ net67 VGND VGND VPWR VPWR game.padded_notes1\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3213_ _0569_ _0574_ _0575_ VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__o21bai_4
X_4193_ game.counter\[18\] _1461_ game.counter\[19\] VGND VGND VPWR VPWR _1465_ sky130_fd_sc_hd__a21oi_1
X_3144_ game.addmisses.a\[13\] game.addmisses.add4.b\[1\] VGND VGND VPWR VPWR _0507_
+ sky130_fd_sc_hd__and2_1
X_3075_ game.addmisses.a\[9\] game.addmisses.add3.b\[1\] VGND VGND VPWR VPWR _0438_
+ sky130_fd_sc_hd__nand2_1
X_3977_ game.scoring_button_2.counts\[9\] game.scoring_button_2.counts\[8\] game.scoring_button_2.counts\[7\]
+ _1291_ VGND VGND VPWR VPWR _1292_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2928_ _0313_ _0327_ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__or2_1
X_5716_ clknet_leaf_22_clk _0006_ net65 VGND VGND VPWR VPWR modetrans.mode\[3\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_18_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2859_ _0163_ _0282_ VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5647_ game.flash_counter\[11\] _2616_ game.flash_counter\[12\] VGND VGND VPWR VPWR
+ _2619_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_103_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5578_ _2577_ VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4529_ _1721_ VGND VGND VPWR VPWR _1727_ sky130_fd_sc_hd__inv_2
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_582 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4880_ _2670_ disp_song.um.drum.next_note2\[30\] VGND VGND VPWR VPWR _1975_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_71_clk clknet_3_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_71_clk sky130_fd_sc_hd__clkbuf_16
X_3900_ game.addhits.add1.b\[1\] game.scoring_button_2.acc\[1\] VGND VGND VPWR VPWR
+ _1230_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3831_ _1068_ _1066_ _1131_ _1164_ _0955_ VGND VGND VPWR VPWR _1181_ sky130_fd_sc_hd__a41o_1
X_3762_ disp_song.mi6.in\[2\] _0926_ VGND VGND VPWR VPWR _1116_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5501_ net140 _2460_ _2462_ net145 VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__a22o_1
X_2713_ _0158_ _0159_ VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__nor2_1
X_3693_ _1046_ _1048_ VGND VGND VPWR VPWR _1049_ sky130_fd_sc_hd__or2_1
X_5432_ _2484_ VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5363_ _2438_ VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4314_ _1558_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_2\[21\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5294_ _0214_ _2377_ VGND VGND VPWR VPWR _2378_ sky130_fd_sc_hd__and2_1
X_4245_ net107 game.scoring_button_2.flash_counter_2\[0\] game.missed_2 VGND VGND
+ VPWR VPWR _1510_ sky130_fd_sc_hd__o21ai_1
X_4176_ _1453_ VGND VGND VPWR VPWR game.scoring_button_2.next_count\[14\] sky130_fd_sc_hd__clkbuf_1
X_3127_ game.addmisses.a\[10\] game.addmisses.add3.b\[2\] VGND VGND VPWR VPWR _0490_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3058_ _0353_ _0425_ _0427_ VGND VGND VPWR VPWR disp_song.um.drum.next_note1\[25\]
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_65_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_62_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_62_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_77_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_608 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_53_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_53_clk sky130_fd_sc_hd__clkbuf_16
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4030_ game.addmisses.add2.b\[1\] _1305_ _1329_ _1339_ _1289_ VGND VGND VPWR VPWR
+ _1340_ sky130_fd_sc_hd__o311a_1
XFILLER_0_47_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5981_ clknet_leaf_25_clk net98 net64 VGND VGND VPWR VPWR game.padded_notes1\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4932_ _2025_ VGND VGND VPWR VPWR _2026_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_44_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_44_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_86_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4863_ disp_song.um.drum.next_idx2\[0\] disp_song.um.drum.next_note2\[24\] _1957_
+ VGND VGND VPWR VPWR _1958_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_86_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4794_ _1917_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_1\[15\]
+ sky130_fd_sc_hd__clkbuf_1
X_3814_ _1066_ _1131_ _1163_ _1164_ _0955_ VGND VGND VPWR VPWR _1165_ sky130_fd_sc_hd__a41o_1
XFILLER_0_104_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3745_ _1098_ _1099_ _0895_ VGND VGND VPWR VPWR _1100_ sky130_fd_sc_hd__o21a_1
X_5415_ _2472_ VGND VGND VPWR VPWR _2473_ sky130_fd_sc_hd__buf_8
X_3676_ _1025_ _1026_ _1031_ VGND VGND VPWR VPWR _1032_ sky130_fd_sc_hd__mux2_2
XFILLER_0_63_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5346_ _0841_ _0847_ highest_score.highest_score\[7\] VGND VGND VPWR VPWR _2424_
+ sky130_fd_sc_hd__a21o_1
X_5277_ _0185_ _2360_ VGND VGND VPWR VPWR _2361_ sky130_fd_sc_hd__or2_1
X_4228_ _1494_ VGND VGND VPWR VPWR _1495_ sky130_fd_sc_hd__inv_2
X_4159_ game.counter\[11\] _1439_ VGND VGND VPWR VPWR _1442_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_35_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_35_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_65_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_26_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_26_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_68_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3530_ _0608_ _0886_ _0888_ VGND VGND VPWR VPWR _0893_ sky130_fd_sc_hd__nor3_1
XFILLER_0_12_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3461_ _0822_ _0823_ VGND VGND VPWR VPWR _0824_ sky130_fd_sc_hd__nor2_2
XFILLER_0_58_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3392_ _0514_ _0523_ VGND VGND VPWR VPWR _0755_ sky130_fd_sc_hd__nand2_1
X_5200_ disp_song.um.drum.next_note1\[11\] _2261_ _0176_ VGND VGND VPWR VPWR _2287_
+ sky130_fd_sc_hd__a21o_1
X_5131_ disp_song.um.drum.next_note1\[20\] disp_song.um.drum.next_note1\[21\] disp_song.um.drum.next_idx1\[0\]
+ VGND VGND VPWR VPWR _2219_ sky130_fd_sc_hd__mux2_1
X_5062_ _2666_ _2085_ _0162_ VGND VGND VPWR VPWR _2153_ sky130_fd_sc_hd__a21o_1
XFILLER_0_74_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4013_ game.addmisses.add1.b\[3\] _1307_ _1323_ _1306_ VGND VGND VPWR VPWR _1325_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5964_ clknet_leaf_34_clk game.scoring_button_1.next_flash_counter_2\[9\] net72 VGND
+ VGND VPWR VPWR game.scoring_button_1.flash_counter_2\[9\] sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_17_clk clknet_3_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_17_clk sky130_fd_sc_hd__clkbuf_16
X_5895_ clknet_leaf_32_clk _0078_ net68 VGND VGND VPWR VPWR game.padded_notes2\[28\]
+ sky130_fd_sc_hd__dfrtp_1
X_4915_ _2664_ _2669_ VGND VGND VPWR VPWR _2009_ sky130_fd_sc_hd__nand2_2
XFILLER_0_47_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4846_ disp_song.um.idx_note2\[1\] _0325_ _0366_ _0179_ VGND VGND VPWR VPWR disp_song.um.next_position\[1\]
+ sky130_fd_sc_hd__o22a_1
XFILLER_0_99_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4777_ game.scoring_button_1.flash_counter_1\[11\] game.scoring_button_1.flash_counter_1\[10\]
+ _1901_ VGND VGND VPWR VPWR _1905_ sky130_fd_sc_hd__and3_1
XFILLER_0_43_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3728_ _1081_ _1080_ VGND VGND VPWR VPWR _1084_ sky130_fd_sc_hd__nor2_1
X_3659_ _0788_ _1014_ VGND VGND VPWR VPWR _1015_ sky130_fd_sc_hd__nand2_1
X_5329_ _0366_ VGND VGND VPWR VPWR disp_song.next_green sky130_fd_sc_hd__inv_2
XFILLER_0_100_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2961_ _0354_ _2661_ _0194_ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__or3b_1
XFILLER_0_8_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4700_ _1852_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_2\[9\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5680_ _2643_ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2892_ _0166_ disp_song.um.idx_note2\[1\] disp_song.um.idx_note2\[0\] VGND VGND VPWR
+ VPWR _0307_ sky130_fd_sc_hd__or3b_1
X_4631_ _1791_ _1436_ VGND VGND VPWR VPWR _1809_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4562_ game.addmisses.a\[9\] _1741_ game.addmisses.a\[10\] VGND VGND VPWR VPWR _1756_
+ sky130_fd_sc_hd__a21oi_1
X_3513_ _0873_ _0875_ VGND VGND VPWR VPWR _0876_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4493_ game.addmisses.a\[1\] _1693_ _1695_ _1691_ VGND VGND VPWR VPWR _1696_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_110_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_6_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_6_clk sky130_fd_sc_hd__clkbuf_16
X_3444_ _0786_ _0789_ VGND VGND VPWR VPWR _0807_ sky130_fd_sc_hd__and2_1
XFILLER_0_40_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6163_ clknet_leaf_21_clk disp_song.um.drum.next_d2\[2\] net61 VGND VGND VPWR VPWR
+ disp_song.display_note2\[2\] sky130_fd_sc_hd__dfrtp_1
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3375_ _0731_ _0737_ VGND VGND VPWR VPWR _0738_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_20_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6094_ clknet_leaf_37_clk disp_song.um.drum.next_note1\[6\] net71 VGND VGND VPWR
+ VPWR disp_song.note1\[6\] sky130_fd_sc_hd__dfstp_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5114_ _2189_ _2198_ _2201_ _0197_ VGND VGND VPWR VPWR _2202_ sky130_fd_sc_hd__o22a_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5045_ disp_song.um.drum.next_note2\[2\] _2134_ _2136_ _1965_ VGND VGND VPWR VPWR
+ _2137_ sky130_fd_sc_hd__a211o_1
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_26_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5947_ clknet_leaf_45_clk game.scoring_button_1.next_flash_counter_1\[15\] net54
+ VGND VGND VPWR VPWR game.scoring_button_1.flash_counter_1\[15\] sky130_fd_sc_hd__dfrtp_1
X_5878_ clknet_leaf_19_clk _0061_ net63 VGND VGND VPWR VPWR game.padded_notes2\[11\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_90_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4829_ _0032_ _1452_ VGND VGND VPWR VPWR _1937_ sky130_fd_sc_hd__and2b_1
XFILLER_0_35_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_577 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_599 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3160_ _0515_ _0520_ _0522_ VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__o21ba_1
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1 disp_song.um.boton2e.sync_b VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__dlygate4sd3_1
X_3091_ _0450_ _0453_ VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__xor2_4
XFILLER_0_9_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5801_ clknet_leaf_55_clk game.scoring_button_2.next_flash_counter_1\[15\] net52
+ VGND VGND VPWR VPWR game.scoring_button_2.flash_counter_1\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5732_ clknet_leaf_73_clk game.scoring_button_2.next_num_misses\[4\] net48 VGND VGND
+ VPWR VPWR game.addmisses.add2.b\[0\] sky130_fd_sc_hd__dfrtp_4
X_3993_ _1305_ _1289_ game.addmisses.add1.b\[0\] VGND VGND VPWR VPWR _1308_ sky130_fd_sc_hd__a21oi_1
X_2944_ _0343_ VGND VGND VPWR VPWR disp_song.um.drum.next_note2\[27\] sky130_fd_sc_hd__inv_2
XFILLER_0_57_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2875_ _0273_ _0294_ VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__nand2_1
X_5663_ _2629_ _2631_ VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__nor2_1
X_4614_ _1800_ VGND VGND VPWR VPWR game.scoring_button_1.next_count\[0\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5594_ disp_song.note1\[29\] game.padded_notes1\[28\] _0209_ VGND VGND VPWR VPWR
+ _2588_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4545_ game.addmisses.a\[8\] _1721_ VGND VGND VPWR VPWR _1741_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4476_ game.scoring_button_1.counts\[0\] game.scoring_button_1.counts\[6\] game.scoring_button_1.counts\[5\]
+ _1679_ VGND VGND VPWR VPWR _1680_ sky130_fd_sc_hd__or4_1
XFILLER_0_13_588 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3427_ _0786_ _0789_ VGND VGND VPWR VPWR _0790_ sky130_fd_sc_hd__nor2_1
X_6146_ clknet_leaf_26_clk net149 net68 VGND VGND VPWR VPWR disp_song.note2\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_3358_ _0714_ _0720_ VGND VGND VPWR VPWR _0721_ sky130_fd_sc_hd__xor2_2
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6077_ clknet_leaf_24_clk disp_song.um.drum.next_idx2\[4\] net64 VGND VGND VPWR VPWR
+ disp_song.um.idx_note2\[4\] sky130_fd_sc_hd__dfstp_2
X_3289_ _0454_ _0460_ _0467_ VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__or3_1
X_5028_ _2067_ _2119_ disp_song.um.drum.next_idx2\[2\] VGND VGND VPWR VPWR _2120_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_441 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_628 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4330_ net176 _1565_ _1568_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_1\[4\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_22_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4261_ game.scoring_button_2.flash_counter_2\[6\] _1518_ VGND VGND VPWR VPWR _1521_
+ sky130_fd_sc_hd__and2_1
X_6000_ clknet_leaf_38_clk _0109_ net66 VGND VGND VPWR VPWR game.padded_notes1\[19\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_66_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3212_ _0570_ _0573_ _0571_ VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__o21ai_1
X_4192_ _1464_ VGND VGND VPWR VPWR game.scoring_button_2.next_count\[18\] sky130_fd_sc_hd__clkbuf_1
X_3143_ game.addmisses.a\[13\] game.addmisses.add4.b\[1\] VGND VGND VPWR VPWR _0506_
+ sky130_fd_sc_hd__or2_1
X_3074_ _0435_ _0436_ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3976_ game.scoring_button_2.counts\[16\] game.scoring_button_2.counts\[15\] game.scoring_button_2.counts\[11\]
+ game.scoring_button_2.counts\[10\] VGND VGND VPWR VPWR _1291_ sky130_fd_sc_hd__or4_1
XFILLER_0_57_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2927_ _0288_ _0330_ _0331_ net191 VGND VGND VPWR VPWR disp_song.um.drum.next_note2\[22\]
+ sky130_fd_sc_hd__a22o_1
X_5715_ clknet_leaf_23_clk _0005_ net65 VGND VGND VPWR VPWR modetrans.mode\[2\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_93_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5646_ net126 _2616_ VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__xor2_1
XFILLER_0_103_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2858_ disp_song.um.idx_note2\[3\] disp_song.um.idx_note2\[4\] _2661_ VGND VGND VPWR
+ VPWR _0282_ sky130_fd_sc_hd__or3b_1
XFILLER_0_60_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5577_ _2576_ game.padded_notes1\[23\] _2472_ VGND VGND VPWR VPWR _2577_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2789_ lvls.level\[1\] lvls.level\[0\] _0200_ VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__mux2_1
X_4528_ _1699_ _1724_ _1726_ VGND VGND VPWR VPWR game.scoring_button_1.next_num_misses\[5\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4459_ game.addhits.a\[15\] _1664_ VGND VGND VPWR VPWR _1666_ sky130_fd_sc_hd__or2_1
X_6129_ clknet_leaf_19_clk disp_song.um.drum.next_note2\[9\] net63 VGND VGND VPWR
+ VPWR disp_song.note2\[9\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_99_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_594 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_99_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3830_ _1046_ _1166_ _0941_ VGND VGND VPWR VPWR _1180_ sky130_fd_sc_hd__o21ai_1
X_3761_ _0925_ _0964_ VGND VGND VPWR VPWR _1115_ sky130_fd_sc_hd__nor2_1
XFILLER_0_109_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2712_ _0156_ _2673_ VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5500_ game.out\[8\] _2460_ _2462_ net140 VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__a22o_1
X_3692_ _0642_ _0638_ _1047_ _1042_ VGND VGND VPWR VPWR _1048_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_42_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5431_ _2483_ net229 _2473_ VGND VGND VPWR VPWR _2484_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5362_ _2437_ highest_score.highest_score\[2\] _2434_ VGND VGND VPWR VPWR _2438_
+ sky130_fd_sc_hd__mux2_1
X_4313_ _1556_ game.missed_2 _1557_ VGND VGND VPWR VPWR _1558_ sky130_fd_sc_hd__and3b_1
XFILLER_0_77_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5293_ _2367_ _2370_ _2371_ _2374_ _2376_ _2216_ VGND VGND VPWR VPWR _2377_ sky130_fd_sc_hd__mux4_1
X_4244_ _1509_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_2\[0\]
+ sky130_fd_sc_hd__clkbuf_1
X_4175_ _1405_ _1452_ VGND VGND VPWR VPWR _1453_ sky130_fd_sc_hd__and2_1
XFILLER_0_97_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3126_ game.addmisses.a\[10\] game.addmisses.add3.b\[2\] VGND VGND VPWR VPWR _0489_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_89_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3057_ _0353_ _0426_ net150 VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_89_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3959_ game.addhits.add4.b\[1\] _1275_ game.addhits.add4.b\[2\] VGND VGND VPWR VPWR
+ _1277_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_60_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5629_ game.flash_counter\[8\] game.flash_counter\[7\] game.flash_counter\[6\] game.flash_counter\[9\]
+ VGND VGND VPWR VPWR _2606_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_13_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_591 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5980_ clknet_leaf_11_clk net95 net61 VGND VGND VPWR VPWR game.scoring_button_1.check_hit.edge_1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4931_ _2009_ _2019_ VGND VGND VPWR VPWR _2025_ sky130_fd_sc_hd__and2_1
X_4862_ _1956_ disp_song.um.drum.next_note2\[25\] VGND VGND VPWR VPWR _1957_ sky130_fd_sc_hd__or2_1
XFILLER_0_74_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3813_ _0633_ _0653_ _0636_ VGND VGND VPWR VPWR _1164_ sky130_fd_sc_hd__or3b_1
XFILLER_0_103_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4793_ _1915_ game.hit_1 _1916_ VGND VGND VPWR VPWR _1917_ sky130_fd_sc_hd__and3b_1
X_3744_ highest_score.highest_score\[1\] highest_score.highest_score\[0\] _0255_ VGND
+ VGND VPWR VPWR _1099_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_12_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3675_ _1028_ _1029_ _1030_ VGND VGND VPWR VPWR _1031_ sky130_fd_sc_hd__or3_4
X_5414_ _2461_ VGND VGND VPWR VPWR _2472_ sky130_fd_sc_hd__buf_8
XFILLER_0_30_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5345_ highest_score.highest_score\[7\] _0841_ _0847_ VGND VGND VPWR VPWR _2423_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_56_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5276_ disp_song.um.drum.next_idx1\[1\] _2323_ VGND VGND VPWR VPWR _2360_ sky130_fd_sc_hd__nor2_1
XFILLER_0_10_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4227_ _1489_ _1493_ VGND VGND VPWR VPWR _1494_ sky130_fd_sc_hd__nor2_1
X_4158_ _1441_ VGND VGND VPWR VPWR game.scoring_button_2.next_count\[10\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_631 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4089_ game.addmisses.add4.b\[1\] _1330_ _1383_ VGND VGND VPWR VPWR _1391_ sky130_fd_sc_hd__and3_1
X_3109_ _0446_ _0470_ _0444_ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__o21a_1
XFILLER_0_77_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3460_ _0763_ _0771_ _0772_ VGND VGND VPWR VPWR _0823_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_110_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3391_ _0738_ _0753_ VGND VGND VPWR VPWR _0754_ sky130_fd_sc_hd__xnor2_1
X_5130_ disp_song.um.drum.next_note1\[22\] disp_song.um.drum.next_note1\[23\] disp_song.um.drum.next_idx1\[0\]
+ VGND VGND VPWR VPWR _2218_ sky130_fd_sc_hd__mux2_1
X_5061_ _2141_ _2148_ _2150_ _2151_ VGND VGND VPWR VPWR _2152_ sky130_fd_sc_hd__o22a_1
X_4012_ _1289_ _1311_ VGND VGND VPWR VPWR _1324_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5963_ clknet_leaf_35_clk game.scoring_button_1.next_flash_counter_2\[8\] net72 VGND
+ VGND VPWR VPWR game.scoring_button_1.flash_counter_2\[8\] sky130_fd_sc_hd__dfrtp_1
X_4914_ _1953_ _1984_ _2008_ VGND VGND VPWR VPWR disp_song.um.drum.next_d2\[0\] sky130_fd_sc_hd__o21a_1
X_5894_ clknet_leaf_32_clk _0077_ net68 VGND VGND VPWR VPWR game.padded_notes2\[27\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_90_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4845_ disp_song.um.idx_note2\[0\] _0325_ _0366_ disp_song.um.idx_note1\[0\] VGND
+ VGND VPWR VPWR disp_song.um.next_position\[0\] sky130_fd_sc_hd__o22a_1
XFILLER_0_28_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4776_ net157 _1901_ _1904_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_1\[10\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_15_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3727_ _1077_ _1082_ VGND VGND VPWR VPWR _1083_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3658_ _0662_ _1013_ VGND VGND VPWR VPWR _1014_ sky130_fd_sc_hd__or2b_1
X_3589_ _0938_ _0942_ _0945_ _0950_ modetrans.mode\[3\] VGND VGND VPWR VPWR _0951_
+ sky130_fd_sc_hd__o311a_1
X_5328_ _2401_ _2402_ _2409_ _0214_ VGND VGND VPWR VPWR disp_song.um.drum.next_d1\[6\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5259_ _2339_ _2341_ _2342_ _2343_ VGND VGND VPWR VPWR _2344_ sky130_fd_sc_hd__o22a_1
XFILLER_0_66_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_626 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2960_ _0352_ _0353_ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2891_ _0306_ VGND VGND VPWR VPWR disp_song.um.drum.next_note2\[12\] sky130_fd_sc_hd__buf_1
XTAP_1192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4630_ _1808_ VGND VGND VPWR VPWR game.scoring_button_1.next_count\[8\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4561_ game.addmisses.a\[10\] game.addmisses.a\[9\] _1741_ VGND VGND VPWR VPWR _1755_
+ sky130_fd_sc_hd__and3_1
X_3512_ game.flash_counter\[13\] game.flash_counter\[10\] _0874_ game.flash_counter\[11\]
+ VGND VGND VPWR VPWR _0875_ sky130_fd_sc_hd__or4b_1
XFILLER_0_12_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4492_ game.addmisses.a\[1\] game.addmisses.a\[0\] VGND VGND VPWR VPWR _1695_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3443_ _0634_ _0805_ _0640_ VGND VGND VPWR VPWR _0806_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_100_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6162_ clknet_leaf_8_clk disp_song.um.drum.next_d2\[1\] net60 VGND VGND VPWR VPWR
+ disp_song.display_note2\[1\] sky130_fd_sc_hd__dfrtp_1
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5113_ _2199_ _2200_ disp_song.um.drum.next_idx1\[1\] VGND VGND VPWR VPWR _2201_
+ sky130_fd_sc_hd__mux2_1
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3374_ _0733_ _0736_ VGND VGND VPWR VPWR _0737_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6093_ clknet_leaf_25_clk disp_song.um.drum.next_note1\[5\] net65 VGND VGND VPWR
+ VPWR disp_song.note1\[5\] sky130_fd_sc_hd__dfrtp_1
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ disp_song.um.drum.next_note2\[0\] _1992_ _2035_ _2135_ disp_song.um.drum.next_note2\[1\]
+ VGND VGND VPWR VPWR _2136_ sky130_fd_sc_hd__a32o_1
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5946_ clknet_leaf_45_clk game.scoring_button_1.next_flash_counter_1\[14\] net53
+ VGND VGND VPWR VPWR game.scoring_button_1.flash_counter_1\[14\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5877_ clknet_leaf_19_clk _0060_ net63 VGND VGND VPWR VPWR game.padded_notes2\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_4828_ _1936_ VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4759_ _1891_ game.hit_1 _1892_ VGND VGND VPWR VPWR _1893_ sky130_fd_sc_hd__and3b_1
XFILLER_0_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_101_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_98_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2 modetrans.u2.sync_pb VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__dlygate4sd3_1
X_3090_ _0451_ _0452_ VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__nand2_2
XFILLER_0_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5800_ clknet_leaf_55_clk game.scoring_button_2.next_flash_counter_1\[14\] net52
+ VGND VGND VPWR VPWR game.scoring_button_2.flash_counter_1\[14\] sky130_fd_sc_hd__dfrtp_1
X_3992_ _0208_ _1306_ VGND VGND VPWR VPWR _1307_ sky130_fd_sc_hd__nor2_2
X_2943_ _2655_ _0279_ _0339_ _0342_ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__o31a_1
X_5731_ clknet_leaf_73_clk game.scoring_button_2.next_num_misses\[3\] net48 VGND VGND
+ VPWR VPWR game.addmisses.add1.b\[3\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_84_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2874_ _2672_ _0158_ VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__nor2_1
X_5662_ _2614_ _2630_ VGND VGND VPWR VPWR _2631_ sky130_fd_sc_hd__nand2_1
X_4613_ game.counter\[0\] game.scoring_button_1.check_hit.in VGND VGND VPWR VPWR _1800_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_32_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5593_ _2587_ VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4544_ game.addmisses.a\[8\] _1721_ VGND VGND VPWR VPWR _1740_ sky130_fd_sc_hd__or2_1
XFILLER_0_40_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4475_ game.scoring_button_1.counts\[1\] game.scoring_button_1.counts\[3\] game.scoring_button_1.counts\[2\]
+ game.scoring_button_1.counts\[4\] VGND VGND VPWR VPWR _1679_ sky130_fd_sc_hd__or4_1
XFILLER_0_0_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3426_ _0787_ _0788_ VGND VGND VPWR VPWR _0789_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6145_ clknet_leaf_27_clk disp_song.um.drum.next_note2\[25\] net68 VGND VGND VPWR
+ VPWR disp_song.note2\[25\] sky130_fd_sc_hd__dfstp_1
X_3357_ _0718_ _0719_ VGND VGND VPWR VPWR _0720_ sky130_fd_sc_hd__nor2_1
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6076_ clknet_leaf_21_clk disp_song.um.drum.next_idx2\[3\] net60 VGND VGND VPWR VPWR
+ disp_song.um.idx_note2\[3\] sky130_fd_sc_hd__dfstp_2
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5027_ disp_song.note2\[3\] disp_song.um.drum.next_idx2\[0\] _2043_ _2064_ VGND VGND
+ VPWR VPWR _2119_ sky130_fd_sc_hd__o211a_1
X_3288_ _0454_ _0468_ _0460_ VGND VGND VPWR VPWR _0651_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_45_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5929_ clknet_leaf_12_clk game.scoring_button_1.next_count\[20\] net58 VGND VGND
+ VPWR VPWR game.scoring_button_1.counts\[20\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_467 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_591 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4260_ _1520_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_2\[5\]
+ sky130_fd_sc_hd__clkbuf_1
X_4191_ _1405_ _1463_ VGND VGND VPWR VPWR _1464_ sky130_fd_sc_hd__and2_1
X_3211_ _0572_ _0573_ VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__xnor2_2
X_3142_ _0437_ _0500_ _0501_ _0435_ VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__a31o_1
X_3073_ game.addmisses.a\[12\] game.addmisses.add4.b\[0\] VGND VGND VPWR VPWR _0436_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_82 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3975_ game.scoring_button_2.counts\[14\] game.scoring_button_2.counts\[13\] game.scoring_button_2.counts\[12\]
+ VGND VGND VPWR VPWR _1290_ sky130_fd_sc_hd__or3_1
X_2926_ _0310_ _0327_ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5714_ clknet_leaf_22_clk _0004_ net59 VGND VGND VPWR VPWR modetrans.mode\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2857_ _0281_ VGND VGND VPWR VPWR disp_song.um.drum.next_note2\[3\] sky130_fd_sc_hd__buf_1
XFILLER_0_17_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5645_ _2618_ VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_478 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5576_ disp_song.note1\[23\] game.padded_notes1\[22\] _2541_ VGND VGND VPWR VPWR
+ _2576_ sky130_fd_sc_hd__mux2_1
X_2788_ _0219_ _0217_ _0218_ net164 VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4527_ game.addmisses.a\[5\] _1691_ _1715_ _1725_ _1675_ VGND VGND VPWR VPWR _1726_
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_111_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4458_ game.addhits.a\[15\] _1664_ VGND VGND VPWR VPWR _1665_ sky130_fd_sc_hd__nand2_1
X_3409_ _0764_ _0770_ _0769_ VGND VGND VPWR VPWR _0772_ sky130_fd_sc_hd__a21o_1
X_6128_ clknet_leaf_19_clk disp_song.um.drum.next_note2\[8\] net63 VGND VGND VPWR
+ VPWR disp_song.note2\[8\] sky130_fd_sc_hd__dfrtp_1
X_4389_ net89 _1607_ game.hit_2 VGND VGND VPWR VPWR _1610_ sky130_fd_sc_hd__o21ai_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6059_ clknet_leaf_14_clk _0015_ net61 VGND VGND VPWR VPWR game.counter\[15\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_68_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3760_ _1077_ VGND VGND VPWR VPWR _1114_ sky130_fd_sc_hd__inv_2
X_2711_ disp_song.um.idx_note2\[4\] _0157_ VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__nor2_2
XFILLER_0_27_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5430_ disp_song.note2\[10\] game.padded_notes2\[9\] _0219_ VGND VGND VPWR VPWR _2483_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3691_ _0649_ _1044_ VGND VGND VPWR VPWR _1047_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5361_ _1021_ _1022_ VGND VGND VPWR VPWR _2437_ sky130_fd_sc_hd__and2_1
XFILLER_0_100_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5292_ _2360_ _2375_ VGND VGND VPWR VPWR _2376_ sky130_fd_sc_hd__or2_1
XFILLER_0_10_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4312_ game.scoring_button_2.flash_counter_2\[21\] _1553_ VGND VGND VPWR VPWR _1557_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_77_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4243_ game.scoring_button_2.flash_counter_2\[0\] _1486_ VGND VGND VPWR VPWR _1509_
+ sky130_fd_sc_hd__and2b_1
X_4174_ _1450_ _1451_ VGND VGND VPWR VPWR _1452_ sky130_fd_sc_hd__nor2_1
X_3125_ _0439_ _0486_ _0438_ VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_96_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3056_ _0194_ _0412_ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__or2_2
XFILLER_0_65_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3958_ _1275_ _1276_ net182 _1227_ VGND VGND VPWR VPWR game.scoring_button_2.next_num_hits\[12\]
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_45_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2909_ _2657_ disp_song.note2\[17\] _0319_ VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3889_ _1222_ VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_1
X_5628_ game.flash_counter\[22\] game.flash_counter\[17\] game.flash_counter\[16\]
+ game.flash_counter\[23\] VGND VGND VPWR VPWR _2605_ sky130_fd_sc_hd__or4b_1
X_5559_ _2564_ net238 _2472_ VGND VGND VPWR VPWR _2565_ sky130_fd_sc_hd__mux2_1
XTAP_1533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4930_ _1956_ _0343_ VGND VGND VPWR VPWR _2024_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4861_ _2669_ VGND VGND VPWR VPWR _1956_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_86_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3812_ _1071_ _1132_ VGND VGND VPWR VPWR _1163_ sky130_fd_sc_hd__nand2_1
X_4792_ game.scoring_button_1.flash_counter_1\[15\] _1912_ VGND VGND VPWR VPWR _1916_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_70_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3743_ highest_score.highest_score\[1\] highest_score.highest_score\[0\] _1054_ VGND
+ VGND VPWR VPWR _1098_ sky130_fd_sc_hd__a21o_1
XFILLER_0_55_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3674_ _0807_ _1017_ net42 VGND VGND VPWR VPWR _1030_ sky130_fd_sc_hd__o21a_1
X_5413_ disp_song.note2\[5\] game.padded_notes2\[4\] _0219_ VGND VGND VPWR VPWR _2471_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5344_ _2421_ VGND VGND VPWR VPWR _2422_ sky130_fd_sc_hd__inv_2
XFILLER_0_100_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5275_ _2195_ _2331_ _2332_ _2359_ _0214_ VGND VGND VPWR VPWR disp_song.um.drum.next_d1\[3\]
+ sky130_fd_sc_hd__o311a_1
XFILLER_0_10_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4226_ _0249_ _1490_ _1491_ _1492_ VGND VGND VPWR VPWR _1493_ sky130_fd_sc_hd__or4_1
X_4157_ _1405_ _1440_ VGND VGND VPWR VPWR _1441_ sky130_fd_sc_hd__and2_1
X_3108_ _0446_ _0470_ VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_69_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4088_ game.addmisses.add4.b\[3\] _1387_ _1389_ VGND VGND VPWR VPWR _1390_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3039_ disp_song.note1\[19\] _0414_ _0410_ _0371_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_46_562 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_104_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_110_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3390_ _0735_ _0746_ _0730_ VGND VGND VPWR VPWR _0753_ sky130_fd_sc_hd__a21boi_1
X_5060_ _1983_ _2005_ _2141_ VGND VGND VPWR VPWR _2151_ sky130_fd_sc_hd__o21ai_1
X_4011_ _1319_ _1322_ VGND VGND VPWR VPWR _1323_ sky130_fd_sc_hd__nor2_1
X_5962_ clknet_leaf_36_clk game.scoring_button_1.next_flash_counter_2\[7\] net72 VGND
+ VGND VPWR VPWR game.scoring_button_1.flash_counter_2\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4913_ _1952_ _2007_ _0214_ _1965_ VGND VGND VPWR VPWR _2008_ sky130_fd_sc_hd__o211a_1
X_5893_ clknet_leaf_26_clk _0076_ net68 VGND VGND VPWR VPWR game.padded_notes2\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_646 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4844_ _1944_ VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4775_ net157 _1901_ game.hit_1 VGND VGND VPWR VPWR _1904_ sky130_fd_sc_hd__a21boi_1
X_3726_ disp_song.mi6.in\[3\] _1081_ VGND VGND VPWR VPWR _1082_ sky130_fd_sc_hd__nand2_2
XFILLER_0_70_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3657_ _0661_ _0665_ VGND VGND VPWR VPWR _1013_ sky130_fd_sc_hd__and2_1
XFILLER_0_2_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3588_ net39 _0948_ _0949_ VGND VGND VPWR VPWR _0950_ sky130_fd_sc_hd__a21o_1
X_5327_ _2404_ _2406_ _2407_ _2408_ disp_song.um.drum.next_idx1\[3\] _0185_ VGND VGND
+ VPWR VPWR _2409_ sky130_fd_sc_hd__mux4_1
X_5258_ _2256_ _2300_ _2339_ VGND VGND VPWR VPWR _2343_ sky130_fd_sc_hd__o21ai_1
X_4209_ game.scoring_button_2.check_hit.in _1477_ VGND VGND VPWR VPWR _1478_ sky130_fd_sc_hd__and2_1
X_5189_ _0415_ _2258_ _2232_ VGND VGND VPWR VPWR _2276_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_3_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2890_ disp_song.note2\[12\] _0269_ _0305_ VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__mux2_1
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4560_ _1675_ _1750_ _1751_ _1754_ VGND VGND VPWR VPWR game.scoring_button_1.next_num_misses\[9\]
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_37_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3511_ game.flash_counter\[15\] game.flash_counter\[12\] game.flash_counter\[14\]
+ game.flash_counter\[22\] VGND VGND VPWR VPWR _0874_ sky130_fd_sc_hd__or4bb_1
X_4491_ game.addmisses.a\[0\] _1675_ _1693_ _1694_ VGND VGND VPWR VPWR game.scoring_button_1.next_num_misses\[0\]
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_100_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3442_ _0544_ _0637_ _0636_ VGND VGND VPWR VPWR _0805_ sky130_fd_sc_hd__and3_1
XFILLER_0_110_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6161_ clknet_leaf_8_clk disp_song.um.drum.next_d2\[0\] net60 VGND VGND VPWR VPWR
+ disp_song.display_note2\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3373_ game.addhits.a\[14\] game.addhits.add4.b\[2\] VGND VGND VPWR VPWR _0736_ sky130_fd_sc_hd__or2_1
X_5112_ disp_song.um.drum.next_note1\[4\] disp_song.um.drum.next_note1\[5\] _0176_
+ VGND VGND VPWR VPWR _2200_ sky130_fd_sc_hd__mux2_1
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6092_ clknet_leaf_42_clk disp_song.um.drum.next_note1\[4\] net64 VGND VGND VPWR
+ VPWR disp_song.note1\[4\] sky130_fd_sc_hd__dfrtp_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5043_ _2009_ _2132_ VGND VGND VPWR VPWR _2135_ sky130_fd_sc_hd__nor2_1
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5945_ clknet_leaf_47_clk game.scoring_button_1.next_flash_counter_1\[13\] net56
+ VGND VGND VPWR VPWR game.scoring_button_1.flash_counter_1\[13\] sky130_fd_sc_hd__dfrtp_1
X_5876_ clknet_leaf_19_clk _0059_ net63 VGND VGND VPWR VPWR game.padded_notes2\[9\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_75_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4827_ _0032_ _1442_ _1443_ VGND VGND VPWR VPWR _1936_ sky130_fd_sc_hd__and3b_1
XFILLER_0_63_627 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4758_ game.scoring_button_1.flash_counter_1\[3\] game.scoring_button_1.flash_counter_1\[4\]
+ _1884_ game.scoring_button_1.flash_counter_1\[5\] VGND VGND VPWR VPWR _1892_ sky130_fd_sc_hd__a31o_1
X_4689_ _1843_ _1830_ _1844_ VGND VGND VPWR VPWR _1845_ sky130_fd_sc_hd__and3b_1
X_3709_ _0633_ _0912_ _1064_ VGND VGND VPWR VPWR _1065_ sky130_fd_sc_hd__or3b_1
XFILLER_0_11_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold3 disp_song.um.boton1e.sync_b VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3991_ _1305_ VGND VGND VPWR VPWR _1306_ sky130_fd_sc_hd__inv_2
X_2942_ _0279_ _0337_ disp_song.note2\[27\] VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_71_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5730_ clknet_leaf_73_clk game.scoring_button_2.next_num_misses\[2\] net48 VGND VGND
+ VPWR VPWR game.addmisses.add1.b\[2\] sky130_fd_sc_hd__dfrtp_2
X_2873_ _0293_ VGND VGND VPWR VPWR disp_song.um.drum.next_note2\[7\] sky130_fd_sc_hd__buf_1
XFILLER_0_84_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5661_ game.flash_counter\[14\] game.flash_counter\[13\] _2623_ game.flash_counter\[15\]
+ VGND VGND VPWR VPWR _2630_ sky130_fd_sc_hd__a31o_1
XFILLER_0_29_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4612_ _0219_ _1791_ _2656_ _1799_ VGND VGND VPWR VPWR game.scoring_button_1.next_good
+ sky130_fd_sc_hd__a31o_1
X_5592_ _2586_ net212 _2472_ VGND VGND VPWR VPWR _2587_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4543_ _1735_ _1736_ _1739_ _1675_ VGND VGND VPWR VPWR game.scoring_button_1.next_num_misses\[7\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4474_ game.scoring_button_1.counts\[22\] game.scoring_button_1.counts\[21\] game.scoring_button_1.counts\[20\]
+ _1677_ VGND VGND VPWR VPWR _1678_ sky130_fd_sc_hd__or4_1
XFILLER_0_40_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3425_ _0661_ _0665_ _0662_ VGND VGND VPWR VPWR _0788_ sky130_fd_sc_hd__a21bo_1
X_6144_ clknet_leaf_28_clk disp_song.um.drum.next_note2\[24\] net68 VGND VGND VPWR
+ VPWR disp_song.note2\[24\] sky130_fd_sc_hd__dfrtp_1
X_3356_ _0716_ _0717_ VGND VGND VPWR VPWR _0719_ sky130_fd_sc_hd__and2_1
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6075_ clknet_leaf_24_clk disp_song.um.drum.next_idx2\[2\] net64 VGND VGND VPWR VPWR
+ disp_song.um.idx_note2\[2\] sky130_fd_sc_hd__dfstp_2
X_3287_ _0460_ _0629_ VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__or2_1
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5026_ _2110_ _2114_ _2116_ _2117_ _2107_ VGND VGND VPWR VPWR _2118_ sky130_fd_sc_hd__o32a_1
XFILLER_0_31_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_75_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5928_ clknet_leaf_12_clk game.scoring_button_1.next_count\[19\] net58 VGND VGND
+ VPWR VPWR game.scoring_button_1.counts\[19\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5859_ clknet_leaf_66_clk game.scoring_button_1.next_num_hits\[8\] net47 VGND VGND
+ VPWR VPWR game.addhits.a\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_109_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_619 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_630 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4190_ game.counter\[18\] _1461_ VGND VGND VPWR VPWR _1463_ sky130_fd_sc_hd__xor2_1
X_3210_ _0564_ _0567_ _0565_ VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__o21a_1
XFILLER_0_66_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3141_ _0502_ _0503_ VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__or2_1
X_3072_ game.addmisses.a\[12\] game.addmisses.add4.b\[0\] VGND VGND VPWR VPWR _0435_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_106_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3974_ _1288_ VGND VGND VPWR VPWR _1289_ sky130_fd_sc_hd__clkbuf_8
X_2925_ disp_song.note2\[21\] _0329_ _0330_ _0285_ VGND VGND VPWR VPWR disp_song.um.drum.next_note2\[21\]
+ sky130_fd_sc_hd__a22o_1
X_5713_ clknet_leaf_5_clk _0003_ net49 VGND VGND VPWR VPWR modetrans.mode\[0\] sky130_fd_sc_hd__dfstp_2
X_2856_ _0269_ disp_song.note2\[3\] _0280_ VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5644_ _2614_ _2615_ _2617_ VGND VGND VPWR VPWR _2618_ sky130_fd_sc_hd__and3_1
XFILLER_0_79_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5575_ _2575_ VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__clkbuf_1
X_2787_ modetrans.mode\[3\] _0217_ _0218_ _0208_ VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4526_ game.addmisses.a\[5\] _1717_ VGND VGND VPWR VPWR _1725_ sky130_fd_sc_hd__nand2_1
X_4457_ game.addhits.a\[13\] _1661_ VGND VGND VPWR VPWR _1664_ sky130_fd_sc_hd__xnor2_1
X_3408_ _0764_ _0770_ VGND VGND VPWR VPWR _0771_ sky130_fd_sc_hd__xor2_4
XFILLER_0_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6127_ clknet_leaf_20_clk disp_song.um.drum.next_note2\[7\] net63 VGND VGND VPWR
+ VPWR disp_song.note2\[7\] sky130_fd_sc_hd__dfstp_1
X_4388_ _1609_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_1\[21\]
+ sky130_fd_sc_hd__clkbuf_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3339_ _0695_ _0701_ VGND VGND VPWR VPWR _0702_ sky130_fd_sc_hd__xor2_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6058_ clknet_leaf_9_clk _0014_ net61 VGND VGND VPWR VPWR game.counter\[14\] sky130_fd_sc_hd__dfrtp_2
X_5009_ _2059_ _2060_ _2026_ VGND VGND VPWR VPWR _2101_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_65_clk clknet_3_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_65_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_68_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_56_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_56_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_86_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2710_ disp_song.um.idx_note2\[3\] _2672_ VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3690_ _1043_ _1045_ VGND VGND VPWR VPWR _1046_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5360_ _2436_ VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__clkbuf_1
X_5291_ disp_song.um.drum.next_idx1\[3\] _2215_ VGND VGND VPWR VPWR _2375_ sky130_fd_sc_hd__and2_1
XFILLER_0_22_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4311_ game.scoring_button_2.flash_counter_2\[21\] _1553_ VGND VGND VPWR VPWR _1556_
+ sky130_fd_sc_hd__and2_1
X_4242_ _1405_ _1495_ _1508_ net135 VGND VGND VPWR VPWR game.scoring_button_2.next_start_count
+ sky130_fd_sc_hd__a22o_1
X_4173_ game.counter\[14\] _1449_ VGND VGND VPWR VPWR _1451_ sky130_fd_sc_hd__and2_1
X_3124_ _0440_ _0486_ VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__xor2_2
XFILLER_0_93_77 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3055_ _0194_ _0410_ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__or2_2
Xclkbuf_leaf_47_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_47_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_92_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3957_ game.addhits.add4.b\[0\] _1268_ _1226_ VGND VGND VPWR VPWR _1276_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_18_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2908_ _0156_ _0297_ _0318_ _0270_ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__or4_1
XFILLER_0_73_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_596 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3888_ _0933_ _1221_ VGND VGND VPWR VPWR _1222_ sky130_fd_sc_hd__and2_1
X_2839_ _0265_ _0266_ disp_song.note2\[0\] VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__o21a_1
XFILLER_0_14_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5627_ game.flash_counter\[21\] game.flash_counter\[20\] VGND VGND VPWR VPWR _2604_
+ sky130_fd_sc_hd__or2b_1
XFILLER_0_103_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5558_ disp_song.note1\[17\] game.padded_notes1\[16\] _2541_ VGND VGND VPWR VPWR
+ _2564_ sky130_fd_sc_hd__mux2_1
X_4509_ _1675_ _1697_ VGND VGND VPWR VPWR _1710_ sky130_fd_sc_hd__nor2_1
X_5489_ disp_song.note2\[29\] game.padded_notes2\[28\] _2497_ VGND VGND VPWR VPWR
+ _2523_ sky130_fd_sc_hd__mux2_1
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_38_clk clknet_3_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_38_clk sky130_fd_sc_hd__clkbuf_16
XTAP_1523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_29_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_29_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_63_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4860_ _1954_ _0343_ disp_song.um.drum.next_idx2\[0\] VGND VGND VPWR VPWR _1955_
+ sky130_fd_sc_hd__mux2_1
X_3811_ _1031_ _1026_ _1091_ VGND VGND VPWR VPWR _1162_ sky130_fd_sc_hd__a21o_1
XFILLER_0_27_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4791_ game.scoring_button_1.flash_counter_1\[15\] _1912_ VGND VGND VPWR VPWR _1915_
+ sky130_fd_sc_hd__and2_1
X_3742_ _1095_ _1096_ _1040_ VGND VGND VPWR VPWR _1097_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_70_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3673_ net42 _0806_ _1016_ VGND VGND VPWR VPWR _1029_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_42_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5412_ _2470_ VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5343_ highest_score.highest_score\[5\] _0840_ _0855_ highest_score.highest_score\[4\]
+ VGND VGND VPWR VPWR _2421_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5274_ _2333_ _2347_ _2358_ _2234_ VGND VGND VPWR VPWR _2359_ sky130_fd_sc_hd__a211o_1
X_4225_ game.counter\[21\] game.counter\[22\] game.counter\[20\] VGND VGND VPWR VPWR
+ _1492_ sky130_fd_sc_hd__or3b_1
X_4156_ _1438_ _1439_ VGND VGND VPWR VPWR _1440_ sky130_fd_sc_hd__nor2_1
X_3107_ _0449_ _0468_ _0469_ _0447_ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__o31a_2
X_4087_ game.addmisses.add4.b\[2\] _1385_ _1388_ VGND VGND VPWR VPWR _1389_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_77_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3038_ _0371_ _0412_ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4989_ _1994_ _2081_ _2667_ VGND VGND VPWR VPWR _2082_ sky130_fd_sc_hd__mux2_1
XFILLER_0_18_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_104_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_110 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4010_ game.addmisses.add1.b\[3\] _1315_ VGND VGND VPWR VPWR _1322_ sky130_fd_sc_hd__nor2_1
X_5961_ clknet_leaf_34_clk game.scoring_button_1.next_flash_counter_2\[6\] net72 VGND
+ VGND VPWR VPWR game.scoring_button_1.flash_counter_2\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4912_ _1998_ _2006_ _1961_ VGND VGND VPWR VPWR _2007_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5892_ clknet_leaf_26_clk _0075_ net68 VGND VGND VPWR VPWR game.padded_notes2\[25\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_47_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4843_ _0032_ _1477_ VGND VGND VPWR VPWR _1944_ sky130_fd_sc_hd__and2b_1
XFILLER_0_47_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4774_ _1903_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_1\[9\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3725_ disp_song.mi6.in\[2\] VGND VGND VPWR VPWR _1081_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_9_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_9_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_3_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3656_ _0806_ VGND VGND VPWR VPWR _1012_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3587_ _0255_ _0258_ VGND VGND VPWR VPWR _0949_ sky130_fd_sc_hd__or2_2
X_5326_ _2325_ _2326_ disp_song.um.drum.next_idx1\[2\] VGND VGND VPWR VPWR _2408_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_474 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5257_ _2254_ _2303_ VGND VGND VPWR VPWR _2342_ sky130_fd_sc_hd__nor2_1
X_4208_ game.counter\[22\] _1474_ VGND VGND VPWR VPWR _1477_ sky130_fd_sc_hd__xnor2_1
X_5188_ _2256_ _2271_ _2273_ _2274_ VGND VGND VPWR VPWR _2275_ sky130_fd_sc_hd__a31o_1
X_4139_ _1405_ _1426_ VGND VGND VPWR VPWR _1427_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_636 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_271 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_3_4__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_4__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_60_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_658 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_84_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3510_ game.flash_counter\[20\] game.flash_counter\[21\] _0871_ _0872_ VGND VGND
+ VPWR VPWR _0873_ sky130_fd_sc_hd__or4_1
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4490_ _1691_ _1675_ game.addmisses.a\[0\] VGND VGND VPWR VPWR _1694_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_100_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3441_ _0781_ _0793_ VGND VGND VPWR VPWR _0804_ sky130_fd_sc_hd__or2_1
XFILLER_0_40_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6160_ clknet_leaf_30_clk net74 net70 VGND VGND VPWR VPWR disp_song.um.boton2e.edge_1
+ sky130_fd_sc_hd__dfrtp_1
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3372_ game.addhits.a\[15\] game.addhits.add4.b\[3\] _0734_ VGND VGND VPWR VPWR _0735_
+ sky130_fd_sc_hd__o21ai_1
X_5111_ disp_song.um.drum.next_note1\[6\] disp_song.um.drum.next_note1\[7\] _0176_
+ VGND VGND VPWR VPWR _2199_ sky130_fd_sc_hd__mux2_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6091_ clknet_leaf_26_clk disp_song.um.drum.next_note1\[3\] net64 VGND VGND VPWR
+ VPWR disp_song.note1\[3\] sky130_fd_sc_hd__dfstp_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5042_ _2133_ VGND VGND VPWR VPWR _2134_ sky130_fd_sc_hd__inv_2
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5944_ clknet_leaf_46_clk game.scoring_button_1.next_flash_counter_1\[12\] net55
+ VGND VGND VPWR VPWR game.scoring_button_1.flash_counter_1\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5875_ clknet_leaf_19_clk _0058_ net63 VGND VGND VPWR VPWR game.padded_notes2\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_4826_ _1935_ VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4757_ game.scoring_button_1.flash_counter_1\[5\] game.scoring_button_1.flash_counter_1\[4\]
+ _1887_ VGND VGND VPWR VPWR _1891_ sky130_fd_sc_hd__and3_1
X_4688_ game.scoring_button_1.flash_counter_2\[6\] _1840_ VGND VGND VPWR VPWR _1844_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_70_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3708_ _0651_ _0652_ VGND VGND VPWR VPWR _1064_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3639_ _0904_ _0996_ _0258_ VGND VGND VPWR VPWR _0997_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5309_ _2247_ _2391_ VGND VGND VPWR VPWR _2392_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_636 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold4 modetrans.u3.sync_pb VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3990_ _1304_ VGND VGND VPWR VPWR _1305_ sky130_fd_sc_hd__clkbuf_4
X_2941_ _2655_ _0340_ _0341_ VGND VGND VPWR VPWR disp_song.um.drum.next_note2\[26\]
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_69_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5660_ _2628_ VGND VGND VPWR VPWR _2629_ sky130_fd_sc_hd__buf_2
XFILLER_0_45_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2872_ _0269_ disp_song.note2\[7\] _0292_ VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__mux2_1
X_4611_ _1792_ _1793_ _1798_ game.hit_1 VGND VGND VPWR VPWR _1799_ sky130_fd_sc_hd__o31a_2
X_5591_ disp_song.note1\[28\] game.padded_notes1\[27\] _0209_ VGND VGND VPWR VPWR
+ _2586_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4542_ _1692_ _1737_ _1738_ _1693_ game.addmisses.a\[7\] VGND VGND VPWR VPWR _1739_
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_111_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4473_ game.scoring_button_1.counts\[19\] game.scoring_button_1.counts\[18\] game.scoring_button_1.counts\[17\]
+ game.scoring_button_1.counts\[16\] VGND VGND VPWR VPWR _1677_ sky130_fd_sc_hd__or4_1
XFILLER_0_40_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3424_ _0661_ _0665_ VGND VGND VPWR VPWR _0787_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6143_ clknet_leaf_30_clk disp_song.um.drum.next_note2\[23\] net69 VGND VGND VPWR
+ VPWR disp_song.note2\[23\] sky130_fd_sc_hd__dfstp_1
X_3355_ _0716_ _0717_ VGND VGND VPWR VPWR _0718_ sky130_fd_sc_hd__nor2_1
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6074_ clknet_leaf_28_clk disp_song.um.drum.next_idx2\[1\] net68 VGND VGND VPWR VPWR
+ disp_song.um.idx_note2\[1\] sky130_fd_sc_hd__dfstp_4
X_3286_ _0552_ _0647_ _0648_ VGND VGND VPWR VPWR _0649_ sky130_fd_sc_hd__a21o_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5025_ _0169_ _2019_ _2679_ VGND VGND VPWR VPWR _2117_ sky130_fd_sc_hd__a21oi_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5927_ clknet_leaf_13_clk game.scoring_button_1.next_count\[18\] net58 VGND VGND
+ VPWR VPWR game.scoring_button_1.counts\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5858_ clknet_leaf_66_clk game.scoring_button_1.next_num_hits\[7\] net46 VGND VGND
+ VPWR VPWR game.addhits.a\[7\] sky130_fd_sc_hd__dfrtp_2
X_5789_ clknet_leaf_54_clk game.scoring_button_2.next_flash_counter_1\[3\] net52 VGND
+ VGND VPWR VPWR game.scoring_button_2.flash_counter_1\[3\] sky130_fd_sc_hd__dfrtp_1
X_4809_ _1926_ game.hit_1 _1927_ VGND VGND VPWR VPWR _1928_ sky130_fd_sc_hd__and3b_1
XFILLER_0_90_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_299 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3140_ _0500_ _0501_ _0437_ VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__a21oi_1
X_3071_ _0402_ _0419_ _0434_ net160 VGND VGND VPWR VPWR disp_song.um.drum.next_note1\[31\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5712_ clknet_leaf_39_clk modetrans.pushed_3 net66 VGND VGND VPWR VPWR modetrans.u2.sync_pb
+ sky130_fd_sc_hd__dfrtp_1
X_3973_ game.scoring_button_2.check_hit.edge_1 _1287_ game.scoring_button_2.hit VGND
+ VGND VPWR VPWR _1288_ sky130_fd_sc_hd__or3_1
X_2924_ disp_song.um.idx_note2\[4\] _0269_ _2675_ disp_song.next_red VGND VGND VPWR
+ VPWR _0330_ sky130_fd_sc_hd__and4_2
X_2855_ _0279_ disp_song.um.idx_note2\[3\] _0161_ VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__or3b_1
X_5643_ _2616_ VGND VGND VPWR VPWR _2617_ sky130_fd_sc_hd__inv_2
XFILLER_0_31_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5574_ _2574_ game.padded_notes1\[22\] _2472_ VGND VGND VPWR VPWR _2575_ sky130_fd_sc_hd__mux2_1
XFILLER_0_60_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2786_ _0219_ _0218_ _0220_ _0217_ VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4525_ _1721_ _1723_ VGND VGND VPWR VPWR _1724_ sky130_fd_sc_hd__xor2_1
XFILLER_0_40_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4456_ game.addhits.a\[13\] _1661_ game.addhits.a\[14\] VGND VGND VPWR VPWR _1663_
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4387_ _1607_ game.hit_2 _1608_ VGND VGND VPWR VPWR _1609_ sky130_fd_sc_hd__and3b_1
X_3407_ _0768_ _0769_ VGND VGND VPWR VPWR _0770_ sky130_fd_sc_hd__nor2_2
X_6126_ clknet_leaf_20_clk disp_song.um.drum.next_note2\[6\] net63 VGND VGND VPWR
+ VPWR disp_song.note2\[6\] sky130_fd_sc_hd__dfrtp_1
X_3338_ _0699_ _0700_ VGND VGND VPWR VPWR _0701_ sky130_fd_sc_hd__nor2_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6057_ clknet_leaf_7_clk _0013_ net59 VGND VGND VPWR VPWR game.counter\[13\] sky130_fd_sc_hd__dfrtp_1
X_3269_ _0624_ _0631_ VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__xnor2_1
X_5008_ disp_song.um.drum.next_idx2\[2\] _2035_ VGND VGND VPWR VPWR _2100_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_95_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_98_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5290_ _2372_ _2373_ _2365_ VGND VGND VPWR VPWR _2374_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4310_ _1555_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_2\[20\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4241_ _0228_ _1496_ _1500_ _1507_ VGND VGND VPWR VPWR _1508_ sky130_fd_sc_hd__and4_1
X_4172_ game.counter\[14\] _1449_ VGND VGND VPWR VPWR _1450_ sky130_fd_sc_hd__nor2_1
X_3123_ _0443_ _0484_ _0485_ _0441_ VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_93_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3054_ _0386_ _0410_ _0424_ VGND VGND VPWR VPWR disp_song.um.drum.next_note1\[24\]
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_65_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3956_ game.addhits.add4.b\[0\] _1268_ VGND VGND VPWR VPWR _1275_ sky130_fd_sc_hd__and2_1
XFILLER_0_85_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2907_ _2654_ _2676_ VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3887_ _0966_ disp_song.display_note2\[6\] _0210_ game.out\[6\] _0208_ VGND VGND
+ VPWR VPWR _1221_ sky130_fd_sc_hd__a221o_2
X_5626_ game.flash_counter\[6\] game.flash_counter\[5\] _2601_ game.flash_counter\[7\]
+ VGND VGND VPWR VPWR _2603_ sky130_fd_sc_hd__a31oi_1
X_2838_ _2661_ _0158_ VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__nand2_1
X_5557_ _2563_ VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__clkbuf_1
X_2769_ _0203_ _0206_ VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5488_ _2522_ VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4508_ _1705_ _1708_ VGND VGND VPWR VPWR _1709_ sky130_fd_sc_hd__nor2_1
X_4439_ game.addhits.a\[8\] _1639_ _1612_ VGND VGND VPWR VPWR _1651_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_111_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6109_ clknet_leaf_38_clk disp_song.um.drum.next_note1\[21\] net67 VGND VGND VPWR
+ VPWR disp_song.note1\[21\] sky130_fd_sc_hd__dfrtp_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_391 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_655 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4790_ _1914_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_1\[14\]
+ sky130_fd_sc_hd__clkbuf_1
X_3810_ _1025_ _1031_ VGND VGND VPWR VPWR _1161_ sky130_fd_sc_hd__and2_1
XFILLER_0_7_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3741_ _0642_ _0638_ net44 VGND VGND VPWR VPWR _1096_ sky130_fd_sc_hd__and3_1
XFILLER_0_70_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_564 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3672_ _0834_ _1027_ net42 VGND VGND VPWR VPWR _1028_ sky130_fd_sc_hd__mux2_2
X_5411_ _2469_ net254 _2462_ VGND VGND VPWR VPWR _2470_ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5342_ highest_score.highest_score\[4\] _0855_ _1024_ highest_score.highest_score\[3\]
+ VGND VGND VPWR VPWR _2420_ sky130_fd_sc_hd__o22a_1
XFILLER_0_2_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5273_ _2333_ _2357_ VGND VGND VPWR VPWR _2358_ sky130_fd_sc_hd__and2b_1
X_4224_ game.counter\[8\] game.counter\[9\] game.counter\[10\] game.counter\[11\]
+ VGND VGND VPWR VPWR _1491_ sky130_fd_sc_hd__or4b_1
X_4155_ game.counter\[10\] _1435_ VGND VGND VPWR VPWR _1439_ sky130_fd_sc_hd__and2_1
X_3106_ _0461_ _0463_ _0465_ VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__nor3_1
X_4086_ game.addmisses.add4.b\[3\] _1387_ VGND VGND VPWR VPWR _1388_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3037_ _0364_ _0410_ _0413_ VGND VGND VPWR VPWR disp_song.um.drum.next_note1\[18\]
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_93_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4988_ _1968_ _1991_ VGND VGND VPWR VPWR _2081_ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3939_ _1256_ _1257_ _1226_ _1252_ _1227_ VGND VGND VPWR VPWR _1263_ sky130_fd_sc_hd__a41o_1
XFILLER_0_33_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_104_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5609_ game.out\[5\] _2460_ _2462_ net93 VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5960_ clknet_leaf_36_clk game.scoring_button_1.next_flash_counter_2\[5\] net72 VGND
+ VGND VPWR VPWR game.scoring_button_1.flash_counter_2\[5\] sky130_fd_sc_hd__dfrtp_1
X_5891_ clknet_leaf_27_clk _0074_ net68 VGND VGND VPWR VPWR game.padded_notes2\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_4911_ _2002_ _2005_ _1983_ VGND VGND VPWR VPWR _2006_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4842_ _1943_ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4773_ _1901_ _1799_ _1902_ VGND VGND VPWR VPWR _1903_ sky130_fd_sc_hd__and3b_1
XFILLER_0_43_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3724_ _1078_ _1079_ VGND VGND VPWR VPWR _1080_ sky130_fd_sc_hd__and2_1
XFILLER_0_7_469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3655_ _0789_ VGND VGND VPWR VPWR _1011_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3586_ _0858_ _0947_ VGND VGND VPWR VPWR _0948_ sky130_fd_sc_hd__nand2_1
X_5325_ _2187_ _2199_ VGND VGND VPWR VPWR _2407_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5256_ _2295_ _2296_ _2256_ VGND VGND VPWR VPWR _2341_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4207_ _1476_ VGND VGND VPWR VPWR game.scoring_button_2.next_count\[21\] sky130_fd_sc_hd__clkbuf_1
X_5187_ _2245_ _2246_ VGND VGND VPWR VPWR _2274_ sky130_fd_sc_hd__nor2_2
X_4138_ game.counter\[6\] _1423_ VGND VGND VPWR VPWR _1426_ sky130_fd_sc_hd__xor2_1
XFILLER_0_97_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4069_ game.addmisses.add3.b\[2\] game.addmisses.add3.b\[1\] game.addmisses.add3.b\[0\]
+ _1357_ VGND VGND VPWR VPWR _1374_ sky130_fd_sc_hd__and4_1
XFILLER_0_78_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire40 net41 VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3440_ _0711_ _0721_ _0802_ VGND VGND VPWR VPWR _0803_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_100_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3371_ _0731_ _0732_ _0733_ VGND VGND VPWR VPWR _0734_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6090_ clknet_leaf_42_clk disp_song.um.drum.next_note1\[2\] net64 VGND VGND VPWR
+ VPWR disp_song.note1\[2\] sky130_fd_sc_hd__dfstp_2
X_5110_ _2193_ _2197_ VGND VGND VPWR VPWR _2198_ sky130_fd_sc_hd__nor2_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5041_ disp_song.um.drum.next_idx2\[1\] _1956_ _2132_ VGND VGND VPWR VPWR _2133_
+ sky130_fd_sc_hd__or3_1
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_87_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5943_ clknet_leaf_52_clk game.scoring_button_1.next_flash_counter_1\[11\] net55
+ VGND VGND VPWR VPWR game.scoring_button_1.flash_counter_1\[11\] sky130_fd_sc_hd__dfrtp_1
X_5874_ clknet_leaf_19_clk _0057_ net63 VGND VGND VPWR VPWR game.padded_notes2\[7\]
+ sky130_fd_sc_hd__dfstp_1
X_4825_ _0032_ _1440_ VGND VGND VPWR VPWR _1935_ sky130_fd_sc_hd__and2b_1
XFILLER_0_47_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4756_ net207 _1887_ _1890_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_1\[4\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_43_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4687_ game.scoring_button_1.flash_counter_2\[6\] _1840_ VGND VGND VPWR VPWR _1843_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_16_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3707_ _1056_ _1062_ _0258_ VGND VGND VPWR VPWR _1063_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3638_ _0943_ _0255_ _0901_ VGND VGND VPWR VPWR _0996_ sky130_fd_sc_hd__and3b_1
X_3569_ _0259_ _0922_ VGND VGND VPWR VPWR _0932_ sky130_fd_sc_hd__nor2_1
X_5308_ _2254_ _2337_ _2390_ _2310_ VGND VGND VPWR VPWR _2391_ sky130_fd_sc_hd__o22a_1
X_5239_ _2203_ _2205_ _2185_ VGND VGND VPWR VPWR _2325_ sky130_fd_sc_hd__mux2_1
XPHY_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_604 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold5 disp_song.um.boton2e.edge_1 VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2940_ _0276_ _0336_ disp_song.note2\[26\] VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_57_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2871_ _0273_ _0291_ VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__nand2_1
XFILLER_0_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4610_ _1794_ _1795_ _1796_ _1797_ VGND VGND VPWR VPWR _1798_ sky130_fd_sc_hd__or4b_1
XFILLER_0_111_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5590_ _2585_ VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4541_ game.addmisses.a\[7\] _1730_ VGND VGND VPWR VPWR _1738_ sky130_fd_sc_hd__or2_1
XFILLER_0_52_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4472_ game.scoring_button_1.counts\[13\] game.scoring_button_1.counts\[12\] game.scoring_button_1.counts\[14\]
+ VGND VGND VPWR VPWR _1676_ sky130_fd_sc_hd__or3_1
XFILLER_0_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3423_ _0660_ _0785_ _0664_ VGND VGND VPWR VPWR _0786_ sky130_fd_sc_hd__a21o_1
XFILLER_0_40_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_110_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_110_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6142_ clknet_leaf_30_clk disp_song.um.drum.next_note2\[22\] net70 VGND VGND VPWR
+ VPWR disp_song.note2\[22\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3354_ _0600_ _0598_ _0492_ VGND VGND VPWR VPWR _0717_ sky130_fd_sc_hd__nand3b_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6073_ clknet_leaf_29_clk disp_song.um.drum.next_idx2\[0\] net69 VGND VGND VPWR VPWR
+ disp_song.um.idx_note2\[0\] sky130_fd_sc_hd__dfstp_4
X_3285_ _0559_ _0553_ VGND VGND VPWR VPWR _0648_ sky130_fd_sc_hd__and2b_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5024_ _2020_ _2017_ _2100_ _2115_ VGND VGND VPWR VPWR _2116_ sky130_fd_sc_hd__o211a_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5926_ clknet_leaf_13_clk game.scoring_button_1.next_count\[17\] net58 VGND VGND
+ VPWR VPWR game.scoring_button_1.counts\[17\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5857_ clknet_leaf_71_clk game.scoring_button_1.next_num_hits\[6\] net46 VGND VGND
+ VPWR VPWR game.addhits.a\[6\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_48_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5788_ clknet_leaf_55_clk game.scoring_button_2.next_flash_counter_1\[2\] net52 VGND
+ VGND VPWR VPWR game.scoring_button_2.flash_counter_1\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_16_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4808_ game.scoring_button_1.flash_counter_1\[19\] game.scoring_button_1.flash_counter_1\[18\]
+ _1919_ game.scoring_button_1.flash_counter_1\[20\] VGND VGND VPWR VPWR _1927_ sky130_fd_sc_hd__a31o_1
XFILLER_0_44_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4739_ _1878_ game.missed_1 _1879_ VGND VGND VPWR VPWR _1880_ sky130_fd_sc_hd__and3b_1
XFILLER_0_50_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_101_255 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_651 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3070_ _0402_ _0421_ VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5711_ clknet_leaf_23_clk net82 net65 VGND VGND VPWR VPWR modetrans.u2.Q2 sky130_fd_sc_hd__dfrtp_1
X_3972_ game.scoring_button_2.check_hit.edge_2 VGND VGND VPWR VPWR _1287_ sky130_fd_sc_hd__inv_2
X_2923_ _0307_ _0327_ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__or2_1
XFILLER_0_72_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2854_ disp_song.um.idx_note2\[1\] disp_song.um.idx_note2\[0\] _0166_ VGND VGND VPWR
+ VPWR _0279_ sky130_fd_sc_hd__nand3_2
X_5642_ game.flash_counter\[10\] game.flash_counter\[9\] game.flash_counter\[8\] _2612_
+ VGND VGND VPWR VPWR _2616_ sky130_fd_sc_hd__and4_1
X_5573_ disp_song.note1\[22\] game.padded_notes1\[21\] _2541_ VGND VGND VPWR VPWR
+ _2574_ sky130_fd_sc_hd__mux2_1
X_2785_ modetrans.mode\[5\] net270 VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4524_ _1720_ _1722_ VGND VGND VPWR VPWR _1723_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4455_ _1661_ _1662_ net189 _1613_ VGND VGND VPWR VPWR game.scoring_button_1.next_num_hits\[12\]
+ sky130_fd_sc_hd__a2bb2o_1
X_3406_ _0766_ _0767_ VGND VGND VPWR VPWR _0769_ sky130_fd_sc_hd__nor2_1
X_4386_ game.scoring_button_2.flash_counter_1\[21\] _1604_ VGND VGND VPWR VPWR _1608_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_40_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6125_ clknet_leaf_24_clk disp_song.um.drum.next_note2\[5\] net64 VGND VGND VPWR
+ VPWR disp_song.note2\[5\] sky130_fd_sc_hd__dfstp_1
X_3337_ _0697_ _0698_ VGND VGND VPWR VPWR _0700_ sky130_fd_sc_hd__nor2_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6056_ clknet_leaf_8_clk _0012_ net60 VGND VGND VPWR VPWR game.counter\[12\] sky130_fd_sc_hd__dfrtp_2
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3268_ _0628_ _0630_ VGND VGND VPWR VPWR _0631_ sky130_fd_sc_hd__nand2_1
X_5007_ _2099_ VGND VGND VPWR VPWR disp_song.um.drum.next_d2\[2\] sky130_fd_sc_hd__clkbuf_1
X_3199_ _0543_ _0560_ _0561_ _0541_ VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_95_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5909_ clknet_leaf_15_clk game.scoring_button_1.next_count\[0\] net62 VGND VGND VPWR
+ VPWR game.scoring_button_1.counts\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_597 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4240_ game.counter\[16\] _0245_ _1502_ _1504_ _1506_ VGND VGND VPWR VPWR _1507_
+ sky130_fd_sc_hd__o2111a_1
XFILLER_0_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4171_ _1443_ _1446_ VGND VGND VPWR VPWR _1449_ sky130_fd_sc_hd__nor2_1
X_3122_ _0477_ _0479_ _0481_ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__nor3_2
X_3053_ _0386_ _0412_ net259 VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_77_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3955_ net219 _1227_ _1274_ _1226_ VGND VGND VPWR VPWR game.scoring_button_2.next_num_hits\[11\]
+ sky130_fd_sc_hd__a22o_1
X_2906_ _2661_ disp_song.um.idx_note2\[4\] _2673_ _0264_ _0317_ VGND VGND VPWR VPWR
+ disp_song.um.drum.next_note2\[16\] sky130_fd_sc_hd__a41o_1
XFILLER_0_45_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3886_ _1220_ VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_1
X_5625_ net142 _2602_ VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2837_ _2654_ _2660_ VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__nand2_2
XFILLER_0_14_621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5556_ _2562_ net226 _2472_ VGND VGND VPWR VPWR _2563_ sky130_fd_sc_hd__mux2_1
X_2768_ pulseout.fin_pulse\[1\] _0204_ _0205_ pulseout.fin_pulse\[0\] VGND VGND VPWR
+ VPWR _0206_ sky130_fd_sc_hd__or4b_4
X_5487_ _2521_ net233 _2515_ VGND VGND VPWR VPWR _2522_ sky130_fd_sc_hd__mux2_1
X_2699_ disp_song.um.idx_note2\[3\] VGND VGND VPWR VPWR _2671_ sky130_fd_sc_hd__inv_2
X_4507_ game.addmisses.a\[3\] _1701_ VGND VGND VPWR VPWR _1708_ sky130_fd_sc_hd__nor2_1
XFILLER_0_13_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4438_ game.addhits.a\[8\] _1639_ VGND VGND VPWR VPWR _1650_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4369_ net174 _1593_ _1413_ VGND VGND VPWR VPWR _1596_ sky130_fd_sc_hd__a21boi_1
X_6108_ clknet_leaf_41_clk disp_song.um.drum.next_note1\[20\] net67 VGND VGND VPWR
+ VPWR disp_song.note1\[20\] sky130_fd_sc_hd__dfrtp_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6039_ clknet_leaf_57_clk _0148_ net50 VGND VGND VPWR VPWR game.flash_counter\[19\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_96_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_645 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_106_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_74_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3740_ _0642_ _0638_ VGND VGND VPWR VPWR _1095_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3671_ _0775_ _0831_ _0790_ _0844_ VGND VGND VPWR VPWR _1027_ sky130_fd_sc_hd__or4_1
X_5410_ disp_song.note2\[4\] game.padded_notes2\[3\] _0219_ VGND VGND VPWR VPWR _2469_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_70_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5341_ highest_score.highest_score\[2\] _2414_ _1024_ highest_score.highest_score\[3\]
+ VGND VGND VPWR VPWR _2419_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5272_ _2352_ _2356_ _2346_ VGND VGND VPWR VPWR _2357_ sky130_fd_sc_hd__mux2_1
X_4223_ _0237_ _0240_ game.counter\[19\] game.counter\[18\] VGND VGND VPWR VPWR _1490_
+ sky130_fd_sc_hd__or4_1
X_4154_ game.counter\[10\] _1435_ VGND VGND VPWR VPWR _1438_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4085_ _1385_ _1386_ VGND VGND VPWR VPWR _1387_ sky130_fd_sc_hd__or2_1
X_3105_ _0461_ _0466_ _0467_ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__o21a_4
X_3036_ _0364_ _0412_ net240 VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4987_ _1986_ _1988_ _2666_ VGND VGND VPWR VPWR _2080_ sky130_fd_sc_hd__mux2_1
X_3938_ _1259_ _1262_ net253 _1227_ VGND VGND VPWR VPWR game.scoring_button_2.next_num_hits\[6\]
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_46_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3869_ _0966_ disp_song.display_note2\[0\] _0211_ game.out\[0\] _0208_ VGND VGND
+ VPWR VPWR _1209_ sky130_fd_sc_hd__a221o_2
XFILLER_0_104_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5608_ net115 _2460_ _2462_ net127 VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5539_ _2551_ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5890_ clknet_leaf_32_clk _0073_ net69 VGND VGND VPWR VPWR game.padded_notes2\[23\]
+ sky130_fd_sc_hd__dfstp_1
X_4910_ _2003_ _2004_ disp_song.um.drum.next_idx2\[1\] VGND VGND VPWR VPWR _2005_
+ sky130_fd_sc_hd__mux2_1
X_4841_ _0032_ _1475_ VGND VGND VPWR VPWR _1943_ sky130_fd_sc_hd__and2b_1
XFILLER_0_74_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4772_ game.scoring_button_1.flash_counter_1\[9\] _1898_ VGND VGND VPWR VPWR _1902_
+ sky130_fd_sc_hd__or2_1
X_3723_ disp_song.mi6.in\[3\] _0926_ VGND VGND VPWR VPWR _1079_ sky130_fd_sc_hd__or2_1
X_3654_ _0930_ _0953_ _1009_ _1010_ _0935_ VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__o41a_2
XFILLER_0_30_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3585_ _0840_ _0946_ VGND VGND VPWR VPWR _0947_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_590 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_100_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5324_ _2317_ _2405_ disp_song.um.drum.next_idx1\[2\] VGND VGND VPWR VPWR _2406_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5255_ _2334_ _2338_ _2339_ VGND VGND VPWR VPWR _2340_ sky130_fd_sc_hd__mux2_1
X_4206_ game.scoring_button_2.check_hit.in _1475_ VGND VGND VPWR VPWR _1476_ sky130_fd_sc_hd__and2_1
XFILLER_0_47_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5186_ _2268_ _2272_ VGND VGND VPWR VPWR _2273_ sky130_fd_sc_hd__or2_1
X_4137_ _1425_ VGND VGND VPWR VPWR game.scoring_button_2.next_count\[5\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4068_ game.addmisses.add3.b\[1\] game.addmisses.add3.b\[0\] _1357_ _1330_ game.addmisses.add3.b\[2\]
+ VGND VGND VPWR VPWR _1373_ sky130_fd_sc_hd__a32o_1
X_3019_ disp_song.um.idx_note1\[0\] disp_song.um.idx_note1\[2\] disp_song.um.idx_note1\[3\]
+ _0179_ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__and4b_2
Xwire41 _0852_ VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3370_ game.addhits.a\[14\] game.addhits.add4.b\[2\] VGND VGND VPWR VPWR _0733_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5040_ _0169_ _1949_ VGND VGND VPWR VPWR _2132_ sky130_fd_sc_hd__or2_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5942_ clknet_leaf_46_clk game.scoring_button_1.next_flash_counter_1\[10\] net55
+ VGND VGND VPWR VPWR game.scoring_button_1.flash_counter_1\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_605 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5873_ clknet_leaf_20_clk _0056_ net63 VGND VGND VPWR VPWR game.padded_notes2\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4824_ _0232_ _0254_ _1436_ VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__o21a_1
XFILLER_0_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4755_ game.scoring_button_1.flash_counter_1\[4\] _1887_ game.hit_1 VGND VGND VPWR
+ VPWR _1890_ sky130_fd_sc_hd__a21boi_1
X_3706_ highest_score.highest_score\[1\] _1057_ _1054_ _1060_ _1061_ VGND VGND VPWR
+ VPWR _1062_ sky130_fd_sc_hd__o311a_1
XFILLER_0_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4686_ _1842_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_2\[5\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3637_ _0891_ _0893_ _0994_ _0941_ VGND VGND VPWR VPWR _0995_ sky130_fd_sc_hd__o31a_1
XFILLER_0_101_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3568_ _0214_ _0928_ _0930_ VGND VGND VPWR VPWR _0931_ sky130_fd_sc_hd__a21o_1
X_5307_ disp_song.note1\[10\] _2232_ _2389_ VGND VGND VPWR VPWR _2390_ sky130_fd_sc_hd__o21a_1
X_3499_ game.flash_counter\[6\] game.flash_counter\[7\] game.flash_counter\[9\] game.flash_counter\[8\]
+ VGND VGND VPWR VPWR _0862_ sky130_fd_sc_hd__o211a_1
X_5238_ _2199_ _2200_ _2185_ VGND VGND VPWR VPWR _2324_ sky130_fd_sc_hd__mux2_1
X_5169_ _2244_ _2252_ VGND VGND VPWR VPWR _2256_ sky130_fd_sc_hd__nor2_4
XPHY_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold6 disp_song.um.boton0e.sync_b VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2870_ disp_song.um.idx_note2\[1\] disp_song.um.idx_note2\[0\] disp_song.um.idx_note2\[2\]
+ VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__and3_1
XFILLER_0_45_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_10_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_10_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4540_ game.addmisses.a\[7\] _1730_ VGND VGND VPWR VPWR _1737_ sky130_fd_sc_hd__nand2_1
X_4471_ _1674_ VGND VGND VPWR VPWR _1675_ sky130_fd_sc_hd__clkbuf_8
X_3422_ _0659_ _0663_ VGND VGND VPWR VPWR _0785_ sky130_fd_sc_hd__nand2_1
X_6141_ clknet_leaf_30_clk disp_song.um.drum.next_note2\[21\] net69 VGND VGND VPWR
+ VPWR disp_song.note2\[21\] sky130_fd_sc_hd__dfstp_1
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3353_ _0590_ _0715_ _0591_ VGND VGND VPWR VPWR _0716_ sky130_fd_sc_hd__a21o_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6072_ clknet_leaf_7_clk _0155_ net59 VGND VGND VPWR VPWR game.scoring_button_1.acc\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_3284_ _0546_ _0560_ VGND VGND VPWR VPWR _0647_ sky130_fd_sc_hd__or2b_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5023_ _2020_ _2015_ VGND VGND VPWR VPWR _2115_ sky130_fd_sc_hd__nand2_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5925_ clknet_leaf_13_clk game.scoring_button_1.next_count\[16\] net58 VGND VGND
+ VPWR VPWR game.scoring_button_1.counts\[16\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5856_ clknet_leaf_66_clk game.scoring_button_1.next_num_hits\[5\] net47 VGND VGND
+ VPWR VPWR game.addhits.a\[5\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_63_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4807_ game.scoring_button_1.flash_counter_1\[19\] game.scoring_button_1.flash_counter_1\[20\]
+ _1922_ VGND VGND VPWR VPWR _1926_ sky130_fd_sc_hd__and3_1
X_2999_ disp_song.um.idx_note1\[3\] _0181_ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__nand2_1
XFILLER_0_63_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5787_ clknet_leaf_55_clk net104 net52 VGND VGND VPWR VPWR game.scoring_button_2.flash_counter_1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4738_ game.scoring_button_1.flash_counter_2\[21\] _1875_ VGND VGND VPWR VPWR _1879_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_9_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4669_ game.scoring_button_1.flash_counter_2\[0\] _1830_ VGND VGND VPWR VPWR _1831_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_3_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_68_clk clknet_3_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_68_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_98_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_59_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_59_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_89_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3971_ game.addhits.add4.b\[3\] _1227_ _1286_ _1226_ VGND VGND VPWR VPWR game.scoring_button_2.next_num_hits\[15\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2922_ _2671_ _0269_ _0164_ _0326_ _0328_ VGND VGND VPWR VPWR disp_song.um.drum.next_note2\[20\]
+ sky130_fd_sc_hd__a41o_1
X_5710_ clknet_leaf_39_clk net75 net66 VGND VGND VPWR VPWR modetrans.u2.Q1 sky130_fd_sc_hd__dfrtp_2
X_2853_ _0278_ VGND VGND VPWR VPWR disp_song.um.drum.next_note2\[2\] sky130_fd_sc_hd__buf_1
X_5641_ game.flash_counter\[9\] game.flash_counter\[8\] _2612_ game.flash_counter\[10\]
+ VGND VGND VPWR VPWR _2615_ sky130_fd_sc_hd__a31o_1
XFILLER_0_38_490 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5572_ _2573_ VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__clkbuf_1
X_2784_ _0209_ VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__buf_8
X_4523_ game.addmisses.a\[5\] _1713_ VGND VGND VPWR VPWR _1722_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4454_ game.addhits.a\[12\] _1654_ _1612_ VGND VGND VPWR VPWR _1662_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_111_576 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4385_ game.scoring_button_2.flash_counter_1\[21\] _1604_ VGND VGND VPWR VPWR _1607_
+ sky130_fd_sc_hd__and2_1
X_3405_ _0766_ _0767_ VGND VGND VPWR VPWR _0768_ sky130_fd_sc_hd__and2_1
X_6124_ clknet_leaf_23_clk disp_song.um.drum.next_note2\[4\] net64 VGND VGND VPWR
+ VPWR disp_song.note2\[4\] sky130_fd_sc_hd__dfrtp_1
X_3336_ _0697_ _0698_ VGND VGND VPWR VPWR _0699_ sky130_fd_sc_hd__and2_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6055_ clknet_leaf_8_clk _0011_ net60 VGND VGND VPWR VPWR game.counter\[11\] sky130_fd_sc_hd__dfrtp_2
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5006_ _0214_ _2098_ VGND VGND VPWR VPWR _2099_ sky130_fd_sc_hd__and2_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3267_ _0460_ _0629_ VGND VGND VPWR VPWR _0630_ sky130_fd_sc_hd__nor2_1
X_3198_ _0553_ _0555_ _0557_ VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__or3_2
XFILLER_0_95_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_95_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5908_ clknet_leaf_10_clk _0089_ net57 VGND VGND VPWR VPWR game.scoring_button_1.hit
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_8_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5839_ clknet_leaf_2_clk game.scoring_button_1.next_num_misses\[4\] net48 VGND VGND
+ VPWR VPWR game.addmisses.a\[4\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_32_600 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_98_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_460 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_110 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_26 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4170_ _1448_ VGND VGND VPWR VPWR game.scoring_button_2.next_count\[13\] sky130_fd_sc_hd__clkbuf_1
X_3121_ _0477_ _0482_ _0483_ VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__o21ba_2
X_3052_ _0384_ _0419_ _0423_ net204 VGND VGND VPWR VPWR disp_song.um.drum.next_note1\[23\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3954_ game.addhits.add3.b\[3\] _1272_ _1268_ VGND VGND VPWR VPWR _1274_ sky130_fd_sc_hd__o21ba_1
X_3885_ _0933_ _1219_ VGND VGND VPWR VPWR _1220_ sky130_fd_sc_hd__and2_1
XFILLER_0_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2905_ _0157_ _0265_ _0316_ disp_song.note2\[16\] VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__o31a_1
X_2836_ _0263_ VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__buf_2
XFILLER_0_73_577 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5624_ game.flash_counter\[5\] _2601_ VGND VGND VPWR VPWR _2602_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5555_ disp_song.note1\[16\] game.padded_notes1\[15\] _2541_ VGND VGND VPWR VPWR
+ _2562_ sky130_fd_sc_hd__mux2_1
X_2767_ pulseout.fin_pulse\[2\] pulseout.fin_pulse\[4\] pulseout.fin_pulse\[3\] VGND
+ VGND VPWR VPWR _0205_ sky130_fd_sc_hd__or3b_1
XFILLER_0_60_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2698_ _2670_ VGND VGND VPWR VPWR disp_song.um.drum.next_idx2\[0\] sky130_fd_sc_hd__clkbuf_8
X_5486_ disp_song.note2\[28\] game.padded_notes2\[27\] _2497_ VGND VGND VPWR VPWR
+ _2521_ sky130_fd_sc_hd__mux2_1
XFILLER_0_77_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4506_ _1675_ _1704_ _1705_ _1707_ VGND VGND VPWR VPWR game.scoring_button_1.next_num_misses\[2\]
+ sky130_fd_sc_hd__o31a_1
X_4437_ _1612_ _1645_ _1649_ net220 VGND VGND VPWR VPWR game.scoring_button_1.next_num_hits\[7\]
+ sky130_fd_sc_hd__a22o_1
X_6107_ clknet_leaf_41_clk disp_song.um.drum.next_note1\[19\] net67 VGND VGND VPWR
+ VPWR disp_song.note1\[19\] sky130_fd_sc_hd__dfstp_1
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4368_ _1595_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_1\[15\]
+ sky130_fd_sc_hd__clkbuf_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3319_ _0674_ _0681_ VGND VGND VPWR VPWR _0682_ sky130_fd_sc_hd__xnor2_2
X_4299_ _1546_ _1486_ _1547_ VGND VGND VPWR VPWR _1548_ sky130_fd_sc_hd__and3b_1
X_6038_ clknet_leaf_57_clk _0147_ net50 VGND VGND VPWR VPWR game.flash_counter\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_603 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3670_ _1021_ _1022_ _1024_ VGND VGND VPWR VPWR _1026_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_36 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5340_ highest_score.highest_score\[2\] _2414_ _2415_ _2416_ _2417_ VGND VGND VPWR
+ VPWR _2418_ sky130_fd_sc_hd__o221a_1
X_5271_ _2339_ _2353_ _2355_ VGND VGND VPWR VPWR _2356_ sky130_fd_sc_hd__o21ba_1
X_4222_ game.counter\[13\] game.counter\[12\] _1487_ _1488_ VGND VGND VPWR VPWR _1489_
+ sky130_fd_sc_hd__or4_1
X_4153_ _1437_ VGND VGND VPWR VPWR game.scoring_button_2.next_count\[9\] sky130_fd_sc_hd__clkbuf_1
X_4084_ game.addmisses.add4.b\[1\] _1379_ VGND VGND VPWR VPWR _1386_ sky130_fd_sc_hd__nor2_1
X_3104_ _0462_ _0465_ _0463_ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__o21a_1
X_3035_ _0411_ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_77_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4986_ _0169_ _2074_ _2078_ VGND VGND VPWR VPWR _2079_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3937_ _1253_ _1254_ _1258_ _1261_ VGND VGND VPWR VPWR _1262_ sky130_fd_sc_hd__a31o_1
XFILLER_0_46_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3868_ _1208_ VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_1
X_2819_ game.counter\[4\] game.counter\[17\] VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5607_ game.out\[3\] _2460_ _2462_ net115 VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3799_ _1049_ _1150_ _1137_ _0896_ VGND VGND VPWR VPWR _1151_ sky130_fd_sc_hd__a31o_1
XFILLER_0_103_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5538_ _2550_ game.padded_notes1\[10\] _2515_ VGND VGND VPWR VPWR _2551_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_111_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5469_ _2509_ VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__clkbuf_1
XTAP_1323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_522 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_544 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_476 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_558 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4840_ _1942_ VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4771_ game.scoring_button_1.flash_counter_1\[9\] _1898_ VGND VGND VPWR VPWR _1901_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_55_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3722_ disp_song.mi6.in\[3\] _0926_ VGND VGND VPWR VPWR _1078_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3653_ _0259_ _1007_ VGND VGND VPWR VPWR _1010_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_399 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5323_ _2221_ _2223_ disp_song.um.drum.next_idx1\[1\] VGND VGND VPWR VPWR _2405_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3584_ net40 _0854_ _0830_ _0834_ VGND VGND VPWR VPWR _0946_ sky130_fd_sc_hd__a2bb2o_1
X_5254_ _0175_ _2187_ _2252_ disp_song.um.drum.next_idx1\[2\] VGND VGND VPWR VPWR
+ _2339_ sky130_fd_sc_hd__o22a_2
X_4205_ _1473_ _1474_ VGND VGND VPWR VPWR _1475_ sky130_fd_sc_hd__and2_1
X_5185_ disp_song.um.drum.next_note1\[17\] _2191_ VGND VGND VPWR VPWR _2272_ sky130_fd_sc_hd__and2_1
X_4136_ _1405_ _0027_ VGND VGND VPWR VPWR _1425_ sky130_fd_sc_hd__and2_1
X_4067_ _1364_ _1371_ _1369_ game.addmisses.add3.b\[3\] VGND VGND VPWR VPWR _1372_
+ sky130_fd_sc_hd__a2bb2o_1
X_3018_ _0380_ _0398_ _0399_ net246 VGND VGND VPWR VPWR disp_song.um.drum.next_note1\[13\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4969_ disp_song.note2\[1\] disp_song.um.drum.next_note2\[0\] disp_song.um.drum.next_idx2\[0\]
+ VGND VGND VPWR VPWR _2063_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_100_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5941_ clknet_leaf_52_clk game.scoring_button_1.next_flash_counter_1\[9\] net55 VGND
+ VGND VPWR VPWR game.scoring_button_1.flash_counter_1\[9\] sky130_fd_sc_hd__dfrtp_1
X_5872_ clknet_leaf_29_clk _0055_ net69 VGND VGND VPWR VPWR game.padded_notes2\[5\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_75_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4823_ _0232_ _0254_ _1432_ VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__o21a_1
XFILLER_0_90_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4754_ _1889_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_1\[3\]
+ sky130_fd_sc_hd__clkbuf_1
X_3705_ highest_score.highest_score\[3\] highest_score.highest_score\[2\] _1052_ VGND
+ VGND VPWR VPWR _1061_ sky130_fd_sc_hd__or3_1
X_4685_ _1840_ game.missed_1 _1841_ VGND VGND VPWR VPWR _1842_ sky130_fd_sc_hd__and3b_1
XFILLER_0_31_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3636_ _0608_ _0675_ _0671_ _0886_ VGND VGND VPWR VPWR _0994_ sky130_fd_sc_hd__a31o_1
XFILLER_0_3_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3567_ _0352_ _0929_ VGND VGND VPWR VPWR _0930_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5306_ disp_song.um.drum.next_note1\[11\] _2191_ disp_song.um.drum.next_idx1\[1\]
+ VGND VGND VPWR VPWR _2389_ sky130_fd_sc_hd__a21o_1
X_3498_ _0840_ _0859_ _0860_ VGND VGND VPWR VPWR _0861_ sky130_fd_sc_hd__o21ai_1
X_5237_ _0191_ _0197_ VGND VGND VPWR VPWR _2323_ sky130_fd_sc_hd__nand2_1
X_5168_ _2249_ _2251_ _2254_ VGND VGND VPWR VPWR _2255_ sky130_fd_sc_hd__mux2_1
X_4119_ game.scoring_button_2.check_hit.in _0248_ _1415_ VGND VGND VPWR VPWR _1416_
+ sky130_fd_sc_hd__and3_1
X_5099_ disp_song.um.drum.next_idx1\[2\] disp_song.um.drum.next_idx1\[1\] VGND VGND
+ VPWR VPWR _2187_ sky130_fd_sc_hd__nand2_2
XFILLER_0_39_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_506 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_580 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold7 modetrans.u3.Q1 VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_108 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4470_ game.scoring_button_1.hit _1673_ VGND VGND VPWR VPWR _1674_ sky130_fd_sc_hd__or2_1
X_3421_ _0782_ _0783_ VGND VGND VPWR VPWR _0784_ sky130_fd_sc_hd__nor2_1
X_6140_ clknet_leaf_28_clk disp_song.um.drum.next_note2\[20\] net68 VGND VGND VPWR
+ VPWR disp_song.note2\[20\] sky130_fd_sc_hd__dfrtp_1
X_3352_ _0585_ _0592_ VGND VGND VPWR VPWR _0715_ sky130_fd_sc_hd__or2b_1
XFILLER_0_21_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3283_ _0640_ _0645_ _0643_ VGND VGND VPWR VPWR _0646_ sky130_fd_sc_hd__o21ai_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6071_ clknet_leaf_10_clk _0154_ net61 VGND VGND VPWR VPWR game.scoring_button_1.acc\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_5022_ _2020_ _2111_ _2105_ _2113_ VGND VGND VPWR VPWR _2114_ sky130_fd_sc_hd__o211a_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5924_ clknet_leaf_13_clk game.scoring_button_1.next_count\[15\] net58 VGND VGND
+ VPWR VPWR game.scoring_button_1.counts\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5855_ clknet_3_1__leaf_clk game.scoring_button_1.next_num_hits\[4\] net48 VGND VGND
+ VPWR VPWR game.addhits.a\[4\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_63_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4806_ net172 _1922_ _1925_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_1\[19\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_35_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2998_ _0380_ _0384_ _0385_ net268 VGND VGND VPWR VPWR disp_song.um.drum.next_note1\[7\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5786_ clknet_leaf_55_clk game.scoring_button_2.next_flash_counter_1\[0\] net52 VGND
+ VGND VPWR VPWR game.scoring_button_2.flash_counter_1\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_56_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4737_ game.scoring_button_1.flash_counter_2\[21\] _1875_ VGND VGND VPWR VPWR _1878_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_71_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4668_ _1791_ _1495_ _1508_ net127 VGND VGND VPWR VPWR game.scoring_button_1.next_start_count
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3619_ _0259_ _0977_ VGND VGND VPWR VPWR _0979_ sky130_fd_sc_hd__nor2_1
X_4599_ _1784_ _1787_ game.addmisses.a\[15\] VGND VGND VPWR VPWR _1788_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3970_ _1283_ _1285_ VGND VGND VPWR VPWR _1286_ sky130_fd_sc_hd__nor2_1
X_2921_ _0163_ _0327_ disp_song.note2\[20\] VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__o21a_1
XFILLER_0_57_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2852_ _0269_ disp_song.note2\[2\] _0277_ VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__mux2_1
X_5640_ _2602_ _2604_ _2605_ _2609_ VGND VGND VPWR VPWR _2614_ sky130_fd_sc_hd__or4_2
XFILLER_0_5_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5571_ _2572_ net225 _2472_ VGND VGND VPWR VPWR _2573_ sky130_fd_sc_hd__mux2_1
X_2783_ _0214_ _0217_ _0218_ modetrans.mode\[5\] VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__a22o_1
X_4522_ game.addmisses.a\[6\] _1720_ game.addmisses.a\[7\] VGND VGND VPWR VPWR _1721_
+ sky130_fd_sc_hd__o21a_2
XFILLER_0_53_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_111_511 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4453_ game.addhits.a\[12\] _1654_ VGND VGND VPWR VPWR _1661_ sky130_fd_sc_hd__and2_1
XFILLER_0_111_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3404_ _0512_ _0524_ _0527_ VGND VGND VPWR VPWR _0767_ sky130_fd_sc_hd__or3b_2
X_4384_ _1606_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_1\[20\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6123_ clknet_leaf_22_clk disp_song.um.drum.next_note2\[3\] net60 VGND VGND VPWR
+ VPWR disp_song.note2\[3\] sky130_fd_sc_hd__dfstp_1
X_3335_ _0600_ _0598_ VGND VGND VPWR VPWR _0698_ sky130_fd_sc_hd__nor2_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6054_ clknet_leaf_8_clk _0010_ net60 VGND VGND VPWR VPWR game.counter\[10\] sky130_fd_sc_hd__dfrtp_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3266_ _0454_ _0468_ VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__xnor2_4
X_5005_ _2087_ _2096_ _2097_ VGND VGND VPWR VPWR _2098_ sky130_fd_sc_hd__mux2_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3197_ _0553_ _0558_ _0559_ VGND VGND VPWR VPWR _0560_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_76_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5907_ clknet_leaf_45_clk game.scoring_button_1.next_good net54 VGND VGND VPWR VPWR
+ game.hit_1 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_48_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5838_ clknet_leaf_2_clk game.scoring_button_1.next_num_misses\[3\] net49 VGND VGND
+ VPWR VPWR game.addmisses.a\[3\] sky130_fd_sc_hd__dfrtp_4
X_5769_ clknet_leaf_17_clk game.scoring_button_2.next_count\[6\] net62 VGND VGND VPWR
+ VPWR game.scoring_button_2.counts\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_612 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_98_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_472 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_38 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3120_ _0478_ _0481_ _0479_ VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_93_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3051_ _0384_ _0421_ VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3953_ _1226_ _1271_ _1273_ _1227_ net198 VGND VGND VPWR VPWR game.scoring_button_2.next_num_hits\[10\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_42_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2904_ _2661_ disp_song.um.idx_note2\[4\] VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__nand2_1
X_3884_ _0966_ disp_song.display_note2\[5\] _0210_ game.out\[5\] _0208_ VGND VGND
+ VPWR VPWR _1219_ sky130_fd_sc_hd__a221o_2
XFILLER_0_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2835_ modetrans.mode\[2\] _2658_ _2659_ VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__and3_1
X_5623_ _0868_ _2595_ VGND VGND VPWR VPWR _2601_ sky130_fd_sc_hd__and2_1
X_5554_ _2561_ VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__clkbuf_1
X_2766_ pulseout.fin_pulse\[5\] VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__inv_2
XFILLER_0_14_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2697_ _2669_ VGND VGND VPWR VPWR _2670_ sky130_fd_sc_hd__inv_2
X_5485_ _2520_ VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_486 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4505_ game.addmisses.a\[2\] _1693_ _1706_ _1699_ VGND VGND VPWR VPWR _1707_ sky130_fd_sc_hd__a211o_1
XFILLER_0_111_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4436_ _1642_ _1643_ _1612_ _1638_ _1613_ VGND VGND VPWR VPWR _1649_ sky130_fd_sc_hd__a41o_1
XFILLER_0_1_583 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4367_ _1593_ game.hit_2 _1594_ VGND VGND VPWR VPWR _1595_ sky130_fd_sc_hd__and3b_1
X_6106_ clknet_leaf_38_clk disp_song.um.drum.next_note1\[18\] net67 VGND VGND VPWR
+ VPWR disp_song.note1\[18\] sky130_fd_sc_hd__dfstp_1
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3318_ _0678_ _0677_ VGND VGND VPWR VPWR _0681_ sky130_fd_sc_hd__and2b_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4298_ game.scoring_button_2.flash_counter_2\[15\] game.scoring_button_2.flash_counter_2\[16\]
+ _1539_ game.scoring_button_2.flash_counter_2\[17\] VGND VGND VPWR VPWR _1547_ sky130_fd_sc_hd__a31o_1
X_6037_ clknet_leaf_58_clk _0146_ net50 VGND VGND VPWR VPWR game.flash_counter\[17\]
+ sky130_fd_sc_hd__dfrtp_2
X_3249_ _0471_ VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__inv_2
XTAP_1505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_615 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_523 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_48 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5270_ _2254_ _2277_ _2339_ _2354_ VGND VGND VPWR VPWR _2355_ sky130_fd_sc_hd__o211a_1
X_4221_ game.counter\[4\] game.counter\[16\] game.counter\[17\] game.counter\[5\]
+ VGND VGND VPWR VPWR _1488_ sky130_fd_sc_hd__or4b_1
X_4152_ _1405_ _1436_ VGND VGND VPWR VPWR _1437_ sky130_fd_sc_hd__and2_1
X_4083_ game.addmisses.add4.b\[0\] game.addmisses.add4.b\[1\] _1363_ VGND VGND VPWR
+ VPWR _1385_ sky130_fd_sc_hd__and3_2
X_3103_ _0464_ _0465_ VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__xnor2_4
X_3034_ _2661_ _0265_ _0357_ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__or3_1
XFILLER_0_53_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4985_ disp_song.um.drum.next_idx2\[2\] _1962_ _2077_ VGND VGND VPWR VPWR _2078_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3936_ _1226_ _1260_ VGND VGND VPWR VPWR _1261_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3867_ _0933_ _1207_ VGND VGND VPWR VPWR _1208_ sky130_fd_sc_hd__and2_1
XFILLER_0_33_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2818_ game.counter\[3\] game.counter\[2\] _0248_ VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__or3_1
X_5606_ net101 _2460_ _2462_ game.out\[3\] VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__a22o_1
X_3798_ _1125_ VGND VGND VPWR VPWR _1150_ sky130_fd_sc_hd__inv_2
X_5537_ disp_song.note1\[10\] game.padded_notes1\[9\] _2541_ VGND VGND VPWR VPWR _2550_
+ sky130_fd_sc_hd__mux2_1
X_2749_ _0191_ VGND VGND VPWR VPWR disp_song.um.drum.next_idx1\[2\] sky130_fd_sc_hd__clkinv_4
XFILLER_0_103_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5468_ _2508_ net211 _2473_ VGND VGND VPWR VPWR _2509_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5399_ _2461_ VGND VGND VPWR VPWR _2462_ sky130_fd_sc_hd__buf_6
XFILLER_0_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4419_ _1612_ _1632_ _1635_ _1613_ net202 VGND VGND VPWR VPWR game.scoring_button_1.next_num_hits\[3\]
+ sky130_fd_sc_hd__a32o_1
XTAP_1302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_74_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_662 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4770_ _1900_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_1\[8\]
+ sky130_fd_sc_hd__clkbuf_1
X_3721_ disp_song.mi6.in\[0\] VGND VGND VPWR VPWR _1077_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_15_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_334 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3652_ _1003_ _0991_ _1008_ _0211_ net38 VGND VGND VPWR VPWR _1009_ sky130_fd_sc_hd__o221a_1
X_3583_ _0258_ _0944_ VGND VGND VPWR VPWR _0945_ sky130_fd_sc_hd__nor2_1
X_5322_ _2318_ _2403_ _0191_ VGND VGND VPWR VPWR _2404_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5253_ _2335_ _2337_ _2254_ VGND VGND VPWR VPWR _2338_ sky130_fd_sc_hd__mux2_1
X_4204_ game.counter\[21\] _1470_ VGND VGND VPWR VPWR _1474_ sky130_fd_sc_hd__nand2_1
X_5184_ _0175_ disp_song.um.drum.next_note1\[16\] VGND VGND VPWR VPWR _2271_ sky130_fd_sc_hd__or2_1
X_4135_ _1423_ _1424_ VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__nor2_1
X_4066_ _1369_ _1370_ VGND VGND VPWR VPWR _1371_ sky130_fd_sc_hd__or2_1
X_3017_ _0382_ _0398_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4968_ _2057_ _2061_ _2034_ VGND VGND VPWR VPWR _2062_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_640 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4899_ _1956_ disp_song.um.drum.next_note2\[13\] _1993_ VGND VGND VPWR VPWR _1994_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_80_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3919_ _1246_ _1247_ VGND VGND VPWR VPWR _1248_ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_406 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5940_ clknet_leaf_46_clk game.scoring_button_1.next_flash_counter_1\[8\] net55 VGND
+ VGND VPWR VPWR game.scoring_button_1.flash_counter_1\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_618 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5871_ clknet_leaf_22_clk _0054_ net64 VGND VGND VPWR VPWR game.padded_notes2\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4822_ _1934_ VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4753_ _1887_ game.hit_1 _1888_ VGND VGND VPWR VPWR _1889_ sky130_fd_sc_hd__and3b_1
XFILLER_0_50_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3704_ _0255_ _1059_ VGND VGND VPWR VPWR _1060_ sky130_fd_sc_hd__and2_1
XFILLER_0_50_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4684_ game.scoring_button_1.flash_counter_2\[3\] game.scoring_button_1.flash_counter_2\[4\]
+ _1833_ game.scoring_button_1.flash_counter_2\[5\] VGND VGND VPWR VPWR _1841_ sky130_fd_sc_hd__a31o_1
XFILLER_0_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3635_ _0919_ _0970_ _0992_ _0915_ VGND VGND VPWR VPWR _0993_ sky130_fd_sc_hd__a211o_1
XFILLER_0_11_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3566_ disp_song.mi6.in\[3\] disp_song.mi6.in\[2\] _0925_ VGND VGND VPWR VPWR _0929_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_11_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3497_ _0855_ _0835_ _0840_ VGND VGND VPWR VPWR _0860_ sky130_fd_sc_hd__or3b_1
X_5305_ _2383_ _2386_ _2387_ VGND VGND VPWR VPWR _2388_ sky130_fd_sc_hd__mux2_1
X_5236_ _0191_ _0197_ _2317_ _2319_ _2321_ VGND VGND VPWR VPWR _2322_ sky130_fd_sc_hd__o311a_1
XFILLER_0_52_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5167_ _2253_ VGND VGND VPWR VPWR _2254_ sky130_fd_sc_hd__buf_4
XFILLER_0_98_507 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4118_ game.counter\[1\] game.counter\[0\] VGND VGND VPWR VPWR _1415_ sky130_fd_sc_hd__nand2_1
X_5098_ disp_song.um.drum.next_idx1\[2\] disp_song.um.drum.next_idx1\[3\] VGND VGND
+ VPWR VPWR _2186_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4049_ _1355_ VGND VGND VPWR VPWR _1356_ sky130_fd_sc_hd__inv_2
XPHY_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_640 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_104_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_584 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold8 game.scoring_button_1.check_hit.edge_1 VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_57_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_651 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3420_ _0673_ _0672_ _0665_ VGND VGND VPWR VPWR _0783_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_52_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3351_ _0712_ _0709_ _0713_ VGND VGND VPWR VPWR _0714_ sky130_fd_sc_hd__a21o_1
XFILLER_0_0_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3282_ _0643_ _0644_ VGND VGND VPWR VPWR _0645_ sky130_fd_sc_hd__nand2_1
X_6070_ clknet_leaf_62_clk highest_score.nxt_mode\[1\] net53 VGND VGND VPWR VPWR highest_score.score_mode\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5021_ _2028_ _2112_ _2042_ VGND VGND VPWR VPWR _2113_ sky130_fd_sc_hd__a21o_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5923_ clknet_leaf_8_clk game.scoring_button_1.next_count\[14\] net60 VGND VGND VPWR
+ VPWR game.scoring_button_1.counts\[14\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_40 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5854_ clknet_leaf_4_clk game.scoring_button_1.next_num_hits\[3\] net49 VGND VGND
+ VPWR VPWR game.addhits.a\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4805_ net172 _1922_ _1799_ VGND VGND VPWR VPWR _1925_ sky130_fd_sc_hd__a21boi_1
X_2997_ _0382_ _0384_ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__nand2_1
X_5785_ clknet_leaf_11_clk game.scoring_button_2.next_count\[22\] net57 VGND VGND
+ VPWR VPWR game.scoring_button_2.counts\[22\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4736_ _1877_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_2\[20\]
+ sky130_fd_sc_hd__clkbuf_1
X_4667_ _1791_ _1689_ _1830_ VGND VGND VPWR VPWR game.scoring_button_1.next_missed
+ sky130_fd_sc_hd__o21bai_1
XFILLER_0_9_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3618_ _0879_ _0977_ VGND VGND VPWR VPWR _0978_ sky130_fd_sc_hd__nand2_1
XFILLER_0_101_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4598_ game.addmisses.a\[14\] game.addmisses.a\[13\] _1765_ VGND VGND VPWR VPWR _1787_
+ sky130_fd_sc_hd__or3_1
X_3549_ _0717_ _0767_ _0911_ _0504_ VGND VGND VPWR VPWR _0912_ sky130_fd_sc_hd__or4b_4
XFILLER_0_86_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5219_ _2293_ _2305_ _2280_ VGND VGND VPWR VPWR _2306_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_610 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2920_ disp_song.um.idx_note2\[4\] _2660_ _2675_ disp_song.next_red VGND VGND VPWR
+ VPWR _0327_ sky130_fd_sc_hd__nand4_2
XFILLER_0_9_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2851_ _0276_ disp_song.um.idx_note2\[3\] _0161_ VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__or3b_1
XFILLER_0_110_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5570_ disp_song.note1\[21\] game.padded_notes1\[20\] _2541_ VGND VGND VPWR VPWR
+ _2572_ sky130_fd_sc_hd__mux2_1
X_2782_ _0217_ _0203_ _0206_ VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__nor3b_2
XFILLER_0_26_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4521_ game.addmisses.a\[5\] _1713_ VGND VGND VPWR VPWR _1720_ sky130_fd_sc_hd__or2_1
X_4452_ net228 _1613_ _1660_ _1612_ VGND VGND VPWR VPWR game.scoring_button_1.next_num_hits\[11\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_111_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3403_ _0765_ _0739_ _0745_ VGND VGND VPWR VPWR _0766_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4383_ _1604_ game.hit_2 _1605_ VGND VGND VPWR VPWR _1606_ sky130_fd_sc_hd__and3b_1
XFILLER_0_21_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6122_ clknet_leaf_22_clk disp_song.um.drum.next_note2\[2\] net60 VGND VGND VPWR
+ VPWR disp_song.note2\[2\] sky130_fd_sc_hd__dfrtp_1
X_3334_ _0579_ _0696_ VGND VGND VPWR VPWR _0697_ sky130_fd_sc_hd__xnor2_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6053_ clknet_leaf_15_clk _0031_ net63 VGND VGND VPWR VPWR game.counter\[9\] sky130_fd_sc_hd__dfrtp_4
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3265_ _0466_ _0626_ _0627_ VGND VGND VPWR VPWR _0628_ sky130_fd_sc_hd__a21o_1
X_5004_ _1960_ _2085_ VGND VGND VPWR VPWR _2097_ sky130_fd_sc_hd__nor2_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3196_ _0554_ _0557_ _0555_ VGND VGND VPWR VPWR _0559_ sky130_fd_sc_hd__o21a_1
XFILLER_0_88_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5906_ clknet_leaf_25_clk game.scoring_button_1.next_missed net64 VGND VGND VPWR
+ VPWR game.missed_1 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_48_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5837_ clknet_leaf_73_clk game.scoring_button_1.next_num_misses\[2\] net49 VGND VGND
+ VPWR VPWR game.addmisses.a\[2\] sky130_fd_sc_hd__dfrtp_2
X_5768_ clknet_leaf_17_clk game.scoring_button_2.next_count\[5\] net62 VGND VGND VPWR
+ VPWR game.scoring_button_2.counts\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4719_ _1864_ game.missed_1 _1865_ VGND VGND VPWR VPWR _1866_ sky130_fd_sc_hd__and3b_1
XFILLER_0_71_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5699_ clknet_leaf_62_clk _0035_ net53 VGND VGND VPWR VPWR highest_score.highest_score\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_102_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_99_602 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_98_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_93_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3050_ _0381_ _0419_ _0422_ net205 VGND VGND VPWR VPWR disp_song.um.drum.next_note1\[22\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3952_ _1269_ game.addhits.add3.b\[3\] _1272_ VGND VGND VPWR VPWR _1273_ sky130_fd_sc_hd__mux2_1
X_2903_ _0315_ VGND VGND VPWR VPWR disp_song.um.drum.next_note2\[15\] sky130_fd_sc_hd__buf_1
X_3883_ _1218_ VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_1
X_5622_ net146 _2600_ VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__xnor2_1
X_2834_ _0256_ _0262_ VGND VGND VPWR VPWR highest_score.nxt_mode\[1\] sky130_fd_sc_hd__xnor2_1
X_5553_ _2560_ game.padded_notes1\[15\] _2472_ VGND VGND VPWR VPWR _2561_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2765_ modetrans.u3.Q2 modetrans.u3.Q1 VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__and2b_1
XFILLER_0_14_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4504_ _1691_ _1703_ VGND VGND VPWR VPWR _1706_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5484_ _2519_ game.padded_notes2\[27\] _2515_ VGND VGND VPWR VPWR _2520_ sky130_fd_sc_hd__mux2_1
X_2696_ disp_song.um.idx_note2\[0\] _2662_ _2668_ VGND VGND VPWR VPWR _2669_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_13_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4435_ _1645_ _1648_ net257 _1613_ VGND VGND VPWR VPWR game.scoring_button_1.next_num_hits\[6\]
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_41_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_595 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4366_ game.scoring_button_2.flash_counter_1\[15\] _1590_ VGND VGND VPWR VPWR _1594_
+ sky130_fd_sc_hd__or2_1
X_6105_ clknet_leaf_42_clk disp_song.um.drum.next_note1\[17\] net67 VGND VGND VPWR
+ VPWR disp_song.note1\[17\] sky130_fd_sc_hd__dfrtp_2
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3317_ _0622_ _0679_ VGND VGND VPWR VPWR _0680_ sky130_fd_sc_hd__xor2_2
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4297_ game.scoring_button_2.flash_counter_2\[17\] game.scoring_button_2.flash_counter_2\[16\]
+ _1542_ VGND VGND VPWR VPWR _1546_ sky130_fd_sc_hd__and3_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6036_ clknet_leaf_58_clk _0145_ net50 VGND VGND VPWR VPWR game.flash_counter\[16\]
+ sky130_fd_sc_hd__dfrtp_4
X_3248_ _0483_ VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__inv_2
X_3179_ game.addhits.a\[4\] game.addhits.add2.b\[0\] VGND VGND VPWR VPWR _0542_ sky130_fd_sc_hd__nor2_1
XTAP_1506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_107_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_107_648 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_535 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4220_ game.counter\[6\] game.counter\[7\] VGND VGND VPWR VPWR _1487_ sky130_fd_sc_hd__nand2_1
X_4151_ _1434_ _1435_ VGND VGND VPWR VPWR _1436_ sky130_fd_sc_hd__nor2_1
XFILLER_0_37_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4082_ _1289_ _1379_ _1380_ _1384_ VGND VGND VPWR VPWR game.scoring_button_2.next_num_misses\[12\]
+ sky130_fd_sc_hd__o31ai_1
X_3102_ _0456_ _0457_ _0458_ VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__o21a_2
X_3033_ _0264_ _0409_ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__nand2_2
X_4984_ _2075_ _2076_ _2667_ VGND VGND VPWR VPWR _2077_ sky130_fd_sc_hd__mux2_1
X_3935_ game.addhits.add2.b\[1\] game.addhits.add2.b\[0\] _1244_ game.addhits.add2.b\[2\]
+ VGND VGND VPWR VPWR _1260_ sky130_fd_sc_hd__a31o_1
XFILLER_0_46_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5605_ net119 _2460_ _2462_ net101 VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3866_ _0966_ disp_song.display_note1\[6\] _0211_ game.out\[13\] _0208_ VGND VGND
+ VPWR VPWR _1207_ sky130_fd_sc_hd__a221o_2
X_2817_ game.counter\[1\] game.counter\[0\] VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__or2_1
XFILLER_0_82_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3797_ _1142_ _1149_ _0935_ VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__o21a_1
X_5536_ _2549_ VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__clkbuf_1
X_2748_ _0190_ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__buf_4
X_5467_ disp_song.note2\[22\] game.padded_notes2\[21\] _2497_ VGND VGND VPWR VPWR
+ _2508_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4418_ _1621_ _1627_ _1629_ VGND VGND VPWR VPWR _1635_ sky130_fd_sc_hd__o21ai_1
X_5398_ _2458_ _2460_ VGND VGND VPWR VPWR _2461_ sky130_fd_sc_hd__nor2_1
X_4349_ net156 _1579_ game.hit_2 VGND VGND VPWR VPWR _1582_ sky130_fd_sc_hd__a21boi_1
X_6019_ clknet_leaf_5_clk net94 net60 VGND VGND VPWR VPWR game.out\[6\] sky130_fd_sc_hd__dfrtp_1
XTAP_1303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3720_ lvls.level\[2\] lvls.level\[1\] modetrans.mode\[5\] VGND VGND VPWR VPWR _1076_
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_99_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_40_clk clknet_3_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_40_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_15_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3651_ _1007_ VGND VGND VPWR VPWR _1008_ sky130_fd_sc_hd__inv_2
X_3582_ highest_score.highest_score\[5\] highest_score.highest_score\[4\] _0255_ _0943_
+ VGND VGND VPWR VPWR _0944_ sky130_fd_sc_hd__o211a_1
X_5321_ _2228_ _2364_ disp_song.um.drum.next_idx1\[1\] VGND VGND VPWR VPWR _2403_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5252_ disp_song.um.drum.next_idx1\[0\] disp_song.um.drum.next_note1\[9\] _2290_
+ _2336_ VGND VGND VPWR VPWR _2337_ sky130_fd_sc_hd__o211a_1
X_4203_ game.counter\[21\] _1470_ VGND VGND VPWR VPWR _1473_ sky130_fd_sc_hd__or2_1
X_5183_ _2267_ _2269_ _2254_ VGND VGND VPWR VPWR _2270_ sky130_fd_sc_hd__mux2_1
X_4134_ game.counter\[4\] _1418_ game.counter\[5\] VGND VGND VPWR VPWR _1424_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4065_ game.addmisses.add3.b\[1\] _1355_ game.addmisses.add3.b\[2\] VGND VGND VPWR
+ VPWR _1370_ sky130_fd_sc_hd__a21oi_1
X_3016_ _0179_ disp_song.um.idx_note1\[3\] disp_song.um.idx_note1\[2\] disp_song.um.idx_note1\[0\]
+ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__and4b_1
XFILLER_0_93_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4967_ _2059_ _2060_ _2020_ VGND VGND VPWR VPWR _2061_ sky130_fd_sc_hd__mux2_1
XFILLER_0_93_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_31_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_31_clk sky130_fd_sc_hd__clkbuf_16
X_4898_ _2670_ disp_song.um.drum.next_note2\[12\] VGND VGND VPWR VPWR _1993_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3918_ _1237_ _1244_ _1240_ VGND VGND VPWR VPWR _1247_ sky130_fd_sc_hd__a21o_1
XFILLER_0_61_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3849_ _0933_ _1195_ VGND VGND VPWR VPWR _1196_ sky130_fd_sc_hd__and2_1
XFILLER_0_104_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5519_ _2537_ net218 _2515_ VGND VGND VPWR VPWR _2538_ sky130_fd_sc_hd__mux2_1
XFILLER_0_89_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_621 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_641 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_22_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_22_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_25_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_110_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5870_ clknet_leaf_22_clk _0053_ net60 VGND VGND VPWR VPWR game.padded_notes2\[3\]
+ sky130_fd_sc_hd__dfstp_1
X_4821_ _0032_ _1430_ VGND VGND VPWR VPWR _1934_ sky130_fd_sc_hd__and2b_1
XFILLER_0_47_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_13_clk clknet_3_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_13_clk sky130_fd_sc_hd__clkbuf_16
X_4752_ game.scoring_button_1.flash_counter_1\[3\] _1884_ VGND VGND VPWR VPWR _1888_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4683_ game.scoring_button_1.flash_counter_2\[5\] game.scoring_button_1.flash_counter_2\[4\]
+ _1836_ VGND VGND VPWR VPWR _1840_ sky130_fd_sc_hd__and3_1
XFILLER_0_43_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3703_ _1055_ _1058_ VGND VGND VPWR VPWR _1059_ sky130_fd_sc_hd__nand2_1
X_3634_ _0667_ _0969_ _0914_ VGND VGND VPWR VPWR _0992_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_50_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3565_ _0925_ _0927_ VGND VGND VPWR VPWR _0928_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3496_ _0857_ _0858_ _0847_ VGND VGND VPWR VPWR _0859_ sky130_fd_sc_hd__or3b_1
X_5304_ _0197_ _2246_ VGND VGND VPWR VPWR _2387_ sky130_fd_sc_hd__xnor2_2
X_5235_ disp_song.um.drum.next_idx1\[2\] _2320_ disp_song.um.drum.next_idx1\[3\] VGND
+ VGND VPWR VPWR _2321_ sky130_fd_sc_hd__a21o_1
XFILLER_0_45_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5166_ _2244_ _2252_ VGND VGND VPWR VPWR _2253_ sky130_fd_sc_hd__or2_1
XFILLER_0_98_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4117_ _1414_ VGND VGND VPWR VPWR game.scoring_button_2.next_count\[0\] sky130_fd_sc_hd__clkbuf_1
X_5097_ _0199_ VGND VGND VPWR VPWR _2185_ sky130_fd_sc_hd__buf_6
X_4048_ game.addmisses.add3.b\[0\] _1335_ VGND VGND VPWR VPWR _1355_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5999_ clknet_leaf_38_clk _0108_ net66 VGND VGND VPWR VPWR game.padded_notes1\[18\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_93_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_652 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold9 modetrans.u2.Q1 VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_108_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_110_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3350_ _0704_ _0707_ VGND VGND VPWR VPWR _0713_ sky130_fd_sc_hd__and2_1
XFILLER_0_21_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5020_ disp_song.um.drum.next_note2\[25\] _1968_ _2667_ VGND VGND VPWR VPWR _2112_
+ sky130_fd_sc_hd__a21o_1
X_3281_ _0628_ _0629_ _0642_ VGND VGND VPWR VPWR _0644_ sky130_fd_sc_hd__a21o_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_2_clk clknet_3_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_2_clk sky130_fd_sc_hd__clkbuf_16
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5922_ clknet_leaf_8_clk game.scoring_button_1.next_count\[13\] net60 VGND VGND VPWR
+ VPWR game.scoring_button_1.counts\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5853_ clknet_leaf_4_clk game.scoring_button_1.next_num_hits\[2\] net49 VGND VGND
+ VPWR VPWR game.addhits.a\[2\] sky130_fd_sc_hd__dfrtp_2
X_5784_ clknet_leaf_11_clk game.scoring_button_2.next_count\[21\] net57 VGND VGND
+ VPWR VPWR game.scoring_button_2.counts\[21\] sky130_fd_sc_hd__dfrtp_1
X_4804_ _1924_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_1\[18\]
+ sky130_fd_sc_hd__clkbuf_1
X_4735_ _1875_ game.missed_1 _1876_ VGND VGND VPWR VPWR _1877_ sky130_fd_sc_hd__and3b_1
X_2996_ disp_song.um.idx_note1\[0\] disp_song.um.idx_note1\[2\] _0177_ _0179_ VGND
+ VGND VPWR VPWR _0384_ sky130_fd_sc_hd__and4_1
XFILLER_0_8_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4666_ _1823_ _1824_ _1829_ game.missed_1 VGND VGND VPWR VPWR _1830_ sky130_fd_sc_hd__o31a_2
XFILLER_0_31_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4597_ _1786_ VGND VGND VPWR VPWR game.scoring_button_1.next_num_misses\[14\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3617_ _0972_ _0974_ _0976_ _0921_ VGND VGND VPWR VPWR _0977_ sky130_fd_sc_hd__a31o_1
XFILLER_0_43_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_101_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3548_ _0617_ _0910_ _0597_ VGND VGND VPWR VPWR _0911_ sky130_fd_sc_hd__a21o_1
XFILLER_0_12_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_86_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3479_ _0762_ _0824_ _0825_ _0826_ VGND VGND VPWR VPWR _0842_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_86_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5218_ _2247_ _2297_ _2301_ _2304_ VGND VGND VPWR VPWR _2305_ sky130_fd_sc_hd__o22a_1
XFILLER_0_98_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5149_ _2185_ _2236_ VGND VGND VPWR VPWR _2237_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_79_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2850_ disp_song.um.idx_note2\[0\] disp_song.um.idx_note2\[2\] disp_song.um.idx_note2\[1\]
+ VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__or3b_2
XFILLER_0_72_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2781_ _0207_ _0215_ _0208_ _0217_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_31_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4520_ _1712_ _1714_ _1719_ _1675_ VGND VGND VPWR VPWR game.scoring_button_1.next_num_misses\[4\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4451_ game.addhits.a\[11\] _1658_ _1654_ VGND VGND VPWR VPWR _1660_ sky130_fd_sc_hd__o21ba_1
X_3402_ _0738_ _0730_ _0747_ VGND VGND VPWR VPWR _0765_ sky130_fd_sc_hd__a21o_1
XFILLER_0_40_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_111_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6121_ clknet_leaf_22_clk disp_song.um.drum.next_note2\[1\] net60 VGND VGND VPWR
+ VPWR disp_song.note2\[1\] sky130_fd_sc_hd__dfstp_1
X_4382_ game.scoring_button_2.flash_counter_1\[19\] game.scoring_button_2.flash_counter_1\[18\]
+ _1597_ game.scoring_button_2.flash_counter_1\[20\] VGND VGND VPWR VPWR _1605_ sky130_fd_sc_hd__a31o_1
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3333_ _0591_ _0592_ VGND VGND VPWR VPWR _0696_ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6052_ clknet_leaf_14_clk _0030_ net58 VGND VGND VPWR VPWR game.counter\[8\] sky130_fd_sc_hd__dfrtp_2
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3264_ _0461_ _0466_ VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5003_ _2092_ _2095_ _2086_ VGND VGND VPWR VPWR _2096_ sky130_fd_sc_hd__mux2_1
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3195_ _0556_ _0557_ VGND VGND VPWR VPWR _0558_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_76_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_72_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5905_ clknet_leaf_44_clk _0088_ net54 VGND VGND VPWR VPWR game.out\[13\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5836_ clknet_leaf_0_clk game.scoring_button_1.next_num_misses\[1\] net49 VGND VGND
+ VPWR VPWR game.addmisses.a\[1\] sky130_fd_sc_hd__dfrtp_4
X_5767_ clknet_leaf_15_clk game.scoring_button_2.next_count\[4\] net62 VGND VGND VPWR
+ VPWR game.scoring_button_2.counts\[4\] sky130_fd_sc_hd__dfrtp_1
X_2979_ disp_song.um.idx_note1\[3\] _0370_ VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4718_ game.scoring_button_1.flash_counter_2\[15\] _1861_ VGND VGND VPWR VPWR _1865_
+ sky130_fd_sc_hd__or2_1
X_5698_ clknet_leaf_1_clk _0034_ net48 VGND VGND VPWR VPWR game.scoring_button_2.acc\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_4649_ _1791_ _1463_ VGND VGND VPWR VPWR _1818_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_97_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3951_ game.addhits.add3.b\[2\] _1267_ VGND VGND VPWR VPWR _1272_ sky130_fd_sc_hd__and2_1
X_2902_ disp_song.note2\[15\] _2657_ _0314_ VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3882_ _0933_ _1217_ VGND VGND VPWR VPWR _1218_ sky130_fd_sc_hd__and2_1
X_5621_ net96 _2597_ _2600_ VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__o21a_1
X_2833_ _0259_ _0261_ VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__nor2_1
X_5552_ disp_song.note1\[15\] game.padded_notes1\[14\] _2541_ VGND VGND VPWR VPWR
+ _2560_ sky130_fd_sc_hd__mux2_1
X_2764_ _0202_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4503_ game.addmisses.a\[3\] _1701_ VGND VGND VPWR VPWR _1705_ sky130_fd_sc_hd__and2_1
XFILLER_0_111_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5483_ disp_song.note2\[27\] game.padded_notes2\[26\] _2497_ VGND VGND VPWR VPWR
+ _2519_ sky130_fd_sc_hd__mux2_1
X_2695_ _2654_ _2663_ VGND VGND VPWR VPWR _2668_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4434_ _1639_ _1640_ _1644_ _1647_ VGND VGND VPWR VPWR _1648_ sky130_fd_sc_hd__a31o_1
XFILLER_0_111_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4365_ game.scoring_button_2.flash_counter_1\[15\] _1590_ VGND VGND VPWR VPWR _1593_
+ sky130_fd_sc_hd__and2_1
X_6104_ clknet_leaf_25_clk disp_song.um.drum.next_note1\[16\] net65 VGND VGND VPWR
+ VPWR disp_song.note1\[16\] sky130_fd_sc_hd__dfrtp_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3316_ _0674_ _0677_ _0678_ VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__a21oi_2
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6035_ clknet_leaf_57_clk _0144_ net51 VGND VGND VPWR VPWR game.flash_counter\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_4296_ net185 _1542_ _1545_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_2\[16\]
+ sky130_fd_sc_hd__o21a_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3247_ _0471_ _0476_ VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__nand2_1
X_3178_ game.addhits.a\[4\] game.addhits.add2.b\[0\] VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__and2_1
XFILLER_0_95_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5819_ clknet_leaf_50_clk game.scoring_button_2.next_flash_counter_2\[10\] net55
+ VGND VGND VPWR VPWR game.scoring_button_2.flash_counter_2\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_639 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_103_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_105_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4150_ game.counter\[8\] game.counter\[9\] _1429_ VGND VGND VPWR VPWR _1435_ sky130_fd_sc_hd__and3_1
X_3101_ _0462_ _0463_ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__or2b_2
X_4081_ net45 _1358_ _1382_ _1383_ VGND VGND VPWR VPWR _1384_ sky130_fd_sc_hd__or4b_1
X_3032_ _2661_ _0357_ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4983_ _1992_ _1976_ VGND VGND VPWR VPWR _2076_ sky130_fd_sc_hd__or2_1
XFILLER_0_93_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3934_ game.addhits.add2.b\[3\] _1258_ VGND VGND VPWR VPWR _1259_ sky130_fd_sc_hd__nor2_1
X_3865_ _1206_ VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_1
X_2816_ game.counter\[16\] game.counter\[21\] game.counter\[22\] VGND VGND VPWR VPWR
+ _0247_ sky130_fd_sc_hd__a21oi_1
X_5604_ game.out\[0\] _2460_ _2462_ net119 VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3796_ _0949_ _1140_ _1148_ _0966_ _1076_ VGND VGND VPWR VPWR _1149_ sky130_fd_sc_hd__a221o_1
X_5535_ _2548_ net214 _2515_ VGND VGND VPWR VPWR _2549_ sky130_fd_sc_hd__mux2_1
X_2747_ _2654_ _0189_ VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__and2_1
X_5466_ _2507_ VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4417_ net208 _1613_ _1634_ _1612_ VGND VGND VPWR VPWR game.scoring_button_1.next_num_hits\[2\]
+ sky130_fd_sc_hd__a22o_1
X_5397_ _2459_ VGND VGND VPWR VPWR _2460_ sky130_fd_sc_hd__buf_4
XFILLER_0_1_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4348_ _1581_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_1\[9\]
+ sky130_fd_sc_hd__clkbuf_1
X_4279_ _1532_ game.missed_2 _1533_ VGND VGND VPWR VPWR _1534_ sky130_fd_sc_hd__and3b_1
X_6018_ clknet_leaf_5_clk _0127_ net60 VGND VGND VPWR VPWR game.out\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_103_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_99_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3650_ _1004_ _1005_ _1006_ _0921_ VGND VGND VPWR VPWR _1007_ sky130_fd_sc_hd__a31o_1
XFILLER_0_43_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3581_ highest_score.highest_score\[5\] highest_score.highest_score\[4\] _0900_ VGND
+ VGND VPWR VPWR _0943_ sky130_fd_sc_hd__a21oi_1
X_5320_ disp_song.um.drum.next_note1\[5\] _2312_ _2360_ _2211_ _2195_ VGND VGND VPWR
+ VPWR _2402_ sky130_fd_sc_hd__a221o_1
XFILLER_0_23_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5251_ _2208_ _2244_ VGND VGND VPWR VPWR _2336_ sky130_fd_sc_hd__nand2_1
X_4202_ _1472_ VGND VGND VPWR VPWR game.scoring_button_2.next_count\[20\] sky130_fd_sc_hd__clkbuf_1
X_5182_ _0175_ disp_song.um.drum.next_note1\[23\] _2191_ _2268_ disp_song.um.drum.next_note1\[22\]
+ VGND VGND VPWR VPWR _2269_ sky130_fd_sc_hd__a32o_1
X_4133_ game.counter\[5\] game.counter\[4\] _1418_ VGND VGND VPWR VPWR _1423_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4064_ game.addmisses.add3.b\[2\] game.addmisses.add3.b\[1\] _1355_ VGND VGND VPWR
+ VPWR _1369_ sky130_fd_sc_hd__and3_1
X_3015_ disp_song.um.idx_note1\[2\] _0180_ _0394_ _0397_ net183 VGND VGND VPWR VPWR
+ disp_song.um.drum.next_note1\[12\] sky130_fd_sc_hd__a32o_1
XFILLER_0_78_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_93_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4966_ _1956_ disp_song.um.drum.next_note2\[15\] _1965_ _2016_ disp_song.um.drum.next_note2\[14\]
+ VGND VGND VPWR VPWR _2060_ sky130_fd_sc_hd__a32o_1
XFILLER_0_19_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4897_ disp_song.um.drum.next_idx2\[2\] _1949_ VGND VGND VPWR VPWR _1992_ sky130_fd_sc_hd__nor2_4
X_3917_ _1243_ _1241_ VGND VGND VPWR VPWR _1246_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3848_ _0966_ disp_song.display_note1\[0\] _0211_ game.out\[7\] _0208_ VGND VGND
+ VPWR VPWR _1195_ sky130_fd_sc_hd__a221o_2
X_3779_ _0633_ _0653_ _1131_ VGND VGND VPWR VPWR _1132_ sky130_fd_sc_hd__o21a_1
X_5518_ disp_song.note1\[4\] game.padded_notes1\[3\] _2497_ VGND VGND VPWR VPWR _2537_
+ sky130_fd_sc_hd__mux2_1
X_5449_ _2495_ net261 _2473_ VGND VGND VPWR VPWR _2496_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4820_ _0232_ _0254_ _1426_ VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__o21a_1
X_4751_ game.scoring_button_1.flash_counter_1\[3\] _1884_ VGND VGND VPWR VPWR _1887_
+ sky130_fd_sc_hd__and2_1
X_4682_ net177 _1836_ _1839_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_2\[4\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_28_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3702_ _1053_ _1052_ _1057_ highest_score.highest_score\[3\] VGND VGND VPWR VPWR
+ _1058_ sky130_fd_sc_hd__a31o_1
XFILLER_0_43_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3633_ _0835_ _0990_ _0848_ VGND VGND VPWR VPWR _0991_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_70_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3564_ disp_song.mi6.in\[2\] _0926_ disp_song.mi6.in\[3\] VGND VGND VPWR VPWR _0927_
+ sky130_fd_sc_hd__o21a_1
X_3495_ _0830_ _0834_ _0821_ _0828_ VGND VGND VPWR VPWR _0858_ sky130_fd_sc_hd__o2bb2a_1
X_5303_ _2255_ _2385_ _2274_ VGND VGND VPWR VPWR _2386_ sky130_fd_sc_hd__mux2_1
X_5234_ _2227_ _2228_ _2185_ VGND VGND VPWR VPWR _2320_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5165_ _0175_ _2185_ VGND VGND VPWR VPWR _2252_ sky130_fd_sc_hd__nor2_4
X_4116_ game.counter\[0\] game.scoring_button_2.check_hit.in VGND VGND VPWR VPWR _1414_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5096_ _2173_ _2175_ _0214_ _2184_ VGND VGND VPWR VPWR disp_song.um.drum.next_d2\[6\]
+ sky130_fd_sc_hd__o211a_1
X_4047_ game.addmisses.add3.b\[0\] _1335_ VGND VGND VPWR VPWR _1354_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5998_ clknet_leaf_38_clk _0107_ net66 VGND VGND VPWR VPWR game.padded_notes1\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_4949_ _1992_ _2042_ VGND VGND VPWR VPWR _2043_ sky130_fd_sc_hd__nand2_4
XFILLER_0_93_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_520 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_575 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_97_597 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_92_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3280_ _0633_ _0641_ _0642_ VGND VGND VPWR VPWR _0643_ sky130_fd_sc_hd__or3b_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5921_ clknet_leaf_8_clk game.scoring_button_1.next_count\[12\] net60 VGND VGND VPWR
+ VPWR game.scoring_button_1.counts\[12\] sky130_fd_sc_hd__dfrtp_1
X_5852_ clknet_leaf_4_clk game.scoring_button_1.next_num_hits\[1\] net49 VGND VGND
+ VPWR VPWR game.addhits.a\[1\] sky130_fd_sc_hd__dfrtp_4
X_5783_ clknet_leaf_11_clk game.scoring_button_2.next_count\[20\] net57 VGND VGND
+ VPWR VPWR game.scoring_button_2.counts\[20\] sky130_fd_sc_hd__dfrtp_1
X_4803_ _1922_ _1799_ _1923_ VGND VGND VPWR VPWR _1924_ sky130_fd_sc_hd__and3b_1
X_4734_ game.scoring_button_1.flash_counter_2\[19\] game.scoring_button_1.flash_counter_2\[18\]
+ _1868_ game.scoring_button_1.flash_counter_2\[20\] VGND VGND VPWR VPWR _1876_ sky130_fd_sc_hd__a31o_1
XFILLER_0_90_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2995_ _0380_ _0381_ _0383_ net262 VGND VGND VPWR VPWR disp_song.um.drum.next_note1\[6\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_569 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4665_ _1825_ _1826_ _1827_ _1828_ VGND VGND VPWR VPWR _1829_ sky130_fd_sc_hd__or4b_1
XFILLER_0_43_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4596_ _1782_ _1785_ _1699_ VGND VGND VPWR VPWR _1786_ sky130_fd_sc_hd__mux2_1
X_3616_ _0907_ _0975_ _0258_ VGND VGND VPWR VPWR _0976_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3547_ _0667_ _0633_ _0650_ _0615_ VGND VGND VPWR VPWR _0910_ sky130_fd_sc_hd__a31o_1
X_3478_ _0830_ _0834_ VGND VGND VPWR VPWR _0841_ sky130_fd_sc_hd__nand2_1
X_5217_ _2256_ _2303_ VGND VGND VPWR VPWR _2304_ sky130_fd_sc_hd__nor2_1
X_5148_ disp_song.um.drum.next_note1\[24\] disp_song.um.drum.next_note1\[25\] disp_song.um.drum.next_idx1\[0\]
+ VGND VGND VPWR VPWR _2236_ sky130_fd_sc_hd__mux2_1
X_5079_ _2157_ _2168_ _2155_ VGND VGND VPWR VPWR _2169_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_106_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2780_ _0216_ VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_5_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_108_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4450_ _1612_ _1657_ _1659_ _1613_ net196 VGND VGND VPWR VPWR game.scoring_button_1.next_num_hits\[10\]
+ sky130_fd_sc_hd__a32o_1
XFILLER_0_41_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3401_ _0758_ _0761_ _0759_ VGND VGND VPWR VPWR _0764_ sky130_fd_sc_hd__o21ai_4
X_4381_ game.scoring_button_2.flash_counter_1\[19\] game.scoring_button_2.flash_counter_1\[20\]
+ _1600_ VGND VGND VPWR VPWR _1604_ sky130_fd_sc_hd__and3_1
XFILLER_0_111_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6120_ clknet_leaf_23_clk disp_song.um.drum.next_note2\[0\] net64 VGND VGND VPWR
+ VPWR disp_song.note2\[0\] sky130_fd_sc_hd__dfrtp_1
X_3332_ _0606_ _0693_ _0694_ VGND VGND VPWR VPWR _0695_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6051_ clknet_leaf_14_clk _0029_ net58 VGND VGND VPWR VPWR game.counter\[7\] sky130_fd_sc_hd__dfrtp_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3263_ _0461_ _0467_ VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__or2_1
X_5002_ _2093_ _2094_ _0169_ VGND VGND VPWR VPWR _2095_ sky130_fd_sc_hd__mux2_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3194_ _0548_ _0549_ _0550_ VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__o21a_1
Xclkbuf_3_5__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_5__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_72_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5904_ clknet_leaf_44_clk net136 net54 VGND VGND VPWR VPWR game.out\[12\] sky130_fd_sc_hd__dfrtp_1
X_5835_ clknet_leaf_0_clk game.scoring_button_1.next_num_misses\[0\] net49 VGND VGND
+ VPWR VPWR game.addmisses.a\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_76_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5766_ clknet_leaf_16_clk game.scoring_button_2.next_count\[3\] net62 VGND VGND VPWR
+ VPWR game.scoring_button_2.counts\[3\] sky130_fd_sc_hd__dfrtp_1
X_2978_ disp_song.um.idx_note1\[0\] _0178_ _0179_ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__nand3_2
X_4717_ game.scoring_button_1.flash_counter_2\[15\] _1861_ VGND VGND VPWR VPWR _1864_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_71_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5697_ clknet_leaf_0_clk _0033_ net48 VGND VGND VPWR VPWR game.scoring_button_2.acc\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_4648_ _1817_ VGND VGND VPWR VPWR game.scoring_button_1.next_count\[17\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_648 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_497 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4579_ _1675_ _1765_ _1766_ _1770_ VGND VGND VPWR VPWR game.scoring_button_1.next_num_misses\[12\]
+ sky130_fd_sc_hd__o31ai_1
XFILLER_0_97_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_94_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold90 disp_song.note1\[20\] VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3950_ game.addhits.add3.b\[2\] _1267_ VGND VGND VPWR VPWR _1271_ sky130_fd_sc_hd__or2_1
X_2901_ _0313_ _0298_ VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__nor2_1
XFILLER_0_58_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3881_ _0966_ disp_song.display_note2\[4\] _0210_ game.out\[4\] _0208_ VGND VGND
+ VPWR VPWR _1217_ sky130_fd_sc_hd__a221o_1
X_5620_ _0868_ _2595_ VGND VGND VPWR VPWR _2600_ sky130_fd_sc_hd__nand2_1
X_2832_ _0260_ VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__buf_2
X_5551_ _2559_ VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2763_ lvls.level\[2\] lvls.level\[1\] _0200_ VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4502_ _1698_ _1703_ VGND VGND VPWR VPWR _1704_ sky130_fd_sc_hd__nor2_1
XFILLER_0_53_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2694_ _2667_ VGND VGND VPWR VPWR disp_song.um.drum.next_idx2\[1\] sky130_fd_sc_hd__clkbuf_8
X_5482_ _2518_ VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4433_ _1612_ _1646_ VGND VGND VPWR VPWR _1647_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4364_ _1592_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_1\[14\]
+ sky130_fd_sc_hd__clkbuf_1
X_6103_ clknet_leaf_38_clk disp_song.um.drum.next_note1\[15\] net67 VGND VGND VPWR
+ VPWR disp_song.note1\[15\] sky130_fd_sc_hd__dfstp_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3315_ _0675_ _0676_ VGND VGND VPWR VPWR _0678_ sky130_fd_sc_hd__and2_1
X_4295_ game.scoring_button_2.flash_counter_2\[16\] _1542_ _1486_ VGND VGND VPWR VPWR
+ _1545_ sky130_fd_sc_hd__a21boi_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6034_ clknet_leaf_56_clk _0143_ net51 VGND VGND VPWR VPWR game.flash_counter\[14\]
+ sky130_fd_sc_hd__dfrtp_2
X_3246_ _0471_ _0484_ VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__xnor2_2
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3177_ _0538_ _0539_ VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__nand2_2
XTAP_1519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5818_ clknet_leaf_50_clk game.scoring_button_2.next_flash_counter_2\[9\] net55 VGND
+ VGND VPWR VPWR game.scoring_button_2.flash_counter_2\[9\] sky130_fd_sc_hd__dfrtp_1
X_5749_ clknet_leaf_3_clk game.scoring_button_2.next_num_hits\[5\] net49 VGND VGND
+ VPWR VPWR game.addhits.add2.b\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_99_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_353 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3100_ game.addmisses.a\[3\] game.addmisses.add1.b\[3\] VGND VGND VPWR VPWR _0463_
+ sky130_fd_sc_hd__nand2_1
X_4080_ game.addmisses.add4.b\[0\] _1381_ VGND VGND VPWR VPWR _1383_ sky130_fd_sc_hd__nand2_1
X_3031_ _0269_ _0407_ _0408_ disp_song.note1\[17\] VGND VGND VPWR VPWR disp_song.um.drum.next_note1\[17\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4982_ _1973_ VGND VGND VPWR VPWR _2075_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3933_ _1256_ _1257_ _1252_ VGND VGND VPWR VPWR _1258_ sky130_fd_sc_hd__or3_1
XFILLER_0_46_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3864_ _0933_ _1205_ VGND VGND VPWR VPWR _1206_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2815_ game.counter\[16\] _0245_ game.counter\[22\] VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__o21a_1
X_5603_ game.padded_notes1\[31\] _2460_ _2462_ net138 VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3795_ _1143_ _1144_ _1147_ VGND VGND VPWR VPWR _1148_ sky130_fd_sc_hd__o21ai_1
X_5534_ disp_song.note1\[9\] game.padded_notes1\[8\] _2541_ VGND VGND VPWR VPWR _2548_
+ sky130_fd_sc_hd__mux2_1
X_2746_ disp_song.um.idx_note1\[2\] _0170_ _0188_ VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_5_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5465_ _2506_ game.padded_notes2\[21\] _2473_ VGND VGND VPWR VPWR _2507_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4416_ _1632_ _1633_ VGND VGND VPWR VPWR _1634_ sky130_fd_sc_hd__nand2_1
X_5396_ game.beat_clk _0209_ VGND VGND VPWR VPWR _2459_ sky130_fd_sc_hd__and2_1
X_4347_ _1579_ _1413_ _1580_ VGND VGND VPWR VPWR _1581_ sky130_fd_sc_hd__and3b_1
X_4278_ game.scoring_button_2.flash_counter_2\[9\] game.scoring_button_2.flash_counter_2\[10\]
+ _1525_ game.scoring_button_2.flash_counter_2\[11\] VGND VGND VPWR VPWR _1533_ sky130_fd_sc_hd__a31o_1
XFILLER_0_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6017_ clknet_leaf_5_clk net116 net60 VGND VGND VPWR VPWR game.out\[4\] sky130_fd_sc_hd__dfrtp_1
X_3229_ _0586_ _0589_ _0587_ VGND VGND VPWR VPWR _0592_ sky130_fd_sc_hd__o21ai_2
XTAP_1305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_629 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_615 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3580_ _0890_ _0940_ _0941_ VGND VGND VPWR VPWR _0942_ sky130_fd_sc_hd__o21a_1
X_5250_ _2288_ VGND VGND VPWR VPWR _2335_ sky130_fd_sc_hd__inv_2
X_4201_ game.scoring_button_2.check_hit.in _1471_ VGND VGND VPWR VPWR _1472_ sky130_fd_sc_hd__and2_1
X_5181_ _0175_ _2230_ VGND VGND VPWR VPWR _2268_ sky130_fd_sc_hd__nor2_1
X_4132_ _1422_ VGND VGND VPWR VPWR game.scoring_button_2.next_count\[4\] sky130_fd_sc_hd__clkbuf_1
X_4063_ _1289_ _1364_ _1365_ _1368_ VGND VGND VPWR VPWR game.scoring_button_2.next_num_misses\[9\]
+ sky130_fd_sc_hd__o31a_1
X_3014_ _0374_ _0392_ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__or2b_1
XFILLER_0_78_437 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4965_ _1956_ disp_song.um.drum.next_note2\[12\] _1968_ _2058_ VGND VGND VPWR VPWR
+ _2059_ sky130_fd_sc_hd__o211a_1
XFILLER_0_74_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3916_ game.addhits.add1.b\[1\] _1227_ _1245_ _1226_ VGND VGND VPWR VPWR game.scoring_button_2.next_num_hits\[1\]
+ sky130_fd_sc_hd__a22o_1
X_4896_ disp_song.um.drum.next_note2\[14\] disp_song.um.drum.next_note2\[15\] _2670_
+ VGND VGND VPWR VPWR _1991_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_654 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_142 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3847_ _1193_ _1194_ _0933_ VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__o21a_1
XFILLER_0_14_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3778_ _0633_ _0630_ _0912_ VGND VGND VPWR VPWR _1131_ sky130_fd_sc_hd__a21oi_1
X_5517_ _2536_ VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__clkbuf_1
X_2729_ _2654_ _0173_ VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_595 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5448_ disp_song.note2\[16\] game.padded_notes2\[15\] _0219_ VGND VGND VPWR VPWR
+ _2495_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5379_ net179 net123 _2448_ VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__o21a_1
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_64_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_103_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_632 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4750_ _1886_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_1\[2\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4681_ net177 _1836_ game.missed_1 VGND VGND VPWR VPWR _1839_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_71_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3701_ highest_score.highest_score\[0\] VGND VGND VPWR VPWR _1057_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3632_ _0840_ _0855_ VGND VGND VPWR VPWR _0990_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3563_ disp_song.mi6.in\[1\] VGND VGND VPWR VPWR _0926_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5302_ _2254_ _2349_ _2384_ _2310_ VGND VGND VPWR VPWR _2385_ sky130_fd_sc_hd__o22a_1
XFILLER_0_59_86 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3494_ _0830_ _0834_ VGND VGND VPWR VPWR _0857_ sky130_fd_sc_hd__and2_1
X_5233_ disp_song.um.drum.next_idx1\[2\] _2318_ disp_song.um.drum.next_idx1\[4\] VGND
+ VGND VPWR VPWR _2319_ sky130_fd_sc_hd__o21a_1
X_5164_ _0175_ disp_song.um.drum.next_note1\[30\] _2195_ _2250_ VGND VGND VPWR VPWR
+ _2251_ sky130_fd_sc_hd__o211a_1
X_4115_ _0219_ _1405_ _2658_ _1413_ VGND VGND VPWR VPWR game.scoring_button_2.next_good
+ sky130_fd_sc_hd__a31o_1
X_5095_ _2677_ _2179_ _2183_ _1950_ VGND VGND VPWR VPWR _2184_ sky130_fd_sc_hd__a211o_1
X_4046_ _1349_ _1350_ _1353_ _1289_ VGND VGND VPWR VPWR game.scoring_button_2.next_num_misses\[7\]
+ sky130_fd_sc_hd__a22o_1
XPHY_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_78_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5997_ clknet_leaf_38_clk _0106_ net66 VGND VGND VPWR VPWR game.padded_notes1\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4948_ _2667_ _2669_ VGND VGND VPWR VPWR _2042_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4879_ disp_song.um.drum.next_idx2\[1\] _1968_ _1973_ VGND VGND VPWR VPWR _1974_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_61_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_621 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_111_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_635 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5920_ clknet_leaf_9_clk game.scoring_button_1.next_count\[11\] net60 VGND VGND VPWR
+ VPWR game.scoring_button_1.counts\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5851_ clknet_leaf_4_clk game.scoring_button_1.next_num_hits\[0\] net49 VGND VGND
+ VPWR VPWR game.addhits.a\[0\] sky130_fd_sc_hd__dfrtp_4
X_2994_ _0382_ _0381_ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__nand2_1
X_5782_ clknet_leaf_11_clk game.scoring_button_2.next_count\[19\] net57 VGND VGND
+ VPWR VPWR game.scoring_button_2.counts\[19\] sky130_fd_sc_hd__dfrtp_1
X_4802_ game.scoring_button_1.flash_counter_1\[18\] _1919_ VGND VGND VPWR VPWR _1923_
+ sky130_fd_sc_hd__or2_1
X_4733_ game.scoring_button_1.flash_counter_2\[19\] game.scoring_button_1.flash_counter_2\[20\]
+ _1871_ VGND VGND VPWR VPWR _1875_ sky130_fd_sc_hd__and3_1
XFILLER_0_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4664_ game.scoring_button_1.flash_counter_2\[17\] game.scoring_button_1.flash_counter_2\[16\]
+ game.scoring_button_1.flash_counter_2\[19\] game.scoring_button_1.flash_counter_2\[18\]
+ VGND VGND VPWR VPWR _1828_ sky130_fd_sc_hd__and4_1
X_4595_ game.addmisses.a\[15\] _1783_ _1784_ VGND VGND VPWR VPWR _1785_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3615_ highest_score.highest_score\[4\] _0902_ VGND VGND VPWR VPWR _0975_ sky130_fd_sc_hd__or2_1
XFILLER_0_101_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3546_ _0612_ _0482_ _0611_ _0613_ VGND VGND VPWR VPWR _0909_ sky130_fd_sc_hd__a31o_2
X_3477_ _0838_ _0839_ _0830_ _0834_ VGND VGND VPWR VPWR _0840_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_50_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5216_ disp_song.note1\[2\] _2232_ _2302_ VGND VGND VPWR VPWR _2303_ sky130_fd_sc_hd__o21ai_1
X_5147_ _0173_ _2231_ _2233_ _2234_ _2185_ VGND VGND VPWR VPWR _2235_ sky130_fd_sc_hd__o221a_1
XFILLER_0_98_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5078_ _2057_ _2061_ _2013_ VGND VGND VPWR VPWR _2168_ sky130_fd_sc_hd__mux2_1
X_4029_ game.addmisses.add2.b\[1\] _1331_ VGND VGND VPWR VPWR _1339_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_109_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_100_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_97_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_284 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4380_ net171 _1600_ _1603_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_1\[19\]
+ sky130_fd_sc_hd__o21a_1
X_3400_ _0762_ _0752_ VGND VGND VPWR VPWR _0763_ sky130_fd_sc_hd__nand2_2
XFILLER_0_0_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3331_ _0605_ _0597_ _0601_ VGND VGND VPWR VPWR _0694_ sky130_fd_sc_hd__or3_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6050_ clknet_leaf_14_clk _0028_ net58 VGND VGND VPWR VPWR game.counter\[6\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_0_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3262_ _0624_ VGND VGND VPWR VPWR _0625_ sky130_fd_sc_hd__inv_2
X_5001_ _2003_ _2004_ _2666_ VGND VGND VPWR VPWR _2094_ sky130_fd_sc_hd__mux2_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3193_ _0554_ _0555_ VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__or2b_1
X_5903_ clknet_leaf_44_clk net118 net53 VGND VGND VPWR VPWR game.out\[11\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5834_ clknet_leaf_11_clk net90 net57 VGND VGND VPWR VPWR game.scoring_button_2.check_hit.edge_1
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5765_ clknet_leaf_16_clk game.scoring_button_2.next_count\[2\] net62 VGND VGND VPWR
+ VPWR game.scoring_button_2.counts\[2\] sky130_fd_sc_hd__dfrtp_1
X_2977_ _0364_ _0367_ _0369_ VGND VGND VPWR VPWR disp_song.um.drum.next_note1\[2\]
+ sky130_fd_sc_hd__o21ai_2
XFILLER_0_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4716_ _1863_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_2\[14\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5696_ _2653_ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4647_ _1791_ _0017_ VGND VGND VPWR VPWR _1817_ sky130_fd_sc_hd__and2_1
XFILLER_0_102_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4578_ _1699_ _1744_ _1768_ _1769_ VGND VGND VPWR VPWR _1770_ sky130_fd_sc_hd__or4b_1
X_3529_ _0675_ _0889_ _0891_ VGND VGND VPWR VPWR _0892_ sky130_fd_sc_hd__a21o_1
XFILLER_0_110_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold91 modetrans.mode\[4\] VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__dlygate4sd3_1
Xhold80 game.addhits.add2.b\[3\] VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2900_ disp_song.um.idx_note2\[1\] disp_song.um.idx_note2\[0\] disp_song.um.idx_note2\[2\]
+ VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__nand3_1
XFILLER_0_97_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3880_ _1216_ VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_70_clk clknet_3_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_70_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_45_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2831_ _0255_ _0258_ VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__and2_1
X_5550_ _2558_ game.padded_notes1\[14\] _2472_ VGND VGND VPWR VPWR _2559_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2762_ _0201_ VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__clkbuf_1
X_5481_ _2517_ net239 _2515_ VGND VGND VPWR VPWR _2518_ sky130_fd_sc_hd__mux2_1
X_4501_ _1701_ _1702_ VGND VGND VPWR VPWR _1703_ sky130_fd_sc_hd__or2_1
X_2693_ _2666_ VGND VGND VPWR VPWR _2667_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4432_ game.addhits.a\[5\] game.addhits.a\[4\] _1630_ game.addhits.a\[6\] VGND VGND
+ VPWR VPWR _1646_ sky130_fd_sc_hd__a31o_1
XFILLER_0_111_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4363_ _1590_ _1413_ _1591_ VGND VGND VPWR VPWR _1592_ sky130_fd_sc_hd__and3b_1
X_6102_ clknet_leaf_37_clk disp_song.um.drum.next_note1\[14\] net67 VGND VGND VPWR
+ VPWR disp_song.note1\[14\] sky130_fd_sc_hd__dfstp_1
XFILLER_0_67_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3314_ _0675_ _0676_ VGND VGND VPWR VPWR _0677_ sky130_fd_sc_hd__or2_1
X_4294_ _1544_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_2\[15\]
+ sky130_fd_sc_hd__clkbuf_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6033_ clknet_leaf_60_clk _0142_ net51 VGND VGND VPWR VPWR game.flash_counter\[13\]
+ sky130_fd_sc_hd__dfrtp_2
X_3245_ _0569_ _0575_ _0607_ _0568_ VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__a22o_2
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3176_ game.addhits.a\[5\] game.addhits.add2.b\[1\] VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_107_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_61_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_61_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_49_579 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_91_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5817_ clknet_leaf_50_clk game.scoring_button_2.next_flash_counter_2\[8\] net55 VGND
+ VGND VPWR VPWR game.scoring_button_2.flash_counter_2\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5748_ clknet_leaf_3_clk game.scoring_button_2.next_num_hits\[4\] net49 VGND VGND
+ VPWR VPWR game.addhits.add2.b\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_106_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5679_ _2614_ _2641_ _2642_ VGND VGND VPWR VPWR _2643_ sky130_fd_sc_hd__and3_1
XFILLER_0_102_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_192 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_52_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_52_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_103_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3030_ _2660_ _0407_ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_619 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4981_ _1955_ _1958_ _2666_ VGND VGND VPWR VPWR _2074_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_43_clk clknet_3_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_43_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_58_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3932_ game.addhits.add2.b\[1\] VGND VGND VPWR VPWR _1257_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3863_ _0966_ disp_song.display_note1\[5\] _0211_ game.out\[12\] _0208_ VGND VGND
+ VPWR VPWR _1205_ sky130_fd_sc_hd__a221o_1
X_2814_ lvls.level\[0\] _0242_ VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__nor2_1
X_5602_ _2593_ VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5533_ _2547_ VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__clkbuf_1
X_3794_ disp_song.mi6.in\[2\] _1145_ _1146_ _1077_ _0925_ VGND VGND VPWR VPWR _1147_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2745_ _0186_ _0187_ _0170_ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__a21oi_1
X_5464_ disp_song.note2\[21\] game.padded_notes2\[20\] _2497_ VGND VGND VPWR VPWR
+ _2506_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5395_ _0209_ modetrans.mode\[5\] VGND VGND VPWR VPWR _2458_ sky130_fd_sc_hd__and2b_1
X_4415_ _1623_ _1630_ _1626_ VGND VGND VPWR VPWR _1633_ sky130_fd_sc_hd__a21o_1
X_4346_ game.scoring_button_2.flash_counter_1\[9\] _1576_ VGND VGND VPWR VPWR _1580_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_111_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4277_ game.scoring_button_2.flash_counter_2\[11\] game.scoring_button_2.flash_counter_2\[10\]
+ _1528_ VGND VGND VPWR VPWR _1532_ sky130_fd_sc_hd__and3_1
X_6016_ clknet_leaf_5_clk net102 net59 VGND VGND VPWR VPWR game.out\[3\] sky130_fd_sc_hd__dfrtp_1
X_3228_ _0585_ _0590_ VGND VGND VPWR VPWR _0591_ sky130_fd_sc_hd__nor2_2
X_3159_ _0521_ _0516_ _0517_ VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_96_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_34_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_34_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_91_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_25_clk clknet_3_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_25_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_28_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_644 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4200_ _1469_ _1470_ VGND VGND VPWR VPWR _1471_ sky130_fd_sc_hd__nor2_1
X_5180_ _2230_ _2266_ disp_song.note1\[20\] disp_song.um.drum.next_idx1\[0\] VGND
+ VGND VPWR VPWR _2267_ sky130_fd_sc_hd__a2bb2o_1
X_4131_ _1405_ _0026_ VGND VGND VPWR VPWR _1422_ sky130_fd_sc_hd__and2_1
X_4062_ game.addmisses.add3.b\[1\] _1330_ _1366_ _1367_ VGND VGND VPWR VPWR _1368_
+ sky130_fd_sc_hd__a31o_1
X_3013_ _0396_ VGND VGND VPWR VPWR disp_song.um.drum.next_note1\[11\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_64_32 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4964_ disp_song.um.drum.next_idx2\[0\] disp_song.um.drum.next_note2\[13\] VGND VGND
+ VPWR VPWR _2058_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_16_clk clknet_3_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_16_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_19_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3915_ _1235_ _1244_ _1237_ VGND VGND VPWR VPWR _1245_ sky130_fd_sc_hd__mux2_1
X_4895_ _1962_ _1989_ VGND VGND VPWR VPWR _1990_ sky130_fd_sc_hd__nor2_1
XFILLER_0_80_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3846_ modetrans.mode\[3\] _0255_ disp_song.toggle_red _0214_ VGND VGND VPWR VPWR
+ _1194_ sky130_fd_sc_hd__a22o_1
XFILLER_0_73_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3777_ _1034_ _1032_ VGND VGND VPWR VPWR _1130_ sky130_fd_sc_hd__and2b_1
X_5516_ _2535_ game.padded_notes1\[3\] _2515_ VGND VGND VPWR VPWR _2536_ sky130_fd_sc_hd__mux2_1
X_2728_ _0171_ _0172_ VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_498 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5447_ _2494_ VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_585 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_100_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5378_ net179 _2447_ VGND VGND VPWR VPWR _2448_ sky130_fd_sc_hd__nand2_1
X_4329_ net176 _1565_ game.hit_2 VGND VGND VPWR VPWR _1568_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_69_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_107_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_571 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_107_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_100_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3700_ _1052_ _1054_ _1055_ VGND VGND VPWR VPWR _1056_ sky130_fd_sc_hd__o21a_1
XFILLER_0_50_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4680_ _1838_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_2\[3\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_625 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3631_ _0953_ _0987_ _0989_ _0935_ VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__o31a_1
XFILLER_0_43_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3562_ disp_song.mi6.in\[4\] VGND VGND VPWR VPWR _0925_ sky130_fd_sc_hd__buf_4
XFILLER_0_3_413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5301_ _2185_ _2231_ disp_song.note1\[26\] _2232_ VGND VGND VPWR VPWR _2384_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_51_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3493_ _0840_ _0850_ _0855_ VGND VGND VPWR VPWR _0856_ sky130_fd_sc_hd__and3_1
XFILLER_0_51_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5232_ _2218_ _2219_ _2185_ VGND VGND VPWR VPWR _2318_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_5_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_5_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_59_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5163_ _0176_ disp_song.um.drum.next_note1\[31\] VGND VGND VPWR VPWR _2250_ sky130_fd_sc_hd__or2_1
X_4114_ _1406_ _1407_ _1412_ game.hit_2 VGND VGND VPWR VPWR _1413_ sky130_fd_sc_hd__o31a_4
X_5094_ _2677_ _2182_ VGND VGND VPWR VPWR _2183_ sky130_fd_sc_hd__nor2_1
X_4045_ _1306_ _1351_ _1352_ _1307_ game.addmisses.add2.b\[3\] VGND VGND VPWR VPWR
+ _1353_ sky130_fd_sc_hd__a32o_1
XFILLER_0_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5996_ clknet_leaf_38_clk _0105_ net66 VGND VGND VPWR VPWR game.padded_notes1\[15\]
+ sky130_fd_sc_hd__dfstp_1
X_4947_ _2037_ _2040_ _2026_ VGND VGND VPWR VPWR _2041_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4878_ disp_song.um.drum.next_note2\[28\] disp_song.um.drum.next_note2\[29\] _2670_
+ VGND VGND VPWR VPWR _1973_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3829_ _1173_ _1179_ _0935_ VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__o21a_1
XFILLER_0_61_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_108_510 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_614 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_103_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5850_ clknet_leaf_68_clk game.scoring_button_1.next_num_misses\[15\] net46 VGND
+ VGND VPWR VPWR game.addmisses.a\[15\] sky130_fd_sc_hd__dfrtp_4
X_2993_ _0359_ _0366_ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__nor2_2
X_5781_ clknet_leaf_11_clk game.scoring_button_2.next_count\[18\] net57 VGND VGND
+ VPWR VPWR game.scoring_button_2.counts\[18\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4801_ game.scoring_button_1.flash_counter_1\[18\] _1919_ VGND VGND VPWR VPWR _1922_
+ sky130_fd_sc_hd__and2_1
X_4732_ net181 _1871_ _1874_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_2\[19\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_28_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4663_ game.scoring_button_1.flash_counter_2\[21\] game.scoring_button_1.flash_counter_2\[20\]
+ game.scoring_button_1.flash_counter_2\[22\] VGND VGND VPWR VPWR _1827_ sky130_fd_sc_hd__or3_1
XFILLER_0_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3614_ _0894_ _0973_ _0896_ VGND VGND VPWR VPWR _0974_ sky130_fd_sc_hd__a21o_1
XFILLER_0_12_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4594_ game.addmisses.a\[14\] _1771_ VGND VGND VPWR VPWR _1784_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3545_ _0902_ _0907_ _0258_ VGND VGND VPWR VPWR _0908_ sky130_fd_sc_hd__a21o_1
X_3476_ _0762_ _0824_ _0825_ _0826_ _0792_ VGND VGND VPWR VPWR _0839_ sky130_fd_sc_hd__o311a_1
X_5215_ _0373_ _2258_ _2232_ VGND VGND VPWR VPWR _2302_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_86_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5146_ _0185_ _0197_ _2187_ VGND VGND VPWR VPWR _2234_ sky130_fd_sc_hd__and3_1
X_5077_ _2013_ _2166_ VGND VGND VPWR VPWR _2167_ sky130_fd_sc_hd__nor2_1
X_4028_ _1335_ _1337_ VGND VGND VPWR VPWR _1338_ sky130_fd_sc_hd__xor2_1
X_5979_ clknet_leaf_10_clk net81 net61 VGND VGND VPWR VPWR game.scoring_button_1.check_hit.edge_2
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_105_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_97_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_85_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_547 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_105 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_111_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3330_ _0683_ _0691_ _0692_ VGND VGND VPWR VPWR _0693_ sky130_fd_sc_hd__o21ba_2
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ _1999_ _2001_ _2667_ VGND VGND VPWR VPWR _2093_ sky130_fd_sc_hd__mux2_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3261_ _0553_ _0623_ _0558_ VGND VGND VPWR VPWR _0624_ sky130_fd_sc_hd__mux2_1
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3192_ game.addhits.a\[3\] game.addhits.add1.b\[3\] VGND VGND VPWR VPWR _0555_ sky130_fd_sc_hd__nand2_1
XFILLER_0_88_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5902_ clknet_leaf_44_clk _0085_ net53 VGND VGND VPWR VPWR game.out\[10\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5833_ clknet_leaf_0_clk net84 net48 VGND VGND VPWR VPWR game.scoring_button_2.check_hit.edge_2
+ sky130_fd_sc_hd__dfrtp_1
X_5764_ clknet_leaf_16_clk game.scoring_button_2.next_count\[1\] net62 VGND VGND VPWR
+ VPWR game.scoring_button_2.counts\[1\] sky130_fd_sc_hd__dfrtp_1
X_2976_ _0368_ _0364_ disp_song.note1\[2\] VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_29_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4715_ _1861_ _1830_ _1862_ VGND VGND VPWR VPWR _1863_ sky130_fd_sc_hd__and3b_1
X_5695_ game.scoring_button_1.acc\[2\] _2529_ VGND VGND VPWR VPWR _2653_ sky130_fd_sc_hd__and2_1
X_4646_ _1816_ VGND VGND VPWR VPWR game.scoring_button_1.next_count\[16\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4577_ net248 _1767_ VGND VGND VPWR VPWR _1769_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_97_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3528_ _0675_ _0890_ VGND VGND VPWR VPWR _0891_ sky130_fd_sc_hd__nor2_1
X_3459_ _0752_ VGND VGND VPWR VPWR _0822_ sky130_fd_sc_hd__inv_2
XFILLER_0_99_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5129_ _2202_ _2214_ _2216_ VGND VGND VPWR VPWR _2217_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_109_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold81 disp_song.note1\[26\] VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 disp_song.note1\[29\] VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__dlygate4sd3_1
Xhold70 game.out\[8\] VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2830_ _0255_ _0258_ VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__nor2_4
XFILLER_0_45_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_455 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2761_ lvls.level\[0\] lvls.level\[2\] _0200_ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__mux2_1
X_5480_ disp_song.note2\[26\] game.padded_notes2\[25\] _2497_ VGND VGND VPWR VPWR
+ _2517_ sky130_fd_sc_hd__mux2_1
X_2692_ _2665_ VGND VGND VPWR VPWR _2666_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_13_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4500_ game.addmisses.a\[1\] game.addmisses.a\[0\] game.addmisses.a\[2\] VGND VGND
+ VPWR VPWR _1702_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_53_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_1 _1201_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_101_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4431_ game.addhits.a\[7\] _1644_ VGND VGND VPWR VPWR _1645_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4362_ game.scoring_button_2.flash_counter_1\[13\] game.scoring_button_2.flash_counter_1\[12\]
+ _1583_ game.scoring_button_2.flash_counter_1\[14\] VGND VGND VPWR VPWR _1591_ sky130_fd_sc_hd__a31o_1
X_6101_ clknet_leaf_37_clk disp_song.um.drum.next_note1\[13\] net71 VGND VGND VPWR
+ VPWR disp_song.note1\[13\] sky130_fd_sc_hd__dfrtp_1
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3313_ _0617_ _0609_ VGND VGND VPWR VPWR _0676_ sky130_fd_sc_hd__nor2_1
X_4293_ _1542_ game.missed_2 _1543_ VGND VGND VPWR VPWR _1544_ sky130_fd_sc_hd__and3b_1
XFILLER_0_67_76 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6032_ clknet_leaf_60_clk _0141_ net51 VGND VGND VPWR VPWR game.flash_counter\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_3244_ _0563_ _0576_ VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__or2b_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3175_ game.addhits.a\[5\] game.addhits.add2.b\[1\] VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__nand2_1
XFILLER_0_107_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5816_ clknet_leaf_49_clk game.scoring_button_2.next_flash_counter_2\[7\] net56 VGND
+ VGND VPWR VPWR game.scoring_button_2.flash_counter_2\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2959_ disp_song.um.idx_note1\[2\] _0179_ disp_song.um.idx_note1\[0\] VGND VGND VPWR
+ VPWR _0353_ sky130_fd_sc_hd__or3b_2
XFILLER_0_17_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5747_ clknet_leaf_3_clk game.scoring_button_2.next_num_hits\[3\] net49 VGND VGND
+ VPWR VPWR game.addhits.add1.b\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5678_ game.flash_counter\[20\] _2640_ VGND VGND VPWR VPWR _2642_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4629_ _1791_ _1432_ VGND VGND VPWR VPWR _1808_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_99_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_99_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_642 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4980_ _2011_ _2051_ _2073_ _0352_ VGND VGND VPWR VPWR disp_song.um.drum.next_d2\[1\]
+ sky130_fd_sc_hd__a211oi_1
XFILLER_0_58_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3931_ game.addhits.add2.b\[2\] VGND VGND VPWR VPWR _1256_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3862_ _1204_ VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_1
X_2813_ _0240_ _0241_ _0243_ game.counter\[21\] VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__a22o_1
X_5601_ _2592_ game.padded_notes1\[31\] _2472_ VGND VGND VPWR VPWR _2593_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5532_ _2546_ net224 _2515_ VGND VGND VPWR VPWR _2547_ sky130_fd_sc_hd__mux2_1
X_3793_ disp_song.mi6.in\[2\] _0926_ _1082_ VGND VGND VPWR VPWR _1146_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_5_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2744_ _0178_ _0180_ VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5463_ _2505_ VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_78_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4414_ _1629_ _1627_ VGND VGND VPWR VPWR _1632_ sky130_fd_sc_hd__or2_1
X_5394_ game.scoring_button_2.check_hit.edge_1 _1287_ net131 _2411_ VGND VGND VPWR
+ VPWR _0049_ sky130_fd_sc_hd__o22a_1
XFILLER_0_111_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4345_ game.scoring_button_2.flash_counter_1\[9\] _1576_ VGND VGND VPWR VPWR _1579_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_94_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4276_ net166 _1528_ _1531_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_2\[10\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_94_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6015_ clknet_leaf_6_clk _0124_ net59 VGND VGND VPWR VPWR game.out\[2\] sky130_fd_sc_hd__dfrtp_1
X_3227_ _0588_ _0589_ VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__xnor2_1
X_3158_ game.addmisses.a\[15\] game.addmisses.add4.b\[3\] VGND VGND VPWR VPWR _0521_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_96_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3089_ game.addmisses.a\[1\] game.addmisses.add1.b\[1\] VGND VGND VPWR VPWR _0452_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_92_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_103_611 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_586 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_102_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_656 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_594 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4130_ net168 _1418_ VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__xor2_1
X_4061_ game.addmisses.add3.b\[1\] _1366_ _1289_ VGND VGND VPWR VPWR _1367_ sky130_fd_sc_hd__o21ai_1
X_3012_ disp_song.um.idx_note1\[0\] _0178_ _0179_ _0394_ _0395_ VGND VGND VPWR VPWR
+ _0396_ sky130_fd_sc_hd__a41o_1
XFILLER_0_64_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_55 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4963_ _2056_ VGND VGND VPWR VPWR _2057_ sky130_fd_sc_hd__inv_2
XFILLER_0_80_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3914_ _1235_ _1242_ _1243_ VGND VGND VPWR VPWR _1244_ sky130_fd_sc_hd__o21ai_2
X_4894_ _1986_ _1988_ disp_song.um.drum.next_idx2\[1\] VGND VGND VPWR VPWR _1989_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3845_ game.missed_1 game.missed_2 _0211_ VGND VGND VPWR VPWR _1193_ sky130_fd_sc_hd__o21a_1
XFILLER_0_13_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_104_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3776_ _1119_ _1128_ _1129_ _0935_ VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__o31a_2
X_5515_ disp_song.note1\[3\] game.padded_notes1\[2\] _2497_ VGND VGND VPWR VPWR _2535_
+ sky130_fd_sc_hd__mux2_1
X_2727_ disp_song.um.idx_note1\[0\] _0170_ VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5446_ _2493_ game.padded_notes2\[15\] _2473_ VGND VGND VPWR VPWR _2494_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5377_ game.beat_clk _0206_ VGND VGND VPWR VPWR _2447_ sky130_fd_sc_hd__or2b_1
X_4328_ _1567_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_1\[3\]
+ sky130_fd_sc_hd__clkbuf_1
X_4259_ _1518_ game.missed_2 _1519_ VGND VGND VPWR VPWR _1520_ sky130_fd_sc_hd__and3b_1
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_130 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_623 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_100_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3630_ _0214_ _0988_ _0986_ _0211_ VGND VGND VPWR VPWR _0989_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3561_ _0849_ _0856_ _0861_ net39 _0923_ VGND VGND VPWR VPWR _0924_ sky130_fd_sc_hd__o311a_1
XFILLER_0_36_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5300_ _2270_ _2382_ _2274_ VGND VGND VPWR VPWR _2383_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3492_ _0830_ _0834_ net40 _0854_ VGND VGND VPWR VPWR _0855_ sky130_fd_sc_hd__o2bb2a_2
X_5231_ _2236_ _2316_ disp_song.um.drum.next_idx1\[1\] VGND VGND VPWR VPWR _2317_
+ sky130_fd_sc_hd__mux2_1
X_5162_ _0175_ disp_song.um.drum.next_note1\[28\] _2191_ _2248_ VGND VGND VPWR VPWR
+ _2249_ sky130_fd_sc_hd__o211a_1
X_5093_ _2180_ _2181_ _0162_ VGND VGND VPWR VPWR _2182_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4113_ _1408_ _1409_ _1410_ _1411_ VGND VGND VPWR VPWR _1412_ sky130_fd_sc_hd__or4b_1
X_4044_ game.addmisses.add2.b\[3\] _1344_ VGND VGND VPWR VPWR _1352_ sky130_fd_sc_hd__or2_1
XPHY_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5995_ clknet_leaf_37_clk _0104_ net71 VGND VGND VPWR VPWR game.padded_notes1\[14\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_59_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4946_ _2038_ _2039_ disp_song.note2\[20\] disp_song.um.drum.next_idx2\[0\] VGND
+ VGND VPWR VPWR _2040_ sky130_fd_sc_hd__a2bb2o_1
X_4877_ _1959_ _1963_ _1971_ _1961_ VGND VGND VPWR VPWR _1972_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_19_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3828_ _0259_ _1171_ _1178_ _0214_ VGND VGND VPWR VPWR _1179_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_61_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3759_ _1103_ _1113_ _0935_ VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__o21a_1
XFILLER_0_30_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5429_ _2482_ VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_97_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_111_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_103_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_589 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4800_ _1921_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_1\[17\]
+ sky130_fd_sc_hd__clkbuf_1
X_2992_ disp_song.um.idx_note1\[0\] disp_song.um.idx_note1\[2\] _0177_ _0179_ VGND
+ VGND VPWR VPWR _0381_ sky130_fd_sc_hd__and4b_1
X_5780_ clknet_leaf_11_clk game.scoring_button_2.next_count\[17\] net57 VGND VGND
+ VPWR VPWR game.scoring_button_2.counts\[17\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4731_ net181 _1871_ _1830_ VGND VGND VPWR VPWR _1874_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_61_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4662_ game.scoring_button_1.flash_counter_2\[8\] game.scoring_button_1.flash_counter_2\[11\]
+ game.scoring_button_1.flash_counter_2\[10\] game.scoring_button_1.flash_counter_2\[9\]
+ VGND VGND VPWR VPWR _1826_ sky130_fd_sc_hd__or4b_1
XFILLER_0_16_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3613_ _0887_ _0939_ VGND VGND VPWR VPWR _0973_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_659 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4593_ game.addmisses.a\[14\] _1771_ _1774_ VGND VGND VPWR VPWR _1783_ sky130_fd_sc_hd__o21a_1
XFILLER_0_9_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3544_ _0255_ _0904_ _0905_ _0906_ VGND VGND VPWR VPWR _0907_ sky130_fd_sc_hd__and4_1
XFILLER_0_12_578 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3475_ _0775_ _0776_ _0811_ _0837_ VGND VGND VPWR VPWR _0838_ sky130_fd_sc_hd__and4b_1
X_5214_ _2254_ _2300_ _2247_ VGND VGND VPWR VPWR _2301_ sky130_fd_sc_hd__o21ai_1
X_5145_ _2232_ disp_song.um.drum.next_note1\[26\] VGND VGND VPWR VPWR _2233_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5076_ _2119_ _2165_ _2026_ VGND VGND VPWR VPWR _2166_ sky130_fd_sc_hd__mux2_1
X_4027_ _1334_ _1336_ VGND VGND VPWR VPWR _1337_ sky130_fd_sc_hd__nand2_1
X_5978_ clknet_leaf_10_clk game.scoring_button_1.next_start_count net57 VGND VGND
+ VPWR VPWR game.scoring_button_1.check_hit.in sky130_fd_sc_hd__dfrtp_4
XFILLER_0_19_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4929_ _1956_ disp_song.um.drum.next_note2\[26\] VGND VGND VPWR VPWR _2023_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_105_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_100_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_106_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_108_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_607 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3260_ _0553_ _0559_ VGND VGND VPWR VPWR _0623_ sky130_fd_sc_hd__nor2_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3191_ game.addhits.a\[3\] game.addhits.add1.b\[3\] VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5901_ clknet_leaf_44_clk net141 net53 VGND VGND VPWR VPWR game.out\[9\] sky130_fd_sc_hd__dfrtp_1
X_5832_ clknet_leaf_10_clk game.scoring_button_2.next_start_count net57 VGND VGND
+ VPWR VPWR game.scoring_button_2.check_hit.in sky130_fd_sc_hd__dfrtp_4
X_5763_ clknet_leaf_16_clk game.scoring_button_2.next_count\[0\] net62 VGND VGND VPWR
+ VPWR game.scoring_button_2.counts\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4714_ game.scoring_button_1.flash_counter_2\[13\] game.scoring_button_1.flash_counter_2\[12\]
+ _1854_ game.scoring_button_1.flash_counter_2\[14\] VGND VGND VPWR VPWR _1862_ sky130_fd_sc_hd__a31o_1
XFILLER_0_84_570 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2975_ _0359_ _0366_ VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__or2_2
X_5694_ _2652_ VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__clkbuf_1
X_4645_ _1791_ _1458_ VGND VGND VPWR VPWR _1816_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_102_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4576_ game.addmisses.a\[12\] _1767_ VGND VGND VPWR VPWR _1768_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3527_ _0886_ _0608_ VGND VGND VPWR VPWR _0890_ sky130_fd_sc_hd__or2b_1
X_3458_ _0775_ _0776_ net43 _0820_ VGND VGND VPWR VPWR _0821_ sky130_fd_sc_hd__and4b_1
X_3389_ _0725_ _0751_ VGND VGND VPWR VPWR _0752_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_99_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5128_ _2187_ _2215_ VGND VGND VPWR VPWR _2216_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5059_ disp_song.um.drum.next_idx2\[1\] _1992_ _2149_ _2000_ _1983_ VGND VGND VPWR
+ VPWR _2150_ sky130_fd_sc_hd__o311a_1
XFILLER_0_109_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_109_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_105_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold71 game.counter\[12\] VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 game.scoring_button_1.flash_counter_1\[13\] VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__dlygate4sd3_1
Xhold60 game.out\[7\] VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__dlygate4sd3_1
Xhold93 game.scoring_button_2.flash_counter_2\[10\] VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_109_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2760_ modetrans.mode\[5\] _2658_ VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__and2_1
X_2691_ _2654_ _2664_ VGND VGND VPWR VPWR _2665_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_2 _1209_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4430_ _1642_ _1643_ _1638_ VGND VGND VPWR VPWR _1644_ sky130_fd_sc_hd__or3_1
X_6100_ clknet_leaf_37_clk disp_song.um.drum.next_note1\[12\] net67 VGND VGND VPWR
+ VPWR disp_song.note1\[12\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_1_567 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4361_ game.scoring_button_2.flash_counter_1\[13\] game.scoring_button_2.flash_counter_1\[14\]
+ _1586_ VGND VGND VPWR VPWR _1590_ sky130_fd_sc_hd__and3_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3312_ _0563_ _0576_ VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__xor2_4
X_4292_ game.scoring_button_2.flash_counter_2\[15\] _1539_ VGND VGND VPWR VPWR _1543_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_67_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3243_ _0597_ _0601_ _0605_ VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__o21a_1
X_6031_ clknet_leaf_60_clk _0140_ net51 VGND VGND VPWR VPWR game.flash_counter\[11\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3174_ _0535_ _0536_ VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_526 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5815_ clknet_leaf_49_clk game.scoring_button_2.next_flash_counter_2\[6\] net56 VGND
+ VGND VPWR VPWR game.scoring_button_2.flash_counter_2\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_609 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2958_ modetrans.mode\[2\] VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__clkinv_4
XFILLER_0_32_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5746_ clknet_leaf_3_clk game.scoring_button_2.next_num_hits\[2\] net49 VGND VGND
+ VPWR VPWR game.addhits.add1.b\[2\] sky130_fd_sc_hd__dfrtp_2
X_5677_ game.flash_counter\[20\] _2640_ VGND VGND VPWR VPWR _2641_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2889_ _0163_ _0298_ VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__nor2_1
X_4628_ _1807_ VGND VGND VPWR VPWR game.scoring_button_1.next_count\[7\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4559_ game.addmisses.a\[9\] _1716_ _1752_ _1753_ VGND VGND VPWR VPWR _1754_ sky130_fd_sc_hd__a31o_1
XFILLER_0_12_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_492 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_94_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_581 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_101_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_610 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3930_ game.addhits.add2.b\[1\] _1227_ _1255_ _1226_ VGND VGND VPWR VPWR game.scoring_button_2.next_num_hits\[5\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3861_ _0933_ _1203_ VGND VGND VPWR VPWR _1204_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2812_ lvls.level\[0\] _0242_ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__or2_1
X_3792_ _1077_ _1078_ _1110_ VGND VGND VPWR VPWR _1145_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_26_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5600_ disp_song.note1\[31\] game.padded_notes1\[30\] _0209_ VGND VGND VPWR VPWR
+ _2592_ sky130_fd_sc_hd__mux2_1
X_5531_ disp_song.note1\[8\] game.padded_notes1\[7\] _2541_ VGND VGND VPWR VPWR _2546_
+ sky130_fd_sc_hd__mux2_1
X_2743_ _0178_ _0180_ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__nand2_1
XFILLER_0_6_637 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_448 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_147 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5462_ _2504_ net251 _2473_ VGND VGND VPWR VPWR _2505_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5393_ _2456_ _0204_ _2454_ _2457_ _0206_ VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__o311a_1
X_4413_ game.addhits.a\[1\] _1613_ _1631_ _1612_ VGND VGND VPWR VPWR game.scoring_button_1.next_num_hits\[1\]
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4344_ _1578_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_1\[8\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6014_ clknet_leaf_22_clk net120 net59 VGND VGND VPWR VPWR game.out\[1\] sky130_fd_sc_hd__dfrtp_1
X_4275_ net166 _1528_ game.missed_2 VGND VGND VPWR VPWR _1531_ sky130_fd_sc_hd__a21boi_1
X_3226_ _0580_ _0581_ _0582_ VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__o21a_1
XFILLER_0_94_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3157_ _0516_ _0519_ VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__xnor2_1
XTAP_1319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_470 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3088_ game.addmisses.a\[1\] game.addmisses.add1.b\[1\] VGND VGND VPWR VPWR _0451_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_613 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_107_428 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_76_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_573 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5729_ clknet_leaf_0_clk game.scoring_button_2.next_num_misses\[1\] net48 VGND VGND
+ VPWR VPWR game.addmisses.add1.b\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_45_584 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_102_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_102_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_99_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_82_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_629 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4060_ game.addmisses.add3.b\[0\] _1357_ VGND VGND VPWR VPWR _1366_ sky130_fd_sc_hd__nand2_1
X_3011_ _0194_ _0359_ _0366_ _0370_ disp_song.note1\[11\] VGND VGND VPWR VPWR _0395_
+ sky130_fd_sc_hd__o41a_1
XFILLER_0_64_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire38 net39 VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__buf_2
X_4962_ _2020_ _2052_ _2053_ _2055_ _1950_ VGND VGND VPWR VPWR _2056_ sky130_fd_sc_hd__o32a_1
X_4893_ _1956_ disp_song.um.drum.next_note2\[9\] _1987_ VGND VGND VPWR VPWR _1988_
+ sky130_fd_sc_hd__o21ai_1
X_3913_ game.addhits.add1.b\[3\] _1234_ VGND VGND VPWR VPWR _1243_ sky130_fd_sc_hd__nand2_1
XFILLER_0_80_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3844_ _1192_ VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3775_ modetrans.mode\[5\] _0952_ _1121_ _0211_ VGND VGND VPWR VPWR _1129_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5514_ _2534_ VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__clkbuf_1
X_2726_ disp_song.um.idx_note1\[0\] _0170_ VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5445_ disp_song.note2\[15\] game.padded_notes2\[14\] _0219_ VGND VGND VPWR VPWR
+ _2493_ sky130_fd_sc_hd__mux2_1
XFILLER_0_42_576 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5376_ _0848_ _2434_ _0899_ VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__o21ai_1
X_4327_ _1565_ game.hit_2 _1566_ VGND VGND VPWR VPWR _1567_ sky130_fd_sc_hd__and3b_1
X_4258_ game.scoring_button_2.flash_counter_2\[3\] game.scoring_button_2.flash_counter_2\[4\]
+ _1511_ game.scoring_button_2.flash_counter_2\[5\] VGND VGND VPWR VPWR _1519_ sky130_fd_sc_hd__a31o_1
X_3209_ _0570_ _0571_ VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__or2b_1
X_4189_ _1462_ VGND VGND VPWR VPWR game.scoring_button_2.next_count\[17\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold190 game.flash_counter\[18\] VGND VGND VPWR VPWR net263 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_16 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_624 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_95_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3560_ _0879_ _0922_ VGND VGND VPWR VPWR _0923_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5230_ _2232_ _0430_ _2233_ VGND VGND VPWR VPWR _2316_ sky130_fd_sc_hd__o21ai_1
X_3491_ _0762_ _0824_ _0825_ _0826_ _0853_ VGND VGND VPWR VPWR _0854_ sky130_fd_sc_hd__o311a_1
X_5161_ _0176_ disp_song.um.drum.next_note1\[29\] VGND VGND VPWR VPWR _2248_ sky130_fd_sc_hd__or2_1
X_5092_ _2082_ _2080_ _0169_ VGND VGND VPWR VPWR _2181_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4112_ game.scoring_button_2.flash_counter_1\[17\] game.scoring_button_2.flash_counter_1\[16\]
+ game.scoring_button_2.flash_counter_1\[19\] game.scoring_button_2.flash_counter_1\[18\]
+ VGND VGND VPWR VPWR _1411_ sky130_fd_sc_hd__and4_1
X_4043_ game.addmisses.add2.b\[3\] _1344_ VGND VGND VPWR VPWR _1351_ sky130_fd_sc_hd__nand2_1
X_5994_ clknet_leaf_37_clk _0103_ net71 VGND VGND VPWR VPWR game.padded_notes1\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4945_ _1956_ disp_song.um.drum.next_note2\[21\] VGND VGND VPWR VPWR _2039_ sky130_fd_sc_hd__nand2_1
X_4876_ _0169_ _1965_ _1966_ _1970_ VGND VGND VPWR VPWR _1971_ sky130_fd_sc_hd__a31o_1
XFILLER_0_6_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3827_ _1174_ _1177_ VGND VGND VPWR VPWR _1178_ sky130_fd_sc_hd__or2b_1
X_3758_ modetrans.mode\[3\] _0949_ _1101_ _1112_ VGND VGND VPWR VPWR _1113_ sky130_fd_sc_hd__a31o_1
X_2709_ disp_song.um.idx_note2\[4\] VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3689_ _0649_ _1044_ _0642_ VGND VGND VPWR VPWR _1045_ sky130_fd_sc_hd__or3b_1
XFILLER_0_42_384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5428_ _2481_ game.padded_notes2\[9\] _2473_ VGND VGND VPWR VPWR _2482_ sky130_fd_sc_hd__mux2_1
X_5359_ _1035_ highest_score.highest_score\[1\] _2434_ VGND VGND VPWR VPWR _2436_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_613 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_77_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_108_589 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_110_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2991_ _0358_ _0366_ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__nor2_2
XFILLER_0_61_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4730_ _1873_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_2\[18\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_657 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_616 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4661_ game.scoring_button_1.flash_counter_2\[13\] game.scoring_button_1.flash_counter_2\[12\]
+ game.scoring_button_1.flash_counter_2\[15\] game.scoring_button_1.flash_counter_2\[14\]
+ VGND VGND VPWR VPWR _1825_ sky130_fd_sc_hd__or4b_1
XFILLER_0_71_424 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3612_ _0916_ _0971_ _0261_ VGND VGND VPWR VPWR _0972_ sky130_fd_sc_hd__o21ai_1
X_4592_ game.addmisses.a\[14\] _1779_ _1781_ VGND VGND VPWR VPWR _1782_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3543_ highest_score.highest_score\[7\] highest_score.highest_score\[6\] _0898_ VGND
+ VGND VPWR VPWR _0906_ sky130_fd_sc_hd__or3_2
XFILLER_0_12_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3474_ _0804_ _0814_ _0836_ VGND VGND VPWR VPWR _0837_ sky130_fd_sc_hd__and3_1
X_5213_ disp_song.um.drum.next_idx1\[0\] _2230_ _2298_ _2299_ VGND VGND VPWR VPWR
+ _2300_ sky130_fd_sc_hd__a211o_1
X_5144_ _0175_ VGND VGND VPWR VPWR _2232_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_19_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5075_ disp_song.note2\[0\] disp_song.um.drum.next_idx2\[1\] disp_song.um.drum.next_idx2\[0\]
+ disp_song.note2\[1\] VGND VGND VPWR VPWR _2165_ sky130_fd_sc_hd__o22a_1
XFILLER_0_79_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4026_ game.addmisses.add2.b\[1\] _1327_ VGND VGND VPWR VPWR _1336_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5977_ clknet_leaf_34_clk game.scoring_button_1.next_flash_counter_2\[22\] net71
+ VGND VGND VPWR VPWR game.scoring_button_1.flash_counter_2\[22\] sky130_fd_sc_hd__dfrtp_1
X_4928_ _2013_ _2021_ VGND VGND VPWR VPWR _2022_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_627 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4859_ disp_song.um.drum.next_note2\[26\] VGND VGND VPWR VPWR _1954_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_573 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_3_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_3_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_15_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_33_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3190_ _0546_ _0552_ VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__nor2_2
X_5900_ clknet_leaf_44_clk _0083_ net53 VGND VGND VPWR VPWR game.out\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_leaf_73_clk clknet_3_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_73_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_76_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5831_ clknet_leaf_52_clk net88 net55 VGND VGND VPWR VPWR game.scoring_button_2.flash_counter_2\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_2974_ _0358_ _0366_ VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__or2_2
XFILLER_0_8_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5762_ clknet_leaf_0_clk net132 net48 VGND VGND VPWR VPWR game.scoring_button_2.hit
+ sky130_fd_sc_hd__dfrtp_1
X_4713_ game.scoring_button_1.flash_counter_2\[13\] game.scoring_button_1.flash_counter_2\[14\]
+ _1857_ VGND VGND VPWR VPWR _1861_ sky130_fd_sc_hd__and3_1
XFILLER_0_84_582 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5693_ net203 _2530_ VGND VGND VPWR VPWR _2652_ sky130_fd_sc_hd__or2_1
X_4644_ _1815_ VGND VGND VPWR VPWR game.scoring_button_1.next_count\[15\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_608 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4575_ game.addmisses.a\[11\] _1743_ _1755_ VGND VGND VPWR VPWR _1767_ sky130_fd_sc_hd__and3_1
XFILLER_0_12_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_587 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3526_ _0608_ _0886_ VGND VGND VPWR VPWR _0889_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3457_ _0814_ _0819_ VGND VGND VPWR VPWR _0820_ sky130_fd_sc_hd__xnor2_1
X_3388_ _0749_ _0750_ VGND VGND VPWR VPWR _0751_ sky130_fd_sc_hd__and2b_1
X_6176_ clknet_leaf_44_clk disp_song.next_green net54 VGND VGND VPWR VPWR disp_song.toggle_green
+ sky130_fd_sc_hd__dfrtp_1
X_5127_ _0191_ _2185_ VGND VGND VPWR VPWR _2215_ sky130_fd_sc_hd__nand2_1
X_5058_ _2001_ VGND VGND VPWR VPWR _2149_ sky130_fd_sc_hd__inv_2
X_4009_ _1289_ _1318_ _1319_ _1321_ VGND VGND VPWR VPWR game.scoring_button_2.next_num_misses\[2\]
+ sky130_fd_sc_hd__o31a_1
XFILLER_0_67_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_64_clk clknet_3_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_64_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_1_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_105_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold50 game.beat_clk VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold83 game.scoring_button_2.flash_counter_1\[10\] VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold61 _0082_ VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 game.out\[10\] VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 game.addhits.add1.b\[2\] VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_55_clk clknet_3_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_55_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_66_560 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2690_ disp_song.um.idx_note2\[1\] _2663_ VGND VGND VPWR VPWR _2664_ sky130_fd_sc_hd__xor2_2
XFILLER_0_41_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_3 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4360_ net173 _1586_ _1589_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_1\[13\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_111_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3311_ _0665_ _0672_ _0673_ VGND VGND VPWR VPWR _0674_ sky130_fd_sc_hd__a21bo_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_579 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4291_ game.scoring_button_2.flash_counter_2\[15\] _1539_ VGND VGND VPWR VPWR _1542_
+ sky130_fd_sc_hd__and2_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3242_ _0604_ VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__inv_2
X_6030_ clknet_leaf_60_clk _0139_ net51 VGND VGND VPWR VPWR game.flash_counter\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3173_ game.addhits.a\[8\] game.addhits.add3.b\[0\] VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__nor2_1
XFILLER_0_107_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_77 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_46_clk clknet_3_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_46_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_49_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5814_ clknet_leaf_50_clk game.scoring_button_2.next_flash_counter_2\[5\] net56 VGND
+ VGND VPWR VPWR game.scoring_button_2.flash_counter_2\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_76_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_106_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2957_ _0351_ VGND VGND VPWR VPWR disp_song.um.drum.next_note1\[0\] sky130_fd_sc_hd__clkbuf_2
XFILLER_0_8_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5745_ clknet_leaf_1_clk game.scoring_button_2.next_num_hits\[1\] net49 VGND VGND
+ VPWR VPWR game.addhits.add1.b\[1\] sky130_fd_sc_hd__dfrtp_4
X_2888_ _0304_ VGND VGND VPWR VPWR disp_song.um.drum.next_note2\[11\] sky130_fd_sc_hd__buf_1
XFILLER_0_96_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5676_ game.flash_counter\[19\] _2636_ VGND VGND VPWR VPWR _2640_ sky130_fd_sc_hd__and2_1
XFILLER_0_32_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4627_ _1791_ _1430_ VGND VGND VPWR VPWR _1807_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4558_ game.addmisses.a\[9\] _1752_ _1675_ VGND VGND VPWR VPWR _1753_ sky130_fd_sc_hd__o21ai_1
X_3509_ game.flash_counter\[17\] game.flash_counter\[16\] game.flash_counter\[6\]
+ game.flash_counter\[7\] VGND VGND VPWR VPWR _0872_ sky130_fd_sc_hd__or4_1
X_4489_ modetrans.mode\[0\] _1692_ VGND VGND VPWR VPWR _1693_ sky130_fd_sc_hd__nor2_2
X_6159_ clknet_leaf_31_clk net78 net70 VGND VGND VPWR VPWR disp_song.um.boton2e.edge_2
+ sky130_fd_sc_hd__dfrtp_1
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_37_clk clknet_3_6__leaf_clk VGND VGND VPWR VPWR clknet_leaf_37_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_94_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_574 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_106_643 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_28_clk clknet_3_7__leaf_clk VGND VGND VPWR VPWR clknet_leaf_28_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_86_622 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_85_187 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3860_ _0966_ disp_song.display_note1\[4\] _0211_ game.out\[11\] _0208_ VGND VGND
+ VPWR VPWR _1203_ sky130_fd_sc_hd__a221o_2
XFILLER_0_73_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2811_ lvls.level\[2\] lvls.level\[1\] VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__nor2_1
X_3791_ _1077_ _0926_ _1082_ _0925_ VGND VGND VPWR VPWR _1144_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_26_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_109_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5530_ _2545_ VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__clkbuf_1
X_2742_ _0185_ VGND VGND VPWR VPWR disp_song.um.drum.next_idx1\[4\] sky130_fd_sc_hd__inv_2
X_5461_ disp_song.note2\[20\] game.padded_notes2\[19\] _2497_ VGND VGND VPWR VPWR
+ _2504_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4412_ _1621_ _1630_ _1623_ VGND VGND VPWR VPWR _1631_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_55 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5392_ pulseout.fin_pulse\[4\] game.beat_clk _2453_ net265 VGND VGND VPWR VPWR _2457_
+ sky130_fd_sc_hd__a31o_1
XFILLER_0_41_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4343_ _1576_ game.hit_2 _1577_ VGND VGND VPWR VPWR _1578_ sky130_fd_sc_hd__and3b_1
XFILLER_0_1_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4274_ _1530_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_2\[9\]
+ sky130_fd_sc_hd__clkbuf_1
X_6013_ clknet_leaf_22_clk net139 net59 VGND VGND VPWR VPWR game.out\[0\] sky130_fd_sc_hd__dfrtp_1
X_3225_ _0586_ _0587_ VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__or2b_1
XFILLER_0_94_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3156_ _0517_ _0518_ VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_19_clk clknet_3_5__leaf_clk VGND VGND VPWR VPWR clknet_leaf_19_clk sky130_fd_sc_hd__clkbuf_16
X_3087_ game.addmisses.add1.b\[0\] game.addmisses.a\[0\] VGND VGND VPWR VPWR _0450_
+ sky130_fd_sc_hd__nand2_2
XTAP_1309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_482 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_346 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_625 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_107_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5728_ clknet_leaf_0_clk game.scoring_button_2.next_num_misses\[0\] net48 VGND VGND
+ VPWR VPWR game.addmisses.add1.b\[0\] sky130_fd_sc_hd__dfrtp_4
X_3989_ _1302_ _1303_ VGND VGND VPWR VPWR _1304_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_596 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_660 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5659_ _0842_ _2622_ _2627_ VGND VGND VPWR VPWR _2628_ sky130_fd_sc_hd__and3_1
XFILLER_0_60_599 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_102_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_99_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3010_ disp_song.note1\[10\] _0393_ _0394_ _0363_ VGND VGND VPWR VPWR disp_song.um.drum.next_note1\[10\]
+ sky130_fd_sc_hd__a22o_1
Xwire39 _0878_ VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__buf_2
X_4961_ _2020_ _2054_ VGND VGND VPWR VPWR _2055_ sky130_fd_sc_hd__nand2_1
XFILLER_0_59_633 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4892_ disp_song.um.drum.next_idx2\[0\] disp_song.um.drum.next_note2\[8\] VGND VGND
+ VPWR VPWR _1987_ sky130_fd_sc_hd__or2_1
X_3912_ _1241_ VGND VGND VPWR VPWR _1242_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3843_ _0933_ _1191_ VGND VGND VPWR VPWR _1192_ sky130_fd_sc_hd__and2_1
XFILLER_0_104_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3774_ _0949_ _1121_ _1127_ modetrans.mode\[3\] VGND VGND VPWR VPWR _1128_ sky130_fd_sc_hd__o211a_1
X_5513_ _2533_ game.padded_notes1\[2\] _2515_ VGND VGND VPWR VPWR _2534_ sky130_fd_sc_hd__mux2_1
X_2725_ _2657_ _2660_ disp_song.toggle_state VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__o21bai_4
X_5444_ _2492_ VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_8_clk clknet_3_4__leaf_clk VGND VGND VPWR VPWR clknet_leaf_8_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_59_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5375_ _2446_ VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__clkbuf_1
X_4326_ game.scoring_button_2.flash_counter_1\[3\] _1562_ VGND VGND VPWR VPWR _1566_
+ sky130_fd_sc_hd__or2_1
X_4257_ game.scoring_button_2.flash_counter_2\[5\] game.scoring_button_2.flash_counter_2\[4\]
+ _1514_ VGND VGND VPWR VPWR _1518_ sky130_fd_sc_hd__and3_1
X_4188_ _1405_ _0017_ VGND VGND VPWR VPWR _1462_ sky130_fd_sc_hd__and2_1
X_3208_ game.addhits.a\[7\] game.addhits.add2.b\[3\] VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__nand2_1
X_3139_ _0437_ _0500_ _0501_ VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__and3_1
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold180 game.addhits.add2.b\[2\] VGND VGND VPWR VPWR net253 sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 _2635_ VGND VGND VPWR VPWR net264 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3490_ _0784_ VGND VGND VPWR VPWR _0853_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5160_ _2245_ _2246_ VGND VGND VPWR VPWR _2247_ sky130_fd_sc_hd__or2_2
X_5091_ _2074_ _2077_ disp_song.um.drum.next_idx2\[2\] VGND VGND VPWR VPWR _2180_
+ sky130_fd_sc_hd__mux2_1
X_4111_ game.scoring_button_2.flash_counter_1\[21\] game.scoring_button_2.flash_counter_1\[20\]
+ game.scoring_button_2.flash_counter_1\[22\] VGND VGND VPWR VPWR _1410_ sky130_fd_sc_hd__or3_1
XFILLER_0_75_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4042_ _1289_ _1335_ VGND VGND VPWR VPWR _1350_ sky130_fd_sc_hd__nor2_1
X_5993_ clknet_leaf_37_clk _0102_ net71 VGND VGND VPWR VPWR game.padded_notes1\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4944_ _2677_ _0162_ _2012_ VGND VGND VPWR VPWR _2038_ sky130_fd_sc_hd__and3_1
XFILLER_0_19_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4875_ disp_song.um.drum.next_idx2\[1\] _1968_ _1969_ VGND VGND VPWR VPWR _1970_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_62_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_74_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3826_ _0925_ _1175_ _1176_ VGND VGND VPWR VPWR _1177_ sky130_fd_sc_hd__or3b_1
XFILLER_0_6_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3757_ _0966_ _1109_ _1111_ _0953_ VGND VGND VPWR VPWR _1112_ sky130_fd_sc_hd__a31o_1
X_2708_ _2679_ VGND VGND VPWR VPWR disp_song.um.drum.next_idx2\[3\] sky130_fd_sc_hd__inv_2
XFILLER_0_42_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3688_ _0625_ net44 VGND VGND VPWR VPWR _1044_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5427_ disp_song.note2\[9\] game.padded_notes2\[8\] _0219_ VGND VGND VPWR VPWR _2481_
+ sky130_fd_sc_hd__mux2_1
X_5358_ _2435_ VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__clkbuf_1
X_4309_ _1553_ game.missed_2 _1554_ VGND VGND VPWR VPWR _1555_ sky130_fd_sc_hd__and3b_1
X_5289_ _2185_ _2221_ _2224_ VGND VGND VPWR VPWR _2373_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_97_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_97_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_606 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_92_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2990_ _0379_ VGND VGND VPWR VPWR disp_song.um.drum.next_note1\[5\] sky130_fd_sc_hd__clkbuf_2
XTAP_1492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4660_ game.scoring_button_1.flash_counter_2\[1\] game.scoring_button_1.flash_counter_2\[0\]
+ game.scoring_button_1.flash_counter_2\[3\] game.scoring_button_1.flash_counter_2\[2\]
+ VGND VGND VPWR VPWR _1824_ sky130_fd_sc_hd__or4_1
XFILLER_0_44_628 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3611_ _0936_ _0970_ _0919_ VGND VGND VPWR VPWR _0971_ sky130_fd_sc_hd__o21a_1
XFILLER_0_43_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_101_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4591_ _1744_ _1780_ VGND VGND VPWR VPWR _1781_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_51 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3542_ _0900_ highest_score.highest_score\[5\] highest_score.highest_score\[4\] VGND
+ VGND VPWR VPWR _0905_ sky130_fd_sc_hd__or3b_1
XFILLER_0_12_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3473_ _0781_ _0791_ _0813_ VGND VGND VPWR VPWR _0836_ sky130_fd_sc_hd__o21ai_1
X_5212_ _2232_ disp_song.um.drum.next_note1\[0\] VGND VGND VPWR VPWR _2299_ sky130_fd_sc_hd__nor2_1
X_5143_ _0430_ _2230_ VGND VGND VPWR VPWR _2231_ sky130_fd_sc_hd__or2_1
X_5074_ _2034_ _2070_ VGND VGND VPWR VPWR _2164_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4025_ game.addmisses.add2.b\[2\] _1334_ game.addmisses.add2.b\[3\] VGND VGND VPWR
+ VPWR _1335_ sky130_fd_sc_hd__o21a_2
XFILLER_0_79_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5976_ clknet_leaf_33_clk game.scoring_button_1.next_flash_counter_2\[21\] net71
+ VGND VGND VPWR VPWR game.scoring_button_1.flash_counter_2\[21\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_260 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4927_ _2015_ _2018_ _2020_ VGND VGND VPWR VPWR _2021_ sky130_fd_sc_hd__mux2_1
X_4858_ _1950_ _1952_ VGND VGND VPWR VPWR _1953_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_617 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_639 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_585 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3809_ _1156_ _1157_ _1160_ _0935_ VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__o31a_2
XFILLER_0_62_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4789_ _1912_ _1799_ _1913_ VGND VGND VPWR VPWR _1914_ sky130_fd_sc_hd__and3b_1
XFILLER_0_42_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_108_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_21_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5830_ clknet_leaf_46_clk game.scoring_button_2.next_flash_counter_2\[21\] net55
+ VGND VGND VPWR VPWR game.scoring_button_2.flash_counter_2\[21\] sky130_fd_sc_hd__dfrtp_1
X_2973_ _0365_ VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__clkbuf_4
X_5761_ clknet_leaf_62_clk game.scoring_button_2.next_good net53 VGND VGND VPWR VPWR
+ game.hit_2 sky130_fd_sc_hd__dfrtp_4
X_4712_ net184 _1857_ _1860_ VGND VGND VPWR VPWR game.scoring_button_1.next_flash_counter_2\[13\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_17_617 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5692_ _2651_ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4643_ _1791_ _1454_ VGND VGND VPWR VPWR _1815_ sky130_fd_sc_hd__and2_1
XFILLER_0_71_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_661 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4574_ game.addmisses.a\[12\] _1749_ VGND VGND VPWR VPWR _1766_ sky130_fd_sc_hd__nor2_1
X_3525_ _0675_ _0671_ VGND VGND VPWR VPWR _0888_ sky130_fd_sc_hd__or2b_1
XFILLER_0_12_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3456_ _0781_ _0818_ VGND VGND VPWR VPWR _0819_ sky130_fd_sc_hd__nor2_1
X_6175_ clknet_leaf_24_clk disp_song.next_red net65 VGND VGND VPWR VPWR disp_song.toggle_red
+ sky130_fd_sc_hd__dfrtp_1
X_3387_ _0527_ _0524_ _0748_ VGND VGND VPWR VPWR _0750_ sky130_fd_sc_hd__a21o_1
XFILLER_0_41_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5126_ _2188_ _2204_ _2206_ _2213_ VGND VGND VPWR VPWR _2214_ sky130_fd_sc_hd__a31o_1
X_5057_ _2147_ _1989_ _1983_ VGND VGND VPWR VPWR _2148_ sky130_fd_sc_hd__mux2_1
X_4008_ game.addmisses.add1.b\[2\] _1307_ _1320_ net45 VGND VGND VPWR VPWR _1321_
+ sky130_fd_sc_hd__a211o_1
XFILLER_0_94_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5959_ clknet_leaf_36_clk game.scoring_button_1.next_flash_counter_2\[4\] net72 VGND
+ VGND VPWR VPWR game.scoring_button_1.flash_counter_2\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_75_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_105_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_101_574 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold40 game.flash_counter\[2\] VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 game.flash_counter\[5\] VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 game.flash_counter\[0\] VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__dlygate4sd3_1
Xhold62 game.out\[12\] VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_98_620 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold95 game.counter\[4\] VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 game.scoring_button_1.flash_counter_1\[10\] VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_85_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_109_641 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_572 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_609 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_108_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_4 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3310_ _0671_ _0667_ _0668_ VGND VGND VPWR VPWR _0673_ sky130_fd_sc_hd__or3_1
XFILLER_0_67_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4290_ _1541_ VGND VGND VPWR VPWR game.scoring_button_2.next_flash_counter_2\[14\]
+ sky130_fd_sc_hd__clkbuf_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3241_ _0602_ _0603_ VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__nor2_1
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3172_ game.addhits.a\[8\] game.addhits.add3.b\[0\] VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__and2_1
XFILLER_0_83_34 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5813_ clknet_leaf_48_clk game.scoring_button_2.next_flash_counter_2\[4\] net56 VGND
+ VGND VPWR VPWR game.scoring_button_2.flash_counter_2\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_8_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2956_ disp_song.note1\[0\] _0349_ _0350_ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__a21bo_1
X_5744_ clknet_leaf_1_clk game.scoring_button_2.next_num_hits\[0\] net48 VGND VGND
+ VPWR VPWR game.addhits.add1.b\[0\] sky130_fd_sc_hd__dfrtp_4
X_2887_ disp_song.note2\[11\] _0269_ _0303_ VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__mux2_1
X_5675_ _2639_ VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__clkbuf_1
X_4626_ _1806_ VGND VGND VPWR VPWR game.scoring_button_1.next_count\[6\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_653 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_102_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4557_ game.addmisses.a\[8\] _1743_ VGND VGND VPWR VPWR _1752_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3508_ game.flash_counter\[19\] game.flash_counter\[18\] VGND VGND VPWR VPWR _0871_
+ sky130_fd_sc_hd__nand2_1
X_4488_ _1691_ VGND VGND VPWR VPWR _1692_ sky130_fd_sc_hd__inv_2
X_3439_ _0722_ _0711_ _0721_ VGND VGND VPWR VPWR _0802_ sky130_fd_sc_hd__a21oi_1
X_6158_ clknet_leaf_30_clk net4 net70 VGND VGND VPWR VPWR disp_song.um.boton2e.sync_b
+ sky130_fd_sc_hd__dfrtp_1
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5109_ _2195_ _2196_ disp_song.um.drum.next_idx1\[1\] VGND VGND VPWR VPWR _2197_
+ sky130_fd_sc_hd__a21oi_1
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6089_ clknet_leaf_43_clk disp_song.um.drum.next_note1\[1\] net64 VGND VGND VPWR
+ VPWR disp_song.note1\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput30 net30 VGND VGND VPWR VPWR top_row[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_101_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_634 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_561 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2810_ _0227_ VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__inv_2
X_3790_ disp_song.mi6.in\[3\] _1116_ _1082_ _0926_ _1077_ VGND VGND VPWR VPWR _1143_
+ sky130_fd_sc_hd__o221a_1
XFILLER_0_54_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2741_ _0170_ _0183_ _0184_ _2654_ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__o211a_4
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5460_ _2503_ VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4411_ _1621_ _1628_ _1629_ VGND VGND VPWR VPWR _1630_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_111_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_78_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5391_ pulseout.fin_pulse\[4\] VGND VGND VPWR VPWR _2456_ sky130_fd_sc_hd__inv_2
XFILLER_0_10_601 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_645 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4342_ game.scoring_button_2.flash_counter_1\[7\] game.scoring_button_2.flash_counter_1\[6\]
+ _1569_ game.scoring_button_2.flash_counter_1\[8\] VGND VGND VPWR VPWR _1577_ sky130_fd_sc_hd__a31o_1
X_4273_ _1528_ _1486_ _1529_ VGND VGND VPWR VPWR _1530_ sky130_fd_sc_hd__and3b_1
X_6012_ clknet_leaf_43_clk _0121_ net65 VGND VGND VPWR VPWR game.padded_notes1\[31\]
+ sky130_fd_sc_hd__dfstp_1
X_3224_ game.addhits.a\[11\] game.addhits.add3.b\[3\] VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__nand2_1
.ends

