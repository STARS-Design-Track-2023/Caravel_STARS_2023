// This is the unpowered netlist.
module sass_synth (cs,
    hwclk,
    n_rst,
    pwm_o,
    seq_led_on,
    seq_play,
    seq_power,
    tempo_select,
    beat_led,
    mode_out,
    multi,
    note1,
    note2,
    note3,
    note4,
    piano_keys);
 input cs;
 input hwclk;
 input n_rst;
 output pwm_o;
 output seq_led_on;
 input seq_play;
 input seq_power;
 input tempo_select;
 output [7:0] beat_led;
 output [1:0] mode_out;
 output [3:0] multi;
 output [3:0] note1;
 output [3:0] note2;
 output [3:0] note3;
 output [3:0] note4;
 input [14:0] piano_keys;

 wire net146;
 wire _0000_;
 wire _0001_;
 wire _0002_;
 wire _0003_;
 wire _0004_;
 wire _0005_;
 wire _0006_;
 wire _0007_;
 wire _0008_;
 wire _0009_;
 wire _0010_;
 wire _0011_;
 wire _0012_;
 wire _0013_;
 wire _0014_;
 wire _0015_;
 wire _0016_;
 wire _0017_;
 wire _0018_;
 wire _0019_;
 wire _0020_;
 wire _0021_;
 wire _0022_;
 wire _0023_;
 wire _0024_;
 wire _0025_;
 wire _0026_;
 wire _0027_;
 wire _0028_;
 wire _0029_;
 wire _0030_;
 wire _0031_;
 wire _0032_;
 wire _0033_;
 wire _0034_;
 wire _0035_;
 wire _0036_;
 wire _0037_;
 wire _0038_;
 wire _0039_;
 wire _0040_;
 wire _0041_;
 wire _0042_;
 wire _0043_;
 wire _0044_;
 wire _0045_;
 wire _0046_;
 wire _0047_;
 wire _0048_;
 wire _0049_;
 wire _0050_;
 wire _0051_;
 wire _0052_;
 wire _0053_;
 wire _0054_;
 wire _0055_;
 wire _0056_;
 wire _0057_;
 wire _0058_;
 wire _0059_;
 wire _0060_;
 wire _0061_;
 wire _0062_;
 wire _0063_;
 wire _0064_;
 wire _0065_;
 wire _0066_;
 wire _0067_;
 wire _0068_;
 wire _0069_;
 wire _0070_;
 wire _0071_;
 wire _0072_;
 wire _0073_;
 wire _0074_;
 wire _0075_;
 wire _0076_;
 wire _0077_;
 wire _0078_;
 wire _0079_;
 wire _0080_;
 wire _0081_;
 wire _0082_;
 wire _0083_;
 wire _0084_;
 wire _0085_;
 wire _0086_;
 wire _0087_;
 wire _0088_;
 wire _0089_;
 wire _0090_;
 wire _0091_;
 wire _0092_;
 wire _0093_;
 wire _0094_;
 wire _0095_;
 wire _0096_;
 wire _0097_;
 wire _0098_;
 wire _0099_;
 wire _0100_;
 wire _0101_;
 wire _0102_;
 wire _0103_;
 wire _0104_;
 wire _0105_;
 wire _0106_;
 wire _0107_;
 wire _0108_;
 wire _0109_;
 wire _0110_;
 wire _0111_;
 wire _0112_;
 wire _0113_;
 wire _0114_;
 wire _0115_;
 wire _0116_;
 wire _0117_;
 wire _0118_;
 wire _0119_;
 wire _0120_;
 wire _0121_;
 wire _0122_;
 wire _0123_;
 wire _0124_;
 wire _0125_;
 wire _0126_;
 wire _0127_;
 wire _0128_;
 wire _0129_;
 wire _0130_;
 wire _0131_;
 wire _0132_;
 wire _0133_;
 wire _0134_;
 wire _0135_;
 wire _0136_;
 wire _0137_;
 wire _0138_;
 wire _0139_;
 wire _0140_;
 wire _0141_;
 wire _0142_;
 wire _0143_;
 wire _0144_;
 wire _0145_;
 wire _0146_;
 wire _0147_;
 wire _0148_;
 wire _0149_;
 wire _0150_;
 wire _0151_;
 wire _0152_;
 wire _0153_;
 wire _0154_;
 wire _0155_;
 wire _0156_;
 wire _0157_;
 wire _0158_;
 wire _0159_;
 wire _0160_;
 wire _0161_;
 wire _0162_;
 wire _0163_;
 wire _0164_;
 wire _0165_;
 wire _0166_;
 wire _0167_;
 wire _0168_;
 wire _0169_;
 wire _0170_;
 wire _0171_;
 wire _0172_;
 wire _0173_;
 wire _0174_;
 wire _0175_;
 wire _0176_;
 wire _0177_;
 wire _0178_;
 wire _0179_;
 wire _0180_;
 wire _0181_;
 wire _0182_;
 wire _0183_;
 wire _0184_;
 wire _0185_;
 wire _0186_;
 wire _0187_;
 wire _0188_;
 wire _0189_;
 wire _0190_;
 wire _0191_;
 wire _0192_;
 wire _0193_;
 wire _0194_;
 wire _0195_;
 wire _0196_;
 wire _0197_;
 wire _0198_;
 wire _0199_;
 wire _0200_;
 wire _0201_;
 wire _0202_;
 wire _0203_;
 wire _0204_;
 wire _0205_;
 wire _0206_;
 wire _0207_;
 wire _0208_;
 wire _0209_;
 wire _0210_;
 wire _0211_;
 wire _0212_;
 wire _0213_;
 wire _0214_;
 wire _0215_;
 wire _0216_;
 wire _0217_;
 wire _0218_;
 wire _0219_;
 wire _0220_;
 wire _0221_;
 wire _0222_;
 wire _0223_;
 wire _0224_;
 wire _0225_;
 wire _0226_;
 wire _0227_;
 wire _0228_;
 wire _0229_;
 wire _0230_;
 wire _0231_;
 wire _0232_;
 wire _0233_;
 wire _0234_;
 wire _0235_;
 wire _0236_;
 wire _0237_;
 wire _0238_;
 wire _0239_;
 wire _0240_;
 wire _0241_;
 wire _0242_;
 wire _0243_;
 wire _0244_;
 wire _0245_;
 wire _0246_;
 wire _0247_;
 wire _0248_;
 wire _0249_;
 wire _0250_;
 wire _0251_;
 wire _0252_;
 wire _0253_;
 wire _0254_;
 wire _0255_;
 wire _0256_;
 wire _0257_;
 wire _0258_;
 wire _0259_;
 wire _0260_;
 wire _0261_;
 wire _0262_;
 wire _0263_;
 wire _0264_;
 wire _0265_;
 wire _0266_;
 wire _0267_;
 wire _0268_;
 wire _0269_;
 wire _0270_;
 wire _0271_;
 wire _0272_;
 wire _0273_;
 wire _0274_;
 wire _0275_;
 wire _0276_;
 wire _0277_;
 wire _0278_;
 wire _0279_;
 wire _0280_;
 wire _0281_;
 wire _0282_;
 wire _0283_;
 wire _0284_;
 wire _0285_;
 wire _0286_;
 wire _0287_;
 wire _0288_;
 wire _0289_;
 wire _0290_;
 wire _0291_;
 wire _0292_;
 wire _0293_;
 wire _0294_;
 wire _0295_;
 wire _0296_;
 wire _0297_;
 wire _0298_;
 wire _0299_;
 wire _0300_;
 wire _0301_;
 wire _0302_;
 wire _0303_;
 wire _0304_;
 wire _0305_;
 wire _0306_;
 wire _0307_;
 wire _0308_;
 wire _0309_;
 wire _0310_;
 wire _0311_;
 wire _0312_;
 wire _0313_;
 wire _0314_;
 wire _0315_;
 wire _0316_;
 wire _0317_;
 wire _0318_;
 wire _0319_;
 wire _0320_;
 wire _0321_;
 wire _0322_;
 wire _0323_;
 wire _0324_;
 wire _0325_;
 wire _0326_;
 wire _0327_;
 wire _0328_;
 wire _0329_;
 wire _0330_;
 wire _0331_;
 wire _0332_;
 wire _0333_;
 wire _0334_;
 wire _0335_;
 wire _0336_;
 wire _0337_;
 wire _0338_;
 wire _0339_;
 wire _0340_;
 wire _0341_;
 wire _0342_;
 wire _0343_;
 wire _0344_;
 wire _0345_;
 wire _0346_;
 wire _0347_;
 wire _0348_;
 wire _0349_;
 wire _0350_;
 wire _0351_;
 wire _0352_;
 wire _0353_;
 wire _0354_;
 wire _0355_;
 wire _0356_;
 wire _0357_;
 wire _0358_;
 wire _0359_;
 wire _0360_;
 wire _0361_;
 wire _0362_;
 wire _0363_;
 wire _0364_;
 wire _0365_;
 wire _0366_;
 wire _0367_;
 wire _0368_;
 wire _0369_;
 wire _0370_;
 wire _0371_;
 wire _0372_;
 wire _0373_;
 wire _0374_;
 wire _0375_;
 wire _0376_;
 wire _0377_;
 wire _0378_;
 wire _0379_;
 wire _0380_;
 wire _0381_;
 wire _0382_;
 wire _0383_;
 wire _0384_;
 wire _0385_;
 wire _0386_;
 wire _0387_;
 wire _0388_;
 wire _0389_;
 wire _0390_;
 wire _0391_;
 wire _0392_;
 wire _0393_;
 wire _0394_;
 wire _0395_;
 wire _0396_;
 wire _0397_;
 wire _0398_;
 wire _0399_;
 wire _0400_;
 wire _0401_;
 wire _0402_;
 wire _0403_;
 wire _0404_;
 wire _0405_;
 wire _0406_;
 wire _0407_;
 wire _0408_;
 wire _0409_;
 wire _0410_;
 wire _0411_;
 wire _0412_;
 wire _0413_;
 wire _0414_;
 wire _0415_;
 wire _0416_;
 wire _0417_;
 wire _0418_;
 wire _0419_;
 wire _0420_;
 wire _0421_;
 wire _0422_;
 wire _0423_;
 wire _0424_;
 wire _0425_;
 wire _0426_;
 wire _0427_;
 wire _0428_;
 wire _0429_;
 wire _0430_;
 wire _0431_;
 wire _0432_;
 wire _0433_;
 wire _0434_;
 wire _0435_;
 wire _0436_;
 wire _0437_;
 wire _0438_;
 wire _0439_;
 wire _0440_;
 wire _0441_;
 wire _0442_;
 wire _0443_;
 wire _0444_;
 wire _0445_;
 wire _0446_;
 wire _0447_;
 wire _0448_;
 wire _0449_;
 wire _0450_;
 wire _0451_;
 wire _0452_;
 wire _0453_;
 wire _0454_;
 wire _0455_;
 wire _0456_;
 wire _0457_;
 wire _0458_;
 wire _0459_;
 wire _0460_;
 wire _0461_;
 wire _0462_;
 wire _0463_;
 wire _0464_;
 wire _0465_;
 wire _0466_;
 wire _0467_;
 wire _0468_;
 wire _0469_;
 wire _0470_;
 wire _0471_;
 wire _0472_;
 wire _0473_;
 wire _0474_;
 wire _0475_;
 wire _0476_;
 wire _0477_;
 wire _0478_;
 wire _0479_;
 wire _0480_;
 wire _0481_;
 wire _0482_;
 wire _0483_;
 wire _0484_;
 wire _0485_;
 wire _0486_;
 wire _0487_;
 wire _0488_;
 wire _0489_;
 wire _0490_;
 wire _0491_;
 wire _0492_;
 wire _0493_;
 wire _0494_;
 wire _0495_;
 wire _0496_;
 wire _0497_;
 wire _0498_;
 wire _0499_;
 wire _0500_;
 wire _0501_;
 wire _0502_;
 wire _0503_;
 wire _0504_;
 wire _0505_;
 wire _0506_;
 wire _0507_;
 wire _0508_;
 wire _0509_;
 wire _0510_;
 wire _0511_;
 wire _0512_;
 wire _0513_;
 wire _0514_;
 wire _0515_;
 wire _0516_;
 wire _0517_;
 wire _0518_;
 wire _0519_;
 wire _0520_;
 wire _0521_;
 wire _0522_;
 wire _0523_;
 wire _0524_;
 wire _0525_;
 wire _0526_;
 wire _0527_;
 wire _0528_;
 wire _0529_;
 wire _0530_;
 wire _0531_;
 wire _0532_;
 wire _0533_;
 wire _0534_;
 wire _0535_;
 wire _0536_;
 wire _0537_;
 wire _0538_;
 wire _0539_;
 wire _0540_;
 wire _0541_;
 wire _0542_;
 wire _0543_;
 wire _0544_;
 wire _0545_;
 wire _0546_;
 wire _0547_;
 wire _0548_;
 wire _0549_;
 wire _0550_;
 wire _0551_;
 wire _0552_;
 wire _0553_;
 wire _0554_;
 wire _0555_;
 wire _0556_;
 wire _0557_;
 wire _0558_;
 wire _0559_;
 wire _0560_;
 wire _0561_;
 wire _0562_;
 wire _0563_;
 wire _0564_;
 wire _0565_;
 wire _0566_;
 wire _0567_;
 wire _0568_;
 wire _0569_;
 wire _0570_;
 wire _0571_;
 wire _0572_;
 wire _0573_;
 wire _0574_;
 wire _0575_;
 wire _0576_;
 wire _0577_;
 wire _0578_;
 wire _0579_;
 wire _0580_;
 wire _0581_;
 wire _0582_;
 wire _0583_;
 wire _0584_;
 wire _0585_;
 wire _0586_;
 wire _0587_;
 wire _0588_;
 wire _0589_;
 wire _0590_;
 wire _0591_;
 wire _0592_;
 wire _0593_;
 wire _0594_;
 wire _0595_;
 wire _0596_;
 wire _0597_;
 wire _0598_;
 wire _0599_;
 wire _0600_;
 wire _0601_;
 wire _0602_;
 wire _0603_;
 wire _0604_;
 wire _0605_;
 wire _0606_;
 wire _0607_;
 wire _0608_;
 wire _0609_;
 wire _0610_;
 wire _0611_;
 wire _0612_;
 wire _0613_;
 wire _0614_;
 wire _0615_;
 wire _0616_;
 wire _0617_;
 wire _0618_;
 wire _0619_;
 wire _0620_;
 wire _0621_;
 wire _0622_;
 wire _0623_;
 wire _0624_;
 wire _0625_;
 wire _0626_;
 wire _0627_;
 wire _0628_;
 wire _0629_;
 wire _0630_;
 wire _0631_;
 wire _0632_;
 wire _0633_;
 wire _0634_;
 wire _0635_;
 wire _0636_;
 wire _0637_;
 wire _0638_;
 wire _0639_;
 wire _0640_;
 wire _0641_;
 wire _0642_;
 wire _0643_;
 wire _0644_;
 wire _0645_;
 wire _0646_;
 wire _0647_;
 wire _0648_;
 wire _0649_;
 wire _0650_;
 wire _0651_;
 wire _0652_;
 wire _0653_;
 wire _0654_;
 wire _0655_;
 wire _0656_;
 wire _0657_;
 wire _0658_;
 wire _0659_;
 wire _0660_;
 wire _0661_;
 wire _0662_;
 wire _0663_;
 wire _0664_;
 wire _0665_;
 wire _0666_;
 wire _0667_;
 wire _0668_;
 wire _0669_;
 wire _0670_;
 wire _0671_;
 wire _0672_;
 wire _0673_;
 wire _0674_;
 wire _0675_;
 wire _0676_;
 wire _0677_;
 wire _0678_;
 wire _0679_;
 wire _0680_;
 wire _0681_;
 wire _0682_;
 wire _0683_;
 wire _0684_;
 wire _0685_;
 wire _0686_;
 wire _0687_;
 wire _0688_;
 wire _0689_;
 wire _0690_;
 wire _0691_;
 wire _0692_;
 wire _0693_;
 wire _0694_;
 wire _0695_;
 wire _0696_;
 wire _0697_;
 wire _0698_;
 wire _0699_;
 wire _0700_;
 wire _0701_;
 wire _0702_;
 wire _0703_;
 wire _0704_;
 wire _0705_;
 wire _0706_;
 wire _0707_;
 wire _0708_;
 wire _0709_;
 wire _0710_;
 wire _0711_;
 wire _0712_;
 wire _0713_;
 wire _0714_;
 wire _0715_;
 wire _0716_;
 wire _0717_;
 wire _0718_;
 wire _0719_;
 wire _0720_;
 wire _0721_;
 wire _0722_;
 wire _0723_;
 wire _0724_;
 wire _0725_;
 wire _0726_;
 wire _0727_;
 wire _0728_;
 wire _0729_;
 wire _0730_;
 wire _0731_;
 wire _0732_;
 wire _0733_;
 wire _0734_;
 wire _0735_;
 wire _0736_;
 wire _0737_;
 wire _0738_;
 wire _0739_;
 wire _0740_;
 wire _0741_;
 wire _0742_;
 wire _0743_;
 wire _0744_;
 wire _0745_;
 wire _0746_;
 wire _0747_;
 wire _0748_;
 wire _0749_;
 wire _0750_;
 wire _0751_;
 wire _0752_;
 wire _0753_;
 wire _0754_;
 wire _0755_;
 wire _0756_;
 wire _0757_;
 wire _0758_;
 wire _0759_;
 wire _0760_;
 wire _0761_;
 wire _0762_;
 wire _0763_;
 wire _0764_;
 wire _0765_;
 wire _0766_;
 wire _0767_;
 wire _0768_;
 wire _0769_;
 wire _0770_;
 wire _0771_;
 wire _0772_;
 wire _0773_;
 wire _0774_;
 wire _0775_;
 wire _0776_;
 wire _0777_;
 wire _0778_;
 wire _0779_;
 wire _0780_;
 wire _0781_;
 wire _0782_;
 wire _0783_;
 wire _0784_;
 wire _0785_;
 wire _0786_;
 wire _0787_;
 wire _0788_;
 wire _0789_;
 wire _0790_;
 wire _0791_;
 wire _0792_;
 wire _0793_;
 wire _0794_;
 wire _0795_;
 wire _0796_;
 wire _0797_;
 wire _0798_;
 wire _0799_;
 wire _0800_;
 wire _0801_;
 wire _0802_;
 wire _0803_;
 wire _0804_;
 wire _0805_;
 wire _0806_;
 wire _0807_;
 wire _0808_;
 wire _0809_;
 wire _0810_;
 wire _0811_;
 wire _0812_;
 wire _0813_;
 wire _0814_;
 wire _0815_;
 wire _0816_;
 wire _0817_;
 wire _0818_;
 wire _0819_;
 wire _0820_;
 wire _0821_;
 wire _0822_;
 wire _0823_;
 wire _0824_;
 wire _0825_;
 wire _0826_;
 wire _0827_;
 wire _0828_;
 wire _0829_;
 wire _0830_;
 wire _0831_;
 wire _0832_;
 wire _0833_;
 wire _0834_;
 wire _0835_;
 wire _0836_;
 wire _0837_;
 wire _0838_;
 wire _0839_;
 wire _0840_;
 wire _0841_;
 wire _0842_;
 wire _0843_;
 wire _0844_;
 wire _0845_;
 wire _0846_;
 wire _0847_;
 wire _0848_;
 wire _0849_;
 wire _0850_;
 wire _0851_;
 wire _0852_;
 wire _0853_;
 wire _0854_;
 wire _0855_;
 wire _0856_;
 wire _0857_;
 wire _0858_;
 wire _0859_;
 wire _0860_;
 wire _0861_;
 wire _0862_;
 wire _0863_;
 wire _0864_;
 wire _0865_;
 wire _0866_;
 wire _0867_;
 wire _0868_;
 wire _0869_;
 wire _0870_;
 wire _0871_;
 wire _0872_;
 wire _0873_;
 wire _0874_;
 wire _0875_;
 wire _0876_;
 wire _0877_;
 wire _0878_;
 wire _0879_;
 wire _0880_;
 wire _0881_;
 wire _0882_;
 wire _0883_;
 wire _0884_;
 wire _0885_;
 wire _0886_;
 wire _0887_;
 wire _0888_;
 wire _0889_;
 wire _0890_;
 wire _0891_;
 wire _0892_;
 wire _0893_;
 wire _0894_;
 wire _0895_;
 wire _0896_;
 wire _0897_;
 wire _0898_;
 wire _0899_;
 wire _0900_;
 wire _0901_;
 wire _0902_;
 wire _0903_;
 wire _0904_;
 wire _0905_;
 wire _0906_;
 wire _0907_;
 wire _0908_;
 wire _0909_;
 wire _0910_;
 wire _0911_;
 wire _0912_;
 wire _0913_;
 wire _0914_;
 wire _0915_;
 wire _0916_;
 wire _0917_;
 wire _0918_;
 wire _0919_;
 wire _0920_;
 wire _0921_;
 wire _0922_;
 wire _0923_;
 wire _0924_;
 wire _0925_;
 wire _0926_;
 wire _0927_;
 wire _0928_;
 wire _0929_;
 wire _0930_;
 wire _0931_;
 wire _0932_;
 wire _0933_;
 wire _0934_;
 wire _0935_;
 wire _0936_;
 wire _0937_;
 wire _0938_;
 wire _0939_;
 wire _0940_;
 wire _0941_;
 wire _0942_;
 wire _0943_;
 wire _0944_;
 wire _0945_;
 wire _0946_;
 wire _0947_;
 wire _0948_;
 wire _0949_;
 wire _0950_;
 wire _0951_;
 wire _0952_;
 wire _0953_;
 wire _0954_;
 wire _0955_;
 wire _0956_;
 wire _0957_;
 wire _0958_;
 wire _0959_;
 wire _0960_;
 wire _0961_;
 wire _0962_;
 wire _0963_;
 wire _0964_;
 wire _0965_;
 wire _0966_;
 wire _0967_;
 wire _0968_;
 wire _0969_;
 wire _0970_;
 wire _0971_;
 wire _0972_;
 wire _0973_;
 wire _0974_;
 wire _0975_;
 wire _0976_;
 wire _0977_;
 wire _0978_;
 wire _0979_;
 wire _0980_;
 wire _0981_;
 wire _0982_;
 wire _0983_;
 wire _0984_;
 wire _0985_;
 wire _0986_;
 wire _0987_;
 wire _0988_;
 wire _0989_;
 wire _0990_;
 wire _0991_;
 wire _0992_;
 wire _0993_;
 wire _0994_;
 wire _0995_;
 wire _0996_;
 wire _0997_;
 wire _0998_;
 wire _0999_;
 wire _1000_;
 wire _1001_;
 wire _1002_;
 wire _1003_;
 wire _1004_;
 wire _1005_;
 wire _1006_;
 wire _1007_;
 wire _1008_;
 wire _1009_;
 wire _1010_;
 wire _1011_;
 wire _1012_;
 wire _1013_;
 wire _1014_;
 wire _1015_;
 wire _1016_;
 wire _1017_;
 wire _1018_;
 wire _1019_;
 wire _1020_;
 wire _1021_;
 wire _1022_;
 wire _1023_;
 wire _1024_;
 wire _1025_;
 wire _1026_;
 wire _1027_;
 wire _1028_;
 wire _1029_;
 wire _1030_;
 wire _1031_;
 wire _1032_;
 wire _1033_;
 wire _1034_;
 wire _1035_;
 wire _1036_;
 wire _1037_;
 wire _1038_;
 wire _1039_;
 wire _1040_;
 wire _1041_;
 wire _1042_;
 wire _1043_;
 wire _1044_;
 wire _1045_;
 wire _1046_;
 wire _1047_;
 wire _1048_;
 wire _1049_;
 wire _1050_;
 wire _1051_;
 wire _1052_;
 wire _1053_;
 wire _1054_;
 wire _1055_;
 wire _1056_;
 wire _1057_;
 wire _1058_;
 wire _1059_;
 wire _1060_;
 wire _1061_;
 wire _1062_;
 wire _1063_;
 wire _1064_;
 wire _1065_;
 wire _1066_;
 wire _1067_;
 wire _1068_;
 wire _1069_;
 wire _1070_;
 wire _1071_;
 wire _1072_;
 wire _1073_;
 wire _1074_;
 wire _1075_;
 wire _1076_;
 wire _1077_;
 wire _1078_;
 wire _1079_;
 wire _1080_;
 wire _1081_;
 wire _1082_;
 wire _1083_;
 wire _1084_;
 wire _1085_;
 wire _1086_;
 wire _1087_;
 wire _1088_;
 wire _1089_;
 wire _1090_;
 wire _1091_;
 wire _1092_;
 wire _1093_;
 wire _1094_;
 wire _1095_;
 wire _1096_;
 wire _1097_;
 wire _1098_;
 wire _1099_;
 wire _1100_;
 wire _1101_;
 wire _1102_;
 wire _1103_;
 wire _1104_;
 wire _1105_;
 wire _1106_;
 wire _1107_;
 wire _1108_;
 wire _1109_;
 wire _1110_;
 wire _1111_;
 wire _1112_;
 wire _1113_;
 wire _1114_;
 wire _1115_;
 wire _1116_;
 wire _1117_;
 wire _1118_;
 wire _1119_;
 wire _1120_;
 wire _1121_;
 wire _1122_;
 wire _1123_;
 wire _1124_;
 wire _1125_;
 wire _1126_;
 wire _1127_;
 wire _1128_;
 wire _1129_;
 wire _1130_;
 wire _1131_;
 wire _1132_;
 wire _1133_;
 wire _1134_;
 wire _1135_;
 wire _1136_;
 wire _1137_;
 wire _1138_;
 wire _1139_;
 wire _1140_;
 wire _1141_;
 wire _1142_;
 wire _1143_;
 wire _1144_;
 wire _1145_;
 wire _1146_;
 wire _1147_;
 wire _1148_;
 wire _1149_;
 wire _1150_;
 wire _1151_;
 wire _1152_;
 wire _1153_;
 wire _1154_;
 wire _1155_;
 wire _1156_;
 wire _1157_;
 wire _1158_;
 wire _1159_;
 wire _1160_;
 wire _1161_;
 wire _1162_;
 wire _1163_;
 wire _1164_;
 wire _1165_;
 wire _1166_;
 wire _1167_;
 wire _1168_;
 wire _1169_;
 wire _1170_;
 wire _1171_;
 wire _1172_;
 wire _1173_;
 wire _1174_;
 wire _1175_;
 wire _1176_;
 wire _1177_;
 wire _1178_;
 wire _1179_;
 wire _1180_;
 wire _1181_;
 wire _1182_;
 wire _1183_;
 wire _1184_;
 wire _1185_;
 wire _1186_;
 wire _1187_;
 wire _1188_;
 wire _1189_;
 wire _1190_;
 wire _1191_;
 wire _1192_;
 wire _1193_;
 wire _1194_;
 wire _1195_;
 wire _1196_;
 wire _1197_;
 wire _1198_;
 wire _1199_;
 wire _1200_;
 wire _1201_;
 wire _1202_;
 wire _1203_;
 wire _1204_;
 wire _1205_;
 wire _1206_;
 wire _1207_;
 wire _1208_;
 wire _1209_;
 wire _1210_;
 wire _1211_;
 wire _1212_;
 wire _1213_;
 wire _1214_;
 wire _1215_;
 wire _1216_;
 wire _1217_;
 wire _1218_;
 wire _1219_;
 wire _1220_;
 wire _1221_;
 wire _1222_;
 wire _1223_;
 wire _1224_;
 wire _1225_;
 wire _1226_;
 wire _1227_;
 wire _1228_;
 wire _1229_;
 wire _1230_;
 wire _1231_;
 wire _1232_;
 wire _1233_;
 wire _1234_;
 wire _1235_;
 wire _1236_;
 wire _1237_;
 wire _1238_;
 wire _1239_;
 wire _1240_;
 wire _1241_;
 wire _1242_;
 wire _1243_;
 wire _1244_;
 wire _1245_;
 wire _1246_;
 wire _1247_;
 wire _1248_;
 wire _1249_;
 wire _1250_;
 wire _1251_;
 wire _1252_;
 wire _1253_;
 wire _1254_;
 wire _1255_;
 wire _1256_;
 wire _1257_;
 wire _1258_;
 wire _1259_;
 wire _1260_;
 wire _1261_;
 wire _1262_;
 wire _1263_;
 wire _1264_;
 wire _1265_;
 wire _1266_;
 wire _1267_;
 wire _1268_;
 wire _1269_;
 wire _1270_;
 wire _1271_;
 wire _1272_;
 wire _1273_;
 wire _1274_;
 wire _1275_;
 wire _1276_;
 wire _1277_;
 wire _1278_;
 wire _1279_;
 wire _1280_;
 wire _1281_;
 wire _1282_;
 wire _1283_;
 wire _1284_;
 wire _1285_;
 wire _1286_;
 wire _1287_;
 wire _1288_;
 wire _1289_;
 wire _1290_;
 wire _1291_;
 wire _1292_;
 wire _1293_;
 wire _1294_;
 wire _1295_;
 wire _1296_;
 wire _1297_;
 wire _1298_;
 wire _1299_;
 wire _1300_;
 wire _1301_;
 wire _1302_;
 wire _1303_;
 wire _1304_;
 wire _1305_;
 wire _1306_;
 wire _1307_;
 wire _1308_;
 wire _1309_;
 wire _1310_;
 wire _1311_;
 wire _1312_;
 wire _1313_;
 wire _1314_;
 wire _1315_;
 wire _1316_;
 wire _1317_;
 wire _1318_;
 wire _1319_;
 wire _1320_;
 wire _1321_;
 wire _1322_;
 wire _1323_;
 wire _1324_;
 wire _1325_;
 wire _1326_;
 wire _1327_;
 wire _1328_;
 wire _1329_;
 wire _1330_;
 wire _1331_;
 wire _1332_;
 wire _1333_;
 wire _1334_;
 wire _1335_;
 wire _1336_;
 wire _1337_;
 wire _1338_;
 wire _1339_;
 wire _1340_;
 wire _1341_;
 wire _1342_;
 wire _1343_;
 wire _1344_;
 wire _1345_;
 wire _1346_;
 wire _1347_;
 wire _1348_;
 wire _1349_;
 wire _1350_;
 wire _1351_;
 wire _1352_;
 wire _1353_;
 wire _1354_;
 wire _1355_;
 wire _1356_;
 wire _1357_;
 wire _1358_;
 wire _1359_;
 wire _1360_;
 wire _1361_;
 wire _1362_;
 wire _1363_;
 wire _1364_;
 wire _1365_;
 wire _1366_;
 wire _1367_;
 wire _1368_;
 wire _1369_;
 wire _1370_;
 wire _1371_;
 wire _1372_;
 wire _1373_;
 wire _1374_;
 wire _1375_;
 wire _1376_;
 wire _1377_;
 wire _1378_;
 wire _1379_;
 wire _1380_;
 wire _1381_;
 wire _1382_;
 wire _1383_;
 wire _1384_;
 wire _1385_;
 wire _1386_;
 wire _1387_;
 wire _1388_;
 wire _1389_;
 wire _1390_;
 wire _1391_;
 wire _1392_;
 wire _1393_;
 wire _1394_;
 wire _1395_;
 wire _1396_;
 wire _1397_;
 wire _1398_;
 wire _1399_;
 wire _1400_;
 wire _1401_;
 wire _1402_;
 wire _1403_;
 wire _1404_;
 wire _1405_;
 wire _1406_;
 wire _1407_;
 wire _1408_;
 wire _1409_;
 wire _1410_;
 wire _1411_;
 wire _1412_;
 wire _1413_;
 wire _1414_;
 wire _1415_;
 wire _1416_;
 wire _1417_;
 wire _1418_;
 wire _1419_;
 wire _1420_;
 wire _1421_;
 wire _1422_;
 wire _1423_;
 wire _1424_;
 wire _1425_;
 wire _1426_;
 wire _1427_;
 wire _1428_;
 wire _1429_;
 wire _1430_;
 wire _1431_;
 wire _1432_;
 wire _1433_;
 wire _1434_;
 wire _1435_;
 wire _1436_;
 wire _1437_;
 wire _1438_;
 wire _1439_;
 wire _1440_;
 wire _1441_;
 wire _1442_;
 wire _1443_;
 wire _1444_;
 wire _1445_;
 wire _1446_;
 wire _1447_;
 wire _1448_;
 wire _1449_;
 wire _1450_;
 wire _1451_;
 wire _1452_;
 wire _1453_;
 wire _1454_;
 wire _1455_;
 wire _1456_;
 wire _1457_;
 wire _1458_;
 wire _1459_;
 wire _1460_;
 wire _1461_;
 wire _1462_;
 wire _1463_;
 wire _1464_;
 wire _1465_;
 wire _1466_;
 wire _1467_;
 wire _1468_;
 wire _1469_;
 wire _1470_;
 wire _1471_;
 wire _1472_;
 wire _1473_;
 wire _1474_;
 wire _1475_;
 wire _1476_;
 wire _1477_;
 wire _1478_;
 wire _1479_;
 wire _1480_;
 wire _1481_;
 wire _1482_;
 wire _1483_;
 wire _1484_;
 wire _1485_;
 wire _1486_;
 wire _1487_;
 wire _1488_;
 wire _1489_;
 wire _1490_;
 wire _1491_;
 wire _1492_;
 wire _1493_;
 wire _1494_;
 wire _1495_;
 wire _1496_;
 wire _1497_;
 wire _1498_;
 wire _1499_;
 wire _1500_;
 wire _1501_;
 wire _1502_;
 wire _1503_;
 wire _1504_;
 wire _1505_;
 wire _1506_;
 wire _1507_;
 wire _1508_;
 wire _1509_;
 wire _1510_;
 wire _1511_;
 wire _1512_;
 wire _1513_;
 wire _1514_;
 wire _1515_;
 wire _1516_;
 wire _1517_;
 wire _1518_;
 wire _1519_;
 wire _1520_;
 wire _1521_;
 wire _1522_;
 wire _1523_;
 wire _1524_;
 wire _1525_;
 wire _1526_;
 wire _1527_;
 wire _1528_;
 wire _1529_;
 wire _1530_;
 wire _1531_;
 wire _1532_;
 wire _1533_;
 wire _1534_;
 wire _1535_;
 wire _1536_;
 wire _1537_;
 wire _1538_;
 wire _1539_;
 wire _1540_;
 wire _1541_;
 wire _1542_;
 wire _1543_;
 wire _1544_;
 wire _1545_;
 wire _1546_;
 wire _1547_;
 wire _1548_;
 wire _1549_;
 wire _1550_;
 wire _1551_;
 wire _1552_;
 wire _1553_;
 wire _1554_;
 wire _1555_;
 wire _1556_;
 wire _1557_;
 wire _1558_;
 wire _1559_;
 wire _1560_;
 wire _1561_;
 wire _1562_;
 wire _1563_;
 wire _1564_;
 wire _1565_;
 wire _1566_;
 wire _1567_;
 wire _1568_;
 wire _1569_;
 wire _1570_;
 wire _1571_;
 wire _1572_;
 wire _1573_;
 wire _1574_;
 wire _1575_;
 wire _1576_;
 wire _1577_;
 wire _1578_;
 wire _1579_;
 wire _1580_;
 wire _1581_;
 wire _1582_;
 wire _1583_;
 wire _1584_;
 wire _1585_;
 wire _1586_;
 wire _1587_;
 wire _1588_;
 wire _1589_;
 wire _1590_;
 wire _1591_;
 wire _1592_;
 wire _1593_;
 wire _1594_;
 wire _1595_;
 wire _1596_;
 wire _1597_;
 wire _1598_;
 wire _1599_;
 wire _1600_;
 wire _1601_;
 wire _1602_;
 wire _1603_;
 wire _1604_;
 wire _1605_;
 wire _1606_;
 wire _1607_;
 wire _1608_;
 wire _1609_;
 wire _1610_;
 wire _1611_;
 wire _1612_;
 wire _1613_;
 wire _1614_;
 wire _1615_;
 wire _1616_;
 wire _1617_;
 wire _1618_;
 wire _1619_;
 wire _1620_;
 wire _1621_;
 wire _1622_;
 wire _1623_;
 wire _1624_;
 wire _1625_;
 wire _1626_;
 wire _1627_;
 wire _1628_;
 wire _1629_;
 wire _1630_;
 wire _1631_;
 wire _1632_;
 wire _1633_;
 wire _1634_;
 wire _1635_;
 wire _1636_;
 wire _1637_;
 wire _1638_;
 wire _1639_;
 wire _1640_;
 wire _1641_;
 wire _1642_;
 wire _1643_;
 wire _1644_;
 wire _1645_;
 wire _1646_;
 wire _1647_;
 wire _1648_;
 wire _1649_;
 wire _1650_;
 wire _1651_;
 wire _1652_;
 wire _1653_;
 wire _1654_;
 wire _1655_;
 wire _1656_;
 wire _1657_;
 wire _1658_;
 wire _1659_;
 wire _1660_;
 wire _1661_;
 wire _1662_;
 wire _1663_;
 wire _1664_;
 wire _1665_;
 wire _1666_;
 wire _1667_;
 wire _1668_;
 wire _1669_;
 wire _1670_;
 wire _1671_;
 wire _1672_;
 wire _1673_;
 wire _1674_;
 wire _1675_;
 wire _1676_;
 wire _1677_;
 wire _1678_;
 wire _1679_;
 wire _1680_;
 wire _1681_;
 wire _1682_;
 wire _1683_;
 wire _1684_;
 wire _1685_;
 wire _1686_;
 wire _1687_;
 wire _1688_;
 wire _1689_;
 wire _1690_;
 wire _1691_;
 wire _1692_;
 wire _1693_;
 wire _1694_;
 wire _1695_;
 wire _1696_;
 wire _1697_;
 wire _1698_;
 wire _1699_;
 wire _1700_;
 wire _1701_;
 wire _1702_;
 wire _1703_;
 wire _1704_;
 wire _1705_;
 wire _1706_;
 wire _1707_;
 wire _1708_;
 wire _1709_;
 wire _1710_;
 wire _1711_;
 wire _1712_;
 wire _1713_;
 wire _1714_;
 wire _1715_;
 wire _1716_;
 wire _1717_;
 wire _1718_;
 wire _1719_;
 wire _1720_;
 wire _1721_;
 wire _1722_;
 wire _1723_;
 wire _1724_;
 wire _1725_;
 wire _1726_;
 wire _1727_;
 wire _1728_;
 wire _1729_;
 wire _1730_;
 wire _1731_;
 wire _1732_;
 wire _1733_;
 wire _1734_;
 wire _1735_;
 wire _1736_;
 wire _1737_;
 wire _1738_;
 wire _1739_;
 wire _1740_;
 wire _1741_;
 wire _1742_;
 wire _1743_;
 wire _1744_;
 wire _1745_;
 wire _1746_;
 wire _1747_;
 wire _1748_;
 wire _1749_;
 wire _1750_;
 wire _1751_;
 wire _1752_;
 wire _1753_;
 wire _1754_;
 wire _1755_;
 wire _1756_;
 wire _1757_;
 wire _1758_;
 wire _1759_;
 wire _1760_;
 wire _1761_;
 wire _1762_;
 wire _1763_;
 wire _1764_;
 wire _1765_;
 wire _1766_;
 wire _1767_;
 wire _1768_;
 wire _1769_;
 wire _1770_;
 wire _1771_;
 wire _1772_;
 wire _1773_;
 wire _1774_;
 wire _1775_;
 wire _1776_;
 wire _1777_;
 wire _1778_;
 wire _1779_;
 wire _1780_;
 wire _1781_;
 wire _1782_;
 wire _1783_;
 wire _1784_;
 wire _1785_;
 wire _1786_;
 wire _1787_;
 wire _1788_;
 wire _1789_;
 wire _1790_;
 wire _1791_;
 wire _1792_;
 wire _1793_;
 wire _1794_;
 wire _1795_;
 wire _1796_;
 wire _1797_;
 wire _1798_;
 wire _1799_;
 wire _1800_;
 wire _1801_;
 wire _1802_;
 wire _1803_;
 wire _1804_;
 wire _1805_;
 wire _1806_;
 wire _1807_;
 wire _1808_;
 wire _1809_;
 wire _1810_;
 wire _1811_;
 wire _1812_;
 wire _1813_;
 wire _1814_;
 wire _1815_;
 wire _1816_;
 wire _1817_;
 wire _1818_;
 wire _1819_;
 wire _1820_;
 wire _1821_;
 wire _1822_;
 wire _1823_;
 wire _1824_;
 wire _1825_;
 wire _1826_;
 wire _1827_;
 wire _1828_;
 wire _1829_;
 wire _1830_;
 wire _1831_;
 wire _1832_;
 wire _1833_;
 wire _1834_;
 wire _1835_;
 wire _1836_;
 wire _1837_;
 wire _1838_;
 wire _1839_;
 wire _1840_;
 wire _1841_;
 wire _1842_;
 wire _1843_;
 wire _1844_;
 wire _1845_;
 wire _1846_;
 wire _1847_;
 wire _1848_;
 wire _1849_;
 wire _1850_;
 wire _1851_;
 wire _1852_;
 wire _1853_;
 wire _1854_;
 wire _1855_;
 wire _1856_;
 wire _1857_;
 wire _1858_;
 wire _1859_;
 wire _1860_;
 wire _1861_;
 wire _1862_;
 wire _1863_;
 wire _1864_;
 wire _1865_;
 wire _1866_;
 wire _1867_;
 wire _1868_;
 wire _1869_;
 wire _1870_;
 wire _1871_;
 wire _1872_;
 wire _1873_;
 wire _1874_;
 wire _1875_;
 wire _1876_;
 wire _1877_;
 wire _1878_;
 wire _1879_;
 wire _1880_;
 wire _1881_;
 wire _1882_;
 wire _1883_;
 wire _1884_;
 wire _1885_;
 wire _1886_;
 wire _1887_;
 wire _1888_;
 wire _1889_;
 wire _1890_;
 wire _1891_;
 wire _1892_;
 wire _1893_;
 wire _1894_;
 wire _1895_;
 wire _1896_;
 wire _1897_;
 wire _1898_;
 wire _1899_;
 wire _1900_;
 wire _1901_;
 wire _1902_;
 wire _1903_;
 wire _1904_;
 wire _1905_;
 wire _1906_;
 wire _1907_;
 wire _1908_;
 wire _1909_;
 wire _1910_;
 wire _1911_;
 wire _1912_;
 wire _1913_;
 wire _1914_;
 wire _1915_;
 wire _1916_;
 wire _1917_;
 wire _1918_;
 wire _1919_;
 wire _1920_;
 wire _1921_;
 wire _1922_;
 wire _1923_;
 wire _1924_;
 wire _1925_;
 wire _1926_;
 wire _1927_;
 wire _1928_;
 wire _1929_;
 wire _1930_;
 wire _1931_;
 wire _1932_;
 wire _1933_;
 wire _1934_;
 wire _1935_;
 wire _1936_;
 wire _1937_;
 wire _1938_;
 wire _1939_;
 wire _1940_;
 wire _1941_;
 wire _1942_;
 wire _1943_;
 wire _1944_;
 wire _1945_;
 wire _1946_;
 wire _1947_;
 wire _1948_;
 wire _1949_;
 wire _1950_;
 wire _1951_;
 wire _1952_;
 wire _1953_;
 wire _1954_;
 wire _1955_;
 wire _1956_;
 wire _1957_;
 wire _1958_;
 wire _1959_;
 wire _1960_;
 wire _1961_;
 wire _1962_;
 wire _1963_;
 wire _1964_;
 wire _1965_;
 wire _1966_;
 wire _1967_;
 wire _1968_;
 wire _1969_;
 wire _1970_;
 wire _1971_;
 wire _1972_;
 wire _1973_;
 wire _1974_;
 wire _1975_;
 wire _1976_;
 wire _1977_;
 wire _1978_;
 wire _1979_;
 wire _1980_;
 wire _1981_;
 wire _1982_;
 wire _1983_;
 wire _1984_;
 wire _1985_;
 wire _1986_;
 wire _1987_;
 wire _1988_;
 wire _1989_;
 wire _1990_;
 wire _1991_;
 wire _1992_;
 wire _1993_;
 wire _1994_;
 wire _1995_;
 wire _1996_;
 wire _1997_;
 wire _1998_;
 wire _1999_;
 wire _2000_;
 wire _2001_;
 wire _2002_;
 wire _2003_;
 wire _2004_;
 wire _2005_;
 wire _2006_;
 wire _2007_;
 wire _2008_;
 wire _2009_;
 wire _2010_;
 wire _2011_;
 wire _2012_;
 wire _2013_;
 wire _2014_;
 wire _2015_;
 wire _2016_;
 wire _2017_;
 wire _2018_;
 wire _2019_;
 wire _2020_;
 wire _2021_;
 wire _2022_;
 wire _2023_;
 wire _2024_;
 wire _2025_;
 wire _2026_;
 wire _2027_;
 wire _2028_;
 wire _2029_;
 wire _2030_;
 wire _2031_;
 wire _2032_;
 wire _2033_;
 wire _2034_;
 wire _2035_;
 wire _2036_;
 wire _2037_;
 wire _2038_;
 wire _2039_;
 wire _2040_;
 wire _2041_;
 wire _2042_;
 wire _2043_;
 wire _2044_;
 wire _2045_;
 wire _2046_;
 wire _2047_;
 wire _2048_;
 wire _2049_;
 wire _2050_;
 wire _2051_;
 wire _2052_;
 wire _2053_;
 wire _2054_;
 wire _2055_;
 wire _2056_;
 wire _2057_;
 wire _2058_;
 wire _2059_;
 wire _2060_;
 wire _2061_;
 wire _2062_;
 wire _2063_;
 wire _2064_;
 wire _2065_;
 wire _2066_;
 wire _2067_;
 wire _2068_;
 wire _2069_;
 wire _2070_;
 wire _2071_;
 wire _2072_;
 wire _2073_;
 wire _2074_;
 wire _2075_;
 wire _2076_;
 wire _2077_;
 wire _2078_;
 wire _2079_;
 wire _2080_;
 wire _2081_;
 wire _2082_;
 wire _2083_;
 wire _2084_;
 wire _2085_;
 wire _2086_;
 wire _2087_;
 wire _2088_;
 wire _2089_;
 wire _2090_;
 wire _2091_;
 wire _2092_;
 wire _2093_;
 wire _2094_;
 wire _2095_;
 wire _2096_;
 wire _2097_;
 wire _2098_;
 wire _2099_;
 wire _2100_;
 wire _2101_;
 wire _2102_;
 wire _2103_;
 wire _2104_;
 wire _2105_;
 wire _2106_;
 wire _2107_;
 wire _2108_;
 wire _2109_;
 wire _2110_;
 wire _2111_;
 wire _2112_;
 wire _2113_;
 wire _2114_;
 wire _2115_;
 wire _2116_;
 wire _2117_;
 wire _2118_;
 wire _2119_;
 wire _2120_;
 wire _2121_;
 wire _2122_;
 wire _2123_;
 wire _2124_;
 wire _2125_;
 wire _2126_;
 wire _2127_;
 wire _2128_;
 wire _2129_;
 wire _2130_;
 wire _2131_;
 wire _2132_;
 wire _2133_;
 wire _2134_;
 wire _2135_;
 wire _2136_;
 wire _2137_;
 wire _2138_;
 wire _2139_;
 wire _2140_;
 wire _2141_;
 wire _2142_;
 wire _2143_;
 wire _2144_;
 wire _2145_;
 wire _2146_;
 wire _2147_;
 wire _2148_;
 wire _2149_;
 wire _2150_;
 wire _2151_;
 wire _2152_;
 wire _2153_;
 wire _2154_;
 wire _2155_;
 wire _2156_;
 wire _2157_;
 wire _2158_;
 wire _2159_;
 wire _2160_;
 wire _2161_;
 wire _2162_;
 wire _2163_;
 wire _2164_;
 wire _2165_;
 wire _2166_;
 wire _2167_;
 wire _2168_;
 wire _2169_;
 wire _2170_;
 wire _2171_;
 wire _2172_;
 wire _2173_;
 wire _2174_;
 wire _2175_;
 wire _2176_;
 wire _2177_;
 wire _2178_;
 wire _2179_;
 wire _2180_;
 wire _2181_;
 wire _2182_;
 wire _2183_;
 wire _2184_;
 wire _2185_;
 wire _2186_;
 wire _2187_;
 wire _2188_;
 wire _2189_;
 wire _2190_;
 wire _2191_;
 wire _2192_;
 wire _2193_;
 wire _2194_;
 wire _2195_;
 wire _2196_;
 wire _2197_;
 wire _2198_;
 wire _2199_;
 wire _2200_;
 wire _2201_;
 wire _2202_;
 wire _2203_;
 wire _2204_;
 wire _2205_;
 wire _2206_;
 wire _2207_;
 wire _2208_;
 wire _2209_;
 wire _2210_;
 wire _2211_;
 wire _2212_;
 wire _2213_;
 wire _2214_;
 wire _2215_;
 wire _2216_;
 wire _2217_;
 wire _2218_;
 wire _2219_;
 wire _2220_;
 wire _2221_;
 wire _2222_;
 wire _2223_;
 wire _2224_;
 wire _2225_;
 wire _2226_;
 wire _2227_;
 wire _2228_;
 wire _2229_;
 wire _2230_;
 wire _2231_;
 wire _2232_;
 wire _2233_;
 wire _2234_;
 wire _2235_;
 wire _2236_;
 wire _2237_;
 wire _2238_;
 wire _2239_;
 wire _2240_;
 wire _2241_;
 wire _2242_;
 wire _2243_;
 wire _2244_;
 wire _2245_;
 wire _2246_;
 wire _2247_;
 wire _2248_;
 wire _2249_;
 wire _2250_;
 wire _2251_;
 wire _2252_;
 wire _2253_;
 wire _2254_;
 wire _2255_;
 wire _2256_;
 wire _2257_;
 wire _2258_;
 wire _2259_;
 wire _2260_;
 wire _2261_;
 wire _2262_;
 wire _2263_;
 wire _2264_;
 wire _2265_;
 wire _2266_;
 wire _2267_;
 wire _2268_;
 wire _2269_;
 wire _2270_;
 wire _2271_;
 wire _2272_;
 wire _2273_;
 wire _2274_;
 wire _2275_;
 wire _2276_;
 wire _2277_;
 wire _2278_;
 wire _2279_;
 wire _2280_;
 wire _2281_;
 wire _2282_;
 wire _2283_;
 wire _2284_;
 wire _2285_;
 wire _2286_;
 wire _2287_;
 wire _2288_;
 wire _2289_;
 wire _2290_;
 wire _2291_;
 wire _2292_;
 wire _2293_;
 wire _2294_;
 wire _2295_;
 wire _2296_;
 wire _2297_;
 wire _2298_;
 wire _2299_;
 wire _2300_;
 wire _2301_;
 wire _2302_;
 wire _2303_;
 wire _2304_;
 wire _2305_;
 wire _2306_;
 wire _2307_;
 wire _2308_;
 wire _2309_;
 wire _2310_;
 wire _2311_;
 wire _2312_;
 wire _2313_;
 wire _2314_;
 wire _2315_;
 wire _2316_;
 wire _2317_;
 wire _2318_;
 wire _2319_;
 wire _2320_;
 wire _2321_;
 wire _2322_;
 wire _2323_;
 wire _2324_;
 wire _2325_;
 wire _2326_;
 wire _2327_;
 wire _2328_;
 wire _2329_;
 wire _2330_;
 wire _2331_;
 wire _2332_;
 wire _2333_;
 wire _2334_;
 wire _2335_;
 wire _2336_;
 wire _2337_;
 wire _2338_;
 wire _2339_;
 wire _2340_;
 wire _2341_;
 wire _2342_;
 wire _2343_;
 wire _2344_;
 wire _2345_;
 wire _2346_;
 wire _2347_;
 wire _2348_;
 wire _2349_;
 wire _2350_;
 wire _2351_;
 wire _2352_;
 wire _2353_;
 wire _2354_;
 wire _2355_;
 wire _2356_;
 wire _2357_;
 wire _2358_;
 wire _2359_;
 wire _2360_;
 wire _2361_;
 wire _2362_;
 wire _2363_;
 wire _2364_;
 wire _2365_;
 wire _2366_;
 wire _2367_;
 wire _2368_;
 wire _2369_;
 wire _2370_;
 wire _2371_;
 wire _2372_;
 wire _2373_;
 wire _2374_;
 wire _2375_;
 wire _2376_;
 wire _2377_;
 wire _2378_;
 wire _2379_;
 wire _2380_;
 wire _2381_;
 wire _2382_;
 wire _2383_;
 wire _2384_;
 wire _2385_;
 wire _2386_;
 wire _2387_;
 wire _2388_;
 wire _2389_;
 wire _2390_;
 wire _2391_;
 wire _2392_;
 wire _2393_;
 wire _2394_;
 wire _2395_;
 wire _2396_;
 wire _2397_;
 wire _2398_;
 wire _2399_;
 wire _2400_;
 wire _2401_;
 wire _2402_;
 wire _2403_;
 wire _2404_;
 wire _2405_;
 wire _2406_;
 wire _2407_;
 wire _2408_;
 wire _2409_;
 wire _2410_;
 wire _2411_;
 wire _2412_;
 wire _2413_;
 wire _2414_;
 wire _2415_;
 wire _2416_;
 wire _2417_;
 wire _2418_;
 wire _2419_;
 wire _2420_;
 wire _2421_;
 wire _2422_;
 wire _2423_;
 wire _2424_;
 wire _2425_;
 wire _2426_;
 wire _2427_;
 wire _2428_;
 wire _2429_;
 wire _2430_;
 wire _2431_;
 wire _2432_;
 wire _2433_;
 wire _2434_;
 wire _2435_;
 wire _2436_;
 wire _2437_;
 wire _2438_;
 wire _2439_;
 wire _2440_;
 wire _2441_;
 wire _2442_;
 wire _2443_;
 wire _2444_;
 wire _2445_;
 wire _2446_;
 wire _2447_;
 wire _2448_;
 wire _2449_;
 wire _2450_;
 wire _2451_;
 wire _2452_;
 wire _2453_;
 wire _2454_;
 wire _2455_;
 wire _2456_;
 wire _2457_;
 wire _2458_;
 wire _2459_;
 wire _2460_;
 wire _2461_;
 wire _2462_;
 wire _2463_;
 wire _2464_;
 wire _2465_;
 wire _2466_;
 wire _2467_;
 wire _2468_;
 wire _2469_;
 wire _2470_;
 wire _2471_;
 wire _2472_;
 wire _2473_;
 wire _2474_;
 wire _2475_;
 wire _2476_;
 wire _2477_;
 wire _2478_;
 wire _2479_;
 wire _2480_;
 wire _2481_;
 wire _2482_;
 wire _2483_;
 wire _2484_;
 wire _2485_;
 wire _2486_;
 wire _2487_;
 wire _2488_;
 wire _2489_;
 wire _2490_;
 wire _2491_;
 wire _2492_;
 wire _2493_;
 wire _2494_;
 wire _2495_;
 wire _2496_;
 wire _2497_;
 wire _2498_;
 wire _2499_;
 wire _2500_;
 wire _2501_;
 wire _2502_;
 wire _2503_;
 wire _2504_;
 wire _2505_;
 wire _2506_;
 wire _2507_;
 wire _2508_;
 wire _2509_;
 wire _2510_;
 wire _2511_;
 wire _2512_;
 wire _2513_;
 wire _2514_;
 wire _2515_;
 wire _2516_;
 wire _2517_;
 wire _2518_;
 wire _2519_;
 wire _2520_;
 wire _2521_;
 wire _2522_;
 wire _2523_;
 wire _2524_;
 wire _2525_;
 wire _2526_;
 wire _2527_;
 wire _2528_;
 wire _2529_;
 wire _2530_;
 wire _2531_;
 wire _2532_;
 wire _2533_;
 wire _2534_;
 wire _2535_;
 wire _2536_;
 wire _2537_;
 wire _2538_;
 wire _2539_;
 wire _2540_;
 wire _2541_;
 wire _2542_;
 wire _2543_;
 wire _2544_;
 wire _2545_;
 wire _2546_;
 wire _2547_;
 wire _2548_;
 wire _2549_;
 wire _2550_;
 wire _2551_;
 wire _2552_;
 wire _2553_;
 wire _2554_;
 wire _2555_;
 wire _2556_;
 wire _2557_;
 wire _2558_;
 wire _2559_;
 wire _2560_;
 wire _2561_;
 wire _2562_;
 wire _2563_;
 wire _2564_;
 wire _2565_;
 wire _2566_;
 wire _2567_;
 wire _2568_;
 wire _2569_;
 wire _2570_;
 wire _2571_;
 wire _2572_;
 wire _2573_;
 wire _2574_;
 wire _2575_;
 wire _2576_;
 wire _2577_;
 wire _2578_;
 wire _2579_;
 wire _2580_;
 wire _2581_;
 wire _2582_;
 wire _2583_;
 wire _2584_;
 wire _2585_;
 wire _2586_;
 wire _2587_;
 wire _2588_;
 wire _2589_;
 wire _2590_;
 wire _2591_;
 wire _2592_;
 wire _2593_;
 wire _2594_;
 wire _2595_;
 wire _2596_;
 wire _2597_;
 wire _2598_;
 wire _2599_;
 wire _2600_;
 wire _2601_;
 wire _2602_;
 wire _2603_;
 wire _2604_;
 wire _2605_;
 wire _2606_;
 wire _2607_;
 wire _2608_;
 wire _2609_;
 wire _2610_;
 wire _2611_;
 wire _2612_;
 wire _2613_;
 wire _2614_;
 wire _2615_;
 wire _2616_;
 wire _2617_;
 wire _2618_;
 wire _2619_;
 wire _2620_;
 wire _2621_;
 wire _2622_;
 wire _2623_;
 wire _2624_;
 wire _2625_;
 wire _2626_;
 wire _2627_;
 wire _2628_;
 wire _2629_;
 wire _2630_;
 wire _2631_;
 wire _2632_;
 wire _2633_;
 wire _2634_;
 wire _2635_;
 wire _2636_;
 wire _2637_;
 wire _2638_;
 wire _2639_;
 wire _2640_;
 wire _2641_;
 wire _2642_;
 wire _2643_;
 wire _2644_;
 wire _2645_;
 wire _2646_;
 wire _2647_;
 wire _2648_;
 wire _2649_;
 wire _2650_;
 wire _2651_;
 wire _2652_;
 wire _2653_;
 wire _2654_;
 wire _2655_;
 wire _2656_;
 wire _2657_;
 wire _2658_;
 wire _2659_;
 wire _2660_;
 wire _2661_;
 wire _2662_;
 wire _2663_;
 wire _2664_;
 wire _2665_;
 wire _2666_;
 wire _2667_;
 wire _2668_;
 wire _2669_;
 wire _2670_;
 wire _2671_;
 wire _2672_;
 wire _2673_;
 wire _2674_;
 wire _2675_;
 wire _2676_;
 wire _2677_;
 wire _2678_;
 wire _2679_;
 wire _2680_;
 wire _2681_;
 wire _2682_;
 wire _2683_;
 wire _2684_;
 wire _2685_;
 wire _2686_;
 wire _2687_;
 wire _2688_;
 wire _2689_;
 wire _2690_;
 wire _2691_;
 wire _2692_;
 wire _2693_;
 wire _2694_;
 wire _2695_;
 wire _2696_;
 wire _2697_;
 wire _2698_;
 wire _2699_;
 wire _2700_;
 wire _2701_;
 wire _2702_;
 wire _2703_;
 wire _2704_;
 wire _2705_;
 wire _2706_;
 wire _2707_;
 wire _2708_;
 wire _2709_;
 wire _2710_;
 wire _2711_;
 wire _2712_;
 wire _2713_;
 wire _2714_;
 wire _2715_;
 wire _2716_;
 wire _2717_;
 wire _2718_;
 wire _2719_;
 wire _2720_;
 wire _2721_;
 wire _2722_;
 wire _2723_;
 wire _2724_;
 wire _2725_;
 wire _2726_;
 wire _2727_;
 wire _2728_;
 wire _2729_;
 wire _2730_;
 wire _2731_;
 wire _2732_;
 wire _2733_;
 wire _2734_;
 wire _2735_;
 wire _2736_;
 wire _2737_;
 wire _2738_;
 wire _2739_;
 wire _2740_;
 wire _2741_;
 wire _2742_;
 wire _2743_;
 wire _2744_;
 wire _2745_;
 wire _2746_;
 wire _2747_;
 wire _2748_;
 wire _2749_;
 wire _2750_;
 wire _2751_;
 wire _2752_;
 wire _2753_;
 wire _2754_;
 wire _2755_;
 wire _2756_;
 wire _2757_;
 wire _2758_;
 wire _2759_;
 wire _2760_;
 wire _2761_;
 wire _2762_;
 wire _2763_;
 wire _2764_;
 wire _2765_;
 wire _2766_;
 wire _2767_;
 wire _2768_;
 wire _2769_;
 wire _2770_;
 wire _2771_;
 wire _2772_;
 wire _2773_;
 wire _2774_;
 wire _2775_;
 wire _2776_;
 wire _2777_;
 wire _2778_;
 wire _2779_;
 wire _2780_;
 wire _2781_;
 wire _2782_;
 wire _2783_;
 wire _2784_;
 wire _2785_;
 wire _2786_;
 wire _2787_;
 wire _2788_;
 wire _2789_;
 wire _2790_;
 wire _2791_;
 wire _2792_;
 wire _2793_;
 wire _2794_;
 wire _2795_;
 wire _2796_;
 wire _2797_;
 wire _2798_;
 wire _2799_;
 wire _2800_;
 wire _2801_;
 wire _2802_;
 wire _2803_;
 wire _2804_;
 wire _2805_;
 wire _2806_;
 wire _2807_;
 wire _2808_;
 wire _2809_;
 wire _2810_;
 wire _2811_;
 wire _2812_;
 wire _2813_;
 wire _2814_;
 wire _2815_;
 wire _2816_;
 wire _2817_;
 wire _2818_;
 wire _2819_;
 wire _2820_;
 wire _2821_;
 wire _2822_;
 wire _2823_;
 wire _2824_;
 wire _2825_;
 wire _2826_;
 wire _2827_;
 wire _2828_;
 wire _2829_;
 wire _2830_;
 wire _2831_;
 wire _2832_;
 wire _2833_;
 wire _2834_;
 wire _2835_;
 wire _2836_;
 wire _2837_;
 wire _2838_;
 wire _2839_;
 wire _2840_;
 wire _2841_;
 wire _2842_;
 wire _2843_;
 wire _2844_;
 wire _2845_;
 wire _2846_;
 wire _2847_;
 wire _2848_;
 wire _2849_;
 wire _2850_;
 wire _2851_;
 wire _2852_;
 wire _2853_;
 wire _2854_;
 wire _2855_;
 wire _2856_;
 wire _2857_;
 wire _2858_;
 wire _2859_;
 wire _2860_;
 wire _2861_;
 wire _2862_;
 wire _2863_;
 wire _2864_;
 wire _2865_;
 wire _2866_;
 wire _2867_;
 wire _2868_;
 wire _2869_;
 wire _2870_;
 wire _2871_;
 wire _2872_;
 wire _2873_;
 wire _2874_;
 wire _2875_;
 wire _2876_;
 wire _2877_;
 wire _2878_;
 wire _2879_;
 wire _2880_;
 wire _2881_;
 wire _2882_;
 wire _2883_;
 wire _2884_;
 wire _2885_;
 wire _2886_;
 wire _2887_;
 wire _2888_;
 wire _2889_;
 wire _2890_;
 wire _2891_;
 wire _2892_;
 wire _2893_;
 wire _2894_;
 wire _2895_;
 wire _2896_;
 wire _2897_;
 wire _2898_;
 wire _2899_;
 wire _2900_;
 wire _2901_;
 wire _2902_;
 wire _2903_;
 wire _2904_;
 wire _2905_;
 wire _2906_;
 wire _2907_;
 wire _2908_;
 wire _2909_;
 wire _2910_;
 wire _2911_;
 wire _2912_;
 wire _2913_;
 wire _2914_;
 wire _2915_;
 wire _2916_;
 wire _2917_;
 wire _2918_;
 wire _2919_;
 wire _2920_;
 wire _2921_;
 wire _2922_;
 wire _2923_;
 wire _2924_;
 wire _2925_;
 wire _2926_;
 wire _2927_;
 wire _2928_;
 wire _2929_;
 wire _2930_;
 wire _2931_;
 wire _2932_;
 wire _2933_;
 wire _2934_;
 wire _2935_;
 wire _2936_;
 wire _2937_;
 wire _2938_;
 wire _2939_;
 wire _2940_;
 wire _2941_;
 wire _2942_;
 wire _2943_;
 wire _2944_;
 wire _2945_;
 wire _2946_;
 wire _2947_;
 wire _2948_;
 wire _2949_;
 wire _2950_;
 wire _2951_;
 wire _2952_;
 wire _2953_;
 wire _2954_;
 wire _2955_;
 wire _2956_;
 wire _2957_;
 wire _2958_;
 wire _2959_;
 wire _2960_;
 wire _2961_;
 wire _2962_;
 wire _2963_;
 wire _2964_;
 wire _2965_;
 wire _2966_;
 wire _2967_;
 wire _2968_;
 wire _2969_;
 wire _2970_;
 wire _2971_;
 wire _2972_;
 wire _2973_;
 wire _2974_;
 wire _2975_;
 wire _2976_;
 wire _2977_;
 wire _2978_;
 wire _2979_;
 wire _2980_;
 wire _2981_;
 wire _2982_;
 wire _2983_;
 wire _2984_;
 wire _2985_;
 wire _2986_;
 wire _2987_;
 wire _2988_;
 wire _2989_;
 wire _2990_;
 wire _2991_;
 wire _2992_;
 wire _2993_;
 wire _2994_;
 wire _2995_;
 wire _2996_;
 wire _2997_;
 wire _2998_;
 wire _2999_;
 wire _3000_;
 wire _3001_;
 wire _3002_;
 wire _3003_;
 wire _3004_;
 wire _3005_;
 wire _3006_;
 wire _3007_;
 wire _3008_;
 wire _3009_;
 wire _3010_;
 wire _3011_;
 wire _3012_;
 wire _3013_;
 wire _3014_;
 wire _3015_;
 wire _3016_;
 wire _3017_;
 wire _3018_;
 wire _3019_;
 wire _3020_;
 wire _3021_;
 wire _3022_;
 wire _3023_;
 wire _3024_;
 wire _3025_;
 wire _3026_;
 wire _3027_;
 wire _3028_;
 wire _3029_;
 wire _3030_;
 wire _3031_;
 wire _3032_;
 wire _3033_;
 wire _3034_;
 wire _3035_;
 wire _3036_;
 wire _3037_;
 wire _3038_;
 wire _3039_;
 wire _3040_;
 wire _3041_;
 wire _3042_;
 wire _3043_;
 wire _3044_;
 wire _3045_;
 wire _3046_;
 wire _3047_;
 wire _3048_;
 wire _3049_;
 wire _3050_;
 wire _3051_;
 wire _3052_;
 wire _3053_;
 wire _3054_;
 wire _3055_;
 wire _3056_;
 wire _3057_;
 wire _3058_;
 wire _3059_;
 wire _3060_;
 wire _3061_;
 wire _3062_;
 wire _3063_;
 wire _3064_;
 wire _3065_;
 wire _3066_;
 wire _3067_;
 wire _3068_;
 wire _3069_;
 wire _3070_;
 wire _3071_;
 wire _3072_;
 wire _3073_;
 wire _3074_;
 wire _3075_;
 wire _3076_;
 wire _3077_;
 wire _3078_;
 wire _3079_;
 wire _3080_;
 wire _3081_;
 wire _3082_;
 wire _3083_;
 wire _3084_;
 wire _3085_;
 wire _3086_;
 wire _3087_;
 wire _3088_;
 wire _3089_;
 wire _3090_;
 wire _3091_;
 wire _3092_;
 wire _3093_;
 wire _3094_;
 wire _3095_;
 wire _3096_;
 wire _3097_;
 wire _3098_;
 wire _3099_;
 wire _3100_;
 wire _3101_;
 wire _3102_;
 wire _3103_;
 wire _3104_;
 wire _3105_;
 wire _3106_;
 wire _3107_;
 wire _3108_;
 wire _3109_;
 wire _3110_;
 wire _3111_;
 wire _3112_;
 wire _3113_;
 wire _3114_;
 wire _3115_;
 wire _3116_;
 wire _3117_;
 wire _3118_;
 wire _3119_;
 wire _3120_;
 wire _3121_;
 wire _3122_;
 wire _3123_;
 wire _3124_;
 wire _3125_;
 wire _3126_;
 wire _3127_;
 wire _3128_;
 wire _3129_;
 wire _3130_;
 wire _3131_;
 wire _3132_;
 wire _3133_;
 wire _3134_;
 wire _3135_;
 wire _3136_;
 wire _3137_;
 wire _3138_;
 wire _3139_;
 wire _3140_;
 wire _3141_;
 wire _3142_;
 wire _3143_;
 wire _3144_;
 wire _3145_;
 wire _3146_;
 wire _3147_;
 wire _3148_;
 wire _3149_;
 wire _3150_;
 wire _3151_;
 wire _3152_;
 wire _3153_;
 wire _3154_;
 wire _3155_;
 wire _3156_;
 wire _3157_;
 wire _3158_;
 wire _3159_;
 wire _3160_;
 wire _3161_;
 wire _3162_;
 wire _3163_;
 wire _3164_;
 wire _3165_;
 wire _3166_;
 wire _3167_;
 wire _3168_;
 wire _3169_;
 wire _3170_;
 wire _3171_;
 wire _3172_;
 wire _3173_;
 wire _3174_;
 wire _3175_;
 wire _3176_;
 wire _3177_;
 wire _3178_;
 wire _3179_;
 wire _3180_;
 wire _3181_;
 wire _3182_;
 wire _3183_;
 wire _3184_;
 wire _3185_;
 wire _3186_;
 wire _3187_;
 wire _3188_;
 wire _3189_;
 wire _3190_;
 wire _3191_;
 wire _3192_;
 wire _3193_;
 wire _3194_;
 wire _3195_;
 wire _3196_;
 wire _3197_;
 wire _3198_;
 wire _3199_;
 wire _3200_;
 wire _3201_;
 wire _3202_;
 wire _3203_;
 wire _3204_;
 wire _3205_;
 wire _3206_;
 wire _3207_;
 wire _3208_;
 wire _3209_;
 wire _3210_;
 wire _3211_;
 wire _3212_;
 wire _3213_;
 wire _3214_;
 wire _3215_;
 wire _3216_;
 wire _3217_;
 wire _3218_;
 wire _3219_;
 wire _3220_;
 wire _3221_;
 wire _3222_;
 wire _3223_;
 wire _3224_;
 wire _3225_;
 wire _3226_;
 wire _3227_;
 wire _3228_;
 wire _3229_;
 wire _3230_;
 wire _3231_;
 wire _3232_;
 wire _3233_;
 wire _3234_;
 wire _3235_;
 wire _3236_;
 wire _3237_;
 wire _3238_;
 wire _3239_;
 wire _3240_;
 wire _3241_;
 wire _3242_;
 wire _3243_;
 wire _3244_;
 wire _3245_;
 wire _3246_;
 wire _3247_;
 wire _3248_;
 wire _3249_;
 wire _3250_;
 wire _3251_;
 wire _3252_;
 wire _3253_;
 wire _3254_;
 wire _3255_;
 wire _3256_;
 wire _3257_;
 wire _3258_;
 wire _3259_;
 wire _3260_;
 wire _3261_;
 wire _3262_;
 wire _3263_;
 wire _3264_;
 wire _3265_;
 wire _3266_;
 wire _3267_;
 wire _3268_;
 wire _3269_;
 wire _3270_;
 wire _3271_;
 wire _3272_;
 wire _3273_;
 wire _3274_;
 wire _3275_;
 wire _3276_;
 wire _3277_;
 wire _3278_;
 wire _3279_;
 wire _3280_;
 wire _3281_;
 wire _3282_;
 wire _3283_;
 wire _3284_;
 wire _3285_;
 wire _3286_;
 wire _3287_;
 wire _3288_;
 wire _3289_;
 wire _3290_;
 wire _3291_;
 wire _3292_;
 wire _3293_;
 wire _3294_;
 wire _3295_;
 wire _3296_;
 wire _3297_;
 wire _3298_;
 wire _3299_;
 wire _3300_;
 wire _3301_;
 wire _3302_;
 wire _3303_;
 wire _3304_;
 wire _3305_;
 wire _3306_;
 wire _3307_;
 wire _3308_;
 wire _3309_;
 wire _3310_;
 wire _3311_;
 wire _3312_;
 wire _3313_;
 wire _3314_;
 wire _3315_;
 wire _3316_;
 wire _3317_;
 wire _3318_;
 wire _3319_;
 wire _3320_;
 wire _3321_;
 wire _3322_;
 wire _3323_;
 wire _3324_;
 wire _3325_;
 wire _3326_;
 wire _3327_;
 wire _3328_;
 wire _3329_;
 wire _3330_;
 wire _3331_;
 wire _3332_;
 wire _3333_;
 wire _3334_;
 wire _3335_;
 wire _3336_;
 wire _3337_;
 wire _3338_;
 wire _3339_;
 wire _3340_;
 wire _3341_;
 wire _3342_;
 wire _3343_;
 wire _3344_;
 wire _3345_;
 wire _3346_;
 wire _3347_;
 wire _3348_;
 wire _3349_;
 wire _3350_;
 wire _3351_;
 wire _3352_;
 wire _3353_;
 wire _3354_;
 wire _3355_;
 wire _3356_;
 wire _3357_;
 wire _3358_;
 wire _3359_;
 wire _3360_;
 wire _3361_;
 wire _3362_;
 wire _3363_;
 wire _3364_;
 wire _3365_;
 wire _3366_;
 wire _3367_;
 wire _3368_;
 wire _3369_;
 wire _3370_;
 wire _3371_;
 wire _3372_;
 wire _3373_;
 wire _3374_;
 wire _3375_;
 wire _3376_;
 wire _3377_;
 wire _3378_;
 wire _3379_;
 wire _3380_;
 wire _3381_;
 wire _3382_;
 wire _3383_;
 wire _3384_;
 wire _3385_;
 wire _3386_;
 wire _3387_;
 wire _3388_;
 wire _3389_;
 wire _3390_;
 wire _3391_;
 wire _3392_;
 wire _3393_;
 wire _3394_;
 wire _3395_;
 wire _3396_;
 wire _3397_;
 wire _3398_;
 wire _3399_;
 wire _3400_;
 wire _3401_;
 wire _3402_;
 wire _3403_;
 wire _3404_;
 wire _3405_;
 wire _3406_;
 wire _3407_;
 wire _3408_;
 wire _3409_;
 wire _3410_;
 wire _3411_;
 wire _3412_;
 wire _3413_;
 wire _3414_;
 wire _3415_;
 wire _3416_;
 wire _3417_;
 wire _3418_;
 wire _3419_;
 wire _3420_;
 wire _3421_;
 wire _3422_;
 wire _3423_;
 wire _3424_;
 wire _3425_;
 wire _3426_;
 wire _3427_;
 wire _3428_;
 wire _3429_;
 wire _3430_;
 wire _3431_;
 wire _3432_;
 wire _3433_;
 wire _3434_;
 wire _3435_;
 wire _3436_;
 wire _3437_;
 wire _3438_;
 wire _3439_;
 wire _3440_;
 wire _3441_;
 wire _3442_;
 wire _3443_;
 wire _3444_;
 wire _3445_;
 wire _3446_;
 wire _3447_;
 wire _3448_;
 wire _3449_;
 wire _3450_;
 wire _3451_;
 wire _3452_;
 wire _3453_;
 wire _3454_;
 wire _3455_;
 wire _3456_;
 wire _3457_;
 wire _3458_;
 wire _3459_;
 wire _3460_;
 wire _3461_;
 wire _3462_;
 wire _3463_;
 wire _3464_;
 wire _3465_;
 wire _3466_;
 wire _3467_;
 wire _3468_;
 wire _3469_;
 wire _3470_;
 wire _3471_;
 wire _3472_;
 wire _3473_;
 wire _3474_;
 wire _3475_;
 wire _3476_;
 wire _3477_;
 wire _3478_;
 wire _3479_;
 wire _3480_;
 wire _3481_;
 wire _3482_;
 wire _3483_;
 wire _3484_;
 wire _3485_;
 wire _3486_;
 wire _3487_;
 wire _3488_;
 wire _3489_;
 wire _3490_;
 wire _3491_;
 wire _3492_;
 wire _3493_;
 wire _3494_;
 wire _3495_;
 wire _3496_;
 wire _3497_;
 wire _3498_;
 wire _3499_;
 wire _3500_;
 wire _3501_;
 wire _3502_;
 wire _3503_;
 wire _3504_;
 wire _3505_;
 wire _3506_;
 wire _3507_;
 wire _3508_;
 wire _3509_;
 wire _3510_;
 wire _3511_;
 wire _3512_;
 wire _3513_;
 wire _3514_;
 wire _3515_;
 wire _3516_;
 wire _3517_;
 wire _3518_;
 wire _3519_;
 wire _3520_;
 wire _3521_;
 wire _3522_;
 wire _3523_;
 wire _3524_;
 wire _3525_;
 wire _3526_;
 wire _3527_;
 wire _3528_;
 wire _3529_;
 wire _3530_;
 wire _3531_;
 wire _3532_;
 wire _3533_;
 wire _3534_;
 wire _3535_;
 wire _3536_;
 wire _3537_;
 wire _3538_;
 wire _3539_;
 wire _3540_;
 wire _3541_;
 wire _3542_;
 wire _3543_;
 wire _3544_;
 wire _3545_;
 wire _3546_;
 wire _3547_;
 wire _3548_;
 wire _3549_;
 wire _3550_;
 wire _3551_;
 wire _3552_;
 wire _3553_;
 wire _3554_;
 wire _3555_;
 wire _3556_;
 wire _3557_;
 wire _3558_;
 wire _3559_;
 wire _3560_;
 wire _3561_;
 wire _3562_;
 wire _3563_;
 wire _3564_;
 wire _3565_;
 wire _3566_;
 wire _3567_;
 wire _3568_;
 wire _3569_;
 wire _3570_;
 wire _3571_;
 wire _3572_;
 wire _3573_;
 wire _3574_;
 wire _3575_;
 wire _3576_;
 wire _3577_;
 wire _3578_;
 wire _3579_;
 wire _3580_;
 wire _3581_;
 wire _3582_;
 wire _3583_;
 wire _3584_;
 wire _3585_;
 wire _3586_;
 wire _3587_;
 wire _3588_;
 wire _3589_;
 wire _3590_;
 wire _3591_;
 wire _3592_;
 wire _3593_;
 wire _3594_;
 wire _3595_;
 wire _3596_;
 wire _3597_;
 wire _3598_;
 wire _3599_;
 wire _3600_;
 wire _3601_;
 wire _3602_;
 wire _3603_;
 wire _3604_;
 wire _3605_;
 wire _3606_;
 wire _3607_;
 wire _3608_;
 wire _3609_;
 wire _3610_;
 wire _3611_;
 wire _3612_;
 wire _3613_;
 wire _3614_;
 wire _3615_;
 wire _3616_;
 wire _3617_;
 wire _3618_;
 wire _3619_;
 wire _3620_;
 wire _3621_;
 wire _3622_;
 wire _3623_;
 wire _3624_;
 wire _3625_;
 wire _3626_;
 wire _3627_;
 wire _3628_;
 wire _3629_;
 wire _3630_;
 wire _3631_;
 wire _3632_;
 wire _3633_;
 wire _3634_;
 wire _3635_;
 wire _3636_;
 wire _3637_;
 wire _3638_;
 wire _3639_;
 wire _3640_;
 wire _3641_;
 wire _3642_;
 wire _3643_;
 wire _3644_;
 wire _3645_;
 wire _3646_;
 wire _3647_;
 wire _3648_;
 wire _3649_;
 wire _3650_;
 wire _3651_;
 wire _3652_;
 wire _3653_;
 wire _3654_;
 wire _3655_;
 wire _3656_;
 wire _3657_;
 wire _3658_;
 wire _3659_;
 wire _3660_;
 wire _3661_;
 wire _3662_;
 wire _3663_;
 wire _3664_;
 wire _3665_;
 wire _3666_;
 wire _3667_;
 wire _3668_;
 wire _3669_;
 wire _3670_;
 wire _3671_;
 wire _3672_;
 wire _3673_;
 wire _3674_;
 wire _3675_;
 wire _3676_;
 wire _3677_;
 wire _3678_;
 wire _3679_;
 wire _3680_;
 wire _3681_;
 wire _3682_;
 wire _3683_;
 wire _3684_;
 wire _3685_;
 wire _3686_;
 wire _3687_;
 wire _3688_;
 wire _3689_;
 wire _3690_;
 wire _3691_;
 wire _3692_;
 wire _3693_;
 wire _3694_;
 wire _3695_;
 wire _3696_;
 wire _3697_;
 wire _3698_;
 wire _3699_;
 wire _3700_;
 wire _3701_;
 wire _3702_;
 wire _3703_;
 wire _3704_;
 wire _3705_;
 wire _3706_;
 wire _3707_;
 wire _3708_;
 wire _3709_;
 wire _3710_;
 wire _3711_;
 wire _3712_;
 wire _3713_;
 wire _3714_;
 wire _3715_;
 wire _3716_;
 wire _3717_;
 wire _3718_;
 wire _3719_;
 wire _3720_;
 wire _3721_;
 wire _3722_;
 wire _3723_;
 wire _3724_;
 wire _3725_;
 wire _3726_;
 wire _3727_;
 wire _3728_;
 wire _3729_;
 wire _3730_;
 wire _3731_;
 wire _3732_;
 wire _3733_;
 wire _3734_;
 wire _3735_;
 wire _3736_;
 wire _3737_;
 wire _3738_;
 wire _3739_;
 wire _3740_;
 wire _3741_;
 wire _3742_;
 wire _3743_;
 wire _3744_;
 wire _3745_;
 wire _3746_;
 wire _3747_;
 wire _3748_;
 wire _3749_;
 wire _3750_;
 wire _3751_;
 wire _3752_;
 wire _3753_;
 wire _3754_;
 wire _3755_;
 wire _3756_;
 wire \inputcont.INTERNAL_MODE ;
 wire \inputcont.INTERNAL_OCTAVE_INPUT ;
 wire \inputcont.INTERNAL_SYNCED_I[0] ;
 wire \inputcont.INTERNAL_SYNCED_I[10] ;
 wire \inputcont.INTERNAL_SYNCED_I[11] ;
 wire \inputcont.INTERNAL_SYNCED_I[12] ;
 wire \inputcont.INTERNAL_SYNCED_I[1] ;
 wire \inputcont.INTERNAL_SYNCED_I[2] ;
 wire \inputcont.INTERNAL_SYNCED_I[3] ;
 wire \inputcont.INTERNAL_SYNCED_I[4] ;
 wire \inputcont.INTERNAL_SYNCED_I[5] ;
 wire \inputcont.INTERNAL_SYNCED_I[6] ;
 wire \inputcont.INTERNAL_SYNCED_I[7] ;
 wire \inputcont.INTERNAL_SYNCED_I[8] ;
 wire \inputcont.INTERNAL_SYNCED_I[9] ;
 wire \inputcont.u1.ff_intermediate[0] ;
 wire \inputcont.u1.ff_intermediate[10] ;
 wire \inputcont.u1.ff_intermediate[11] ;
 wire \inputcont.u1.ff_intermediate[12] ;
 wire \inputcont.u1.ff_intermediate[13] ;
 wire \inputcont.u1.ff_intermediate[14] ;
 wire \inputcont.u1.ff_intermediate[1] ;
 wire \inputcont.u1.ff_intermediate[2] ;
 wire \inputcont.u1.ff_intermediate[3] ;
 wire \inputcont.u1.ff_intermediate[4] ;
 wire \inputcont.u1.ff_intermediate[5] ;
 wire \inputcont.u1.ff_intermediate[6] ;
 wire \inputcont.u1.ff_intermediate[7] ;
 wire \inputcont.u1.ff_intermediate[8] ;
 wire \inputcont.u1.ff_intermediate[9] ;
 wire \inputcont.u2.next_in ;
 wire \inputcont.u3.next_in ;
 wire net1;
 wire net10;
 wire net100;
 wire net101;
 wire net102;
 wire net103;
 wire net104;
 wire net105;
 wire net106;
 wire net107;
 wire net108;
 wire net109;
 wire net11;
 wire net110;
 wire net111;
 wire net112;
 wire net113;
 wire net114;
 wire net115;
 wire net116;
 wire net117;
 wire net118;
 wire net119;
 wire net12;
 wire net120;
 wire net121;
 wire net122;
 wire net123;
 wire net124;
 wire net125;
 wire net126;
 wire net127;
 wire net128;
 wire net129;
 wire net13;
 wire net130;
 wire net131;
 wire net132;
 wire net133;
 wire net134;
 wire net135;
 wire net136;
 wire net137;
 wire net138;
 wire net139;
 wire net14;
 wire net140;
 wire net141;
 wire net142;
 wire net143;
 wire net144;
 wire net145;
 wire net147;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net88;
 wire net89;
 wire net9;
 wire net90;
 wire net91;
 wire net92;
 wire net93;
 wire net94;
 wire net95;
 wire net96;
 wire net97;
 wire net98;
 wire net99;
 wire \oct.next_state[0] ;
 wire \oct.next_state[1] ;
 wire \oct.next_state[2] ;
 wire \oct.state[0] ;
 wire \oct.state[1] ;
 wire \oct.state[2] ;
 wire \pm.count[0] ;
 wire \pm.count[1] ;
 wire \pm.count[2] ;
 wire \pm.count[3] ;
 wire \pm.count[4] ;
 wire \pm.count[5] ;
 wire \pm.count[6] ;
 wire \pm.count[7] ;
 wire \pm.count[8] ;
 wire \pm.current_waveform[0] ;
 wire \pm.current_waveform[1] ;
 wire \pm.current_waveform[2] ;
 wire \pm.current_waveform[3] ;
 wire \pm.current_waveform[4] ;
 wire \pm.current_waveform[5] ;
 wire \pm.current_waveform[6] ;
 wire \pm.current_waveform[7] ;
 wire \pm.current_waveform[8] ;
 wire \pm.next_count[0] ;
 wire \pm.next_count[1] ;
 wire \pm.next_count[2] ;
 wire \pm.next_count[3] ;
 wire \pm.next_count[4] ;
 wire \pm.next_count[5] ;
 wire \pm.next_count[6] ;
 wire \pm.next_count[7] ;
 wire \pm.next_count[8] ;
 wire \pm.next_pwm_o ;
 wire \pm.pwm_o ;
 wire \rate_clk.count[0] ;
 wire \rate_clk.count[1] ;
 wire \rate_clk.count[2] ;
 wire \rate_clk.count[3] ;
 wire \rate_clk.count[4] ;
 wire \rate_clk.count[5] ;
 wire \rate_clk.count[6] ;
 wire \rate_clk.count[7] ;
 wire \rate_clk.next_count[0] ;
 wire \rate_clk.next_count[1] ;
 wire \rate_clk.next_count[2] ;
 wire \rate_clk.next_count[3] ;
 wire \rate_clk.next_count[4] ;
 wire \rate_clk.next_count[5] ;
 wire \rate_clk.next_count[6] ;
 wire \rate_clk.next_count[7] ;
 wire \select1.sequencer_on ;
 wire \seq.beat[0] ;
 wire \seq.beat[1] ;
 wire \seq.beat[2] ;
 wire \seq.beat[3] ;
 wire \seq.clk_div.count[0] ;
 wire \seq.clk_div.count[10] ;
 wire \seq.clk_div.count[11] ;
 wire \seq.clk_div.count[12] ;
 wire \seq.clk_div.count[13] ;
 wire \seq.clk_div.count[14] ;
 wire \seq.clk_div.count[15] ;
 wire \seq.clk_div.count[16] ;
 wire \seq.clk_div.count[17] ;
 wire \seq.clk_div.count[18] ;
 wire \seq.clk_div.count[19] ;
 wire \seq.clk_div.count[1] ;
 wire \seq.clk_div.count[20] ;
 wire \seq.clk_div.count[21] ;
 wire \seq.clk_div.count[2] ;
 wire \seq.clk_div.count[3] ;
 wire \seq.clk_div.count[4] ;
 wire \seq.clk_div.count[5] ;
 wire \seq.clk_div.count[6] ;
 wire \seq.clk_div.count[7] ;
 wire \seq.clk_div.count[8] ;
 wire \seq.clk_div.count[9] ;
 wire \seq.clk_div.next_count[0] ;
 wire \seq.clk_div.next_count[10] ;
 wire \seq.clk_div.next_count[11] ;
 wire \seq.clk_div.next_count[12] ;
 wire \seq.clk_div.next_count[13] ;
 wire \seq.clk_div.next_count[14] ;
 wire \seq.clk_div.next_count[15] ;
 wire \seq.clk_div.next_count[16] ;
 wire \seq.clk_div.next_count[17] ;
 wire \seq.clk_div.next_count[18] ;
 wire \seq.clk_div.next_count[19] ;
 wire \seq.clk_div.next_count[1] ;
 wire \seq.clk_div.next_count[20] ;
 wire \seq.clk_div.next_count[21] ;
 wire \seq.clk_div.next_count[2] ;
 wire \seq.clk_div.next_count[3] ;
 wire \seq.clk_div.next_count[4] ;
 wire \seq.clk_div.next_count[5] ;
 wire \seq.clk_div.next_count[6] ;
 wire \seq.clk_div.next_count[7] ;
 wire \seq.clk_div.next_count[8] ;
 wire \seq.clk_div.next_count[9] ;
 wire \seq.encode.inter_keys[0] ;
 wire \seq.encode.inter_keys[10] ;
 wire \seq.encode.inter_keys[1] ;
 wire \seq.encode.keys_edge_det[0] ;
 wire \seq.encode.keys_edge_det[10] ;
 wire \seq.encode.keys_edge_det[1] ;
 wire \seq.encode.keys_edge_det[2] ;
 wire \seq.encode.keys_edge_det[3] ;
 wire \seq.encode.keys_edge_det[4] ;
 wire \seq.encode.keys_edge_det[5] ;
 wire \seq.encode.keys_edge_det[6] ;
 wire \seq.encode.keys_edge_det[7] ;
 wire \seq.encode.keys_edge_det[8] ;
 wire \seq.encode.keys_edge_det[9] ;
 wire \seq.encode.keys_sync[0] ;
 wire \seq.encode.keys_sync[10] ;
 wire \seq.encode.keys_sync[1] ;
 wire \seq.encode.next_play ;
 wire \seq.encode.next_sequencer_on ;
 wire \seq.encode.play ;
 wire \seq.player_1.next_state[0] ;
 wire \seq.player_1.next_state[1] ;
 wire \seq.player_1.next_state[2] ;
 wire \seq.player_1.next_state[3] ;
 wire \seq.player_1.state[0] ;
 wire \seq.player_1.state[1] ;
 wire \seq.player_1.state[2] ;
 wire \seq.player_1.state[3] ;
 wire \seq.player_2.next_state[0] ;
 wire \seq.player_2.next_state[1] ;
 wire \seq.player_2.next_state[2] ;
 wire \seq.player_2.next_state[3] ;
 wire \seq.player_2.state[0] ;
 wire \seq.player_2.state[1] ;
 wire \seq.player_2.state[2] ;
 wire \seq.player_2.state[3] ;
 wire \seq.player_3.next_state[0] ;
 wire \seq.player_3.next_state[1] ;
 wire \seq.player_3.next_state[2] ;
 wire \seq.player_3.next_state[3] ;
 wire \seq.player_3.state[0] ;
 wire \seq.player_3.state[1] ;
 wire \seq.player_3.state[2] ;
 wire \seq.player_3.state[3] ;
 wire \seq.player_4.next_state[0] ;
 wire \seq.player_4.next_state[1] ;
 wire \seq.player_4.next_state[2] ;
 wire \seq.player_4.next_state[3] ;
 wire \seq.player_4.state[0] ;
 wire \seq.player_4.state[1] ;
 wire \seq.player_4.state[2] ;
 wire \seq.player_4.state[3] ;
 wire \seq.player_5.next_state[0] ;
 wire \seq.player_5.next_state[1] ;
 wire \seq.player_5.next_state[2] ;
 wire \seq.player_5.next_state[3] ;
 wire \seq.player_5.state[0] ;
 wire \seq.player_5.state[1] ;
 wire \seq.player_5.state[2] ;
 wire \seq.player_5.state[3] ;
 wire \seq.player_6.next_state[0] ;
 wire \seq.player_6.next_state[1] ;
 wire \seq.player_6.next_state[2] ;
 wire \seq.player_6.next_state[3] ;
 wire \seq.player_6.state[0] ;
 wire \seq.player_6.state[1] ;
 wire \seq.player_6.state[2] ;
 wire \seq.player_6.state[3] ;
 wire \seq.player_7.next_state[0] ;
 wire \seq.player_7.next_state[1] ;
 wire \seq.player_7.next_state[2] ;
 wire \seq.player_7.next_state[3] ;
 wire \seq.player_7.state[0] ;
 wire \seq.player_7.state[1] ;
 wire \seq.player_7.state[2] ;
 wire \seq.player_7.state[3] ;
 wire \seq.player_8.next_state[0] ;
 wire \seq.player_8.next_state[1] ;
 wire \seq.player_8.next_state[2] ;
 wire \seq.player_8.next_state[3] ;
 wire \seq.player_8.state[0] ;
 wire \seq.player_8.state[1] ;
 wire \seq.player_8.state[2] ;
 wire \seq.player_8.state[3] ;
 wire \seq.tempo_select.next_state[0] ;
 wire \seq.tempo_select.next_state[1] ;
 wire \seq.tempo_select.state[0] ;
 wire \seq.tempo_select.state[1] ;
 wire seq_play_on;
 wire seq_power_on;
 wire \sound1.count[0] ;
 wire \sound1.count[10] ;
 wire \sound1.count[11] ;
 wire \sound1.count[12] ;
 wire \sound1.count[13] ;
 wire \sound1.count[14] ;
 wire \sound1.count[15] ;
 wire \sound1.count[16] ;
 wire \sound1.count[17] ;
 wire \sound1.count[18] ;
 wire \sound1.count[1] ;
 wire \sound1.count[2] ;
 wire \sound1.count[3] ;
 wire \sound1.count[4] ;
 wire \sound1.count[5] ;
 wire \sound1.count[6] ;
 wire \sound1.count[7] ;
 wire \sound1.count[8] ;
 wire \sound1.count[9] ;
 wire \sound1.count_m[0] ;
 wire \sound1.count_m[10] ;
 wire \sound1.count_m[11] ;
 wire \sound1.count_m[12] ;
 wire \sound1.count_m[13] ;
 wire \sound1.count_m[14] ;
 wire \sound1.count_m[15] ;
 wire \sound1.count_m[16] ;
 wire \sound1.count_m[17] ;
 wire \sound1.count_m[18] ;
 wire \sound1.count_m[1] ;
 wire \sound1.count_m[2] ;
 wire \sound1.count_m[3] ;
 wire \sound1.count_m[4] ;
 wire \sound1.count_m[5] ;
 wire \sound1.count_m[6] ;
 wire \sound1.count_m[7] ;
 wire \sound1.count_m[8] ;
 wire \sound1.count_m[9] ;
 wire \sound1.divisor_m[0] ;
 wire \sound1.divisor_m[10] ;
 wire \sound1.divisor_m[11] ;
 wire \sound1.divisor_m[12] ;
 wire \sound1.divisor_m[13] ;
 wire \sound1.divisor_m[14] ;
 wire \sound1.divisor_m[15] ;
 wire \sound1.divisor_m[16] ;
 wire \sound1.divisor_m[17] ;
 wire \sound1.divisor_m[18] ;
 wire \sound1.divisor_m[1] ;
 wire \sound1.divisor_m[2] ;
 wire \sound1.divisor_m[3] ;
 wire \sound1.divisor_m[4] ;
 wire \sound1.divisor_m[5] ;
 wire \sound1.divisor_m[6] ;
 wire \sound1.divisor_m[7] ;
 wire \sound1.divisor_m[8] ;
 wire \sound1.divisor_m[9] ;
 wire \sound1.osc.next_count[0] ;
 wire \sound1.osc.next_count[10] ;
 wire \sound1.osc.next_count[11] ;
 wire \sound1.osc.next_count[12] ;
 wire \sound1.osc.next_count[13] ;
 wire \sound1.osc.next_count[14] ;
 wire \sound1.osc.next_count[15] ;
 wire \sound1.osc.next_count[16] ;
 wire \sound1.osc.next_count[17] ;
 wire \sound1.osc.next_count[18] ;
 wire \sound1.osc.next_count[1] ;
 wire \sound1.osc.next_count[2] ;
 wire \sound1.osc.next_count[3] ;
 wire \sound1.osc.next_count[4] ;
 wire \sound1.osc.next_count[5] ;
 wire \sound1.osc.next_count[6] ;
 wire \sound1.osc.next_count[7] ;
 wire \sound1.osc.next_count[8] ;
 wire \sound1.osc.next_count[9] ;
 wire \sound1.sdiv.A[0] ;
 wire \sound1.sdiv.A[10] ;
 wire \sound1.sdiv.A[11] ;
 wire \sound1.sdiv.A[12] ;
 wire \sound1.sdiv.A[13] ;
 wire \sound1.sdiv.A[14] ;
 wire \sound1.sdiv.A[15] ;
 wire \sound1.sdiv.A[16] ;
 wire \sound1.sdiv.A[17] ;
 wire \sound1.sdiv.A[18] ;
 wire \sound1.sdiv.A[19] ;
 wire \sound1.sdiv.A[1] ;
 wire \sound1.sdiv.A[20] ;
 wire \sound1.sdiv.A[21] ;
 wire \sound1.sdiv.A[22] ;
 wire \sound1.sdiv.A[23] ;
 wire \sound1.sdiv.A[24] ;
 wire \sound1.sdiv.A[25] ;
 wire \sound1.sdiv.A[26] ;
 wire \sound1.sdiv.A[2] ;
 wire \sound1.sdiv.A[3] ;
 wire \sound1.sdiv.A[4] ;
 wire \sound1.sdiv.A[5] ;
 wire \sound1.sdiv.A[6] ;
 wire \sound1.sdiv.A[7] ;
 wire \sound1.sdiv.A[8] ;
 wire \sound1.sdiv.A[9] ;
 wire \sound1.sdiv.C[0] ;
 wire \sound1.sdiv.C[1] ;
 wire \sound1.sdiv.C[2] ;
 wire \sound1.sdiv.C[3] ;
 wire \sound1.sdiv.C[4] ;
 wire \sound1.sdiv.C[5] ;
 wire \sound1.sdiv.Q[0] ;
 wire \sound1.sdiv.Q[10] ;
 wire \sound1.sdiv.Q[11] ;
 wire \sound1.sdiv.Q[12] ;
 wire \sound1.sdiv.Q[13] ;
 wire \sound1.sdiv.Q[14] ;
 wire \sound1.sdiv.Q[15] ;
 wire \sound1.sdiv.Q[16] ;
 wire \sound1.sdiv.Q[17] ;
 wire \sound1.sdiv.Q[18] ;
 wire \sound1.sdiv.Q[19] ;
 wire \sound1.sdiv.Q[1] ;
 wire \sound1.sdiv.Q[20] ;
 wire \sound1.sdiv.Q[21] ;
 wire \sound1.sdiv.Q[22] ;
 wire \sound1.sdiv.Q[23] ;
 wire \sound1.sdiv.Q[24] ;
 wire \sound1.sdiv.Q[25] ;
 wire \sound1.sdiv.Q[26] ;
 wire \sound1.sdiv.Q[27] ;
 wire \sound1.sdiv.Q[2] ;
 wire \sound1.sdiv.Q[3] ;
 wire \sound1.sdiv.Q[4] ;
 wire \sound1.sdiv.Q[5] ;
 wire \sound1.sdiv.Q[6] ;
 wire \sound1.sdiv.Q[7] ;
 wire \sound1.sdiv.Q[8] ;
 wire \sound1.sdiv.Q[9] ;
 wire \sound1.sdiv.dived ;
 wire \sound1.sdiv.next_dived ;
 wire \sound1.sdiv.next_start ;
 wire \sound1.sdiv.start ;
 wire \sound2.count[0] ;
 wire \sound2.count[10] ;
 wire \sound2.count[11] ;
 wire \sound2.count[12] ;
 wire \sound2.count[13] ;
 wire \sound2.count[14] ;
 wire \sound2.count[15] ;
 wire \sound2.count[16] ;
 wire \sound2.count[17] ;
 wire \sound2.count[18] ;
 wire \sound2.count[1] ;
 wire \sound2.count[2] ;
 wire \sound2.count[3] ;
 wire \sound2.count[4] ;
 wire \sound2.count[5] ;
 wire \sound2.count[6] ;
 wire \sound2.count[7] ;
 wire \sound2.count[8] ;
 wire \sound2.count[9] ;
 wire \sound2.count_m[0] ;
 wire \sound2.count_m[10] ;
 wire \sound2.count_m[11] ;
 wire \sound2.count_m[12] ;
 wire \sound2.count_m[13] ;
 wire \sound2.count_m[14] ;
 wire \sound2.count_m[15] ;
 wire \sound2.count_m[16] ;
 wire \sound2.count_m[17] ;
 wire \sound2.count_m[18] ;
 wire \sound2.count_m[1] ;
 wire \sound2.count_m[2] ;
 wire \sound2.count_m[3] ;
 wire \sound2.count_m[4] ;
 wire \sound2.count_m[5] ;
 wire \sound2.count_m[6] ;
 wire \sound2.count_m[7] ;
 wire \sound2.count_m[8] ;
 wire \sound2.count_m[9] ;
 wire \sound2.divisor_m[0] ;
 wire \sound2.divisor_m[10] ;
 wire \sound2.divisor_m[11] ;
 wire \sound2.divisor_m[12] ;
 wire \sound2.divisor_m[13] ;
 wire \sound2.divisor_m[14] ;
 wire \sound2.divisor_m[15] ;
 wire \sound2.divisor_m[16] ;
 wire \sound2.divisor_m[17] ;
 wire \sound2.divisor_m[18] ;
 wire \sound2.divisor_m[1] ;
 wire \sound2.divisor_m[2] ;
 wire \sound2.divisor_m[3] ;
 wire \sound2.divisor_m[4] ;
 wire \sound2.divisor_m[5] ;
 wire \sound2.divisor_m[6] ;
 wire \sound2.divisor_m[7] ;
 wire \sound2.divisor_m[8] ;
 wire \sound2.divisor_m[9] ;
 wire \sound2.osc.next_count[0] ;
 wire \sound2.osc.next_count[10] ;
 wire \sound2.osc.next_count[11] ;
 wire \sound2.osc.next_count[12] ;
 wire \sound2.osc.next_count[13] ;
 wire \sound2.osc.next_count[14] ;
 wire \sound2.osc.next_count[15] ;
 wire \sound2.osc.next_count[16] ;
 wire \sound2.osc.next_count[17] ;
 wire \sound2.osc.next_count[18] ;
 wire \sound2.osc.next_count[1] ;
 wire \sound2.osc.next_count[2] ;
 wire \sound2.osc.next_count[3] ;
 wire \sound2.osc.next_count[4] ;
 wire \sound2.osc.next_count[5] ;
 wire \sound2.osc.next_count[6] ;
 wire \sound2.osc.next_count[7] ;
 wire \sound2.osc.next_count[8] ;
 wire \sound2.osc.next_count[9] ;
 wire \sound2.sdiv.A[0] ;
 wire \sound2.sdiv.A[10] ;
 wire \sound2.sdiv.A[11] ;
 wire \sound2.sdiv.A[12] ;
 wire \sound2.sdiv.A[13] ;
 wire \sound2.sdiv.A[14] ;
 wire \sound2.sdiv.A[15] ;
 wire \sound2.sdiv.A[16] ;
 wire \sound2.sdiv.A[17] ;
 wire \sound2.sdiv.A[18] ;
 wire \sound2.sdiv.A[19] ;
 wire \sound2.sdiv.A[1] ;
 wire \sound2.sdiv.A[20] ;
 wire \sound2.sdiv.A[21] ;
 wire \sound2.sdiv.A[22] ;
 wire \sound2.sdiv.A[23] ;
 wire \sound2.sdiv.A[24] ;
 wire \sound2.sdiv.A[25] ;
 wire \sound2.sdiv.A[26] ;
 wire \sound2.sdiv.A[2] ;
 wire \sound2.sdiv.A[3] ;
 wire \sound2.sdiv.A[4] ;
 wire \sound2.sdiv.A[5] ;
 wire \sound2.sdiv.A[6] ;
 wire \sound2.sdiv.A[7] ;
 wire \sound2.sdiv.A[8] ;
 wire \sound2.sdiv.A[9] ;
 wire \sound2.sdiv.C[0] ;
 wire \sound2.sdiv.C[1] ;
 wire \sound2.sdiv.C[2] ;
 wire \sound2.sdiv.C[3] ;
 wire \sound2.sdiv.C[4] ;
 wire \sound2.sdiv.C[5] ;
 wire \sound2.sdiv.Q[0] ;
 wire \sound2.sdiv.Q[10] ;
 wire \sound2.sdiv.Q[11] ;
 wire \sound2.sdiv.Q[12] ;
 wire \sound2.sdiv.Q[13] ;
 wire \sound2.sdiv.Q[14] ;
 wire \sound2.sdiv.Q[15] ;
 wire \sound2.sdiv.Q[16] ;
 wire \sound2.sdiv.Q[17] ;
 wire \sound2.sdiv.Q[18] ;
 wire \sound2.sdiv.Q[19] ;
 wire \sound2.sdiv.Q[1] ;
 wire \sound2.sdiv.Q[20] ;
 wire \sound2.sdiv.Q[21] ;
 wire \sound2.sdiv.Q[22] ;
 wire \sound2.sdiv.Q[23] ;
 wire \sound2.sdiv.Q[24] ;
 wire \sound2.sdiv.Q[25] ;
 wire \sound2.sdiv.Q[26] ;
 wire \sound2.sdiv.Q[27] ;
 wire \sound2.sdiv.Q[2] ;
 wire \sound2.sdiv.Q[3] ;
 wire \sound2.sdiv.Q[4] ;
 wire \sound2.sdiv.Q[5] ;
 wire \sound2.sdiv.Q[6] ;
 wire \sound2.sdiv.Q[7] ;
 wire \sound2.sdiv.Q[8] ;
 wire \sound2.sdiv.Q[9] ;
 wire \sound2.sdiv.dived ;
 wire \sound2.sdiv.next_dived ;
 wire \sound2.sdiv.next_start ;
 wire \sound2.sdiv.start ;
 wire \sound3.count[0] ;
 wire \sound3.count[10] ;
 wire \sound3.count[11] ;
 wire \sound3.count[12] ;
 wire \sound3.count[13] ;
 wire \sound3.count[14] ;
 wire \sound3.count[15] ;
 wire \sound3.count[16] ;
 wire \sound3.count[17] ;
 wire \sound3.count[18] ;
 wire \sound3.count[1] ;
 wire \sound3.count[2] ;
 wire \sound3.count[3] ;
 wire \sound3.count[4] ;
 wire \sound3.count[5] ;
 wire \sound3.count[6] ;
 wire \sound3.count[7] ;
 wire \sound3.count[8] ;
 wire \sound3.count[9] ;
 wire \sound3.count_m[0] ;
 wire \sound3.count_m[10] ;
 wire \sound3.count_m[11] ;
 wire \sound3.count_m[12] ;
 wire \sound3.count_m[13] ;
 wire \sound3.count_m[14] ;
 wire \sound3.count_m[15] ;
 wire \sound3.count_m[16] ;
 wire \sound3.count_m[17] ;
 wire \sound3.count_m[18] ;
 wire \sound3.count_m[1] ;
 wire \sound3.count_m[2] ;
 wire \sound3.count_m[3] ;
 wire \sound3.count_m[4] ;
 wire \sound3.count_m[5] ;
 wire \sound3.count_m[6] ;
 wire \sound3.count_m[7] ;
 wire \sound3.count_m[8] ;
 wire \sound3.count_m[9] ;
 wire \sound3.divisor_m[0] ;
 wire \sound3.divisor_m[10] ;
 wire \sound3.divisor_m[11] ;
 wire \sound3.divisor_m[12] ;
 wire \sound3.divisor_m[13] ;
 wire \sound3.divisor_m[14] ;
 wire \sound3.divisor_m[15] ;
 wire \sound3.divisor_m[16] ;
 wire \sound3.divisor_m[17] ;
 wire \sound3.divisor_m[18] ;
 wire \sound3.divisor_m[1] ;
 wire \sound3.divisor_m[2] ;
 wire \sound3.divisor_m[3] ;
 wire \sound3.divisor_m[4] ;
 wire \sound3.divisor_m[5] ;
 wire \sound3.divisor_m[6] ;
 wire \sound3.divisor_m[7] ;
 wire \sound3.divisor_m[8] ;
 wire \sound3.divisor_m[9] ;
 wire \sound3.osc.next_count[0] ;
 wire \sound3.osc.next_count[10] ;
 wire \sound3.osc.next_count[11] ;
 wire \sound3.osc.next_count[12] ;
 wire \sound3.osc.next_count[13] ;
 wire \sound3.osc.next_count[14] ;
 wire \sound3.osc.next_count[15] ;
 wire \sound3.osc.next_count[16] ;
 wire \sound3.osc.next_count[17] ;
 wire \sound3.osc.next_count[18] ;
 wire \sound3.osc.next_count[1] ;
 wire \sound3.osc.next_count[2] ;
 wire \sound3.osc.next_count[3] ;
 wire \sound3.osc.next_count[4] ;
 wire \sound3.osc.next_count[5] ;
 wire \sound3.osc.next_count[6] ;
 wire \sound3.osc.next_count[7] ;
 wire \sound3.osc.next_count[8] ;
 wire \sound3.osc.next_count[9] ;
 wire \sound3.sdiv.A[0] ;
 wire \sound3.sdiv.A[10] ;
 wire \sound3.sdiv.A[11] ;
 wire \sound3.sdiv.A[12] ;
 wire \sound3.sdiv.A[13] ;
 wire \sound3.sdiv.A[14] ;
 wire \sound3.sdiv.A[15] ;
 wire \sound3.sdiv.A[16] ;
 wire \sound3.sdiv.A[17] ;
 wire \sound3.sdiv.A[18] ;
 wire \sound3.sdiv.A[19] ;
 wire \sound3.sdiv.A[1] ;
 wire \sound3.sdiv.A[20] ;
 wire \sound3.sdiv.A[21] ;
 wire \sound3.sdiv.A[22] ;
 wire \sound3.sdiv.A[23] ;
 wire \sound3.sdiv.A[24] ;
 wire \sound3.sdiv.A[25] ;
 wire \sound3.sdiv.A[26] ;
 wire \sound3.sdiv.A[2] ;
 wire \sound3.sdiv.A[3] ;
 wire \sound3.sdiv.A[4] ;
 wire \sound3.sdiv.A[5] ;
 wire \sound3.sdiv.A[6] ;
 wire \sound3.sdiv.A[7] ;
 wire \sound3.sdiv.A[8] ;
 wire \sound3.sdiv.A[9] ;
 wire \sound3.sdiv.C[0] ;
 wire \sound3.sdiv.C[1] ;
 wire \sound3.sdiv.C[2] ;
 wire \sound3.sdiv.C[3] ;
 wire \sound3.sdiv.C[4] ;
 wire \sound3.sdiv.C[5] ;
 wire \sound3.sdiv.Q[0] ;
 wire \sound3.sdiv.Q[10] ;
 wire \sound3.sdiv.Q[11] ;
 wire \sound3.sdiv.Q[12] ;
 wire \sound3.sdiv.Q[13] ;
 wire \sound3.sdiv.Q[14] ;
 wire \sound3.sdiv.Q[15] ;
 wire \sound3.sdiv.Q[16] ;
 wire \sound3.sdiv.Q[17] ;
 wire \sound3.sdiv.Q[18] ;
 wire \sound3.sdiv.Q[19] ;
 wire \sound3.sdiv.Q[1] ;
 wire \sound3.sdiv.Q[20] ;
 wire \sound3.sdiv.Q[21] ;
 wire \sound3.sdiv.Q[22] ;
 wire \sound3.sdiv.Q[23] ;
 wire \sound3.sdiv.Q[24] ;
 wire \sound3.sdiv.Q[25] ;
 wire \sound3.sdiv.Q[26] ;
 wire \sound3.sdiv.Q[27] ;
 wire \sound3.sdiv.Q[2] ;
 wire \sound3.sdiv.Q[3] ;
 wire \sound3.sdiv.Q[4] ;
 wire \sound3.sdiv.Q[5] ;
 wire \sound3.sdiv.Q[6] ;
 wire \sound3.sdiv.Q[7] ;
 wire \sound3.sdiv.Q[8] ;
 wire \sound3.sdiv.Q[9] ;
 wire \sound3.sdiv.dived ;
 wire \sound3.sdiv.next_dived ;
 wire \sound3.sdiv.next_start ;
 wire \sound3.sdiv.start ;
 wire \sound4.count[0] ;
 wire \sound4.count[10] ;
 wire \sound4.count[11] ;
 wire \sound4.count[12] ;
 wire \sound4.count[13] ;
 wire \sound4.count[14] ;
 wire \sound4.count[15] ;
 wire \sound4.count[16] ;
 wire \sound4.count[17] ;
 wire \sound4.count[18] ;
 wire \sound4.count[1] ;
 wire \sound4.count[2] ;
 wire \sound4.count[3] ;
 wire \sound4.count[4] ;
 wire \sound4.count[5] ;
 wire \sound4.count[6] ;
 wire \sound4.count[7] ;
 wire \sound4.count[8] ;
 wire \sound4.count[9] ;
 wire \sound4.count_m[0] ;
 wire \sound4.count_m[10] ;
 wire \sound4.count_m[11] ;
 wire \sound4.count_m[12] ;
 wire \sound4.count_m[13] ;
 wire \sound4.count_m[14] ;
 wire \sound4.count_m[15] ;
 wire \sound4.count_m[16] ;
 wire \sound4.count_m[17] ;
 wire \sound4.count_m[18] ;
 wire \sound4.count_m[1] ;
 wire \sound4.count_m[2] ;
 wire \sound4.count_m[3] ;
 wire \sound4.count_m[4] ;
 wire \sound4.count_m[5] ;
 wire \sound4.count_m[6] ;
 wire \sound4.count_m[7] ;
 wire \sound4.count_m[8] ;
 wire \sound4.count_m[9] ;
 wire \sound4.divisor_m[0] ;
 wire \sound4.divisor_m[10] ;
 wire \sound4.divisor_m[11] ;
 wire \sound4.divisor_m[12] ;
 wire \sound4.divisor_m[13] ;
 wire \sound4.divisor_m[14] ;
 wire \sound4.divisor_m[15] ;
 wire \sound4.divisor_m[16] ;
 wire \sound4.divisor_m[17] ;
 wire \sound4.divisor_m[18] ;
 wire \sound4.divisor_m[1] ;
 wire \sound4.divisor_m[2] ;
 wire \sound4.divisor_m[3] ;
 wire \sound4.divisor_m[4] ;
 wire \sound4.divisor_m[5] ;
 wire \sound4.divisor_m[6] ;
 wire \sound4.divisor_m[7] ;
 wire \sound4.divisor_m[8] ;
 wire \sound4.divisor_m[9] ;
 wire \sound4.osc.next_count[0] ;
 wire \sound4.osc.next_count[10] ;
 wire \sound4.osc.next_count[11] ;
 wire \sound4.osc.next_count[12] ;
 wire \sound4.osc.next_count[13] ;
 wire \sound4.osc.next_count[14] ;
 wire \sound4.osc.next_count[15] ;
 wire \sound4.osc.next_count[16] ;
 wire \sound4.osc.next_count[17] ;
 wire \sound4.osc.next_count[18] ;
 wire \sound4.osc.next_count[1] ;
 wire \sound4.osc.next_count[2] ;
 wire \sound4.osc.next_count[3] ;
 wire \sound4.osc.next_count[4] ;
 wire \sound4.osc.next_count[5] ;
 wire \sound4.osc.next_count[6] ;
 wire \sound4.osc.next_count[7] ;
 wire \sound4.osc.next_count[8] ;
 wire \sound4.osc.next_count[9] ;
 wire \sound4.sdiv.A[0] ;
 wire \sound4.sdiv.A[10] ;
 wire \sound4.sdiv.A[11] ;
 wire \sound4.sdiv.A[12] ;
 wire \sound4.sdiv.A[13] ;
 wire \sound4.sdiv.A[14] ;
 wire \sound4.sdiv.A[15] ;
 wire \sound4.sdiv.A[16] ;
 wire \sound4.sdiv.A[17] ;
 wire \sound4.sdiv.A[18] ;
 wire \sound4.sdiv.A[19] ;
 wire \sound4.sdiv.A[1] ;
 wire \sound4.sdiv.A[20] ;
 wire \sound4.sdiv.A[21] ;
 wire \sound4.sdiv.A[22] ;
 wire \sound4.sdiv.A[23] ;
 wire \sound4.sdiv.A[24] ;
 wire \sound4.sdiv.A[25] ;
 wire \sound4.sdiv.A[26] ;
 wire \sound4.sdiv.A[2] ;
 wire \sound4.sdiv.A[3] ;
 wire \sound4.sdiv.A[4] ;
 wire \sound4.sdiv.A[5] ;
 wire \sound4.sdiv.A[6] ;
 wire \sound4.sdiv.A[7] ;
 wire \sound4.sdiv.A[8] ;
 wire \sound4.sdiv.A[9] ;
 wire \sound4.sdiv.C[0] ;
 wire \sound4.sdiv.C[1] ;
 wire \sound4.sdiv.C[2] ;
 wire \sound4.sdiv.C[3] ;
 wire \sound4.sdiv.C[4] ;
 wire \sound4.sdiv.C[5] ;
 wire \sound4.sdiv.Q[0] ;
 wire \sound4.sdiv.Q[10] ;
 wire \sound4.sdiv.Q[11] ;
 wire \sound4.sdiv.Q[12] ;
 wire \sound4.sdiv.Q[13] ;
 wire \sound4.sdiv.Q[14] ;
 wire \sound4.sdiv.Q[15] ;
 wire \sound4.sdiv.Q[16] ;
 wire \sound4.sdiv.Q[17] ;
 wire \sound4.sdiv.Q[18] ;
 wire \sound4.sdiv.Q[19] ;
 wire \sound4.sdiv.Q[1] ;
 wire \sound4.sdiv.Q[20] ;
 wire \sound4.sdiv.Q[21] ;
 wire \sound4.sdiv.Q[22] ;
 wire \sound4.sdiv.Q[23] ;
 wire \sound4.sdiv.Q[24] ;
 wire \sound4.sdiv.Q[25] ;
 wire \sound4.sdiv.Q[26] ;
 wire \sound4.sdiv.Q[27] ;
 wire \sound4.sdiv.Q[2] ;
 wire \sound4.sdiv.Q[3] ;
 wire \sound4.sdiv.Q[4] ;
 wire \sound4.sdiv.Q[5] ;
 wire \sound4.sdiv.Q[6] ;
 wire \sound4.sdiv.Q[7] ;
 wire \sound4.sdiv.Q[8] ;
 wire \sound4.sdiv.Q[9] ;
 wire \sound4.sdiv.dived ;
 wire \sound4.sdiv.next_dived ;
 wire \sound4.sdiv.next_start ;
 wire \sound4.sdiv.start ;
 wire tempo_select_on;
 wire \wave.mode[0] ;
 wire \wave.mode[1] ;
 wire \wave.next_state[0] ;
 wire \wave.next_state[1] ;
 wire \wave_comb.u1.A[0] ;
 wire \wave_comb.u1.A[10] ;
 wire \wave_comb.u1.A[1] ;
 wire \wave_comb.u1.A[2] ;
 wire \wave_comb.u1.A[3] ;
 wire \wave_comb.u1.A[4] ;
 wire \wave_comb.u1.A[5] ;
 wire \wave_comb.u1.A[6] ;
 wire \wave_comb.u1.A[7] ;
 wire \wave_comb.u1.A[8] ;
 wire \wave_comb.u1.A[9] ;
 wire \wave_comb.u1.C[0] ;
 wire \wave_comb.u1.C[1] ;
 wire \wave_comb.u1.C[2] ;
 wire \wave_comb.u1.C[3] ;
 wire \wave_comb.u1.C[4] ;
 wire \wave_comb.u1.C[5] ;
 wire \wave_comb.u1.M[0] ;
 wire \wave_comb.u1.M[1] ;
 wire \wave_comb.u1.M[2] ;
 wire \wave_comb.u1.Q[0] ;
 wire \wave_comb.u1.Q[10] ;
 wire \wave_comb.u1.Q[11] ;
 wire \wave_comb.u1.Q[1] ;
 wire \wave_comb.u1.Q[2] ;
 wire \wave_comb.u1.Q[3] ;
 wire \wave_comb.u1.Q[4] ;
 wire \wave_comb.u1.Q[5] ;
 wire \wave_comb.u1.Q[6] ;
 wire \wave_comb.u1.Q[7] ;
 wire \wave_comb.u1.Q[8] ;
 wire \wave_comb.u1.Q[9] ;
 wire \wave_comb.u1.dived ;
 wire \wave_comb.u1.next_dived ;
 wire \wave_comb.u1.next_start ;
 wire \wave_comb.u1.start ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_1111_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(net41));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(net44));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(net58));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(\inputcont.u1.ff_intermediate[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(\inputcont.u1.ff_intermediate[10] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(\inputcont.u1.ff_intermediate[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(\inputcont.u1.ff_intermediate[1] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(\inputcont.u1.ff_intermediate[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(\inputcont.u1.ff_intermediate[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(\inputcont.u1.ff_intermediate[9] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(\inputcont.u1.ff_intermediate[9] ));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_298 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_765 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_241 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_307 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_322 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_396 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_416 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_643 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_100_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_706 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_100_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_100 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_106 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_244 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_35 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_355 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_401 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_418 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_422 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_503 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_549 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_577 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_61 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_647 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_653 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_101_687 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_723 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_101_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_101 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_136 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_175 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_220 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_244 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_289 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_338 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_350 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_433 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_459 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_603 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_708 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_720 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_116 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_128 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_140 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_188 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_228 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_243 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_378 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_391 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_404 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_458 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_656 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_693 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_103_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_103_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_73 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_738 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_103_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_103_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_204 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_212 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_403 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_566 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_602 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_614 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_674 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_71 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_104_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_154 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_187 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_374 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_386 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_411 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_105_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_686 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_707 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_105_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_329 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_352 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_434 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_521 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_576 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_616 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_675 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_690 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_106_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_725 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_133 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_173 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_182 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_218 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_301 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_343 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_510 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_534 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_543 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_551 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_107_682 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_107_89 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_98 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_118 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_271 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_530 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_108_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_568 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_576 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_596 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_618 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_666 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_678 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_690 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_108_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_85 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_216 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_319 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_368 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_492 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_505 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_561 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_608 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_680 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_109_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_109_96 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_115 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_172 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_321 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_377 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_10_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_424 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_448 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_472 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_486 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_10_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_110 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_125 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_188 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_210 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_256 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_327 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_331 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_395 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_399 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_468 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_477 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_621 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_110_628 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_633 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_654 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_675 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_110_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_110_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_110_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_108 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_221 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_254 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_315 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_402 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_452 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_463 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_525 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_584 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_111_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_670 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_111_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_111_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_771 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_172 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_273 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_112_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_361 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_371 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_395 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_444 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_459 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_627 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_635 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_322 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_359 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_461 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_493 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_557 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_670 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_113_676 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_113_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_113_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_114 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_122 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_312 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_507 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_527 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_567 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_649 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_653 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_665 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_114_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_114_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_136 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_184 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_407 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_538 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_610 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_626 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_634 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_115_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_115_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_115_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_109 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_117 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_339 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_351 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_433 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_459 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_116_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_116_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_116_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_116_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_460 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_535 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_117_642 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_117_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_307 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_385 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_414 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_432 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_444 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_545 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_118_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_118_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_13 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_25 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_261 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_293 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_317 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_37 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_373 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_479 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_49 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_119_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_552 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_124 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_156 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_181 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_193 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_264 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_372 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_411 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_476 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_11 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_341 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_417 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_487 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_515 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_556 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_564 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_120_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_761 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_120_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_337 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_490 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_552 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_121_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_578 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_121_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_338 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_353 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_379 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_450 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_122_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_551 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_563 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_122_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_354 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_366 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_372 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_380 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_455 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_486 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_123_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_123_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_577 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_123_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_177 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_346 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_562 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_582 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_611 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_124_635 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_124_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_125_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_125_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_358 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_438 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_460 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_495 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_499 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_126_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_556 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_126_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_341 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_353 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_357 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_416 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_447 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_487 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_495 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_127_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_532 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_127_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_610 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_127_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_155 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_190 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_345 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_483 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_543 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_563 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_568 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_574 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_128_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_728 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_740 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_128_752 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_128_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_129_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_457 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_469 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_129_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_129_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_129_770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_186 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_204 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_216 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_324 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_336 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_418 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_421 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_12_453 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_12_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_12_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_289 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_301 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_44 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_517 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_531 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_537 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_651 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_697 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_718 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_753 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_762 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_130_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_130_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_151 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_179 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_301 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_349 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_493 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_13_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_172 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_194 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_201 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_14_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_326 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_433 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_14_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_493 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_509 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_14_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_123 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_135 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_162 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_214 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_284 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_357 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_458 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_494 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_15_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_579 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_151 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_195 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_206 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_259 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_264 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_276 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_303 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_307 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_325 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_16_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_475 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_525 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_570 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_574 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_599 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_16_634 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_16_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_108 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_145 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_166 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_173 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_179 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_257 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_269 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_277 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_423 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_494 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_509 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_600 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_612 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_17_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_96 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_107 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_119 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_394 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_442 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_474 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_492 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_504 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_18_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_553 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_570 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_63 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_18_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_18_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_131 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_143 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_176 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_188 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_293 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_330 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_348 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_501 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_19_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_650 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_662 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_19_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_709 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_71 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_174 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_182 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_206 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_257 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_396 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_408 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_430 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_462 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_1_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_530 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_534 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_559 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_1_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_753 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_1_765 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_102 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_157 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_213 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_20_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_389 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_432 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_444 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_468 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_20_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_508 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_581 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_618 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_665 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_20_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_136 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_390 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_407 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_415 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_446 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_46 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_502 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_21_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_21_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_685 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_73 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_156 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_317 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_328 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_341 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_37 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_452 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_513 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_524 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_551 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_22_563 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_573 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_586 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_22_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_713 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_22_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_116 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_143 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_278 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_316 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_328 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_405 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_420 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_456 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_464 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_484 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_493 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_503 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_629 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_23_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_661 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_75 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_82 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_23_94 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_107 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_197 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_209 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_265 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_389 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_428 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_515 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_549 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_553 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_565 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_24_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_593 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_614 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_757 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_82 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_140 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_164 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_179 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_202 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_263 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_431 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_443 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_447 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_458 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_25_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_485 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_497 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_520 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_573 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_659 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_765 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_164 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_220 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_232 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_251 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_260 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_287 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_347 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_373 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_395 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_450 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_489 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_500 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_530 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_630 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_26_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_26_769 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_26_90 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_98 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_147 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_152 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_185 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_215 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_302 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_314 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_33 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_331 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_357 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_473 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_27_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_321 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_360 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_397 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_490 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_630 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_757 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_28_76 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_28_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_108 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_132 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_186 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_198 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_210 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_223 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_233 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_264 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_417 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_445 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_455 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_492 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_585 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_596 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_604 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_765 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_29_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_121 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_129 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_134 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_158 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_304 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_323 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_359 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_374 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_2_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_455 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_468 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_491 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_521 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_2_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_108 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_128 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_235 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_386 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_398 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_419 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_469 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_522 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_553 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_602 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_638 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_30_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_30_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_160 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_175 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_213 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_266 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_291 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_299 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_346 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_350 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_374 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_386 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_409 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_469 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_481 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_509 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_552 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_637 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_708 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_720 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_735 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_31_738 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_80 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_94 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_186 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_194 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_215 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_223 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_454 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_496 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_508 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_587 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_607 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_615 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_32_640 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_82 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_100 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_118 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_126 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_182 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_190 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_220 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_265 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_33_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_35 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_406 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_411 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_465 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_526 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_639 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_647 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_33_670 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_702 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_714 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_79 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_104 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_114 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_152 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_170 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_274 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_283 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_342 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_34_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_566 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_599 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_621 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_627 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_34_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_687 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_707 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_34_714 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_91 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_207 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_247 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_308 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_429 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_461 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_48 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_525 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_589 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_615 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_66 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_671 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_683 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_687 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_701 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_35_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_741 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_751 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_35_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_87 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_159 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_171 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_188 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_224 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_283 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_321 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_351 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_38 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_473 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_536 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_542 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_568 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_36_610 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_617 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_745 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_36_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_95 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_144 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_194 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_332 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_354 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_376 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_388 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_432 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_438 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_467 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_487 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_511 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_37_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_569 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_590 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_600 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_689 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_708 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_756 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_76 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_760 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_95 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_122 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_128 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_231 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_244 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_285 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_402 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_414 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_429 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_470 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_488 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_524 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_545 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_563 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_60 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_612 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_624 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_656 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_38_679 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_745 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_38_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_103 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_120 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_149 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_166 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_188 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_196 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_239 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_257 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_305 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_317 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_323 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_349 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_436 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_490 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_498 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_505 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_537 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_549 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_593 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_640 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_656 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_660 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_703 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_727 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_746 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_139 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_155 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_162 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_187 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_401 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_407 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_411 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_3_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_480 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_487 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_3_502 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_525 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_3_534 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_195 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_212 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_277 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_342 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_352 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_391 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_403 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_462 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_474 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_490 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_518 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_531 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_536 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_587 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_593 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_614 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_620 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_648 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_662 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_677 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_40_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_85 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_119 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_199 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_237 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_286 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_316 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_335 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_341 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_381 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_404 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_416 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_424 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_440 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_465 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_483 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_559 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_567 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_574 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_598 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_610 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_634 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_41_642 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_647 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_716 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_41_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_120 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_132 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_166 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_174 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_193 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_206 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_239 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_292 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_309 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_336 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_356 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_378 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_436 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_481 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_495 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_52 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_546 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_564 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_595 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_60 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_616 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_623 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_633 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_66 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_42_665 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_685 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_694 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_710 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_714 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_737 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_749 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_42_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_96 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_150 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_176 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_193 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_207 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_305 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_334 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_413 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_441 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_465 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_534 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_596 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_624 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_648 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_43_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_660 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_678 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_693 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_717 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_43_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_742 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_751 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_763 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_771 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_127 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_173 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_181 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_185 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_208 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_277 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_317 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_347 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_355 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_379 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_445 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_467 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_481 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_488 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_500 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_508 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_537 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_543 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_642 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_67 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_44_698 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_705 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_44_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_744 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_757 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_183 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_211 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_247 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_401 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_532 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_625 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_129 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_235 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_251 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_307 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_334 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_340 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_348 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_399 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_424 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_494 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_506 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_518 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_527 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_531 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_616 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_46_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_677 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_724 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_736 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_46_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_11 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_142 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_154 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_207 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_214 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_222 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_254 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_293 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_317 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_370 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_388 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_415 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_427 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_458 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_479 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_483 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_495 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_511 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_519 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_597 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_612 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_652 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_664 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_709 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_768 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_103 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_115 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_159 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_183 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_224 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_228 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_241 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_249 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_278 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_318 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_338 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_376 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_388 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_399 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_407 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_466 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_474 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_506 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_516 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_533 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_571 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_587 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_641 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_645 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_663 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_672 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_684 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_48_696 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_70 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_727 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_739 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_745 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_48_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_140 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_144 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_152 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_207 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_245 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_272 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_320 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_332 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_359 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_371 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_383 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_42 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_439 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_447 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_456 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_484 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_517 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_529 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_561 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_577 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_598 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_6 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_605 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_649 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_65 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_677 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_49_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_707 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_721 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_49_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_129 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_133 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_174 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_182 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_194 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_233 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_297 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_306 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_313 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_320 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_332 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_339 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_412 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_421 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_435 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_459 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_471 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_480 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_504 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_4_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_579 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_699 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_4_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_107 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_126 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_130 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_195 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_205 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_229 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_295 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_307 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_334 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_342 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_375 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_454 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_472 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_552 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_568 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_580 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_601 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_613 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_636 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_677 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_754 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_50_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_85 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_50_99 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_104 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_125 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_144 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_193 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_205 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_258 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_310 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_322 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_330 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_348 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_417 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_51_425 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_460 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_488 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_494 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_50 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_51_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_515 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_581 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_593 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_684 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_689 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_713 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_741 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_764 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_123 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_157 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_174 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_217 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_258 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_270 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_282 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_455 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_467 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_495 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_507 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_542 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_612 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_624 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_636 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_664 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_725 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_737 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_743 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_52_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_52_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_156 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_192 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_242 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_263 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_267 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_288 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_327 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_351 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_375 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_437 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_470 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_482 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_513 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_558 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_612 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_630 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_634 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_681 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_705 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_717 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_164 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_202 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_318 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_344 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_362 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_383 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_412 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_475 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_541 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_601 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_622 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_657 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_669 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_726 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_54_738 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_54_769 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_54_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_113 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_169 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_174 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_178 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_184 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_203 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_211 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_218 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_238 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_281 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_311 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_335 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_348 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_356 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_364 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_381 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_422 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_556 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_585 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_593 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_612 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_627 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_633 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_639 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_658 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_704 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_712 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_55_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_729 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_761 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_767 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_161 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_185 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_215 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_229 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_291 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_304 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_327 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_333 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_457 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_468 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_502 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_525 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_580 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_611 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_623 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_669 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_681 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_699 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_709 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_56_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_56_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_150 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_314 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_367 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_376 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_380 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_400 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_423 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_435 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_517 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_591 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_629 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_641 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_649 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_683 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_748 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_121 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_174 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_185 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_197 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_204 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_225 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_259 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_273 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_305 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_58_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_392 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_475 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_589 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_683 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_58_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_134 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_234 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_284 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_308 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_328 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_353 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_431 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_461 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_546 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_556 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_615 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_59_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_683 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_687 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_719 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_749 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_151 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_167 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_176 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_237 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_289 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_312 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_324 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_356 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_360 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_381 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_432 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_446 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_483 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_5_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_510 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_522 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_5_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_112 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_120 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_175 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_187 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_222 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_288 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_339 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_377 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_385 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_437 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_498 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_609 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_60_621 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_643 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_666 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_678 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_688 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_698 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_701 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_724 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_730 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_764 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_181 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_213 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_223 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_229 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_238 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_256 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_279 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_286 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_292 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_61_311 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_369 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_430 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_442 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_461 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_473 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_502 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_543 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_576 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_588 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_606 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_632 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_644 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_652 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_673 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_692 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_696 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_61_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_228 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_240 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_259 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_330 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_342 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_350 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_360 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_381 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_419 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_439 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_451 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_463 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_475 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_477 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_557 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_59 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_62_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_652 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_664 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_676 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_688 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_720 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_62_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_754 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_766 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_162 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_178 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_265 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_302 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_319 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_330 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_47 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_481 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_503 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_539 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_552 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_587 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_599 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_669 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_673 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_63_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_706 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_722 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_63_750 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_768 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_128 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_215 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_309 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_332 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_361 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_384 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_403 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_415 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_450 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_462 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_64_501 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_516 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_524 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_64_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_653 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_678 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_701 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_744 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_75 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_148 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_200 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_249 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_279 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_335 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_353 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_368 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_387 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_511 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_523 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_535 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_547 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_559 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_592 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_65_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_65_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_629 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_657 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_661 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_697 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_703 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_750 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_767 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_103 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_113 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_131 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_179 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_200 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_216 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_220 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_244 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_286 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_389 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_401 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_414 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_446 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_454 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_485 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_507 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_519 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_531 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_536 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_547 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_553 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_565 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_604 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_616 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_624 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_645 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_674 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_698 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_70 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_721 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_66_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_755 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_66_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_95 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_196 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_262 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_274 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_290 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_306 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_315 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_337 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_360 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_372 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_401 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_468 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_476 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_520 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_67_528 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_559 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_687 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_705 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_720 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_729 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_109 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_203 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_211 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_219 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_237 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_251 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_253 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_268 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_276 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_287 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_352 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_360 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_382 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_429 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_441 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_453 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_465 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_506 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_533 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_545 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_553 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_575 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_597 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_609 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_621 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_633 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_64 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_669 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_675 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_699 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_68_710 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_732 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_740 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_68_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_136 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_193 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_205 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_237 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_281 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_306 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_318 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_324 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_361 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_384 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_42 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_425 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_449 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_469 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_516 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_544 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_553 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_558 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_567 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_614 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_654 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_666 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_714 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_725 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_138 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_141 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_168 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_18 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_184 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_203 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_215 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_227 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_300 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_309 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_353 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_371 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_387 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_394 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_424 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_441 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_482 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_486 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_492 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_522 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_6_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_701 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_6_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_120 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_132 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_136 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_154 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_171 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_184 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_203 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_21 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_238 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_250 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_253 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_37 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_388 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_396 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_405 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_437 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_454 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_473 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_485 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_494 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_506 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_52 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_577 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_70_586 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_589 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_626 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_630 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_649 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_70_725 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_733 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_747 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_96 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_135 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_147 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_190 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_223 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_242 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_246 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_366 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_378 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_382 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_429 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_444 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_458 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_466 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_476 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_488 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_536 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_585 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_613 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_635 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_646 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_673 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_726 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_737 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_71_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_112 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_128 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_150 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_162 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_214 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_23 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_230 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_274 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_282 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_290 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_300 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_338 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_362 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_380 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_392 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_400 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_407 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_437 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_450 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_462 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_47 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_477 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_489 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_512 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_523 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_554 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_596 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_608 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_61 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_620 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_72_628 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_643 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_650 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_658 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_675 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_707 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_736 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_748 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_72_768 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_102 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_165 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_186 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_198 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_210 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_222 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_240 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_261 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_279 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_318 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_330 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_35 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_354 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_373 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_405 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_42 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_440 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_466 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_478 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_502 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_528 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_540 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_548 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_555 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_577 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_608 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_641 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_647 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_694 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_702 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_725 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_73_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_752 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_764 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_172 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_209 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_231 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_258 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_266 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_276 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_288 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_300 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_329 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_341 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_353 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_373 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_417 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_424 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_432 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_464 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_472 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_531 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_566 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_586 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_619 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_62 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_648 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_660 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_672 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_684 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_690 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_74_698 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_74_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_102 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_108 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_155 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_185 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_221 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_241 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_249 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_277 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_281 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_285 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_303 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_320 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_334 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_349 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_357 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_374 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_408 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_420 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_424 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_441 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_517 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_549 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_564 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_572 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_583 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_595 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_608 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_626 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_638 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_644 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_652 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_664 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_668 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_695 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_771 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_75_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_75_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_100 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_112 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_120 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_150 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_162 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_180 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_192 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_221 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_233 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_250 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_260 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_316 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_324 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_343 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_363 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_365 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_397 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_444 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_452 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_477 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_481 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_485 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_492 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_500 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_514 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_568 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_58 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_601 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_633 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_666 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_70 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_734 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_754 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_765 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_76_82 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_88 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_100 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_120 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_128 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_138 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_144 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_208 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_213 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_317 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_329 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_357 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_380 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_428 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_440 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_469 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_481 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_513 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_521 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_554 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_592 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_623 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_632 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_644 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_678 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_690 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_702 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_714 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_77_726 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_77_769 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_101 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_107 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_119 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_166 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_170 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_178 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_197 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_204 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_240 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_246 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_284 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_318 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_330 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_342 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_362 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_377 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_404 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_429 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_437 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_44 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_453 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_459 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_490 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_502 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_508 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_545 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_569 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_581 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_589 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_618 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_640 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_743 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_78_769 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_121 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_155 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_181 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_218 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_259 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_271 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_279 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_298 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_306 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_346 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_359 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_363 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_382 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_400 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_412 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_426 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_447 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_47 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_501 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_517 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_537 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_569 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_577 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_588 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_594 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_602 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_653 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_66 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_671 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_673 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_79_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_719 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_74 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_771 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_90 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_79_98 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_143 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_164 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_175 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_237 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_285 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_297 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_335 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_366 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_378 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_390 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_399 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_40 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_406 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_415 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_427 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_446 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_7_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_464 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_487 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_512 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_52 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_538 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_558 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_570 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_582 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_594 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_606 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_7_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_123 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_132 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_156 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_221 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_227 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_253 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_265 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_274 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_304 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_315 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_332 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_344 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_352 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_358 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_369 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_378 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_390 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_394 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_414 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_430 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_436 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_461 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_470 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_499 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_515 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_554 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_558 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_564 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_580 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_608 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_61 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_620 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_630 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_648 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_652 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_683 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_69 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_695 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_701 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_716 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_742 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_97 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_110 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_124 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_142 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_201 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_220 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_231 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_255 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_267 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_301 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_313 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_325 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_337 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_349 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_373 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_405 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_447 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_45 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_484 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_492 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_510 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_516 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_524 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_532 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_536 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_577 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_583 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_615 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_617 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_658 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_670 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_711 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_723 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_81_770 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_105 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_129 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_137 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_197 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_230 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_250 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_271 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_283 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_295 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_307 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_345 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_363 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_374 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_386 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_390 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_397 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_409 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_421 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_433 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_443 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_451 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_513 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_525 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_531 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_541 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_565 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_622 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_629 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_650 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_67 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_701 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_721 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_737 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_82_746 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_754 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_82_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_113 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_125 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_129 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_133 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_145 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_169 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_212 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_225 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_248 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_252 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_28 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_304 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_360 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_364 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_40 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_414 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_423 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_431 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_472 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_496 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_505 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_52 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_532 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_573 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_585 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_593 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_604 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_83_610 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_626 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_638 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_646 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_680 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_692 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_704 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_711 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_719 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_83_736 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_83_744 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_83_749 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_137 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_149 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_172 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_209 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_221 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_233 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_239 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_246 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_312 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_327 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_333 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_369 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_386 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_398 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_427 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_439 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_45 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_451 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_463 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_498 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_520 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_529 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_546 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_558 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_566 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_586 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_641 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_655 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_689 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_697 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_718 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_722 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_84_753 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_763 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_771 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_84_82 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_158 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_178 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_190 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_233 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_256 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_268 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_281 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_356 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_386 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_393 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_405 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_417 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_434 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_446 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_456 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_468 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_480 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_85_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_512 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_524 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_536 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_548 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_561 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_570 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_580 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_588 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_614 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_85_625 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_645 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_671 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_673 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_696 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_729 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_741 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_764 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_85_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_90 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_109 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_130 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_138 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_190 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_231 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_253 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_261 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_276 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_288 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_29 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_304 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_344 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_397 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_486 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_498 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_515 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_519 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_540 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_560 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_572 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_584 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_596 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_600 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_608 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_620 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_626 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_633 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_86_657 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_675 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_713 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_86_738 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_86_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_104 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_119 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_127 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_154 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_162 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_177 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_183 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_225 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_23 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_237 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_242 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_249 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_257 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_334 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_343 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_365 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_377 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_416 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_428 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_436 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_445 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_449 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_459 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_50 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_503 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_511 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_523 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_544 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_559 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_569 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_581 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_593 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_601 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_607 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_617 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_645 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_657 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_662 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_87_670 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_685 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_713 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_729 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_87_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_749 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_83 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_114 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_126 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_158 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_170 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_184 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_191 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_209 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_239 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_278 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_290 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_300 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_331 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_343 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_362 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_373 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_383 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_457 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_477 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_489 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_497 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_52 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_530 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_545 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_557 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_565 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_581 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_88_596 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_605 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_618 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_64 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_88_640 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_652 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_679 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_691 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_699 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_709 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_721 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_733 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_739 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_764 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_93 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_102 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_125 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_164 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_189 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_202 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_222 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_225 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_232 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_266 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_305 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_313 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_325 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_342 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_354 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_366 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_377 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_382 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_390 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_413 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_440 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_449 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_470 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_476 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_498 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_511 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_527 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_549 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_561 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_569 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_575 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_587 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_599 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_611 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_629 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_645 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_673 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_685 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_693 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_713 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_72 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_729 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_756 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_89_768 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_84 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_96 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_118 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_177 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_195 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_211 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_235 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_247 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_251 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_277 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_284 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_296 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_333 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_398 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_410 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_418 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_433 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_457 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_469 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_475 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_489 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_526 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_54 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_546 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_559 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_563 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_584 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_643 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_657 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_681 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_693 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_699 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_715 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_739 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_8_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_769 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_97 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_101 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_109 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_122 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_135 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_139 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_141 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_155 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_163 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_168 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_180 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_195 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_202 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_213 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_230 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_253 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_265 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_276 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_280 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_302 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_309 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_321 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_356 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_389 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_401 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_413 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_419 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_434 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_44 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_452 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_464 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_484 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_496 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_504 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_522 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_530 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_533 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_551 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_56 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_563 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_601 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_613 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_622 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_90_630 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_657 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_682 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_708 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_716 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_737 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_745 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_751 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_761 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_90_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_90_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_107 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_111 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_119 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_152 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_164 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_199 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_211 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_219 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_228 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_236 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_245 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_301 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_328 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_337 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_375 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_391 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_393 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_408 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_420 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_428 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_436 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_442 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_46 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_462 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_470 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_500 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_517 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_529 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_91_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_567 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_579 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_587 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_613 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_617 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_647 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_91_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_668 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_91_693 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_712 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_724 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_91_758 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_95 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_12 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_122 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_134 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_150 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_160 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_209 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_221 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_24 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_251 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_258 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_269 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_281 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_293 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_305 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_333 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_345 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_351 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_363 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_365 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_371 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_379 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_419 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_433 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_445 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_474 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_489 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_501 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_513 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_528 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_542 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_555 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_589 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_620 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_632 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_668 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_686 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_698 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_712 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_724 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_92_736 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_740 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_749 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_755 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_762 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_77 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_92_770 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_91 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_99 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_111 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_113 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_124 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_160 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_175 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_223 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_253 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_264 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_276 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_315 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_345 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_356 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_368 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_385 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_445 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_457 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_461 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_485 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_518 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_530 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_542 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_93_557 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_569 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_595 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_607 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_617 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_642 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_646 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_656 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_668 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_682 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_713 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_93_726 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_755 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_93_771 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_99 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_106 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_119 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_131 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_141 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_153 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_165 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_182 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_188 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_192 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_197 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_23 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_231 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_239 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_248 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_263 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_287 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_299 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_307 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_309 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_313 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_346 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_358 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_365 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_387 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_393 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_402 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_410 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_417 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_425 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_43 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_470 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_500 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_512 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_520 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_533 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_541 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_552 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_576 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_627 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_639 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_643 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_658 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_670 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_694 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_708 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_94_716 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_732 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_744 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_94_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_116 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_124 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_130 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_140 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_152 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_157 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_190 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_202 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_208 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_232 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_244 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_251 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_263 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_273 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_279 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_310 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_314 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_320 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_346 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_357 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_369 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_383 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_391 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_425 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_449 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_483 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_491 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_503 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_505 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_544 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_556 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_567 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_579 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_591 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_615 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_627 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_639 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_647 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_655 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_663 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_679 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_691 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_703 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_715 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_724 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_729 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_737 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_747 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_753 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_767 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_95_82 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_90 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_109 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_117 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_141 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_156 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_168 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_175 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_195 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_209 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_217 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_222 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_234 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_242 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_250 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_265 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_306 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_309 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_321 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_325 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_354 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_362 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_385 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_397 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_421 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_443 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_456 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_468 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_477 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_514 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_541 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_554 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_578 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_586 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_589 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_597 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_603 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_619 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_96_624 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_628 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_685 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_697 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_706 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_732 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_740 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_96_757 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_766 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_96_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_97 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_102 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_110 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_127 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_146 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_186 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_198 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_206 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_225 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_236 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_246 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_252 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_272 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_281 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_305 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_357 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_361 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_365 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_377 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_387 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_393 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_401 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_413 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_429 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_441 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_447 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_457 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_465 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_491 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_503 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_97_516 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_539 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_547 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_553 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_559 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_561 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_573 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_594 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_602 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_97_614 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_97_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_682 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_694 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_715 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_727 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_747 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_759 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_771 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_102 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_114 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_126 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_138 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_165 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_180 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_197 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_210 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_218 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_224 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_234 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_246 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_253 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_270 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_278 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_321 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_333 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_355 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_363 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_365 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_399 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_411 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_419 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_421 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_442 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_446 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_475 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_489 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_501 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_528 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_545 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_564 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_576 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_601 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_625 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_637 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_643 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_98_645 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_651 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_660 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_672 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_678 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_68 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_699 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_704 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_716 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_728 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_98_740 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_746 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_755 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_757 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_769 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_85 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_101 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_110 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_113 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_147 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_159 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_232 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_244 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_261 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_281 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_293 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_326 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_334 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_337 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_345 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_369 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_377 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_416 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_425 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_437 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_453 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_460 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_472 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_478 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_505 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_51 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_526 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_538 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_550 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_558 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_571 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_583 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_595 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_62 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_631 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_650 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_99_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_671 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_693 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_99_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_74 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_99_741 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_762 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_99_766 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_86 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_113 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_123 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_131 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_143 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_161 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_178 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_205 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_217 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_233 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_245 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_260 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_272 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_277 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_286 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_294 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_301 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_319 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_331 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_335 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_337 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_349 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_387 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_391 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_393 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_410 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_414 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_435 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_447 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_449 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_478 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_503 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_9_525 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_541 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_554 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_573 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_597 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_609 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_615 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_629 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_653 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_665 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_709 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_721 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_727 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_741 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_753 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_765 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_771 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1057 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1058 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1059 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1060 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1061 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1062 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1063 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1064 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1065 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1066 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1067 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1068 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1069 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1070 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1071 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1072 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1073 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1074 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1075 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1076 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1077 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1078 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1079 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1080 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1081 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1082 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1083 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1084 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1085 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1086 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1087 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1088 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1089 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1090 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1091 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1092 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1093 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1094 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1095 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1096 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1097 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1098 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1099 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1100 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1101 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1102 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1103 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1104 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1105 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1106 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1107 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1108 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1109 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1110 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1111 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1112 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1113 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1114 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1115 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1116 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1117 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1118 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1119 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1120 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1121 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1122 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1123 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1124 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1125 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1126 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1127 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1128 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1129 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1130 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1131 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1132 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1133 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1134 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1135 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1136 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1137 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1138 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1139 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1140 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1141 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1142 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1143 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1144 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1145 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1146 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1147 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1148 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1149 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1150 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1151 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1152 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1153 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1154 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1155 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1156 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1157 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1158 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1159 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1160 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1161 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1162 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1163 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1164 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1165 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_1999 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2000 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2001 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2002 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2003 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2004 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2005 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2006 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2007 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2008 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2009 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2010 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2011 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2012 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2013 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2014 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2015 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2016 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2017 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2018 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2019 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2020 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2021 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2022 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2023 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2024 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2025 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2026 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2027 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2028 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2029 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2030 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2031 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2032 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2033 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2034 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2035 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2036 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2037 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2038 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2039 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2040 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2041 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2042 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2043 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2044 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2045 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2046 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2047 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2048 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2049 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2050 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2051 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2052 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2053 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2054 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2055 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_2056 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_628 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_629 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_630 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_631 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_632 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_633 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_634 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_635 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_636 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_637 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_638 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_639 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_640 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_641 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_642 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_643 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_644 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_645 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_646 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_647 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_648 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_649 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_650 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_651 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_652 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_653 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_654 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_655 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_656 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_657 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_658 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_659 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_660 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_661 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_662 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_663 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_664 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_665 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_666 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_667 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_668 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_669 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_670 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_671 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_672 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_673 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_674 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_675 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_676 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_677 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_678 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_679 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_680 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_681 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_682 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_683 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_684 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_685 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_686 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_687 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_688 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_689 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_690 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_691 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_692 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_693 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_694 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_695 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_696 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_697 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_698 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_699 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_700 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_701 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_702 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_703 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_704 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_705 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_706 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_707 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_708 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_709 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_710 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_711 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_712 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_713 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_714 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_715 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_716 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_717 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_718 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_719 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_720 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_721 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_722 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_723 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_724 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_725 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_726 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_727 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_728 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_729 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_730 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_731 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_732 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_733 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_734 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_735 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_736 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_737 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_738 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_739 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_740 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_741 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_742 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_743 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_744 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_745 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_746 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_747 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_748 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_749 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_750 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_751 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_752 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_753 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_754 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_755 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_756 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_757 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_758 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_759 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_760 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_761 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_762 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_763 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_764 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_765 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_766 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_767 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_768 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_769 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_770 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_771 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_772 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_773 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_774 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_775 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_776 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_777 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_778 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_779 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_780 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_781 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_782 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_783 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_784 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_785 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_786 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_787 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_788 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_789 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_790 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_791 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_792 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_793 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_794 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_795 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_796 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_797 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_798 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_799 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_800 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_801 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_802 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_803 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_804 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_805 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_806 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_807 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_808 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_809 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_810 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_811 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_812 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_813 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_814 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_815 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_816 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_817 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_818 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_819 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_820 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_821 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_822 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_823 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_824 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_825 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_826 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_827 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_828 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_829 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_830 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_831 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_832 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_833 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_834 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_835 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_836 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_837 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_838 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_839 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_840 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_841 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_842 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_843 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_844 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_845 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_846 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_847 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_848 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_849 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_850 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_851 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_852 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_853 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_854 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_855 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_856 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_857 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_858 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_859 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_860 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_861 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_862 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_863 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_864 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_865 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_866 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_867 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_868 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_869 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_870 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_871 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_872 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_873 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_874 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_875 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_876 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_877 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_878 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_879 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_880 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_881 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_882 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_883 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_884 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_885 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_886 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_887 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_888 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_889 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_890 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_891 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_892 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_893 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_894 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_895 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_896 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_897 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_898 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_899 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_900 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_901 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_902 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_903 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_904 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_905 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_906 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_907 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_908 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_909 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_910 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_911 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_912 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_913 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_914 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_915 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_916 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_917 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_918 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_919 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_920 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_921 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_922 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_923 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_924 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_925 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_926 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_927 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_928 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_929 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_930 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_931 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_932 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_933 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_934 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_935 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_936 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_937 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_938 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_939 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_940 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_941 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_942 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_943 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_944 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_945 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_946 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_947 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_948 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_949 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_950 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_951 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_952 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_953 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_954 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_955 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_956 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_957 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_958 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_959 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_960 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_961 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_962 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_963 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_964 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_965 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_966 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_967 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_968 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_969 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_970 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_971 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_972 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_973 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_974 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_975 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_976 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_977 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_978 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_979 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_980 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_981 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_982 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_983 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_984 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_985 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_986 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_987 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_988 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_989 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_990 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_991 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_992 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_993 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_994 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_995 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_996 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_997 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_998 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_999 ();
 sky130_fd_sc_hd__inv_2 _3757_ (.A(\inputcont.INTERNAL_SYNCED_I[10] ),
    .Y(_0441_));
 sky130_fd_sc_hd__or4_1 _3758_ (.A(\inputcont.INTERNAL_SYNCED_I[0] ),
    .B(\inputcont.INTERNAL_SYNCED_I[1] ),
    .C(\inputcont.INTERNAL_SYNCED_I[3] ),
    .D(\inputcont.INTERNAL_SYNCED_I[2] ),
    .X(_0442_));
 sky130_fd_sc_hd__clkbuf_8 _3759_ (.A(_0442_),
    .X(_0443_));
 sky130_fd_sc_hd__or4_4 _3760_ (.A(\inputcont.INTERNAL_SYNCED_I[5] ),
    .B(\inputcont.INTERNAL_SYNCED_I[4] ),
    .C(\inputcont.INTERNAL_SYNCED_I[7] ),
    .D(\inputcont.INTERNAL_SYNCED_I[6] ),
    .X(_0444_));
 sky130_fd_sc_hd__or4_4 _3761_ (.A(\inputcont.INTERNAL_SYNCED_I[9] ),
    .B(\inputcont.INTERNAL_SYNCED_I[8] ),
    .C(_0443_),
    .D(_0444_),
    .X(_0445_));
 sky130_fd_sc_hd__inv_2 _3762_ (.A(\inputcont.INTERNAL_SYNCED_I[12] ),
    .Y(_0446_));
 sky130_fd_sc_hd__or4_2 _3763_ (.A(_0446_),
    .B(\inputcont.INTERNAL_SYNCED_I[11] ),
    .C(\inputcont.INTERNAL_SYNCED_I[10] ),
    .D(_0445_),
    .X(_0447_));
 sky130_fd_sc_hd__nor2_1 _3764_ (.A(_0443_),
    .B(_0444_),
    .Y(_0448_));
 sky130_fd_sc_hd__inv_2 _3765_ (.A(\inputcont.INTERNAL_SYNCED_I[1] ),
    .Y(_0449_));
 sky130_fd_sc_hd__inv_2 _3766_ (.A(_0443_),
    .Y(_0450_));
 sky130_fd_sc_hd__a221o_1 _3767_ (.A1(_0449_),
    .A2(\inputcont.INTERNAL_SYNCED_I[2] ),
    .B1(\inputcont.INTERNAL_SYNCED_I[4] ),
    .B2(_0450_),
    .C1(\inputcont.INTERNAL_SYNCED_I[0] ),
    .X(_0451_));
 sky130_fd_sc_hd__a21oi_1 _3768_ (.A1(\inputcont.INTERNAL_SYNCED_I[8] ),
    .A2(_0448_),
    .B1(_0451_),
    .Y(_0452_));
 sky130_fd_sc_hd__or4b_2 _3769_ (.A(\inputcont.INTERNAL_SYNCED_I[5] ),
    .B(_0443_),
    .C(\inputcont.INTERNAL_SYNCED_I[4] ),
    .D_N(\inputcont.INTERNAL_SYNCED_I[6] ),
    .X(_0453_));
 sky130_fd_sc_hd__o2111ai_4 _3770_ (.A1(_0441_),
    .A2(_0445_),
    .B1(_0447_),
    .C1(_0452_),
    .D1(_0453_),
    .Y(net35));
 sky130_fd_sc_hd__or3_1 _3771_ (.A(\inputcont.INTERNAL_SYNCED_I[8] ),
    .B(_0443_),
    .C(_0444_),
    .X(_0454_));
 sky130_fd_sc_hd__o21ba_1 _3772_ (.A1(\inputcont.INTERNAL_SYNCED_I[9] ),
    .A2(\inputcont.INTERNAL_SYNCED_I[10] ),
    .B1_N(_0454_),
    .X(_0455_));
 sky130_fd_sc_hd__inv_2 _3773_ (.A(\inputcont.INTERNAL_SYNCED_I[5] ),
    .Y(_0456_));
 sky130_fd_sc_hd__nor2_1 _3774_ (.A(\inputcont.INTERNAL_SYNCED_I[1] ),
    .B(\inputcont.INTERNAL_SYNCED_I[2] ),
    .Y(_0457_));
 sky130_fd_sc_hd__o32a_1 _3775_ (.A1(_0456_),
    .A2(\inputcont.INTERNAL_SYNCED_I[4] ),
    .A3(_0443_),
    .B1(_0457_),
    .B2(\inputcont.INTERNAL_SYNCED_I[0] ),
    .X(_0458_));
 sky130_fd_sc_hd__nand3b_2 _3776_ (.A_N(_0455_),
    .B(_0458_),
    .C(_0453_),
    .Y(net36));
 sky130_fd_sc_hd__or2_1 _3777_ (.A(\inputcont.INTERNAL_SYNCED_I[0] ),
    .B(\inputcont.INTERNAL_SYNCED_I[1] ),
    .X(_0459_));
 sky130_fd_sc_hd__nor2_1 _3778_ (.A(\inputcont.INTERNAL_SYNCED_I[2] ),
    .B(_0459_),
    .Y(_0460_));
 sky130_fd_sc_hd__or3b_1 _3779_ (.A(\inputcont.INTERNAL_SYNCED_I[10] ),
    .B(_0445_),
    .C_N(\inputcont.INTERNAL_SYNCED_I[11] ),
    .X(_0461_));
 sky130_fd_sc_hd__nand2_1 _3780_ (.A(_0447_),
    .B(_0461_),
    .Y(_0462_));
 sky130_fd_sc_hd__or2_2 _3781_ (.A(\inputcont.INTERNAL_SYNCED_I[5] ),
    .B(\inputcont.INTERNAL_SYNCED_I[4] ),
    .X(_0463_));
 sky130_fd_sc_hd__o21a_1 _3782_ (.A1(\inputcont.INTERNAL_SYNCED_I[6] ),
    .A2(_0463_),
    .B1(_0450_),
    .X(_0464_));
 sky130_fd_sc_hd__a211o_1 _3783_ (.A1(\inputcont.INTERNAL_SYNCED_I[3] ),
    .A2(_0460_),
    .B1(_0462_),
    .C1(_0464_),
    .X(net37));
 sky130_fd_sc_hd__or4b_1 _3784_ (.A(\inputcont.INTERNAL_SYNCED_I[6] ),
    .B(_0443_),
    .C(_0463_),
    .D_N(\inputcont.INTERNAL_SYNCED_I[7] ),
    .X(_0465_));
 sky130_fd_sc_hd__inv_2 _3785_ (.A(_0465_),
    .Y(_0466_));
 sky130_fd_sc_hd__a211o_1 _3786_ (.A1(\inputcont.INTERNAL_SYNCED_I[8] ),
    .A2(_0448_),
    .B1(_0455_),
    .C1(_0466_),
    .X(_0467_));
 sky130_fd_sc_hd__or2_1 _3787_ (.A(_0462_),
    .B(_0467_),
    .X(_0468_));
 sky130_fd_sc_hd__clkbuf_4 _3788_ (.A(_0468_),
    .X(net38));
 sky130_fd_sc_hd__and2b_1 _3789_ (.A_N(net1),
    .B(\wave.mode[0] ),
    .X(_0469_));
 sky130_fd_sc_hd__clkbuf_4 _3790_ (.A(_0469_),
    .X(net30));
 sky130_fd_sc_hd__or3b_1 _3791_ (.A(_0464_),
    .B(_0443_),
    .C_N(_0461_),
    .X(_0470_));
 sky130_fd_sc_hd__o21a_1 _3792_ (.A1(_0467_),
    .A2(_0470_),
    .B1(\inputcont.INTERNAL_SYNCED_I[12] ),
    .X(_0471_));
 sky130_fd_sc_hd__inv_2 _3793_ (.A(_0471_),
    .Y(_0472_));
 sky130_fd_sc_hd__nand2_1 _3794_ (.A(\inputcont.INTERNAL_SYNCED_I[11] ),
    .B(_0461_),
    .Y(_0473_));
 sky130_fd_sc_hd__o21a_1 _3795_ (.A1(_0443_),
    .A2(_0444_),
    .B1(\inputcont.INTERNAL_SYNCED_I[8] ),
    .X(_0474_));
 sky130_fd_sc_hd__o31a_2 _3796_ (.A1(\inputcont.INTERNAL_SYNCED_I[8] ),
    .A2(_0443_),
    .A3(_0444_),
    .B1(\inputcont.INTERNAL_SYNCED_I[9] ),
    .X(_0475_));
 sky130_fd_sc_hd__o31a_1 _3797_ (.A1(\inputcont.INTERNAL_SYNCED_I[6] ),
    .A2(_0443_),
    .A3(_0463_),
    .B1(\inputcont.INTERNAL_SYNCED_I[7] ),
    .X(_0476_));
 sky130_fd_sc_hd__a2111o_1 _3798_ (.A1(\inputcont.INTERNAL_SYNCED_I[10] ),
    .A2(_0445_),
    .B1(_0474_),
    .C1(_0475_),
    .D1(_0476_),
    .X(_0477_));
 sky130_fd_sc_hd__o21ai_4 _3799_ (.A1(\inputcont.INTERNAL_SYNCED_I[4] ),
    .A2(_0443_),
    .B1(\inputcont.INTERNAL_SYNCED_I[5] ),
    .Y(_0478_));
 sky130_fd_sc_hd__o21ai_4 _3800_ (.A1(_0443_),
    .A2(_0463_),
    .B1(\inputcont.INTERNAL_SYNCED_I[6] ),
    .Y(_0479_));
 sky130_fd_sc_hd__o31ai_4 _3801_ (.A1(\inputcont.INTERNAL_SYNCED_I[0] ),
    .A2(\inputcont.INTERNAL_SYNCED_I[1] ),
    .A3(\inputcont.INTERNAL_SYNCED_I[2] ),
    .B1(\inputcont.INTERNAL_SYNCED_I[3] ),
    .Y(_0480_));
 sky130_fd_sc_hd__nand2_2 _3802_ (.A(\inputcont.INTERNAL_SYNCED_I[0] ),
    .B(\inputcont.INTERNAL_SYNCED_I[1] ),
    .Y(_0481_));
 sky130_fd_sc_hd__o21ai_4 _3803_ (.A1(\inputcont.INTERNAL_SYNCED_I[0] ),
    .A2(\inputcont.INTERNAL_SYNCED_I[1] ),
    .B1(\inputcont.INTERNAL_SYNCED_I[2] ),
    .Y(_0482_));
 sky130_fd_sc_hd__o41ai_1 _3804_ (.A1(\inputcont.INTERNAL_SYNCED_I[0] ),
    .A2(\inputcont.INTERNAL_SYNCED_I[1] ),
    .A3(\inputcont.INTERNAL_SYNCED_I[3] ),
    .A4(\inputcont.INTERNAL_SYNCED_I[2] ),
    .B1(\inputcont.INTERNAL_SYNCED_I[4] ),
    .Y(_0483_));
 sky130_fd_sc_hd__and4_1 _3805_ (.A(_0480_),
    .B(_0481_),
    .C(_0482_),
    .D(net67),
    .X(_0484_));
 sky130_fd_sc_hd__buf_2 _3806_ (.A(_0484_),
    .X(_0485_));
 sky130_fd_sc_hd__and4b_1 _3807_ (.A_N(_0477_),
    .B(_0478_),
    .C(_0479_),
    .D(_0485_),
    .X(_0486_));
 sky130_fd_sc_hd__nand2_1 _3808_ (.A(_0473_),
    .B(_0486_),
    .Y(_0487_));
 sky130_fd_sc_hd__nor2_1 _3809_ (.A(_0474_),
    .B(_0475_),
    .Y(_0488_));
 sky130_fd_sc_hd__o31ai_2 _3810_ (.A1(\inputcont.INTERNAL_SYNCED_I[6] ),
    .A2(_0443_),
    .A3(_0463_),
    .B1(\inputcont.INTERNAL_SYNCED_I[7] ),
    .Y(_0489_));
 sky130_fd_sc_hd__and4_1 _3811_ (.A(_0479_),
    .B(_0478_),
    .C(_0485_),
    .D(_0489_),
    .X(_0490_));
 sky130_fd_sc_hd__clkbuf_4 _3812_ (.A(_0490_),
    .X(_0491_));
 sky130_fd_sc_hd__and4_1 _3813_ (.A(\inputcont.INTERNAL_SYNCED_I[10] ),
    .B(_0445_),
    .C(_0488_),
    .D(_0491_),
    .X(_0492_));
 sky130_fd_sc_hd__or2b_1 _3814_ (.A(_0479_),
    .B_N(_0478_),
    .X(_0493_));
 sky130_fd_sc_hd__nand2_1 _3815_ (.A(_0483_),
    .B(_0493_),
    .Y(_0494_));
 sky130_fd_sc_hd__and3_1 _3816_ (.A(_0480_),
    .B(_0481_),
    .C(_0482_),
    .X(_0495_));
 sky130_fd_sc_hd__and3_1 _3817_ (.A(\inputcont.INTERNAL_SYNCED_I[2] ),
    .B(_0459_),
    .C(_0481_),
    .X(_0496_));
 sky130_fd_sc_hd__a221o_1 _3818_ (.A1(_0474_),
    .A2(_0491_),
    .B1(_0494_),
    .B2(_0495_),
    .C1(_0496_),
    .X(_0497_));
 sky130_fd_sc_hd__or2_1 _3819_ (.A(_0492_),
    .B(_0497_),
    .X(_0498_));
 sky130_fd_sc_hd__o21ba_4 _3820_ (.A1(_0472_),
    .A2(_0487_),
    .B1_N(_0498_),
    .X(_0499_));
 sky130_fd_sc_hd__clkinv_4 _3821_ (.A(_0499_),
    .Y(net39));
 sky130_fd_sc_hd__o21ai_4 _3822_ (.A1(_0443_),
    .A2(_0444_),
    .B1(\inputcont.INTERNAL_SYNCED_I[8] ),
    .Y(_0500_));
 sky130_fd_sc_hd__nand2_1 _3823_ (.A(_0479_),
    .B(_0478_),
    .Y(_0501_));
 sky130_fd_sc_hd__nand2_2 _3824_ (.A(_0481_),
    .B(_0482_),
    .Y(_0502_));
 sky130_fd_sc_hd__a211o_1 _3825_ (.A1(_0485_),
    .A2(_0501_),
    .B1(_0492_),
    .C1(_0502_),
    .X(_0503_));
 sky130_fd_sc_hd__a31oi_4 _3826_ (.A1(_0500_),
    .A2(_0475_),
    .A3(_0491_),
    .B1(_0503_),
    .Y(_0504_));
 sky130_fd_sc_hd__inv_2 _3827_ (.A(_0504_),
    .Y(net40));
 sky130_fd_sc_hd__a21boi_1 _3828_ (.A1(_0472_),
    .A2(_0473_),
    .B1_N(_0486_),
    .Y(_0505_));
 sky130_fd_sc_hd__a41o_1 _3829_ (.A1(_0479_),
    .A2(_0478_),
    .A3(_0480_),
    .A4(net67),
    .B1(_0502_),
    .X(_0506_));
 sky130_fd_sc_hd__nor2b_2 _3830_ (.A(_0505_),
    .B_N(_0506_),
    .Y(_0507_));
 sky130_fd_sc_hd__inv_2 _3831_ (.A(_0507_),
    .Y(net41));
 sky130_fd_sc_hd__and3_1 _3832_ (.A(_0479_),
    .B(_0478_),
    .C(_0485_),
    .X(_0508_));
 sky130_fd_sc_hd__a21o_2 _3833_ (.A1(_0508_),
    .A2(_0477_),
    .B1(_0505_),
    .X(net42));
 sky130_fd_sc_hd__and2b_1 _3834_ (.A_N(net1),
    .B(\wave.mode[1] ),
    .X(_0509_));
 sky130_fd_sc_hd__buf_4 _3835_ (.A(_0509_),
    .X(net31));
 sky130_fd_sc_hd__nand2_1 _3836_ (.A(_0471_),
    .B(_0487_),
    .Y(_0510_));
 sky130_fd_sc_hd__and3_1 _3837_ (.A(\inputcont.INTERNAL_SYNCED_I[0] ),
    .B(\inputcont.INTERNAL_SYNCED_I[1] ),
    .C(\inputcont.INTERNAL_SYNCED_I[2] ),
    .X(_0511_));
 sky130_fd_sc_hd__buf_2 _3838_ (.A(_0511_),
    .X(_0512_));
 sky130_fd_sc_hd__a31oi_4 _3839_ (.A1(_0480_),
    .A2(_0481_),
    .A3(_0482_),
    .B1(net67),
    .Y(_0513_));
 sky130_fd_sc_hd__a211o_1 _3840_ (.A1(\inputcont.INTERNAL_SYNCED_I[3] ),
    .A2(_0502_),
    .B1(_0512_),
    .C1(_0513_),
    .X(_0514_));
 sky130_fd_sc_hd__nor2_2 _3841_ (.A(_0500_),
    .B(_0491_),
    .Y(_0515_));
 sky130_fd_sc_hd__nor2_1 _3842_ (.A(_0478_),
    .B(_0485_),
    .Y(_0516_));
 sky130_fd_sc_hd__a21oi_1 _3843_ (.A1(_0478_),
    .A2(_0485_),
    .B1(_0479_),
    .Y(_0517_));
 sky130_fd_sc_hd__a31oi_2 _3844_ (.A1(_0479_),
    .A2(_0478_),
    .A3(_0485_),
    .B1(_0489_),
    .Y(_0518_));
 sky130_fd_sc_hd__or4_2 _3845_ (.A(_0514_),
    .B(_0516_),
    .C(_0517_),
    .D(_0518_),
    .X(_0519_));
 sky130_fd_sc_hd__nor2_1 _3846_ (.A(_0515_),
    .B(_0519_),
    .Y(_0520_));
 sky130_fd_sc_hd__a21boi_4 _3847_ (.A1(_0500_),
    .A2(_0491_),
    .B1_N(_0475_),
    .Y(_0521_));
 sky130_fd_sc_hd__nor2_1 _3848_ (.A(\inputcont.INTERNAL_SYNCED_I[9] ),
    .B(_0454_),
    .Y(_0522_));
 sky130_fd_sc_hd__a211oi_4 _3849_ (.A1(_0488_),
    .A2(_0491_),
    .B1(_0441_),
    .C1(_0522_),
    .Y(_0523_));
 sky130_fd_sc_hd__nor4_1 _3850_ (.A(_0473_),
    .B(_0486_),
    .C(_0521_),
    .D(_0523_),
    .Y(_0524_));
 sky130_fd_sc_hd__or2_2 _3851_ (.A(_0478_),
    .B(_0485_),
    .X(_0525_));
 sky130_fd_sc_hd__a21o_1 _3852_ (.A1(_0478_),
    .A2(_0485_),
    .B1(_0479_),
    .X(_0526_));
 sky130_fd_sc_hd__and3b_1 _3853_ (.A_N(_0514_),
    .B(_0525_),
    .C(_0526_),
    .X(_0527_));
 sky130_fd_sc_hd__o41a_1 _3854_ (.A1(_0515_),
    .A2(_0518_),
    .A3(_0521_),
    .A4(_0523_),
    .B1(_0527_),
    .X(_0528_));
 sky130_fd_sc_hd__inv_2 _3855_ (.A(_0513_),
    .Y(_0529_));
 sky130_fd_sc_hd__a21oi_1 _3856_ (.A1(\inputcont.INTERNAL_SYNCED_I[3] ),
    .A2(_0502_),
    .B1(_0512_),
    .Y(_0530_));
 sky130_fd_sc_hd__nand2_1 _3857_ (.A(_0525_),
    .B(_0526_),
    .Y(_0531_));
 sky130_fd_sc_hd__and3_1 _3858_ (.A(_0529_),
    .B(_0530_),
    .C(_0531_),
    .X(_0532_));
 sky130_fd_sc_hd__a211o_1 _3859_ (.A1(_0520_),
    .A2(_0524_),
    .B1(_0528_),
    .C1(_0532_),
    .X(_0533_));
 sky130_fd_sc_hd__or3_2 _3860_ (.A(_0510_),
    .B(_0514_),
    .C(_0533_),
    .X(_0534_));
 sky130_fd_sc_hd__or4b_1 _3861_ (.A(_0515_),
    .B(_0519_),
    .C(_0521_),
    .D_N(_0523_),
    .X(_0535_));
 sky130_fd_sc_hd__a21o_1 _3862_ (.A1(_0525_),
    .A2(_0517_),
    .B1(_0513_),
    .X(_0536_));
 sky130_fd_sc_hd__nor3_1 _3863_ (.A(_0500_),
    .B(_0491_),
    .C(_0519_),
    .Y(_0537_));
 sky130_fd_sc_hd__a211oi_1 _3864_ (.A1(_0530_),
    .A2(_0536_),
    .B1(net57),
    .C1(_0512_),
    .Y(_0538_));
 sky130_fd_sc_hd__and3_1 _3865_ (.A(_0534_),
    .B(_0535_),
    .C(_0538_),
    .X(_0539_));
 sky130_fd_sc_hd__buf_4 _3866_ (.A(_0539_),
    .X(_0540_));
 sky130_fd_sc_hd__inv_2 _3867_ (.A(_0540_),
    .Y(net43));
 sky130_fd_sc_hd__or2_1 _3868_ (.A(_0521_),
    .B(_0523_),
    .X(_0541_));
 sky130_fd_sc_hd__a211oi_1 _3869_ (.A1(_0520_),
    .A2(_0541_),
    .B1(_0512_),
    .C1(_0532_),
    .Y(_0542_));
 sky130_fd_sc_hd__inv_2 _3870_ (.A(_0542_),
    .Y(net44));
 sky130_fd_sc_hd__nor2_1 _3871_ (.A(_0513_),
    .B(_0531_),
    .Y(_0543_));
 sky130_fd_sc_hd__a21boi_1 _3872_ (.A1(\inputcont.INTERNAL_SYNCED_I[3] ),
    .A2(_0502_),
    .B1_N(_0543_),
    .Y(_0544_));
 sky130_fd_sc_hd__nand2_1 _3873_ (.A(_0520_),
    .B(_0524_),
    .Y(_0545_));
 sky130_fd_sc_hd__o211a_2 _3874_ (.A1(_0512_),
    .A2(_0544_),
    .B1(_0534_),
    .C1(_0545_),
    .X(_0546_));
 sky130_fd_sc_hd__inv_2 _3875_ (.A(_0546_),
    .Y(net45));
 sky130_fd_sc_hd__a21oi_1 _3876_ (.A1(_0520_),
    .A2(_0541_),
    .B1(net57),
    .Y(_0547_));
 sky130_fd_sc_hd__nand2_1 _3877_ (.A(_0518_),
    .B(_0527_),
    .Y(_0548_));
 sky130_fd_sc_hd__and3_2 _3878_ (.A(_0545_),
    .B(_0547_),
    .C(_0548_),
    .X(_0549_));
 sky130_fd_sc_hd__nand2_4 _3879_ (.A(_0549_),
    .B(_0534_),
    .Y(net46));
 sky130_fd_sc_hd__and3_1 _3880_ (.A(\rate_clk.count[1] ),
    .B(\rate_clk.count[0] ),
    .C(\rate_clk.count[2] ),
    .X(_0550_));
 sky130_fd_sc_hd__and2_1 _3881_ (.A(\rate_clk.count[3] ),
    .B(_0550_),
    .X(_0551_));
 sky130_fd_sc_hd__and3_1 _3882_ (.A(\rate_clk.count[5] ),
    .B(\rate_clk.count[4] ),
    .C(_0551_),
    .X(_0552_));
 sky130_fd_sc_hd__and2_2 _3883_ (.A(\rate_clk.count[6] ),
    .B(_0552_),
    .X(_0553_));
 sky130_fd_sc_hd__nand2_8 _3884_ (.A(\rate_clk.count[7] ),
    .B(_0553_),
    .Y(_0554_));
 sky130_fd_sc_hd__inv_2 _3885_ (.A(\sound4.sdiv.start ),
    .Y(_0555_));
 sky130_fd_sc_hd__a311oi_4 _3886_ (.A1(\sound4.sdiv.C[4] ),
    .A2(\sound4.sdiv.C[3] ),
    .A3(\sound4.sdiv.C[2] ),
    .B1(_0555_),
    .C1(\sound4.sdiv.C[5] ),
    .Y(_0556_));
 sky130_fd_sc_hd__inv_2 _3887_ (.A(_0556_),
    .Y(_0557_));
 sky130_fd_sc_hd__inv_2 _3888_ (.A(\sound2.sdiv.start ),
    .Y(_0558_));
 sky130_fd_sc_hd__a311oi_4 _3889_ (.A1(\sound2.sdiv.C[4] ),
    .A2(\sound2.sdiv.C[3] ),
    .A3(\sound2.sdiv.C[2] ),
    .B1(_0558_),
    .C1(\sound2.sdiv.C[5] ),
    .Y(_0559_));
 sky130_fd_sc_hd__inv_2 _3890_ (.A(_0559_),
    .Y(_0560_));
 sky130_fd_sc_hd__inv_2 _3891_ (.A(\sound3.sdiv.start ),
    .Y(_0561_));
 sky130_fd_sc_hd__a311oi_4 _3892_ (.A1(\sound3.sdiv.C[4] ),
    .A2(\sound3.sdiv.C[3] ),
    .A3(\sound3.sdiv.C[2] ),
    .B1(_0561_),
    .C1(\sound3.sdiv.C[5] ),
    .Y(_0562_));
 sky130_fd_sc_hd__inv_2 _3893_ (.A(_0562_),
    .Y(_0563_));
 sky130_fd_sc_hd__inv_2 _3894_ (.A(\sound1.sdiv.start ),
    .Y(_0564_));
 sky130_fd_sc_hd__a311oi_4 _3895_ (.A1(\sound1.sdiv.C[4] ),
    .A2(\sound1.sdiv.C[3] ),
    .A3(\sound1.sdiv.C[2] ),
    .B1(_0564_),
    .C1(\sound1.sdiv.C[5] ),
    .Y(_0565_));
 sky130_fd_sc_hd__inv_2 _3896_ (.A(net65),
    .Y(_0566_));
 sky130_fd_sc_hd__a22o_1 _3897_ (.A1(\sound3.sdiv.dived ),
    .A2(_0563_),
    .B1(_0566_),
    .B2(\sound1.sdiv.dived ),
    .X(_0567_));
 sky130_fd_sc_hd__a221o_2 _3898_ (.A1(\sound4.sdiv.dived ),
    .A2(_0557_),
    .B1(_0560_),
    .B2(\sound2.sdiv.dived ),
    .C1(_0567_),
    .X(_0568_));
 sky130_fd_sc_hd__nand2_8 _3899_ (.A(_0554_),
    .B(_0568_),
    .Y(_0569_));
 sky130_fd_sc_hd__inv_2 _3900_ (.A(\wave_comb.u1.start ),
    .Y(_0570_));
 sky130_fd_sc_hd__a2111o_4 _3901_ (.A1(\wave_comb.u1.C[3] ),
    .A2(\wave_comb.u1.C[2] ),
    .B1(_0570_),
    .C1(\wave_comb.u1.C[5] ),
    .D1(\wave_comb.u1.C[4] ),
    .X(_0571_));
 sky130_fd_sc_hd__and2_1 _3902_ (.A(_0569_),
    .B(_0571_),
    .X(_0572_));
 sky130_fd_sc_hd__clkbuf_8 _3903_ (.A(_0572_),
    .X(_0573_));
 sky130_fd_sc_hd__inv_2 _3904_ (.A(_0573_),
    .Y(\wave_comb.u1.next_start ));
 sky130_fd_sc_hd__and3_1 _3905_ (.A(\rate_clk.count[6] ),
    .B(\rate_clk.count[7] ),
    .C(_0552_),
    .X(_0574_));
 sky130_fd_sc_hd__clkbuf_16 _3906_ (.A(_0574_),
    .X(_0575_));
 sky130_fd_sc_hd__nor2_4 _3907_ (.A(_0575_),
    .B(_0556_),
    .Y(_0576_));
 sky130_fd_sc_hd__inv_2 _3908_ (.A(_0576_),
    .Y(\sound4.sdiv.next_start ));
 sky130_fd_sc_hd__nor2_8 _3909_ (.A(_0575_),
    .B(net147),
    .Y(_0577_));
 sky130_fd_sc_hd__inv_2 _3910_ (.A(_0577_),
    .Y(\sound3.sdiv.next_start ));
 sky130_fd_sc_hd__nor2_8 _3911_ (.A(_0575_),
    .B(net66),
    .Y(_0578_));
 sky130_fd_sc_hd__inv_2 _3912_ (.A(_0578_),
    .Y(\sound2.sdiv.next_start ));
 sky130_fd_sc_hd__nor2_4 _3913_ (.A(_0575_),
    .B(net65),
    .Y(_0579_));
 sky130_fd_sc_hd__inv_2 _3914_ (.A(_0579_),
    .Y(\sound1.sdiv.next_start ));
 sky130_fd_sc_hd__nor3_1 _3915_ (.A(_0510_),
    .B(_0514_),
    .C(_0533_),
    .Y(_0580_));
 sky130_fd_sc_hd__o311a_1 _3916_ (.A1(_0512_),
    .A2(_0533_),
    .A3(_0580_),
    .B1(_0502_),
    .C1(\inputcont.INTERNAL_SYNCED_I[3] ),
    .X(_0581_));
 sky130_fd_sc_hd__o31a_2 _3917_ (.A1(_0510_),
    .A2(_0513_),
    .A3(_0533_),
    .B1(_0530_),
    .X(_0582_));
 sky130_fd_sc_hd__a21o_1 _3918_ (.A1(_0549_),
    .A2(_0582_),
    .B1(_0529_),
    .X(_0583_));
 sky130_fd_sc_hd__a41o_1 _3919_ (.A1(_0529_),
    .A2(_0525_),
    .A3(_0549_),
    .A4(_0582_),
    .B1(_0526_),
    .X(_0584_));
 sky130_fd_sc_hd__a31o_1 _3920_ (.A1(_0529_),
    .A2(_0549_),
    .A3(_0582_),
    .B1(_0525_),
    .X(_0585_));
 sky130_fd_sc_hd__and4b_1 _3921_ (.A_N(_0581_),
    .B(_0583_),
    .C(_0584_),
    .D(_0585_),
    .X(_0586_));
 sky130_fd_sc_hd__clkbuf_4 _3922_ (.A(_0586_),
    .X(_0587_));
 sky130_fd_sc_hd__or2b_1 _3923_ (.A(_0581_),
    .B_N(_0583_),
    .X(_0588_));
 sky130_fd_sc_hd__a21oi_2 _3924_ (.A1(_0584_),
    .A2(_0585_),
    .B1(_0588_),
    .Y(_0589_));
 sky130_fd_sc_hd__nand3_2 _3925_ (.A(_0548_),
    .B(_0543_),
    .C(_0582_),
    .Y(_0590_));
 sky130_fd_sc_hd__o21ba_1 _3926_ (.A1(_0515_),
    .A2(_0521_),
    .B1_N(_0519_),
    .X(_0591_));
 sky130_fd_sc_hd__o21a_1 _3927_ (.A1(_0590_),
    .A2(_0591_),
    .B1(_0523_),
    .X(_0592_));
 sky130_fd_sc_hd__inv_2 _3928_ (.A(_0545_),
    .Y(_0593_));
 sky130_fd_sc_hd__o31a_1 _3929_ (.A1(_0593_),
    .A2(net57),
    .A3(_0590_),
    .B1(_0521_),
    .X(_0594_));
 sky130_fd_sc_hd__or2_2 _3930_ (.A(_0592_),
    .B(_0594_),
    .X(_0595_));
 sky130_fd_sc_hd__nand2_1 _3931_ (.A(_0515_),
    .B(_0590_),
    .Y(_0596_));
 sky130_fd_sc_hd__a311o_1 _3932_ (.A1(_0545_),
    .A2(_0543_),
    .A3(_0582_),
    .B1(_0489_),
    .C1(_0508_),
    .X(_0597_));
 sky130_fd_sc_hd__and3b_1 _3933_ (.A_N(_0595_),
    .B(_0596_),
    .C(_0597_),
    .X(_0598_));
 sky130_fd_sc_hd__o21ba_1 _3934_ (.A1(_0514_),
    .A2(_0533_),
    .B1_N(_0510_),
    .X(_0599_));
 sky130_fd_sc_hd__inv_2 _3935_ (.A(_0547_),
    .Y(_0600_));
 sky130_fd_sc_hd__nor2_1 _3936_ (.A(_0473_),
    .B(_0486_),
    .Y(_0601_));
 sky130_fd_sc_hd__o21a_1 _3937_ (.A1(_0600_),
    .A2(_0590_),
    .B1(_0601_),
    .X(_0602_));
 sky130_fd_sc_hd__nor2_1 _3938_ (.A(_0599_),
    .B(_0602_),
    .Y(_0603_));
 sky130_fd_sc_hd__and3_1 _3939_ (.A(_0587_),
    .B(_0597_),
    .C(_0596_),
    .X(_0604_));
 sky130_fd_sc_hd__or3b_2 _3940_ (.A(_0603_),
    .B(_0595_),
    .C_N(_0604_),
    .X(_0605_));
 sky130_fd_sc_hd__o31a_2 _3941_ (.A1(_0588_),
    .A2(_0589_),
    .A3(_0598_),
    .B1(_0605_),
    .X(_0606_));
 sky130_fd_sc_hd__nand2_8 _3942_ (.A(_0587_),
    .B(_0606_),
    .Y(net34));
 sky130_fd_sc_hd__inv_2 _3943_ (.A(\inputcont.INTERNAL_SYNCED_I[3] ),
    .Y(_0607_));
 sky130_fd_sc_hd__and2_1 _3944_ (.A(\inputcont.INTERNAL_SYNCED_I[6] ),
    .B(\inputcont.INTERNAL_SYNCED_I[8] ),
    .X(_0608_));
 sky130_fd_sc_hd__nor2_1 _3945_ (.A(\inputcont.INTERNAL_SYNCED_I[6] ),
    .B(\inputcont.INTERNAL_SYNCED_I[8] ),
    .Y(_0609_));
 sky130_fd_sc_hd__nor2_1 _3946_ (.A(_0608_),
    .B(_0609_),
    .Y(_0610_));
 sky130_fd_sc_hd__xnor2_1 _3947_ (.A(\inputcont.INTERNAL_SYNCED_I[10] ),
    .B(_0610_),
    .Y(_0611_));
 sky130_fd_sc_hd__inv_2 _3948_ (.A(\inputcont.INTERNAL_SYNCED_I[4] ),
    .Y(_0612_));
 sky130_fd_sc_hd__a21oi_1 _3949_ (.A1(_0459_),
    .A2(_0481_),
    .B1(\inputcont.INTERNAL_SYNCED_I[2] ),
    .Y(_0613_));
 sky130_fd_sc_hd__or2_1 _3950_ (.A(_0496_),
    .B(_0613_),
    .X(_0614_));
 sky130_fd_sc_hd__nor2_1 _3951_ (.A(_0612_),
    .B(_0614_),
    .Y(_0615_));
 sky130_fd_sc_hd__and2_1 _3952_ (.A(_0612_),
    .B(_0614_),
    .X(_0616_));
 sky130_fd_sc_hd__or2_1 _3953_ (.A(_0615_),
    .B(_0616_),
    .X(_0617_));
 sky130_fd_sc_hd__xor2_1 _3954_ (.A(\inputcont.INTERNAL_SYNCED_I[11] ),
    .B(_0617_),
    .X(_0618_));
 sky130_fd_sc_hd__nor2_1 _3955_ (.A(_0611_),
    .B(_0618_),
    .Y(_0619_));
 sky130_fd_sc_hd__and2_1 _3956_ (.A(_0611_),
    .B(_0618_),
    .X(_0620_));
 sky130_fd_sc_hd__nor2_1 _3957_ (.A(_0619_),
    .B(_0620_),
    .Y(_0621_));
 sky130_fd_sc_hd__and2_1 _3958_ (.A(\inputcont.INTERNAL_SYNCED_I[7] ),
    .B(_0621_),
    .X(_0622_));
 sky130_fd_sc_hd__nor2_1 _3959_ (.A(\inputcont.INTERNAL_SYNCED_I[7] ),
    .B(_0621_),
    .Y(_0623_));
 sky130_fd_sc_hd__nor2_1 _3960_ (.A(_0622_),
    .B(_0623_),
    .Y(_0624_));
 sky130_fd_sc_hd__xnor2_1 _3961_ (.A(\inputcont.INTERNAL_SYNCED_I[9] ),
    .B(_0624_),
    .Y(_0625_));
 sky130_fd_sc_hd__or2_1 _3962_ (.A(_0456_),
    .B(_0625_),
    .X(_0626_));
 sky130_fd_sc_hd__nand2_1 _3963_ (.A(_0456_),
    .B(_0625_),
    .Y(_0627_));
 sky130_fd_sc_hd__nand2_1 _3964_ (.A(_0626_),
    .B(_0627_),
    .Y(_0628_));
 sky130_fd_sc_hd__xnor2_1 _3965_ (.A(_0446_),
    .B(_0628_),
    .Y(_0629_));
 sky130_fd_sc_hd__nor2_2 _3966_ (.A(_0607_),
    .B(_0629_),
    .Y(_0630_));
 sky130_fd_sc_hd__and2_1 _3967_ (.A(_0607_),
    .B(_0629_),
    .X(_0631_));
 sky130_fd_sc_hd__or2_4 _3968_ (.A(_0630_),
    .B(_0631_),
    .X(_0632_));
 sky130_fd_sc_hd__nor2_2 _3969_ (.A(net34),
    .B(_0632_),
    .Y(net32));
 sky130_fd_sc_hd__a21oi_1 _3970_ (.A1(\inputcont.INTERNAL_SYNCED_I[10] ),
    .A2(_0610_),
    .B1(_0608_),
    .Y(_0633_));
 sky130_fd_sc_hd__o2bb2a_1 _3971_ (.A1_N(\inputcont.INTERNAL_SYNCED_I[4] ),
    .A2_N(_0512_),
    .B1(_0615_),
    .B2(_0502_),
    .X(_0634_));
 sky130_fd_sc_hd__inv_2 _3972_ (.A(_0617_),
    .Y(_0635_));
 sky130_fd_sc_hd__a21oi_1 _3973_ (.A1(\inputcont.INTERNAL_SYNCED_I[11] ),
    .A2(_0635_),
    .B1(_0619_),
    .Y(_0636_));
 sky130_fd_sc_hd__xnor2_1 _3974_ (.A(_0634_),
    .B(_0636_),
    .Y(_0637_));
 sky130_fd_sc_hd__xnor2_1 _3975_ (.A(_0633_),
    .B(_0637_),
    .Y(_0638_));
 sky130_fd_sc_hd__a21oi_1 _3976_ (.A1(\inputcont.INTERNAL_SYNCED_I[9] ),
    .A2(_0624_),
    .B1(_0622_),
    .Y(_0639_));
 sky130_fd_sc_hd__xnor2_1 _3977_ (.A(_0638_),
    .B(_0639_),
    .Y(_0640_));
 sky130_fd_sc_hd__o21a_1 _3978_ (.A1(_0446_),
    .A2(_0628_),
    .B1(_0626_),
    .X(_0641_));
 sky130_fd_sc_hd__xnor2_2 _3979_ (.A(_0640_),
    .B(_0641_),
    .Y(_0642_));
 sky130_fd_sc_hd__xnor2_4 _3980_ (.A(_0630_),
    .B(_0642_),
    .Y(_0643_));
 sky130_fd_sc_hd__nor2_2 _3981_ (.A(net34),
    .B(_0643_),
    .Y(net33));
 sky130_fd_sc_hd__and2_1 _3982_ (.A(_0554_),
    .B(_0568_),
    .X(_0644_));
 sky130_fd_sc_hd__buf_4 _3983_ (.A(_0644_),
    .X(_0645_));
 sky130_fd_sc_hd__nor2_2 _3984_ (.A(_0645_),
    .B(_0571_),
    .Y(_0646_));
 sky130_fd_sc_hd__buf_4 _3985_ (.A(_0646_),
    .X(\wave_comb.u1.next_dived ));
 sky130_fd_sc_hd__inv_2 _3986_ (.A(\pm.count[0] ),
    .Y(\pm.next_count[0] ));
 sky130_fd_sc_hd__xor2_1 _3987_ (.A(\pm.count[1] ),
    .B(\pm.count[0] ),
    .X(\pm.next_count[1] ));
 sky130_fd_sc_hd__and3_1 _3988_ (.A(\pm.count[1] ),
    .B(\pm.count[0] ),
    .C(\pm.count[2] ),
    .X(_0647_));
 sky130_fd_sc_hd__a21oi_1 _3989_ (.A1(\pm.count[1] ),
    .A2(\pm.count[0] ),
    .B1(\pm.count[2] ),
    .Y(_0648_));
 sky130_fd_sc_hd__nor2_1 _3990_ (.A(_0647_),
    .B(_0648_),
    .Y(\pm.next_count[2] ));
 sky130_fd_sc_hd__and2_1 _3991_ (.A(\pm.count[3] ),
    .B(_0647_),
    .X(_0649_));
 sky130_fd_sc_hd__nor2_1 _3992_ (.A(\pm.count[3] ),
    .B(_0647_),
    .Y(_0650_));
 sky130_fd_sc_hd__nor2_1 _3993_ (.A(_0649_),
    .B(_0650_),
    .Y(\pm.next_count[3] ));
 sky130_fd_sc_hd__inv_2 _3994_ (.A(\pm.count[4] ),
    .Y(_0651_));
 sky130_fd_sc_hd__xnor2_1 _3995_ (.A(_0651_),
    .B(_0649_),
    .Y(\pm.next_count[4] ));
 sky130_fd_sc_hd__and3_1 _3996_ (.A(\pm.count[5] ),
    .B(\pm.count[4] ),
    .C(_0649_),
    .X(_0652_));
 sky130_fd_sc_hd__a21oi_1 _3997_ (.A1(\pm.count[4] ),
    .A2(_0649_),
    .B1(\pm.count[5] ),
    .Y(_0653_));
 sky130_fd_sc_hd__nor2_1 _3998_ (.A(_0652_),
    .B(_0653_),
    .Y(\pm.next_count[5] ));
 sky130_fd_sc_hd__and2_1 _3999_ (.A(\pm.count[6] ),
    .B(_0652_),
    .X(_0654_));
 sky130_fd_sc_hd__buf_1 _4000_ (.A(_0654_),
    .X(_0655_));
 sky130_fd_sc_hd__nor2_1 _4001_ (.A(\pm.count[6] ),
    .B(_0652_),
    .Y(_0656_));
 sky130_fd_sc_hd__nor2_1 _4002_ (.A(_0655_),
    .B(_0656_),
    .Y(\pm.next_count[6] ));
 sky130_fd_sc_hd__inv_2 _4003_ (.A(\pm.count[7] ),
    .Y(_0657_));
 sky130_fd_sc_hd__xnor2_1 _4004_ (.A(_0657_),
    .B(_0655_),
    .Y(\pm.next_count[7] ));
 sky130_fd_sc_hd__a21boi_1 _4005_ (.A1(\pm.count[7] ),
    .A2(_0655_),
    .B1_N(\pm.count[8] ),
    .Y(\pm.next_count[8] ));
 sky130_fd_sc_hd__inv_2 _4006_ (.A(\inputcont.u3.next_in ),
    .Y(_0658_));
 sky130_fd_sc_hd__and3_1 _4007_ (.A(\wave.mode[0] ),
    .B(\inputcont.INTERNAL_MODE ),
    .C(_0658_),
    .X(_0659_));
 sky130_fd_sc_hd__a21oi_1 _4008_ (.A1(\inputcont.INTERNAL_MODE ),
    .A2(_0658_),
    .B1(\wave.mode[0] ),
    .Y(_0660_));
 sky130_fd_sc_hd__nor2_1 _4009_ (.A(_0659_),
    .B(_0660_),
    .Y(\wave.next_state[0] ));
 sky130_fd_sc_hd__xor2_1 _4010_ (.A(\wave.mode[1] ),
    .B(_0659_),
    .X(\wave.next_state[1] ));
 sky130_fd_sc_hd__inv_2 _4011_ (.A(\seq.encode.keys_sync[10] ),
    .Y(_0661_));
 sky130_fd_sc_hd__o21ai_1 _4012_ (.A1(_0661_),
    .A2(\seq.encode.keys_edge_det[10] ),
    .B1(\seq.tempo_select.state[0] ),
    .Y(_0662_));
 sky130_fd_sc_hd__or3_1 _4013_ (.A(_0661_),
    .B(\seq.encode.keys_edge_det[10] ),
    .C(\seq.tempo_select.state[0] ),
    .X(_0663_));
 sky130_fd_sc_hd__nand2_1 _4014_ (.A(_0662_),
    .B(_0663_),
    .Y(\seq.tempo_select.next_state[0] ));
 sky130_fd_sc_hd__nand2_1 _4015_ (.A(\seq.tempo_select.state[1] ),
    .B(\seq.tempo_select.state[0] ),
    .Y(_0664_));
 sky130_fd_sc_hd__or2_1 _4016_ (.A(\seq.tempo_select.state[1] ),
    .B(\seq.tempo_select.state[0] ),
    .X(_0665_));
 sky130_fd_sc_hd__nand2_1 _4017_ (.A(_0664_),
    .B(_0665_),
    .Y(_0666_));
 sky130_fd_sc_hd__xor2_1 _4018_ (.A(_0662_),
    .B(_0666_),
    .X(\seq.tempo_select.next_state[1] ));
 sky130_fd_sc_hd__nand2_1 _4019_ (.A(_0587_),
    .B(_0597_),
    .Y(_0667_));
 sky130_fd_sc_hd__inv_2 _4020_ (.A(_0599_),
    .Y(_0668_));
 sky130_fd_sc_hd__o21ba_1 _4021_ (.A1(_0668_),
    .A2(_0602_),
    .B1_N(_0592_),
    .X(_0669_));
 sky130_fd_sc_hd__o21a_1 _4022_ (.A1(_0594_),
    .A2(_0669_),
    .B1(_0596_),
    .X(_0670_));
 sky130_fd_sc_hd__or3b_1 _4023_ (.A(_0588_),
    .B(_0584_),
    .C_N(_0585_),
    .X(_0671_));
 sky130_fd_sc_hd__o21a_1 _4024_ (.A1(_0581_),
    .A2(_0583_),
    .B1(_0671_),
    .X(_0672_));
 sky130_fd_sc_hd__o21ai_4 _4025_ (.A1(_0667_),
    .A2(_0670_),
    .B1(_0672_),
    .Y(net47));
 sky130_fd_sc_hd__a21oi_4 _4026_ (.A1(_0604_),
    .A2(_0595_),
    .B1(_0589_),
    .Y(_0673_));
 sky130_fd_sc_hd__inv_2 _4027_ (.A(_0673_),
    .Y(net48));
 sky130_fd_sc_hd__nand2_2 _4028_ (.A(_0587_),
    .B(_0605_),
    .Y(net49));
 sky130_fd_sc_hd__inv_2 _4029_ (.A(_0606_),
    .Y(net50));
 sky130_fd_sc_hd__buf_12 _4030_ (.A(\oct.state[2] ),
    .X(_0674_));
 sky130_fd_sc_hd__inv_4 _4031_ (.A(_0674_),
    .Y(_0675_));
 sky130_fd_sc_hd__buf_12 _4032_ (.A(\oct.state[1] ),
    .X(_0676_));
 sky130_fd_sc_hd__buf_12 _4033_ (.A(\oct.state[0] ),
    .X(_0677_));
 sky130_fd_sc_hd__nand2_8 _4034_ (.A(_0676_),
    .B(_0677_),
    .Y(_0678_));
 sky130_fd_sc_hd__nor2_4 _4035_ (.A(_0675_),
    .B(_0678_),
    .Y(_0679_));
 sky130_fd_sc_hd__inv_8 _4036_ (.A(\oct.state[0] ),
    .Y(_0680_));
 sky130_fd_sc_hd__nor2_4 _4037_ (.A(_0676_),
    .B(_0680_),
    .Y(_0681_));
 sky130_fd_sc_hd__nor2b_4 _4038_ (.A(\inputcont.u2.next_in ),
    .B_N(\inputcont.INTERNAL_OCTAVE_INPUT ),
    .Y(_0682_));
 sky130_fd_sc_hd__nor2_8 _4039_ (.A(_0674_),
    .B(_0678_),
    .Y(_0683_));
 sky130_fd_sc_hd__nor2_8 _4040_ (.A(_0676_),
    .B(\oct.state[0] ),
    .Y(_0684_));
 sky130_fd_sc_hd__buf_12 _4041_ (.A(_0675_),
    .X(_0685_));
 sky130_fd_sc_hd__inv_6 _4042_ (.A(_0676_),
    .Y(_0686_));
 sky130_fd_sc_hd__nor2_8 _4043_ (.A(_0686_),
    .B(_0677_),
    .Y(_0687_));
 sky130_fd_sc_hd__nand2_8 _4044_ (.A(_0685_),
    .B(_0687_),
    .Y(_0688_));
 sky130_fd_sc_hd__nand2_1 _4045_ (.A(_0682_),
    .B(_0688_),
    .Y(_0689_));
 sky130_fd_sc_hd__o32a_1 _4046_ (.A1(_0681_),
    .A2(_0682_),
    .A3(_0683_),
    .B1(_0684_),
    .B2(_0689_),
    .X(_0690_));
 sky130_fd_sc_hd__or2_1 _4047_ (.A(_0679_),
    .B(_0690_),
    .X(_0691_));
 sky130_fd_sc_hd__clkbuf_1 _4048_ (.A(_0691_),
    .X(\oct.next_state[0] ));
 sky130_fd_sc_hd__o32a_1 _4049_ (.A1(_0682_),
    .A2(_0683_),
    .A3(_0687_),
    .B1(_0689_),
    .B2(_0681_),
    .X(_0692_));
 sky130_fd_sc_hd__or2_1 _4050_ (.A(_0679_),
    .B(_0692_),
    .X(_0693_));
 sky130_fd_sc_hd__clkbuf_1 _4051_ (.A(_0693_),
    .X(\oct.next_state[1] ));
 sky130_fd_sc_hd__nor2_2 _4052_ (.A(_0676_),
    .B(_0675_),
    .Y(_0694_));
 sky130_fd_sc_hd__buf_12 _4053_ (.A(_0674_),
    .X(_0695_));
 sky130_fd_sc_hd__nand2_4 _4054_ (.A(_0695_),
    .B(_0687_),
    .Y(_0696_));
 sky130_fd_sc_hd__nor2_1 _4055_ (.A(_0682_),
    .B(_0696_),
    .Y(_0697_));
 sky130_fd_sc_hd__a211o_1 _4056_ (.A1(_0682_),
    .A2(_0683_),
    .B1(_0694_),
    .C1(_0697_),
    .X(\oct.next_state[2] ));
 sky130_fd_sc_hd__buf_8 _4057_ (.A(\select1.sequencer_on ),
    .X(_0698_));
 sky130_fd_sc_hd__inv_4 _4058_ (.A(_0698_),
    .Y(_0699_));
 sky130_fd_sc_hd__buf_12 _4059_ (.A(_0699_),
    .X(_0700_));
 sky130_fd_sc_hd__nor2_8 _4060_ (.A(_0700_),
    .B(net1),
    .Y(net52));
 sky130_fd_sc_hd__or3_4 _4061_ (.A(\seq.beat[1] ),
    .B(\seq.beat[0] ),
    .C(\seq.beat[2] ),
    .X(_0701_));
 sky130_fd_sc_hd__inv_2 _4062_ (.A(\seq.beat[3] ),
    .Y(_0702_));
 sky130_fd_sc_hd__nand2_4 _4063_ (.A(_0702_),
    .B(net52),
    .Y(_0703_));
 sky130_fd_sc_hd__nor2_1 _4064_ (.A(_0701_),
    .B(_0703_),
    .Y(net22));
 sky130_fd_sc_hd__or3b_4 _4065_ (.A(\seq.beat[0] ),
    .B(\seq.beat[2] ),
    .C_N(\seq.beat[1] ),
    .X(_0704_));
 sky130_fd_sc_hd__nor2_1 _4066_ (.A(_0703_),
    .B(_0704_),
    .Y(net23));
 sky130_fd_sc_hd__or3b_4 _4067_ (.A(\seq.beat[1] ),
    .B(\seq.beat[0] ),
    .C_N(\seq.beat[2] ),
    .X(_0705_));
 sky130_fd_sc_hd__nor2_2 _4068_ (.A(_0703_),
    .B(_0705_),
    .Y(net24));
 sky130_fd_sc_hd__nand3b_2 _4069_ (.A_N(\seq.beat[0] ),
    .B(\seq.beat[2] ),
    .C(\seq.beat[1] ),
    .Y(_0706_));
 sky130_fd_sc_hd__nor2_2 _4070_ (.A(_0703_),
    .B(_0706_),
    .Y(net25));
 sky130_fd_sc_hd__nand2_8 _4071_ (.A(\seq.beat[3] ),
    .B(net52),
    .Y(_0707_));
 sky130_fd_sc_hd__nor2_1 _4072_ (.A(_0701_),
    .B(_0707_),
    .Y(net26));
 sky130_fd_sc_hd__nor2_1 _4073_ (.A(_0704_),
    .B(_0707_),
    .Y(net27));
 sky130_fd_sc_hd__nor2_1 _4074_ (.A(_0705_),
    .B(_0707_),
    .Y(net28));
 sky130_fd_sc_hd__nor2_1 _4075_ (.A(_0706_),
    .B(_0707_),
    .Y(net29));
 sky130_fd_sc_hd__and2b_1 _4076_ (.A_N(net1),
    .B(net19),
    .X(_0708_));
 sky130_fd_sc_hd__clkbuf_1 _4077_ (.A(_0708_),
    .X(seq_play_on));
 sky130_fd_sc_hd__and2b_1 _4078_ (.A_N(net1),
    .B(net20),
    .X(_0709_));
 sky130_fd_sc_hd__clkbuf_1 _4079_ (.A(_0709_),
    .X(seq_power_on));
 sky130_fd_sc_hd__and2b_1 _4080_ (.A_N(net1),
    .B(net21),
    .X(_0710_));
 sky130_fd_sc_hd__clkbuf_1 _4081_ (.A(_0710_),
    .X(tempo_select_on));
 sky130_fd_sc_hd__and2b_1 _4082_ (.A_N(net1),
    .B(\pm.pwm_o ),
    .X(_0711_));
 sky130_fd_sc_hd__clkbuf_1 _4083_ (.A(_0711_),
    .X(net51));
 sky130_fd_sc_hd__and2b_1 _4084_ (.A_N(\seq.encode.keys_edge_det[9] ),
    .B(\inputcont.INTERNAL_SYNCED_I[7] ),
    .X(_0712_));
 sky130_fd_sc_hd__and2_1 _4085_ (.A(\seq.player_8.state[0] ),
    .B(_0712_),
    .X(_0713_));
 sky130_fd_sc_hd__a311o_1 _4086_ (.A1(\seq.player_8.state[1] ),
    .A2(\seq.player_8.state[2] ),
    .A3(\seq.player_8.state[3] ),
    .B1(_0713_),
    .C1(_0700_),
    .X(_0714_));
 sky130_fd_sc_hd__o21ba_1 _4087_ (.A1(\seq.player_8.state[0] ),
    .A2(_0712_),
    .B1_N(_0714_),
    .X(\seq.player_8.next_state[0] ));
 sky130_fd_sc_hd__and3_1 _4088_ (.A(\seq.player_8.state[0] ),
    .B(\seq.player_8.state[1] ),
    .C(_0712_),
    .X(_0715_));
 sky130_fd_sc_hd__nor2_1 _4089_ (.A(\seq.player_8.state[1] ),
    .B(_0713_),
    .Y(_0716_));
 sky130_fd_sc_hd__a2111oi_1 _4090_ (.A1(\seq.player_8.state[2] ),
    .A2(\seq.player_8.state[3] ),
    .B1(_0715_),
    .C1(_0716_),
    .D1(_0700_),
    .Y(\seq.player_8.next_state[1] ));
 sky130_fd_sc_hd__nand2_1 _4091_ (.A(\seq.player_8.state[2] ),
    .B(\seq.player_8.state[3] ),
    .Y(_0717_));
 sky130_fd_sc_hd__xor2_1 _4092_ (.A(\seq.player_8.state[2] ),
    .B(_0715_),
    .X(_0718_));
 sky130_fd_sc_hd__clkbuf_8 _4093_ (.A(_0698_),
    .X(_0719_));
 sky130_fd_sc_hd__o211a_1 _4094_ (.A1(_0717_),
    .A2(_0716_),
    .B1(_0718_),
    .C1(_0719_),
    .X(\seq.player_8.next_state[2] ));
 sky130_fd_sc_hd__a31o_1 _4095_ (.A1(\seq.player_8.state[1] ),
    .A2(\seq.player_8.state[2] ),
    .A3(_0713_),
    .B1(\seq.player_8.state[3] ),
    .X(_0720_));
 sky130_fd_sc_hd__o211a_1 _4096_ (.A1(_0717_),
    .A2(_0716_),
    .B1(_0720_),
    .C1(_0719_),
    .X(\seq.player_8.next_state[3] ));
 sky130_fd_sc_hd__and2b_1 _4097_ (.A_N(\seq.encode.keys_edge_det[8] ),
    .B(\inputcont.INTERNAL_SYNCED_I[6] ),
    .X(_0721_));
 sky130_fd_sc_hd__and2_1 _4098_ (.A(\seq.player_7.state[0] ),
    .B(_0721_),
    .X(_0722_));
 sky130_fd_sc_hd__a311o_1 _4099_ (.A1(\seq.player_7.state[1] ),
    .A2(\seq.player_7.state[2] ),
    .A3(\seq.player_7.state[3] ),
    .B1(_0722_),
    .C1(_0700_),
    .X(_0723_));
 sky130_fd_sc_hd__o21ba_1 _4100_ (.A1(\seq.player_7.state[0] ),
    .A2(_0721_),
    .B1_N(_0723_),
    .X(\seq.player_7.next_state[0] ));
 sky130_fd_sc_hd__and3_1 _4101_ (.A(\seq.player_7.state[0] ),
    .B(\seq.player_7.state[1] ),
    .C(_0721_),
    .X(_0724_));
 sky130_fd_sc_hd__nor2_1 _4102_ (.A(\seq.player_7.state[1] ),
    .B(_0722_),
    .Y(_0725_));
 sky130_fd_sc_hd__a2111oi_1 _4103_ (.A1(\seq.player_7.state[2] ),
    .A2(\seq.player_7.state[3] ),
    .B1(_0724_),
    .C1(_0725_),
    .D1(_0700_),
    .Y(\seq.player_7.next_state[1] ));
 sky130_fd_sc_hd__nand2_1 _4104_ (.A(\seq.player_7.state[2] ),
    .B(\seq.player_7.state[3] ),
    .Y(_0726_));
 sky130_fd_sc_hd__xor2_1 _4105_ (.A(\seq.player_7.state[2] ),
    .B(_0724_),
    .X(_0727_));
 sky130_fd_sc_hd__o211a_1 _4106_ (.A1(_0726_),
    .A2(_0725_),
    .B1(_0727_),
    .C1(_0719_),
    .X(\seq.player_7.next_state[2] ));
 sky130_fd_sc_hd__a31o_1 _4107_ (.A1(\seq.player_7.state[1] ),
    .A2(\seq.player_7.state[2] ),
    .A3(_0722_),
    .B1(\seq.player_7.state[3] ),
    .X(_0728_));
 sky130_fd_sc_hd__o211a_1 _4108_ (.A1(_0726_),
    .A2(_0725_),
    .B1(_0728_),
    .C1(_0719_),
    .X(\seq.player_7.next_state[3] ));
 sky130_fd_sc_hd__nor2_1 _4109_ (.A(_0456_),
    .B(\seq.encode.keys_edge_det[7] ),
    .Y(_0729_));
 sky130_fd_sc_hd__and2_1 _4110_ (.A(\seq.player_6.state[0] ),
    .B(_0729_),
    .X(_0730_));
 sky130_fd_sc_hd__a311o_1 _4111_ (.A1(\seq.player_6.state[1] ),
    .A2(\seq.player_6.state[2] ),
    .A3(\seq.player_6.state[3] ),
    .B1(_0730_),
    .C1(_0700_),
    .X(_0731_));
 sky130_fd_sc_hd__o21ba_1 _4112_ (.A1(\seq.player_6.state[0] ),
    .A2(_0729_),
    .B1_N(_0731_),
    .X(\seq.player_6.next_state[0] ));
 sky130_fd_sc_hd__and3_1 _4113_ (.A(\seq.player_6.state[0] ),
    .B(\seq.player_6.state[1] ),
    .C(_0729_),
    .X(_0732_));
 sky130_fd_sc_hd__nor2_1 _4114_ (.A(\seq.player_6.state[1] ),
    .B(_0730_),
    .Y(_0733_));
 sky130_fd_sc_hd__a2111oi_1 _4115_ (.A1(\seq.player_6.state[2] ),
    .A2(\seq.player_6.state[3] ),
    .B1(_0732_),
    .C1(_0733_),
    .D1(_0700_),
    .Y(\seq.player_6.next_state[1] ));
 sky130_fd_sc_hd__nand2_1 _4116_ (.A(\seq.player_6.state[2] ),
    .B(\seq.player_6.state[3] ),
    .Y(_0734_));
 sky130_fd_sc_hd__xor2_1 _4117_ (.A(\seq.player_6.state[2] ),
    .B(_0732_),
    .X(_0735_));
 sky130_fd_sc_hd__o211a_1 _4118_ (.A1(_0734_),
    .A2(_0733_),
    .B1(_0735_),
    .C1(_0719_),
    .X(\seq.player_6.next_state[2] ));
 sky130_fd_sc_hd__a31o_1 _4119_ (.A1(\seq.player_6.state[1] ),
    .A2(\seq.player_6.state[2] ),
    .A3(_0730_),
    .B1(\seq.player_6.state[3] ),
    .X(_0736_));
 sky130_fd_sc_hd__o211a_1 _4120_ (.A1(_0734_),
    .A2(_0733_),
    .B1(_0736_),
    .C1(_0719_),
    .X(\seq.player_6.next_state[3] ));
 sky130_fd_sc_hd__nor2_1 _4121_ (.A(_0612_),
    .B(\seq.encode.keys_edge_det[6] ),
    .Y(_0737_));
 sky130_fd_sc_hd__and2_1 _4122_ (.A(\seq.player_5.state[0] ),
    .B(_0737_),
    .X(_0738_));
 sky130_fd_sc_hd__a311o_1 _4123_ (.A1(\seq.player_5.state[1] ),
    .A2(\seq.player_5.state[2] ),
    .A3(\seq.player_5.state[3] ),
    .B1(_0738_),
    .C1(_0700_),
    .X(_0739_));
 sky130_fd_sc_hd__o21ba_1 _4124_ (.A1(\seq.player_5.state[0] ),
    .A2(_0737_),
    .B1_N(_0739_),
    .X(\seq.player_5.next_state[0] ));
 sky130_fd_sc_hd__and3_1 _4125_ (.A(\seq.player_5.state[0] ),
    .B(\seq.player_5.state[1] ),
    .C(_0737_),
    .X(_0740_));
 sky130_fd_sc_hd__nor2_1 _4126_ (.A(\seq.player_5.state[1] ),
    .B(_0738_),
    .Y(_0741_));
 sky130_fd_sc_hd__a2111oi_1 _4127_ (.A1(\seq.player_5.state[2] ),
    .A2(\seq.player_5.state[3] ),
    .B1(_0740_),
    .C1(_0741_),
    .D1(_0700_),
    .Y(\seq.player_5.next_state[1] ));
 sky130_fd_sc_hd__nand2_1 _4128_ (.A(\seq.player_5.state[2] ),
    .B(\seq.player_5.state[3] ),
    .Y(_0742_));
 sky130_fd_sc_hd__xor2_1 _4129_ (.A(\seq.player_5.state[2] ),
    .B(_0740_),
    .X(_0743_));
 sky130_fd_sc_hd__o211a_1 _4130_ (.A1(_0742_),
    .A2(_0741_),
    .B1(_0743_),
    .C1(_0719_),
    .X(\seq.player_5.next_state[2] ));
 sky130_fd_sc_hd__a31o_1 _4131_ (.A1(\seq.player_5.state[1] ),
    .A2(\seq.player_5.state[2] ),
    .A3(_0738_),
    .B1(\seq.player_5.state[3] ),
    .X(_0744_));
 sky130_fd_sc_hd__o211a_1 _4132_ (.A1(_0742_),
    .A2(_0741_),
    .B1(_0744_),
    .C1(_0719_),
    .X(\seq.player_5.next_state[3] ));
 sky130_fd_sc_hd__nor2_1 _4133_ (.A(_0607_),
    .B(\seq.encode.keys_edge_det[5] ),
    .Y(_0745_));
 sky130_fd_sc_hd__and2_1 _4134_ (.A(\seq.player_4.state[0] ),
    .B(_0745_),
    .X(_0746_));
 sky130_fd_sc_hd__a311o_1 _4135_ (.A1(\seq.player_4.state[1] ),
    .A2(\seq.player_4.state[2] ),
    .A3(\seq.player_4.state[3] ),
    .B1(_0746_),
    .C1(_0700_),
    .X(_0747_));
 sky130_fd_sc_hd__o21ba_1 _4136_ (.A1(\seq.player_4.state[0] ),
    .A2(_0745_),
    .B1_N(_0747_),
    .X(\seq.player_4.next_state[0] ));
 sky130_fd_sc_hd__and3_1 _4137_ (.A(\seq.player_4.state[0] ),
    .B(\seq.player_4.state[1] ),
    .C(_0745_),
    .X(_0748_));
 sky130_fd_sc_hd__nor2_1 _4138_ (.A(\seq.player_4.state[1] ),
    .B(_0746_),
    .Y(_0749_));
 sky130_fd_sc_hd__a2111oi_1 _4139_ (.A1(\seq.player_4.state[2] ),
    .A2(\seq.player_4.state[3] ),
    .B1(_0748_),
    .C1(_0749_),
    .D1(_0700_),
    .Y(\seq.player_4.next_state[1] ));
 sky130_fd_sc_hd__nand2_1 _4140_ (.A(\seq.player_4.state[2] ),
    .B(\seq.player_4.state[3] ),
    .Y(_0750_));
 sky130_fd_sc_hd__xor2_1 _4141_ (.A(\seq.player_4.state[2] ),
    .B(_0748_),
    .X(_0751_));
 sky130_fd_sc_hd__o211a_1 _4142_ (.A1(_0750_),
    .A2(_0749_),
    .B1(_0751_),
    .C1(_0719_),
    .X(\seq.player_4.next_state[2] ));
 sky130_fd_sc_hd__a31o_1 _4143_ (.A1(\seq.player_4.state[1] ),
    .A2(\seq.player_4.state[2] ),
    .A3(_0746_),
    .B1(\seq.player_4.state[3] ),
    .X(_0752_));
 sky130_fd_sc_hd__o211a_1 _4144_ (.A1(_0750_),
    .A2(_0749_),
    .B1(_0752_),
    .C1(_0719_),
    .X(\seq.player_4.next_state[3] ));
 sky130_fd_sc_hd__and2b_1 _4145_ (.A_N(\seq.encode.keys_edge_det[4] ),
    .B(\inputcont.INTERNAL_SYNCED_I[2] ),
    .X(_0753_));
 sky130_fd_sc_hd__and2_1 _4146_ (.A(\seq.player_3.state[0] ),
    .B(_0753_),
    .X(_0754_));
 sky130_fd_sc_hd__a311o_1 _4147_ (.A1(\seq.player_3.state[1] ),
    .A2(\seq.player_3.state[2] ),
    .A3(\seq.player_3.state[3] ),
    .B1(_0754_),
    .C1(_0700_),
    .X(_0755_));
 sky130_fd_sc_hd__o21ba_1 _4148_ (.A1(\seq.player_3.state[0] ),
    .A2(_0753_),
    .B1_N(_0755_),
    .X(\seq.player_3.next_state[0] ));
 sky130_fd_sc_hd__and3_1 _4149_ (.A(\seq.player_3.state[0] ),
    .B(\seq.player_3.state[1] ),
    .C(_0753_),
    .X(_0756_));
 sky130_fd_sc_hd__nor2_1 _4150_ (.A(\seq.player_3.state[1] ),
    .B(_0754_),
    .Y(_0757_));
 sky130_fd_sc_hd__a2111oi_1 _4151_ (.A1(\seq.player_3.state[2] ),
    .A2(\seq.player_3.state[3] ),
    .B1(_0756_),
    .C1(_0757_),
    .D1(_0700_),
    .Y(\seq.player_3.next_state[1] ));
 sky130_fd_sc_hd__nand2_1 _4152_ (.A(\seq.player_3.state[2] ),
    .B(\seq.player_3.state[3] ),
    .Y(_0758_));
 sky130_fd_sc_hd__xor2_1 _4153_ (.A(\seq.player_3.state[2] ),
    .B(_0756_),
    .X(_0759_));
 sky130_fd_sc_hd__o211a_1 _4154_ (.A1(_0758_),
    .A2(_0757_),
    .B1(_0759_),
    .C1(_0719_),
    .X(\seq.player_3.next_state[2] ));
 sky130_fd_sc_hd__a31o_1 _4155_ (.A1(\seq.player_3.state[1] ),
    .A2(\seq.player_3.state[2] ),
    .A3(_0754_),
    .B1(\seq.player_3.state[3] ),
    .X(_0760_));
 sky130_fd_sc_hd__o211a_1 _4156_ (.A1(_0758_),
    .A2(_0757_),
    .B1(_0760_),
    .C1(_0719_),
    .X(\seq.player_3.next_state[3] ));
 sky130_fd_sc_hd__nor2_1 _4157_ (.A(_0449_),
    .B(\seq.encode.keys_edge_det[3] ),
    .Y(_0761_));
 sky130_fd_sc_hd__and2_1 _4158_ (.A(\seq.player_2.state[0] ),
    .B(_0761_),
    .X(_0762_));
 sky130_fd_sc_hd__a311o_1 _4159_ (.A1(\seq.player_2.state[1] ),
    .A2(\seq.player_2.state[2] ),
    .A3(\seq.player_2.state[3] ),
    .B1(_0762_),
    .C1(_0700_),
    .X(_0763_));
 sky130_fd_sc_hd__o21ba_1 _4160_ (.A1(\seq.player_2.state[0] ),
    .A2(_0761_),
    .B1_N(_0763_),
    .X(\seq.player_2.next_state[0] ));
 sky130_fd_sc_hd__and3_1 _4161_ (.A(\seq.player_2.state[0] ),
    .B(\seq.player_2.state[1] ),
    .C(_0761_),
    .X(_0764_));
 sky130_fd_sc_hd__nor2_1 _4162_ (.A(\seq.player_2.state[1] ),
    .B(_0762_),
    .Y(_0765_));
 sky130_fd_sc_hd__a2111oi_1 _4163_ (.A1(\seq.player_2.state[2] ),
    .A2(\seq.player_2.state[3] ),
    .B1(_0764_),
    .C1(_0765_),
    .D1(_0700_),
    .Y(\seq.player_2.next_state[1] ));
 sky130_fd_sc_hd__nand2_1 _4164_ (.A(\seq.player_2.state[2] ),
    .B(\seq.player_2.state[3] ),
    .Y(_0766_));
 sky130_fd_sc_hd__xor2_1 _4165_ (.A(\seq.player_2.state[2] ),
    .B(_0764_),
    .X(_0767_));
 sky130_fd_sc_hd__o211a_1 _4166_ (.A1(_0766_),
    .A2(_0765_),
    .B1(_0767_),
    .C1(_0719_),
    .X(\seq.player_2.next_state[2] ));
 sky130_fd_sc_hd__a31o_1 _4167_ (.A1(\seq.player_2.state[1] ),
    .A2(\seq.player_2.state[2] ),
    .A3(_0762_),
    .B1(\seq.player_2.state[3] ),
    .X(_0768_));
 sky130_fd_sc_hd__o211a_1 _4168_ (.A1(_0766_),
    .A2(_0765_),
    .B1(_0768_),
    .C1(_0719_),
    .X(\seq.player_2.next_state[3] ));
 sky130_fd_sc_hd__and2b_1 _4169_ (.A_N(\seq.encode.keys_edge_det[2] ),
    .B(\inputcont.INTERNAL_SYNCED_I[0] ),
    .X(_0769_));
 sky130_fd_sc_hd__and2_1 _4170_ (.A(\seq.player_1.state[0] ),
    .B(_0769_),
    .X(_0770_));
 sky130_fd_sc_hd__a311o_1 _4171_ (.A1(\seq.player_1.state[1] ),
    .A2(\seq.player_1.state[2] ),
    .A3(\seq.player_1.state[3] ),
    .B1(_0770_),
    .C1(_0700_),
    .X(_0771_));
 sky130_fd_sc_hd__o21ba_1 _4172_ (.A1(\seq.player_1.state[0] ),
    .A2(_0769_),
    .B1_N(_0771_),
    .X(\seq.player_1.next_state[0] ));
 sky130_fd_sc_hd__and3_1 _4173_ (.A(\seq.player_1.state[0] ),
    .B(\seq.player_1.state[1] ),
    .C(_0769_),
    .X(_0772_));
 sky130_fd_sc_hd__nor2_1 _4174_ (.A(\seq.player_1.state[1] ),
    .B(_0770_),
    .Y(_0773_));
 sky130_fd_sc_hd__a2111oi_1 _4175_ (.A1(\seq.player_1.state[2] ),
    .A2(\seq.player_1.state[3] ),
    .B1(_0772_),
    .C1(_0773_),
    .D1(_0700_),
    .Y(\seq.player_1.next_state[1] ));
 sky130_fd_sc_hd__nand2_1 _4176_ (.A(\seq.player_1.state[2] ),
    .B(\seq.player_1.state[3] ),
    .Y(_0774_));
 sky130_fd_sc_hd__xor2_1 _4177_ (.A(\seq.player_1.state[2] ),
    .B(_0772_),
    .X(_0775_));
 sky130_fd_sc_hd__o211a_1 _4178_ (.A1(_0774_),
    .A2(_0773_),
    .B1(_0775_),
    .C1(_0719_),
    .X(\seq.player_1.next_state[2] ));
 sky130_fd_sc_hd__a31o_1 _4179_ (.A1(\seq.player_1.state[1] ),
    .A2(\seq.player_1.state[2] ),
    .A3(_0770_),
    .B1(\seq.player_1.state[3] ),
    .X(_0776_));
 sky130_fd_sc_hd__o211a_1 _4180_ (.A1(_0774_),
    .A2(_0773_),
    .B1(_0776_),
    .C1(_0719_),
    .X(\seq.player_1.next_state[3] ));
 sky130_fd_sc_hd__nor2_1 _4181_ (.A(_0700_),
    .B(\seq.clk_div.count[0] ),
    .Y(\seq.clk_div.next_count[0] ));
 sky130_fd_sc_hd__and2_1 _4182_ (.A(\seq.clk_div.count[1] ),
    .B(\seq.clk_div.count[0] ),
    .X(_0777_));
 sky130_fd_sc_hd__o21ai_1 _4183_ (.A1(\seq.clk_div.count[1] ),
    .A2(\seq.clk_div.count[0] ),
    .B1(_0719_),
    .Y(_0778_));
 sky130_fd_sc_hd__nor2_1 _4184_ (.A(_0777_),
    .B(_0778_),
    .Y(\seq.clk_div.next_count[1] ));
 sky130_fd_sc_hd__inv_2 _4185_ (.A(\seq.clk_div.count[18] ),
    .Y(_0779_));
 sky130_fd_sc_hd__inv_2 _4186_ (.A(\seq.clk_div.count[10] ),
    .Y(_0780_));
 sky130_fd_sc_hd__o2111a_1 _4187_ (.A1(\seq.tempo_select.state[1] ),
    .A2(\seq.clk_div.count[12] ),
    .B1(_0779_),
    .C1(\seq.clk_div.count[6] ),
    .D1(_0780_),
    .X(_0781_));
 sky130_fd_sc_hd__or2b_1 _4188_ (.A(\seq.tempo_select.state[1] ),
    .B_N(\seq.tempo_select.state[0] ),
    .X(_0782_));
 sky130_fd_sc_hd__or4bb_1 _4189_ (.A(\seq.clk_div.count[5] ),
    .B(\seq.clk_div.count[15] ),
    .C_N(\seq.clk_div.count[17] ),
    .D_N(\seq.clk_div.count[3] ),
    .X(_0783_));
 sky130_fd_sc_hd__a21oi_1 _4190_ (.A1(\seq.clk_div.count[19] ),
    .A2(_0782_),
    .B1(_0783_),
    .Y(_0784_));
 sky130_fd_sc_hd__and2b_1 _4191_ (.A_N(\seq.tempo_select.state[0] ),
    .B(\seq.tempo_select.state[1] ),
    .X(_0785_));
 sky130_fd_sc_hd__o22ai_1 _4192_ (.A1(\seq.tempo_select.state[0] ),
    .A2(_0781_),
    .B1(_0784_),
    .B2(_0785_),
    .Y(_0786_));
 sky130_fd_sc_hd__nand2_1 _4193_ (.A(\seq.tempo_select.state[0] ),
    .B(\seq.clk_div.count[4] ),
    .Y(_0787_));
 sky130_fd_sc_hd__or4_1 _4194_ (.A(\seq.clk_div.count[6] ),
    .B(\seq.clk_div.count[12] ),
    .C(\seq.clk_div.count[16] ),
    .D(_0779_),
    .X(_0788_));
 sky130_fd_sc_hd__inv_2 _4195_ (.A(\seq.clk_div.count[2] ),
    .Y(_0789_));
 sky130_fd_sc_hd__a21oi_1 _4196_ (.A1(_0789_),
    .A2(\seq.clk_div.count[14] ),
    .B1(\seq.tempo_select.state[1] ),
    .Y(_0790_));
 sky130_fd_sc_hd__inv_2 _4197_ (.A(\seq.clk_div.count[20] ),
    .Y(_0791_));
 sky130_fd_sc_hd__nand2_1 _4198_ (.A(\seq.tempo_select.state[1] ),
    .B(\seq.clk_div.count[5] ),
    .Y(_0792_));
 sky130_fd_sc_hd__o22a_1 _4199_ (.A1(\seq.tempo_select.state[1] ),
    .A2(_0791_),
    .B1(_0792_),
    .B2(\seq.clk_div.count[12] ),
    .X(_0793_));
 sky130_fd_sc_hd__or3b_1 _4200_ (.A(\seq.tempo_select.state[0] ),
    .B(\seq.clk_div.count[4] ),
    .C_N(\seq.clk_div.count[16] ),
    .X(_0794_));
 sky130_fd_sc_hd__o32a_1 _4201_ (.A1(_0787_),
    .A2(_0788_),
    .A3(_0790_),
    .B1(_0793_),
    .B2(_0794_),
    .X(_0795_));
 sky130_fd_sc_hd__inv_2 _4202_ (.A(\seq.clk_div.count[7] ),
    .Y(_0796_));
 sky130_fd_sc_hd__o22a_1 _4203_ (.A1(\seq.clk_div.count[20] ),
    .A2(_0664_),
    .B1(_0665_),
    .B2(\seq.clk_div.count[21] ),
    .X(_0797_));
 sky130_fd_sc_hd__or4bb_1 _4204_ (.A(\seq.clk_div.count[3] ),
    .B(\seq.clk_div.count[17] ),
    .C_N(_0785_),
    .D_N(\seq.clk_div.count[15] ),
    .X(_0798_));
 sky130_fd_sc_hd__nand2_1 _4205_ (.A(\seq.clk_div.count[11] ),
    .B(\seq.clk_div.count[19] ),
    .Y(_0799_));
 sky130_fd_sc_hd__a2111o_1 _4206_ (.A1(_0782_),
    .A2(_0798_),
    .B1(_0799_),
    .C1(\seq.clk_div.count[21] ),
    .D1(\seq.clk_div.count[20] ),
    .X(_0800_));
 sky130_fd_sc_hd__o21ai_1 _4207_ (.A1(_0796_),
    .A2(_0797_),
    .B1(_0800_),
    .Y(_0801_));
 sky130_fd_sc_hd__inv_2 _4208_ (.A(\seq.clk_div.count[13] ),
    .Y(_0802_));
 sky130_fd_sc_hd__o2bb2a_1 _4209_ (.A1_N(\seq.clk_div.count[7] ),
    .A2_N(\seq.clk_div.count[11] ),
    .B1(_0802_),
    .B2(\seq.clk_div.count[21] ),
    .X(_0803_));
 sky130_fd_sc_hd__o211a_1 _4210_ (.A1(\seq.clk_div.count[10] ),
    .A2(_0779_),
    .B1(_0777_),
    .C1(_0803_),
    .X(_0804_));
 sky130_fd_sc_hd__o21ai_1 _4211_ (.A1(_0789_),
    .A2(\seq.clk_div.count[14] ),
    .B1(_0782_),
    .Y(_0805_));
 sky130_fd_sc_hd__inv_2 _4212_ (.A(\seq.clk_div.count[8] ),
    .Y(_0806_));
 sky130_fd_sc_hd__a211o_1 _4213_ (.A1(\seq.tempo_select.state[0] ),
    .A2(_0802_),
    .B1(\seq.clk_div.count[9] ),
    .C1(_0806_),
    .X(_0807_));
 sky130_fd_sc_hd__nand2_1 _4214_ (.A(\seq.tempo_select.state[1] ),
    .B(_0807_),
    .Y(_0808_));
 sky130_fd_sc_hd__a21o_1 _4215_ (.A1(_0806_),
    .A2(\seq.clk_div.count[9] ),
    .B1(\seq.tempo_select.state[1] ),
    .X(_0809_));
 sky130_fd_sc_hd__and4_1 _4216_ (.A(_0804_),
    .B(_0805_),
    .C(_0808_),
    .D(_0809_),
    .X(_0810_));
 sky130_fd_sc_hd__or4bb_1 _4217_ (.A(_0786_),
    .B(_0795_),
    .C_N(_0801_),
    .D_N(_0810_),
    .X(_0811_));
 sky130_fd_sc_hd__and2_1 _4218_ (.A(_0719_),
    .B(_0811_),
    .X(_0812_));
 sky130_fd_sc_hd__buf_4 _4219_ (.A(_0812_),
    .X(_0813_));
 sky130_fd_sc_hd__o21ai_1 _4220_ (.A1(\seq.clk_div.count[2] ),
    .A2(_0777_),
    .B1(_0813_),
    .Y(_0814_));
 sky130_fd_sc_hd__a21oi_1 _4221_ (.A1(\seq.clk_div.count[2] ),
    .A2(_0777_),
    .B1(_0814_),
    .Y(\seq.clk_div.next_count[2] ));
 sky130_fd_sc_hd__and3_1 _4222_ (.A(\seq.clk_div.count[2] ),
    .B(\seq.clk_div.count[3] ),
    .C(_0777_),
    .X(_0815_));
 sky130_fd_sc_hd__a31o_1 _4223_ (.A1(\seq.clk_div.count[1] ),
    .A2(\seq.clk_div.count[0] ),
    .A3(\seq.clk_div.count[2] ),
    .B1(\seq.clk_div.count[3] ),
    .X(_0816_));
 sky130_fd_sc_hd__and3b_1 _4224_ (.A_N(_0815_),
    .B(_0816_),
    .C(_0813_),
    .X(_0817_));
 sky130_fd_sc_hd__clkbuf_1 _4225_ (.A(_0817_),
    .X(\seq.clk_div.next_count[3] ));
 sky130_fd_sc_hd__o21ai_1 _4226_ (.A1(\seq.clk_div.count[4] ),
    .A2(_0815_),
    .B1(_0813_),
    .Y(_0818_));
 sky130_fd_sc_hd__a21oi_1 _4227_ (.A1(\seq.clk_div.count[4] ),
    .A2(_0815_),
    .B1(_0818_),
    .Y(\seq.clk_div.next_count[4] ));
 sky130_fd_sc_hd__and3_1 _4228_ (.A(\seq.clk_div.count[4] ),
    .B(\seq.clk_div.count[5] ),
    .C(_0815_),
    .X(_0819_));
 sky130_fd_sc_hd__a21o_1 _4229_ (.A1(\seq.clk_div.count[4] ),
    .A2(_0815_),
    .B1(\seq.clk_div.count[5] ),
    .X(_0820_));
 sky130_fd_sc_hd__and3b_1 _4230_ (.A_N(_0819_),
    .B(_0820_),
    .C(_0813_),
    .X(_0821_));
 sky130_fd_sc_hd__clkbuf_1 _4231_ (.A(_0821_),
    .X(\seq.clk_div.next_count[5] ));
 sky130_fd_sc_hd__and2_1 _4232_ (.A(\seq.clk_div.count[6] ),
    .B(_0819_),
    .X(_0822_));
 sky130_fd_sc_hd__o21ai_1 _4233_ (.A1(\seq.clk_div.count[6] ),
    .A2(_0819_),
    .B1(_0813_),
    .Y(_0823_));
 sky130_fd_sc_hd__nor2_1 _4234_ (.A(_0822_),
    .B(_0823_),
    .Y(\seq.clk_div.next_count[6] ));
 sky130_fd_sc_hd__and3_1 _4235_ (.A(\seq.clk_div.count[6] ),
    .B(\seq.clk_div.count[7] ),
    .C(_0819_),
    .X(_0824_));
 sky130_fd_sc_hd__o21ai_1 _4236_ (.A1(\seq.clk_div.count[7] ),
    .A2(_0822_),
    .B1(_0813_),
    .Y(_0825_));
 sky130_fd_sc_hd__nor2_1 _4237_ (.A(_0824_),
    .B(_0825_),
    .Y(\seq.clk_div.next_count[7] ));
 sky130_fd_sc_hd__or2_1 _4238_ (.A(\seq.clk_div.count[8] ),
    .B(_0824_),
    .X(_0826_));
 sky130_fd_sc_hd__nand2_1 _4239_ (.A(\seq.clk_div.count[8] ),
    .B(_0824_),
    .Y(_0827_));
 sky130_fd_sc_hd__and3_1 _4240_ (.A(_0813_),
    .B(_0826_),
    .C(_0827_),
    .X(_0828_));
 sky130_fd_sc_hd__clkbuf_1 _4241_ (.A(_0828_),
    .X(\seq.clk_div.next_count[8] ));
 sky130_fd_sc_hd__and3_1 _4242_ (.A(\seq.clk_div.count[8] ),
    .B(\seq.clk_div.count[9] ),
    .C(_0824_),
    .X(_0829_));
 sky130_fd_sc_hd__a21o_1 _4243_ (.A1(\seq.clk_div.count[8] ),
    .A2(_0824_),
    .B1(\seq.clk_div.count[9] ),
    .X(_0830_));
 sky130_fd_sc_hd__and3b_1 _4244_ (.A_N(_0829_),
    .B(_0813_),
    .C(_0830_),
    .X(_0831_));
 sky130_fd_sc_hd__clkbuf_1 _4245_ (.A(_0831_),
    .X(\seq.clk_div.next_count[9] ));
 sky130_fd_sc_hd__and4_1 _4246_ (.A(\seq.clk_div.count[8] ),
    .B(\seq.clk_div.count[9] ),
    .C(\seq.clk_div.count[10] ),
    .D(_0824_),
    .X(_0832_));
 sky130_fd_sc_hd__or2_1 _4247_ (.A(\seq.clk_div.count[10] ),
    .B(_0829_),
    .X(_0833_));
 sky130_fd_sc_hd__and3b_1 _4248_ (.A_N(_0832_),
    .B(_0813_),
    .C(_0833_),
    .X(_0834_));
 sky130_fd_sc_hd__clkbuf_1 _4249_ (.A(_0834_),
    .X(\seq.clk_div.next_count[10] ));
 sky130_fd_sc_hd__and3_1 _4250_ (.A(\seq.clk_div.count[10] ),
    .B(\seq.clk_div.count[11] ),
    .C(_0829_),
    .X(_0835_));
 sky130_fd_sc_hd__or2_1 _4251_ (.A(\seq.clk_div.count[11] ),
    .B(_0832_),
    .X(_0836_));
 sky130_fd_sc_hd__and3b_1 _4252_ (.A_N(_0835_),
    .B(_0813_),
    .C(_0836_),
    .X(_0837_));
 sky130_fd_sc_hd__clkbuf_1 _4253_ (.A(_0837_),
    .X(\seq.clk_div.next_count[11] ));
 sky130_fd_sc_hd__and2_1 _4254_ (.A(\seq.clk_div.count[12] ),
    .B(_0835_),
    .X(_0838_));
 sky130_fd_sc_hd__or2_1 _4255_ (.A(\seq.clk_div.count[12] ),
    .B(_0835_),
    .X(_0839_));
 sky130_fd_sc_hd__and3b_1 _4256_ (.A_N(_0838_),
    .B(_0813_),
    .C(_0839_),
    .X(_0840_));
 sky130_fd_sc_hd__clkbuf_1 _4257_ (.A(_0840_),
    .X(\seq.clk_div.next_count[12] ));
 sky130_fd_sc_hd__and4_1 _4258_ (.A(\seq.clk_div.count[11] ),
    .B(\seq.clk_div.count[12] ),
    .C(\seq.clk_div.count[13] ),
    .D(_0832_),
    .X(_0841_));
 sky130_fd_sc_hd__or2_1 _4259_ (.A(\seq.clk_div.count[13] ),
    .B(_0838_),
    .X(_0842_));
 sky130_fd_sc_hd__and3b_1 _4260_ (.A_N(_0841_),
    .B(_0813_),
    .C(_0842_),
    .X(_0843_));
 sky130_fd_sc_hd__clkbuf_1 _4261_ (.A(_0843_),
    .X(\seq.clk_div.next_count[13] ));
 sky130_fd_sc_hd__and3_1 _4262_ (.A(\seq.clk_div.count[13] ),
    .B(\seq.clk_div.count[14] ),
    .C(_0838_),
    .X(_0844_));
 sky130_fd_sc_hd__or2_1 _4263_ (.A(\seq.clk_div.count[14] ),
    .B(_0841_),
    .X(_0845_));
 sky130_fd_sc_hd__and3b_1 _4264_ (.A_N(_0844_),
    .B(_0813_),
    .C(_0845_),
    .X(_0846_));
 sky130_fd_sc_hd__clkbuf_1 _4265_ (.A(_0846_),
    .X(\seq.clk_div.next_count[14] ));
 sky130_fd_sc_hd__and3_1 _4266_ (.A(\seq.clk_div.count[14] ),
    .B(\seq.clk_div.count[15] ),
    .C(_0841_),
    .X(_0847_));
 sky130_fd_sc_hd__or2_1 _4267_ (.A(\seq.clk_div.count[15] ),
    .B(_0844_),
    .X(_0848_));
 sky130_fd_sc_hd__and3b_1 _4268_ (.A_N(_0847_),
    .B(_0813_),
    .C(_0848_),
    .X(_0849_));
 sky130_fd_sc_hd__clkbuf_1 _4269_ (.A(_0849_),
    .X(\seq.clk_div.next_count[15] ));
 sky130_fd_sc_hd__and2_1 _4270_ (.A(\seq.clk_div.count[16] ),
    .B(_0847_),
    .X(_0850_));
 sky130_fd_sc_hd__or2_1 _4271_ (.A(\seq.clk_div.count[16] ),
    .B(_0847_),
    .X(_0851_));
 sky130_fd_sc_hd__and3b_1 _4272_ (.A_N(_0850_),
    .B(_0813_),
    .C(_0851_),
    .X(_0852_));
 sky130_fd_sc_hd__clkbuf_1 _4273_ (.A(_0852_),
    .X(\seq.clk_div.next_count[16] ));
 sky130_fd_sc_hd__and4_1 _4274_ (.A(\seq.clk_div.count[15] ),
    .B(\seq.clk_div.count[16] ),
    .C(\seq.clk_div.count[17] ),
    .D(_0844_),
    .X(_0853_));
 sky130_fd_sc_hd__inv_2 _4275_ (.A(_0853_),
    .Y(_0854_));
 sky130_fd_sc_hd__o211a_1 _4276_ (.A1(\seq.clk_div.count[17] ),
    .A2(_0850_),
    .B1(_0854_),
    .C1(_0813_),
    .X(\seq.clk_div.next_count[17] ));
 sky130_fd_sc_hd__and3_1 _4277_ (.A(\seq.clk_div.count[17] ),
    .B(\seq.clk_div.count[18] ),
    .C(_0850_),
    .X(_0855_));
 sky130_fd_sc_hd__or2_1 _4278_ (.A(\seq.clk_div.count[18] ),
    .B(_0853_),
    .X(_0856_));
 sky130_fd_sc_hd__and3b_1 _4279_ (.A_N(_0855_),
    .B(_0813_),
    .C(_0856_),
    .X(_0857_));
 sky130_fd_sc_hd__clkbuf_1 _4280_ (.A(_0857_),
    .X(\seq.clk_div.next_count[18] ));
 sky130_fd_sc_hd__nand3_1 _4281_ (.A(\seq.clk_div.count[18] ),
    .B(\seq.clk_div.count[19] ),
    .C(_0853_),
    .Y(_0858_));
 sky130_fd_sc_hd__o211a_1 _4282_ (.A1(\seq.clk_div.count[19] ),
    .A2(_0855_),
    .B1(_0858_),
    .C1(_0813_),
    .X(\seq.clk_div.next_count[19] ));
 sky130_fd_sc_hd__nor2_1 _4283_ (.A(_0791_),
    .B(_0858_),
    .Y(_0859_));
 sky130_fd_sc_hd__nand2_1 _4284_ (.A(_0791_),
    .B(_0858_),
    .Y(_0860_));
 sky130_fd_sc_hd__and3b_1 _4285_ (.A_N(_0859_),
    .B(_0813_),
    .C(_0860_),
    .X(_0861_));
 sky130_fd_sc_hd__clkbuf_1 _4286_ (.A(_0861_),
    .X(\seq.clk_div.next_count[20] ));
 sky130_fd_sc_hd__o21ai_1 _4287_ (.A1(\seq.clk_div.count[21] ),
    .A2(_0859_),
    .B1(_0813_),
    .Y(_0862_));
 sky130_fd_sc_hd__a21oi_1 _4288_ (.A1(\seq.clk_div.count[21] ),
    .A2(_0859_),
    .B1(_0862_),
    .Y(\seq.clk_div.next_count[21] ));
 sky130_fd_sc_hd__or2b_1 _4289_ (.A(\seq.encode.keys_edge_det[0] ),
    .B_N(\seq.encode.keys_sync[0] ),
    .X(_0863_));
 sky130_fd_sc_hd__xnor2_1 _4290_ (.A(\seq.encode.play ),
    .B(_0863_),
    .Y(\seq.encode.next_play ));
 sky130_fd_sc_hd__and2b_1 _4291_ (.A_N(\seq.encode.keys_edge_det[1] ),
    .B(\seq.encode.keys_sync[1] ),
    .X(_0864_));
 sky130_fd_sc_hd__xnor2_1 _4292_ (.A(_0700_),
    .B(_0864_),
    .Y(\seq.encode.next_sequencer_on ));
 sky130_fd_sc_hd__or2_1 _4293_ (.A(_0575_),
    .B(_0566_),
    .X(_0865_));
 sky130_fd_sc_hd__clkbuf_8 _4294_ (.A(_0865_),
    .X(_0866_));
 sky130_fd_sc_hd__inv_4 _4295_ (.A(_0866_),
    .Y(_0867_));
 sky130_fd_sc_hd__buf_4 _4296_ (.A(_0867_),
    .X(\sound1.sdiv.next_dived ));
 sky130_fd_sc_hd__or2_1 _4297_ (.A(_0674_),
    .B(_0677_),
    .X(_0868_));
 sky130_fd_sc_hd__buf_6 _4298_ (.A(_0868_),
    .X(_0869_));
 sky130_fd_sc_hd__nor3_1 _4299_ (.A(\seq.beat[1] ),
    .B(\seq.beat[0] ),
    .C(\seq.beat[2] ),
    .Y(_0870_));
 sky130_fd_sc_hd__a31o_2 _4300_ (.A1(_0702_),
    .A2(\seq.encode.play ),
    .A3(_0870_),
    .B1(\inputcont.INTERNAL_SYNCED_I[0] ),
    .X(_0871_));
 sky130_fd_sc_hd__o41a_1 _4301_ (.A1(\seq.player_1.state[0] ),
    .A2(\seq.player_1.state[1] ),
    .A3(\seq.player_1.state[2] ),
    .A4(\seq.player_1.state[3] ),
    .B1(_0698_),
    .X(_0872_));
 sky130_fd_sc_hd__nand2_1 _4302_ (.A(_0871_),
    .B(_0872_),
    .Y(_0873_));
 sky130_fd_sc_hd__nor3b_1 _4303_ (.A(\seq.beat[0] ),
    .B(\seq.beat[2] ),
    .C_N(\seq.beat[1] ),
    .Y(_0874_));
 sky130_fd_sc_hd__a31o_1 _4304_ (.A1(_0702_),
    .A2(\seq.encode.play ),
    .A3(_0874_),
    .B1(\inputcont.INTERNAL_SYNCED_I[1] ),
    .X(_0875_));
 sky130_fd_sc_hd__and2_1 _4305_ (.A(\select1.sequencer_on ),
    .B(_0875_),
    .X(_0876_));
 sky130_fd_sc_hd__or4_1 _4306_ (.A(\seq.player_2.state[0] ),
    .B(\seq.player_2.state[1] ),
    .C(\seq.player_2.state[2] ),
    .D(\seq.player_2.state[3] ),
    .X(_0877_));
 sky130_fd_sc_hd__nand2_1 _4307_ (.A(_0876_),
    .B(_0877_),
    .Y(_0878_));
 sky130_fd_sc_hd__nor3b_1 _4308_ (.A(\seq.beat[1] ),
    .B(\seq.beat[0] ),
    .C_N(\seq.beat[2] ),
    .Y(_0879_));
 sky130_fd_sc_hd__a31o_1 _4309_ (.A1(_0702_),
    .A2(\seq.encode.play ),
    .A3(_0879_),
    .B1(\inputcont.INTERNAL_SYNCED_I[2] ),
    .X(_0880_));
 sky130_fd_sc_hd__and2_1 _4310_ (.A(\select1.sequencer_on ),
    .B(_0880_),
    .X(_0881_));
 sky130_fd_sc_hd__or4_1 _4311_ (.A(\seq.player_3.state[0] ),
    .B(\seq.player_3.state[1] ),
    .C(\seq.player_3.state[2] ),
    .D(\seq.player_3.state[3] ),
    .X(_0882_));
 sky130_fd_sc_hd__nand2_1 _4312_ (.A(_0881_),
    .B(_0882_),
    .Y(_0883_));
 sky130_fd_sc_hd__and3b_1 _4313_ (.A_N(\seq.beat[0] ),
    .B(\seq.beat[2] ),
    .C(\seq.beat[1] ),
    .X(_0884_));
 sky130_fd_sc_hd__a31o_1 _4314_ (.A1(_0702_),
    .A2(\seq.encode.play ),
    .A3(_0884_),
    .B1(\inputcont.INTERNAL_SYNCED_I[3] ),
    .X(_0885_));
 sky130_fd_sc_hd__and2_1 _4315_ (.A(\select1.sequencer_on ),
    .B(_0885_),
    .X(_0886_));
 sky130_fd_sc_hd__or4_1 _4316_ (.A(\seq.player_4.state[0] ),
    .B(\seq.player_4.state[1] ),
    .C(\seq.player_4.state[2] ),
    .D(\seq.player_4.state[3] ),
    .X(_0887_));
 sky130_fd_sc_hd__nand2_1 _4317_ (.A(_0886_),
    .B(_0887_),
    .Y(_0888_));
 sky130_fd_sc_hd__a31o_1 _4318_ (.A1(\seq.beat[3] ),
    .A2(\seq.encode.play ),
    .A3(_0870_),
    .B1(\inputcont.INTERNAL_SYNCED_I[4] ),
    .X(_0889_));
 sky130_fd_sc_hd__and2_1 _4319_ (.A(\select1.sequencer_on ),
    .B(_0889_),
    .X(_0890_));
 sky130_fd_sc_hd__or4_1 _4320_ (.A(\seq.player_5.state[0] ),
    .B(\seq.player_5.state[1] ),
    .C(\seq.player_5.state[2] ),
    .D(\seq.player_5.state[3] ),
    .X(_0891_));
 sky130_fd_sc_hd__nand2_1 _4321_ (.A(_0890_),
    .B(_0891_),
    .Y(_0892_));
 sky130_fd_sc_hd__a31o_1 _4322_ (.A1(\seq.beat[3] ),
    .A2(\seq.encode.play ),
    .A3(_0874_),
    .B1(\inputcont.INTERNAL_SYNCED_I[5] ),
    .X(_0893_));
 sky130_fd_sc_hd__and2_1 _4323_ (.A(\select1.sequencer_on ),
    .B(_0893_),
    .X(_0894_));
 sky130_fd_sc_hd__or4_1 _4324_ (.A(\seq.player_6.state[0] ),
    .B(\seq.player_6.state[1] ),
    .C(\seq.player_6.state[2] ),
    .D(\seq.player_6.state[3] ),
    .X(_0895_));
 sky130_fd_sc_hd__nand2_1 _4325_ (.A(_0894_),
    .B(_0895_),
    .Y(_0896_));
 sky130_fd_sc_hd__a31o_1 _4326_ (.A1(\seq.beat[3] ),
    .A2(\seq.encode.play ),
    .A3(_0879_),
    .B1(\inputcont.INTERNAL_SYNCED_I[6] ),
    .X(_0897_));
 sky130_fd_sc_hd__and2_1 _4327_ (.A(\select1.sequencer_on ),
    .B(_0897_),
    .X(_0898_));
 sky130_fd_sc_hd__or4_1 _4328_ (.A(\seq.player_7.state[0] ),
    .B(\seq.player_7.state[1] ),
    .C(\seq.player_7.state[2] ),
    .D(\seq.player_7.state[3] ),
    .X(_0899_));
 sky130_fd_sc_hd__a31oi_1 _4329_ (.A1(\seq.beat[3] ),
    .A2(\seq.encode.play ),
    .A3(_0884_),
    .B1(\inputcont.INTERNAL_SYNCED_I[7] ),
    .Y(_0900_));
 sky130_fd_sc_hd__a31oi_2 _4330_ (.A1(\select1.sequencer_on ),
    .A2(_0897_),
    .A3(_0899_),
    .B1(_0900_),
    .Y(_0901_));
 sky130_fd_sc_hd__a22o_1 _4331_ (.A1(\seq.player_7.state[1] ),
    .A2(_0898_),
    .B1(_0901_),
    .B2(\seq.player_8.state[1] ),
    .X(_0902_));
 sky130_fd_sc_hd__a22o_1 _4332_ (.A1(\seq.player_6.state[1] ),
    .A2(_0894_),
    .B1(_0896_),
    .B2(_0902_),
    .X(_0903_));
 sky130_fd_sc_hd__a22o_1 _4333_ (.A1(\seq.player_5.state[1] ),
    .A2(_0890_),
    .B1(_0892_),
    .B2(_0903_),
    .X(_0904_));
 sky130_fd_sc_hd__a22o_1 _4334_ (.A1(\seq.player_4.state[1] ),
    .A2(_0886_),
    .B1(_0888_),
    .B2(_0904_),
    .X(_0905_));
 sky130_fd_sc_hd__a22o_1 _4335_ (.A1(\seq.player_3.state[1] ),
    .A2(_0881_),
    .B1(_0883_),
    .B2(_0905_),
    .X(_0906_));
 sky130_fd_sc_hd__a22o_1 _4336_ (.A1(\seq.player_2.state[1] ),
    .A2(_0876_),
    .B1(_0878_),
    .B2(_0906_),
    .X(_0907_));
 sky130_fd_sc_hd__a22o_1 _4337_ (.A1(\seq.player_1.state[1] ),
    .A2(_0871_),
    .B1(_0873_),
    .B2(_0907_),
    .X(_0908_));
 sky130_fd_sc_hd__mux2_4 _4338_ (.A0(net36),
    .A1(_0908_),
    .S(_0698_),
    .X(_0909_));
 sky130_fd_sc_hd__a22o_1 _4339_ (.A1(\seq.player_7.state[0] ),
    .A2(_0898_),
    .B1(_0901_),
    .B2(\seq.player_8.state[0] ),
    .X(_0910_));
 sky130_fd_sc_hd__a22o_1 _4340_ (.A1(\seq.player_6.state[0] ),
    .A2(_0894_),
    .B1(_0896_),
    .B2(_0910_),
    .X(_0911_));
 sky130_fd_sc_hd__a22o_1 _4341_ (.A1(\seq.player_5.state[0] ),
    .A2(_0890_),
    .B1(_0892_),
    .B2(_0911_),
    .X(_0912_));
 sky130_fd_sc_hd__a22o_1 _4342_ (.A1(\seq.player_4.state[0] ),
    .A2(_0886_),
    .B1(_0888_),
    .B2(_0912_),
    .X(_0913_));
 sky130_fd_sc_hd__a22o_1 _4343_ (.A1(\seq.player_3.state[0] ),
    .A2(_0881_),
    .B1(_0883_),
    .B2(_0913_),
    .X(_0914_));
 sky130_fd_sc_hd__a22o_1 _4344_ (.A1(\seq.player_2.state[0] ),
    .A2(_0876_),
    .B1(_0878_),
    .B2(_0914_),
    .X(_0915_));
 sky130_fd_sc_hd__a22o_1 _4345_ (.A1(\seq.player_1.state[0] ),
    .A2(_0871_),
    .B1(_0873_),
    .B2(_0915_),
    .X(_0916_));
 sky130_fd_sc_hd__nand2_1 _4346_ (.A(_0698_),
    .B(_0916_),
    .Y(_0917_));
 sky130_fd_sc_hd__a21boi_4 _4347_ (.A1(_0699_),
    .A2(net35),
    .B1_N(_0917_),
    .Y(_0918_));
 sky130_fd_sc_hd__a22o_1 _4348_ (.A1(\seq.player_7.state[2] ),
    .A2(_0898_),
    .B1(_0901_),
    .B2(\seq.player_8.state[2] ),
    .X(_0919_));
 sky130_fd_sc_hd__a22o_1 _4349_ (.A1(\seq.player_6.state[2] ),
    .A2(_0894_),
    .B1(_0896_),
    .B2(_0919_),
    .X(_0920_));
 sky130_fd_sc_hd__a22o_1 _4350_ (.A1(\seq.player_5.state[2] ),
    .A2(_0890_),
    .B1(_0892_),
    .B2(_0920_),
    .X(_0921_));
 sky130_fd_sc_hd__a22o_1 _4351_ (.A1(\seq.player_4.state[2] ),
    .A2(_0886_),
    .B1(_0888_),
    .B2(_0921_),
    .X(_0922_));
 sky130_fd_sc_hd__a22o_1 _4352_ (.A1(\seq.player_3.state[2] ),
    .A2(_0881_),
    .B1(_0883_),
    .B2(_0922_),
    .X(_0923_));
 sky130_fd_sc_hd__a22o_1 _4353_ (.A1(\seq.player_2.state[2] ),
    .A2(_0876_),
    .B1(_0878_),
    .B2(_0923_),
    .X(_0924_));
 sky130_fd_sc_hd__a22o_1 _4354_ (.A1(\seq.player_1.state[2] ),
    .A2(_0871_),
    .B1(_0873_),
    .B2(_0924_),
    .X(_0925_));
 sky130_fd_sc_hd__mux2_2 _4355_ (.A0(net37),
    .A1(_0925_),
    .S(_0698_),
    .X(_0926_));
 sky130_fd_sc_hd__a22o_1 _4356_ (.A1(\seq.player_7.state[3] ),
    .A2(_0897_),
    .B1(_0901_),
    .B2(\seq.player_8.state[3] ),
    .X(_0927_));
 sky130_fd_sc_hd__and3_1 _4357_ (.A(\select1.sequencer_on ),
    .B(_0896_),
    .C(_0927_),
    .X(_0928_));
 sky130_fd_sc_hd__and3_1 _4358_ (.A(\select1.sequencer_on ),
    .B(\seq.player_6.state[3] ),
    .C(_0893_),
    .X(_0929_));
 sky130_fd_sc_hd__o21a_1 _4359_ (.A1(_0928_),
    .A2(_0929_),
    .B1(_0892_),
    .X(_0930_));
 sky130_fd_sc_hd__a22o_1 _4360_ (.A1(_0886_),
    .A2(_0887_),
    .B1(_0890_),
    .B2(\seq.player_5.state[3] ),
    .X(_0931_));
 sky130_fd_sc_hd__o221a_1 _4361_ (.A1(\seq.player_4.state[3] ),
    .A2(_0888_),
    .B1(_0930_),
    .B2(_0931_),
    .C1(_0883_),
    .X(_0932_));
 sky130_fd_sc_hd__a22o_1 _4362_ (.A1(_0876_),
    .A2(_0877_),
    .B1(_0881_),
    .B2(\seq.player_3.state[3] ),
    .X(_0933_));
 sky130_fd_sc_hd__o221a_1 _4363_ (.A1(\seq.player_2.state[3] ),
    .A2(_0878_),
    .B1(_0932_),
    .B2(_0933_),
    .C1(_0873_),
    .X(_0934_));
 sky130_fd_sc_hd__and3_1 _4364_ (.A(_0698_),
    .B(\seq.player_1.state[3] ),
    .C(_0871_),
    .X(_0935_));
 sky130_fd_sc_hd__a211oi_4 _4365_ (.A1(_0699_),
    .A2(net38),
    .B1(_0934_),
    .C1(_0935_),
    .Y(_0936_));
 sky130_fd_sc_hd__nand2_2 _4366_ (.A(_0926_),
    .B(_0936_),
    .Y(_0937_));
 sky130_fd_sc_hd__or3_1 _4367_ (.A(_0909_),
    .B(_0918_),
    .C(_0937_),
    .X(_0938_));
 sky130_fd_sc_hd__clkbuf_8 _4368_ (.A(_0938_),
    .X(_0939_));
 sky130_fd_sc_hd__a21bo_2 _4369_ (.A1(_0699_),
    .A2(net35),
    .B1_N(_0917_),
    .X(_0940_));
 sky130_fd_sc_hd__or2b_1 _4370_ (.A(_0937_),
    .B_N(_0909_),
    .X(_0941_));
 sky130_fd_sc_hd__or2_1 _4371_ (.A(_0940_),
    .B(_0941_),
    .X(_0942_));
 sky130_fd_sc_hd__buf_4 _4372_ (.A(_0942_),
    .X(_0943_));
 sky130_fd_sc_hd__nor2_8 _4373_ (.A(_0674_),
    .B(_0677_),
    .Y(_0944_));
 sky130_fd_sc_hd__nor2_4 _4374_ (.A(_0686_),
    .B(_0680_),
    .Y(_0945_));
 sky130_fd_sc_hd__nor2_8 _4375_ (.A(_0945_),
    .B(net64),
    .Y(_0946_));
 sky130_fd_sc_hd__nor2_4 _4376_ (.A(_0675_),
    .B(_0946_),
    .Y(_0947_));
 sky130_fd_sc_hd__or2_4 _4377_ (.A(_0944_),
    .B(_0947_),
    .X(_0948_));
 sky130_fd_sc_hd__nor2_2 _4378_ (.A(_0926_),
    .B(_0936_),
    .Y(_0949_));
 sky130_fd_sc_hd__nand3_4 _4379_ (.A(_0949_),
    .B(_0909_),
    .C(_0940_),
    .Y(_0950_));
 sky130_fd_sc_hd__nor2_1 _4380_ (.A(_0686_),
    .B(_0675_),
    .Y(_0951_));
 sky130_fd_sc_hd__nor2_8 _4381_ (.A(_0674_),
    .B(_0684_),
    .Y(_0952_));
 sky130_fd_sc_hd__or2_1 _4382_ (.A(_0951_),
    .B(_0952_),
    .X(_0953_));
 sky130_fd_sc_hd__clkbuf_8 _4383_ (.A(_0953_),
    .X(_0954_));
 sky130_fd_sc_hd__nor2b_2 _4384_ (.A(_0926_),
    .B_N(_0936_),
    .Y(_0955_));
 sky130_fd_sc_hd__nand2_1 _4385_ (.A(_0940_),
    .B(_0955_),
    .Y(_0956_));
 sky130_fd_sc_hd__or2_1 _4386_ (.A(_0909_),
    .B(_0956_),
    .X(_0957_));
 sky130_fd_sc_hd__buf_4 _4387_ (.A(_0957_),
    .X(_0958_));
 sky130_fd_sc_hd__buf_8 _4388_ (.A(_0951_),
    .X(_0959_));
 sky130_fd_sc_hd__or2_4 _4389_ (.A(_0959_),
    .B(_0944_),
    .X(_0960_));
 sky130_fd_sc_hd__o22a_1 _4390_ (.A1(_0950_),
    .A2(_0954_),
    .B1(_0958_),
    .B2(_0960_),
    .X(_0961_));
 sky130_fd_sc_hd__o221a_1 _4391_ (.A1(_0869_),
    .A2(_0939_),
    .B1(_0943_),
    .B2(_0948_),
    .C1(_0961_),
    .X(_0962_));
 sky130_fd_sc_hd__or2_1 _4392_ (.A(_0676_),
    .B(\oct.state[0] ),
    .X(_0963_));
 sky130_fd_sc_hd__buf_8 _4393_ (.A(_0963_),
    .X(_0964_));
 sky130_fd_sc_hd__nand2_1 _4394_ (.A(_0909_),
    .B(_0955_),
    .Y(_0965_));
 sky130_fd_sc_hd__or2_1 _4395_ (.A(_0918_),
    .B(_0965_),
    .X(_0966_));
 sky130_fd_sc_hd__clkbuf_4 _4396_ (.A(_0966_),
    .X(_0967_));
 sky130_fd_sc_hd__or2_1 _4397_ (.A(_0918_),
    .B(_0941_),
    .X(_0968_));
 sky130_fd_sc_hd__buf_4 _4398_ (.A(_0968_),
    .X(_0969_));
 sky130_fd_sc_hd__nand2_8 _4399_ (.A(_0686_),
    .B(\oct.state[0] ),
    .Y(_0970_));
 sky130_fd_sc_hd__nor2_8 _4400_ (.A(_0674_),
    .B(_0970_),
    .Y(_0971_));
 sky130_fd_sc_hd__nor2_1 _4401_ (.A(_0675_),
    .B(_0687_),
    .Y(_0972_));
 sky130_fd_sc_hd__or2_4 _4402_ (.A(_0971_),
    .B(_0972_),
    .X(_0973_));
 sky130_fd_sc_hd__or3b_4 _4403_ (.A(_0909_),
    .B(_0936_),
    .C_N(_0926_),
    .X(_0974_));
 sky130_fd_sc_hd__or2_1 _4404_ (.A(_0918_),
    .B(_0974_),
    .X(_0975_));
 sky130_fd_sc_hd__clkbuf_4 _4405_ (.A(_0975_),
    .X(_0976_));
 sky130_fd_sc_hd__nand2_8 _4406_ (.A(_0678_),
    .B(_0964_),
    .Y(_0977_));
 sky130_fd_sc_hd__nor2_4 _4407_ (.A(_0685_),
    .B(_0977_),
    .Y(_0978_));
 sky130_fd_sc_hd__or2_4 _4408_ (.A(_0978_),
    .B(_0971_),
    .X(_0979_));
 sky130_fd_sc_hd__or3b_1 _4409_ (.A(_0918_),
    .B(_0909_),
    .C_N(_0949_),
    .X(_0980_));
 sky130_fd_sc_hd__buf_4 _4410_ (.A(_0980_),
    .X(_0981_));
 sky130_fd_sc_hd__nand2_4 _4411_ (.A(_0676_),
    .B(_0680_),
    .Y(_0982_));
 sky130_fd_sc_hd__nor2_8 _4412_ (.A(_0674_),
    .B(_0982_),
    .Y(_0983_));
 sky130_fd_sc_hd__or2_1 _4413_ (.A(_0983_),
    .B(_0951_),
    .X(_0984_));
 sky130_fd_sc_hd__buf_4 _4414_ (.A(_0984_),
    .X(_0985_));
 sky130_fd_sc_hd__o22a_1 _4415_ (.A1(_0976_),
    .A2(_0979_),
    .B1(_0981_),
    .B2(_0985_),
    .X(_0986_));
 sky130_fd_sc_hd__o221a_1 _4416_ (.A1(_0964_),
    .A2(_0967_),
    .B1(_0969_),
    .B2(_0973_),
    .C1(_0986_),
    .X(_0987_));
 sky130_fd_sc_hd__or2_2 _4417_ (.A(_0909_),
    .B(_0940_),
    .X(_0988_));
 sky130_fd_sc_hd__or3_1 _4418_ (.A(_0926_),
    .B(_0936_),
    .C(_0988_),
    .X(_0989_));
 sky130_fd_sc_hd__clkbuf_8 _4419_ (.A(_0989_),
    .X(_0990_));
 sky130_fd_sc_hd__or2_1 _4420_ (.A(_0988_),
    .B(_0937_),
    .X(_0991_));
 sky130_fd_sc_hd__buf_4 _4421_ (.A(_0991_),
    .X(_0992_));
 sky130_fd_sc_hd__nor2_4 _4422_ (.A(_0674_),
    .B(_0680_),
    .Y(_0993_));
 sky130_fd_sc_hd__nand3_4 _4423_ (.A(_0949_),
    .B(_0909_),
    .C(_0918_),
    .Y(_0994_));
 sky130_fd_sc_hd__nor2_1 _4424_ (.A(_0686_),
    .B(_0674_),
    .Y(_0995_));
 sky130_fd_sc_hd__buf_8 _4425_ (.A(_0995_),
    .X(_0996_));
 sky130_fd_sc_hd__nor2_8 _4426_ (.A(net64),
    .B(_0996_),
    .Y(_0997_));
 sky130_fd_sc_hd__o32a_1 _4427_ (.A1(_0959_),
    .A2(_0992_),
    .A3(_0993_),
    .B1(_0994_),
    .B2(_0997_),
    .X(_0998_));
 sky130_fd_sc_hd__or2_1 _4428_ (.A(_0940_),
    .B(_0974_),
    .X(_0999_));
 sky130_fd_sc_hd__buf_4 _4429_ (.A(_0999_),
    .X(_1000_));
 sky130_fd_sc_hd__nor2_8 _4430_ (.A(_0685_),
    .B(_0680_),
    .Y(_1001_));
 sky130_fd_sc_hd__or2_1 _4431_ (.A(_0940_),
    .B(_0965_),
    .X(_1002_));
 sky130_fd_sc_hd__buf_4 _4432_ (.A(_1002_),
    .X(_1003_));
 sky130_fd_sc_hd__buf_8 _4433_ (.A(_0972_),
    .X(_1004_));
 sky130_fd_sc_hd__nor2_2 _4434_ (.A(_0944_),
    .B(_1004_),
    .Y(_1005_));
 sky130_fd_sc_hd__o22a_1 _4435_ (.A1(_1000_),
    .A2(_1001_),
    .B1(_1003_),
    .B2(_1005_),
    .X(_1006_));
 sky130_fd_sc_hd__o311a_1 _4436_ (.A1(_0990_),
    .A2(_0978_),
    .A3(_0944_),
    .B1(_0998_),
    .C1(_1006_),
    .X(_1007_));
 sky130_fd_sc_hd__nand3_1 _4437_ (.A(_0962_),
    .B(_0987_),
    .C(_1007_),
    .Y(_1008_));
 sky130_fd_sc_hd__xor2_1 _4438_ (.A(\sound1.count[1] ),
    .B(_1008_),
    .X(_1009_));
 sky130_fd_sc_hd__nand2_8 _4439_ (.A(_0685_),
    .B(_0681_),
    .Y(_1010_));
 sky130_fd_sc_hd__or2_4 _4440_ (.A(_0695_),
    .B(_0678_),
    .X(_1011_));
 sky130_fd_sc_hd__nor2_4 _4441_ (.A(_0675_),
    .B(_0970_),
    .Y(_1012_));
 sky130_fd_sc_hd__or2_1 _4442_ (.A(_0944_),
    .B(_1012_),
    .X(_1013_));
 sky130_fd_sc_hd__buf_4 _4443_ (.A(_1013_),
    .X(_1014_));
 sky130_fd_sc_hd__nand2_8 _4444_ (.A(_0695_),
    .B(_0964_),
    .Y(_1015_));
 sky130_fd_sc_hd__nand2_4 _4445_ (.A(_1015_),
    .B(_0869_),
    .Y(_1016_));
 sky130_fd_sc_hd__nor2_2 _4446_ (.A(_0683_),
    .B(_0947_),
    .Y(_1017_));
 sky130_fd_sc_hd__nor2_4 _4447_ (.A(_0674_),
    .B(_0964_),
    .Y(_1018_));
 sky130_fd_sc_hd__nor2_4 _4448_ (.A(_0675_),
    .B(_0945_),
    .Y(_1019_));
 sky130_fd_sc_hd__or2_4 _4449_ (.A(_1018_),
    .B(_1019_),
    .X(_1020_));
 sky130_fd_sc_hd__o22a_1 _4450_ (.A1(_0950_),
    .A2(_1017_),
    .B1(_1020_),
    .B2(_0994_),
    .X(_1021_));
 sky130_fd_sc_hd__o221a_1 _4451_ (.A1(_0979_),
    .A2(_0958_),
    .B1(_0992_),
    .B2(_1016_),
    .C1(_1021_),
    .X(_1022_));
 sky130_fd_sc_hd__o221a_1 _4452_ (.A1(_1011_),
    .A2(_0967_),
    .B1(_1003_),
    .B2(_1014_),
    .C1(_1022_),
    .X(_1023_));
 sky130_fd_sc_hd__nor2_2 _4453_ (.A(_0685_),
    .B(_0681_),
    .Y(_1024_));
 sky130_fd_sc_hd__buf_8 _4454_ (.A(_1024_),
    .X(_1025_));
 sky130_fd_sc_hd__nand2_4 _4455_ (.A(_0695_),
    .B(_0677_),
    .Y(_1026_));
 sky130_fd_sc_hd__nand2_2 _4456_ (.A(_0964_),
    .B(_1026_),
    .Y(_1027_));
 sky130_fd_sc_hd__nor2_8 _4457_ (.A(_0695_),
    .B(_0946_),
    .Y(_1028_));
 sky130_fd_sc_hd__o32a_1 _4458_ (.A1(_0969_),
    .A2(_1025_),
    .A3(_1028_),
    .B1(_1005_),
    .B2(_0943_),
    .X(_1029_));
 sky130_fd_sc_hd__o221a_1 _4459_ (.A1(_1000_),
    .A2(_1025_),
    .B1(_1027_),
    .B2(_0976_),
    .C1(_1029_),
    .X(_1030_));
 sky130_fd_sc_hd__o211a_1 _4460_ (.A1(_0981_),
    .A2(_0997_),
    .B1(_1023_),
    .C1(_1030_),
    .X(_1031_));
 sky130_fd_sc_hd__o221a_2 _4461_ (.A1(_0990_),
    .A2(_0973_),
    .B1(_0939_),
    .B2(_1010_),
    .C1(_1031_),
    .X(_1032_));
 sky130_fd_sc_hd__or2_2 _4462_ (.A(_0679_),
    .B(_0971_),
    .X(_1033_));
 sky130_fd_sc_hd__nor2_2 _4463_ (.A(_0685_),
    .B(_0677_),
    .Y(_1034_));
 sky130_fd_sc_hd__nor2_4 _4464_ (.A(_0952_),
    .B(_1034_),
    .Y(_1035_));
 sky130_fd_sc_hd__a211o_1 _4465_ (.A1(_0940_),
    .A2(_0944_),
    .B1(_1004_),
    .C1(_0974_),
    .X(_1036_));
 sky130_fd_sc_hd__o221a_1 _4466_ (.A1(_0992_),
    .A2(_1033_),
    .B1(_1035_),
    .B2(_0981_),
    .C1(_1036_),
    .X(_1037_));
 sky130_fd_sc_hd__nor2_8 _4467_ (.A(_0676_),
    .B(_0695_),
    .Y(_1038_));
 sky130_fd_sc_hd__or2_4 _4468_ (.A(_1019_),
    .B(_1038_),
    .X(_1039_));
 sky130_fd_sc_hd__nor2_4 _4469_ (.A(_0674_),
    .B(_0977_),
    .Y(_1040_));
 sky130_fd_sc_hd__nor2_8 _4470_ (.A(_1019_),
    .B(net63),
    .Y(_1041_));
 sky130_fd_sc_hd__nor2_2 _4471_ (.A(_0944_),
    .B(_0947_),
    .Y(_1042_));
 sky130_fd_sc_hd__nor2_2 _4472_ (.A(_0679_),
    .B(_0944_),
    .Y(_1043_));
 sky130_fd_sc_hd__o22a_1 _4473_ (.A1(_0958_),
    .A2(_1042_),
    .B1(_1043_),
    .B2(_0967_),
    .X(_1044_));
 sky130_fd_sc_hd__o221a_1 _4474_ (.A1(_1003_),
    .A2(_1039_),
    .B1(_1041_),
    .B2(_0939_),
    .C1(_1044_),
    .X(_1045_));
 sky130_fd_sc_hd__nor2_4 _4475_ (.A(_0674_),
    .B(_0945_),
    .Y(_1046_));
 sky130_fd_sc_hd__o22a_1 _4476_ (.A1(_0950_),
    .A2(_0996_),
    .B1(_1046_),
    .B2(_0994_),
    .X(_1047_));
 sky130_fd_sc_hd__o221a_1 _4477_ (.A1(_0990_),
    .A2(_0996_),
    .B1(_1040_),
    .B2(_0969_),
    .C1(_0943_),
    .X(_1048_));
 sky130_fd_sc_hd__o22a_1 _4478_ (.A1(_1001_),
    .A2(_1047_),
    .B1(_1048_),
    .B2(_0947_),
    .X(_1049_));
 sky130_fd_sc_hd__and3_2 _4479_ (.A(_1037_),
    .B(_1045_),
    .C(_1049_),
    .X(_1050_));
 sky130_fd_sc_hd__a2bb2o_1 _4480_ (.A1_N(\sound1.count[2] ),
    .A2_N(_1032_),
    .B1(_1050_),
    .B2(\sound1.count[11] ),
    .X(_1051_));
 sky130_fd_sc_hd__or2_1 _4481_ (.A(_0944_),
    .B(_0969_),
    .X(_1052_));
 sky130_fd_sc_hd__nor2_4 _4482_ (.A(net64),
    .B(_1001_),
    .Y(_1053_));
 sky130_fd_sc_hd__o32a_1 _4483_ (.A1(_0679_),
    .A2(_0950_),
    .A3(_1040_),
    .B1(_1053_),
    .B2(_0992_),
    .X(_1054_));
 sky130_fd_sc_hd__or2_4 _4484_ (.A(_0676_),
    .B(_0695_),
    .X(_1055_));
 sky130_fd_sc_hd__nand2_2 _4485_ (.A(_0678_),
    .B(_1055_),
    .Y(_1056_));
 sky130_fd_sc_hd__nand2_2 _4486_ (.A(_0695_),
    .B(_0970_),
    .Y(_1057_));
 sky130_fd_sc_hd__nand2_4 _4487_ (.A(_0685_),
    .B(_0977_),
    .Y(_1058_));
 sky130_fd_sc_hd__nor2_2 _4488_ (.A(_1018_),
    .B(_0959_),
    .Y(_1059_));
 sky130_fd_sc_hd__o22a_1 _4489_ (.A1(_0956_),
    .A2(_1026_),
    .B1(_1059_),
    .B2(_0981_),
    .X(_1060_));
 sky130_fd_sc_hd__o221a_1 _4490_ (.A1(_0939_),
    .A2(_1057_),
    .B1(_1058_),
    .B2(_0958_),
    .C1(_1060_),
    .X(_1061_));
 sky130_fd_sc_hd__nand2_4 _4491_ (.A(_0676_),
    .B(_0685_),
    .Y(_1062_));
 sky130_fd_sc_hd__nand2_2 _4492_ (.A(_0964_),
    .B(_1062_),
    .Y(_1063_));
 sky130_fd_sc_hd__a21oi_4 _4493_ (.A1(_0674_),
    .A2(_0684_),
    .B1(_0683_),
    .Y(_1064_));
 sky130_fd_sc_hd__o22a_1 _4494_ (.A1(_0979_),
    .A2(_1003_),
    .B1(_0943_),
    .B2(_0983_),
    .X(_1065_));
 sky130_fd_sc_hd__o221a_1 _4495_ (.A1(_1000_),
    .A2(_1063_),
    .B1(_1064_),
    .B2(_0994_),
    .C1(_1065_),
    .X(_1066_));
 sky130_fd_sc_hd__o211a_1 _4496_ (.A1(_0990_),
    .A2(_1056_),
    .B1(_1061_),
    .C1(_1066_),
    .X(_1067_));
 sky130_fd_sc_hd__o311a_1 _4497_ (.A1(_0677_),
    .A2(_0976_),
    .A3(_1038_),
    .B1(_1054_),
    .C1(_1067_),
    .X(_1068_));
 sky130_fd_sc_hd__nand3b_1 _4498_ (.A_N(_0949_),
    .B(_0937_),
    .C(_0974_),
    .Y(_1069_));
 sky130_fd_sc_hd__a21o_4 _4499_ (.A1(_0988_),
    .A2(_0955_),
    .B1(_1069_),
    .X(_1070_));
 sky130_fd_sc_hd__o211ai_4 _4500_ (.A1(_0676_),
    .A2(_1052_),
    .B1(_1068_),
    .C1(_1070_),
    .Y(_1071_));
 sky130_fd_sc_hd__inv_2 _4501_ (.A(_1071_),
    .Y(_1072_));
 sky130_fd_sc_hd__inv_2 _4502_ (.A(\sound1.count[7] ),
    .Y(_1073_));
 sky130_fd_sc_hd__o22a_1 _4503_ (.A1(_1015_),
    .A2(_0981_),
    .B1(_0969_),
    .B2(_0946_),
    .X(_1074_));
 sky130_fd_sc_hd__o221a_1 _4504_ (.A1(_0688_),
    .A2(_0958_),
    .B1(_0943_),
    .B2(_0971_),
    .C1(_1074_),
    .X(_1075_));
 sky130_fd_sc_hd__or2_1 _4505_ (.A(_0679_),
    .B(_1046_),
    .X(_1076_));
 sky130_fd_sc_hd__buf_4 _4506_ (.A(_1076_),
    .X(_1077_));
 sky130_fd_sc_hd__nand2_2 _4507_ (.A(_0695_),
    .B(_0680_),
    .Y(_1078_));
 sky130_fd_sc_hd__nand2_4 _4508_ (.A(_0970_),
    .B(_0869_),
    .Y(_1079_));
 sky130_fd_sc_hd__o22a_1 _4509_ (.A1(_0956_),
    .A2(_1078_),
    .B1(_1079_),
    .B2(_0992_),
    .X(_1080_));
 sky130_fd_sc_hd__o221a_1 _4510_ (.A1(_0990_),
    .A2(_0960_),
    .B1(_0994_),
    .B2(_1039_),
    .C1(_1080_),
    .X(_1081_));
 sky130_fd_sc_hd__or2_1 _4511_ (.A(_0680_),
    .B(_0976_),
    .X(_1082_));
 sky130_fd_sc_hd__nor2_4 _4512_ (.A(_0694_),
    .B(_0996_),
    .Y(_1083_));
 sky130_fd_sc_hd__or2_1 _4513_ (.A(_0950_),
    .B(_1083_),
    .X(_1084_));
 sky130_fd_sc_hd__nor2_2 _4514_ (.A(_0959_),
    .B(_0952_),
    .Y(_1085_));
 sky130_fd_sc_hd__o22a_1 _4515_ (.A1(_0952_),
    .A2(_1000_),
    .B1(_1003_),
    .B2(_1085_),
    .X(_1086_));
 sky130_fd_sc_hd__and3_1 _4516_ (.A(_1082_),
    .B(_1084_),
    .C(_1086_),
    .X(_1087_));
 sky130_fd_sc_hd__o311a_1 _4517_ (.A1(_0684_),
    .A2(_0939_),
    .A3(_1077_),
    .B1(_1081_),
    .C1(_1087_),
    .X(_1088_));
 sky130_fd_sc_hd__nand2_1 _4518_ (.A(_1075_),
    .B(_1088_),
    .Y(_1089_));
 sky130_fd_sc_hd__or2_1 _4519_ (.A(_0967_),
    .B(_1025_),
    .X(_1090_));
 sky130_fd_sc_hd__a21o_1 _4520_ (.A1(_0976_),
    .A2(_0994_),
    .B1(_0960_),
    .X(_1091_));
 sky130_fd_sc_hd__or3_1 _4521_ (.A(_0993_),
    .B(_0943_),
    .C(_1012_),
    .X(_1092_));
 sky130_fd_sc_hd__a21o_1 _4522_ (.A1(_0992_),
    .A2(_1003_),
    .B1(_0948_),
    .X(_1093_));
 sky130_fd_sc_hd__o2111a_1 _4523_ (.A1(_0996_),
    .A2(_1090_),
    .B1(_1091_),
    .C1(_1092_),
    .D1(_1093_),
    .X(_1094_));
 sky130_fd_sc_hd__nand2_4 _4524_ (.A(_0685_),
    .B(_0677_),
    .Y(_1095_));
 sky130_fd_sc_hd__or2_2 _4525_ (.A(_0983_),
    .B(_0978_),
    .X(_1096_));
 sky130_fd_sc_hd__nor2_2 _4526_ (.A(_0952_),
    .B(_0972_),
    .Y(_1097_));
 sky130_fd_sc_hd__o22a_1 _4527_ (.A1(_0969_),
    .A2(_1096_),
    .B1(_1097_),
    .B2(_1000_),
    .X(_1098_));
 sky130_fd_sc_hd__o221a_1 _4528_ (.A1(_0939_),
    .A2(_1095_),
    .B1(_1056_),
    .B2(_0958_),
    .C1(_1098_),
    .X(_1099_));
 sky130_fd_sc_hd__nor2_1 _4529_ (.A(_0674_),
    .B(_0687_),
    .Y(_1100_));
 sky130_fd_sc_hd__or2_4 _4530_ (.A(_1100_),
    .B(_0959_),
    .X(_1101_));
 sky130_fd_sc_hd__or3_1 _4531_ (.A(_0977_),
    .B(_0950_),
    .C(_0996_),
    .X(_1102_));
 sky130_fd_sc_hd__o221a_1 _4532_ (.A1(_0981_),
    .A2(_1041_),
    .B1(_1101_),
    .B2(_0990_),
    .C1(_1102_),
    .X(_1103_));
 sky130_fd_sc_hd__and3_2 _4533_ (.A(_1094_),
    .B(_1099_),
    .C(_1103_),
    .X(_1104_));
 sky130_fd_sc_hd__a22o_1 _4534_ (.A1(_1073_),
    .A2(_1089_),
    .B1(_1104_),
    .B2(\sound1.count[0] ),
    .X(_1105_));
 sky130_fd_sc_hd__a221o_1 _4535_ (.A1(\sound1.count[2] ),
    .A2(_1032_),
    .B1(_1072_),
    .B2(\sound1.count[6] ),
    .C1(_1105_),
    .X(_1106_));
 sky130_fd_sc_hd__nor2_8 _4536_ (.A(_0685_),
    .B(_0684_),
    .Y(_1107_));
 sky130_fd_sc_hd__o211a_1 _4537_ (.A1(_0683_),
    .A2(_0981_),
    .B1(_0992_),
    .C1(_1052_),
    .X(_1108_));
 sky130_fd_sc_hd__o22a_1 _4538_ (.A1(_0677_),
    .A2(_1084_),
    .B1(_1090_),
    .B2(_0952_),
    .X(_1109_));
 sky130_fd_sc_hd__nor2_2 _4539_ (.A(_0944_),
    .B(_1012_),
    .Y(_1110_));
 sky130_fd_sc_hd__nand2_4 _4540_ (.A(_0685_),
    .B(_0970_),
    .Y(_1111_));
 sky130_fd_sc_hd__nand2_4 _4541_ (.A(_1015_),
    .B(_1111_),
    .Y(_1112_));
 sky130_fd_sc_hd__nand2_2 _4542_ (.A(_1015_),
    .B(_1062_),
    .Y(_1113_));
 sky130_fd_sc_hd__o32a_1 _4543_ (.A1(_0687_),
    .A2(_1001_),
    .A3(_0943_),
    .B1(_0997_),
    .B2(_0939_),
    .X(_1114_));
 sky130_fd_sc_hd__o221a_1 _4544_ (.A1(_0976_),
    .A2(_1112_),
    .B1(_1113_),
    .B2(_1000_),
    .C1(_1114_),
    .X(_1115_));
 sky130_fd_sc_hd__a21oi_4 _4545_ (.A1(_0695_),
    .A2(net64),
    .B1(_1040_),
    .Y(_1116_));
 sky130_fd_sc_hd__o22a_1 _4546_ (.A1(_0990_),
    .A2(_1064_),
    .B1(_1116_),
    .B2(_0994_),
    .X(_1117_));
 sky130_fd_sc_hd__o2111a_1 _4547_ (.A1(_0958_),
    .A2(_1110_),
    .B1(_1115_),
    .C1(_1117_),
    .D1(_1070_),
    .X(_1118_));
 sky130_fd_sc_hd__o311a_1 _4548_ (.A1(_0676_),
    .A2(_1003_),
    .A3(_1034_),
    .B1(_1109_),
    .C1(_1118_),
    .X(_1119_));
 sky130_fd_sc_hd__o21ai_2 _4549_ (.A1(_1107_),
    .A2(_1108_),
    .B1(_1119_),
    .Y(_1120_));
 sky130_fd_sc_hd__nand2_1 _4550_ (.A(\sound1.count[13] ),
    .B(_1120_),
    .Y(_1121_));
 sky130_fd_sc_hd__or2_1 _4551_ (.A(\sound1.count[13] ),
    .B(_1120_),
    .X(_1122_));
 sky130_fd_sc_hd__nor2_2 _4552_ (.A(_0679_),
    .B(_0971_),
    .Y(_1123_));
 sky130_fd_sc_hd__or2_1 _4553_ (.A(_0683_),
    .B(_1034_),
    .X(_1124_));
 sky130_fd_sc_hd__buf_4 _4554_ (.A(_1124_),
    .X(_1125_));
 sky130_fd_sc_hd__nor2_4 _4555_ (.A(_0959_),
    .B(net63),
    .Y(_1126_));
 sky130_fd_sc_hd__nor2_4 _4556_ (.A(_1025_),
    .B(_1038_),
    .Y(_1127_));
 sky130_fd_sc_hd__or2_1 _4557_ (.A(_0995_),
    .B(_0947_),
    .X(_1128_));
 sky130_fd_sc_hd__clkbuf_8 _4558_ (.A(_1128_),
    .X(_1129_));
 sky130_fd_sc_hd__or2_1 _4559_ (.A(_0994_),
    .B(_1129_),
    .X(_1130_));
 sky130_fd_sc_hd__o221a_1 _4560_ (.A1(_0992_),
    .A2(_1126_),
    .B1(_1127_),
    .B2(_0990_),
    .C1(_1130_),
    .X(_1131_));
 sky130_fd_sc_hd__o221a_1 _4561_ (.A1(_0967_),
    .A2(_1123_),
    .B1(_1125_),
    .B2(_0958_),
    .C1(_1131_),
    .X(_1132_));
 sky130_fd_sc_hd__nor2_4 _4562_ (.A(_0674_),
    .B(_0681_),
    .Y(_1133_));
 sky130_fd_sc_hd__nor2_4 _4563_ (.A(_1107_),
    .B(_1133_),
    .Y(_1134_));
 sky130_fd_sc_hd__nor2_2 _4564_ (.A(_1107_),
    .B(net63),
    .Y(_1135_));
 sky130_fd_sc_hd__o22a_1 _4565_ (.A1(_0943_),
    .A2(_1134_),
    .B1(_1135_),
    .B2(_0950_),
    .X(_1136_));
 sky130_fd_sc_hd__o22a_1 _4566_ (.A1(_0696_),
    .A2(_0939_),
    .B1(_1003_),
    .B2(_1041_),
    .X(_1137_));
 sky130_fd_sc_hd__nand2_8 _4567_ (.A(_0685_),
    .B(_0678_),
    .Y(_1138_));
 sky130_fd_sc_hd__nor2_4 _4568_ (.A(_0959_),
    .B(_1028_),
    .Y(_1139_));
 sky130_fd_sc_hd__nor2_4 _4569_ (.A(_0945_),
    .B(_1038_),
    .Y(_1140_));
 sky130_fd_sc_hd__nor2_2 _4570_ (.A(_1038_),
    .B(_1034_),
    .Y(_1141_));
 sky130_fd_sc_hd__o22a_1 _4571_ (.A1(_1000_),
    .A2(_1140_),
    .B1(_1141_),
    .B2(_0976_),
    .X(_1142_));
 sky130_fd_sc_hd__o221a_1 _4572_ (.A1(_0981_),
    .A2(_1138_),
    .B1(_1139_),
    .B2(_0969_),
    .C1(_1142_),
    .X(_1143_));
 sky130_fd_sc_hd__and3_1 _4573_ (.A(_1136_),
    .B(_1137_),
    .C(_1143_),
    .X(_1144_));
 sky130_fd_sc_hd__and3_2 _4574_ (.A(_1070_),
    .B(_1132_),
    .C(_1144_),
    .X(_1145_));
 sky130_fd_sc_hd__or2_4 _4575_ (.A(_0683_),
    .B(_0694_),
    .X(_1146_));
 sky130_fd_sc_hd__or2_1 _4576_ (.A(_0994_),
    .B(_1053_),
    .X(_1147_));
 sky130_fd_sc_hd__o221a_1 _4577_ (.A1(_0983_),
    .A2(_0992_),
    .B1(_1146_),
    .B2(_0990_),
    .C1(_1147_),
    .X(_1148_));
 sky130_fd_sc_hd__o221a_1 _4578_ (.A1(_0943_),
    .A2(_1012_),
    .B1(_1127_),
    .B2(_0969_),
    .C1(_1148_),
    .X(_1149_));
 sky130_fd_sc_hd__o311a_1 _4579_ (.A1(_0680_),
    .A2(_0959_),
    .A3(_0958_),
    .B1(_1149_),
    .C1(_1070_),
    .X(_1150_));
 sky130_fd_sc_hd__nand2_2 _4580_ (.A(_0696_),
    .B(_1055_),
    .Y(_1151_));
 sky130_fd_sc_hd__or3_1 _4581_ (.A(_1107_),
    .B(_1003_),
    .C(_1040_),
    .X(_1152_));
 sky130_fd_sc_hd__o221a_1 _4582_ (.A1(_0939_),
    .A2(_1134_),
    .B1(_1151_),
    .B2(_0981_),
    .C1(_1152_),
    .X(_1153_));
 sky130_fd_sc_hd__or2_4 _4583_ (.A(_1018_),
    .B(_0978_),
    .X(_1154_));
 sky130_fd_sc_hd__o22a_1 _4584_ (.A1(_0950_),
    .A2(_1125_),
    .B1(_1154_),
    .B2(_1000_),
    .X(_1155_));
 sky130_fd_sc_hd__o221a_1 _4585_ (.A1(_0967_),
    .A2(_1095_),
    .B1(_1042_),
    .B2(_0976_),
    .C1(_1155_),
    .X(_1156_));
 sky130_fd_sc_hd__and3_2 _4586_ (.A(_1150_),
    .B(_1153_),
    .C(_1156_),
    .X(_1157_));
 sky130_fd_sc_hd__nor2_4 _4587_ (.A(_0685_),
    .B(_0982_),
    .Y(_1158_));
 sky130_fd_sc_hd__or2_2 _4588_ (.A(_1100_),
    .B(_1158_),
    .X(_1159_));
 sky130_fd_sc_hd__o22a_1 _4589_ (.A1(_0685_),
    .A2(_0981_),
    .B1(_0939_),
    .B2(_1159_),
    .X(_1160_));
 sky130_fd_sc_hd__o221a_1 _4590_ (.A1(_0680_),
    .A2(_0958_),
    .B1(_1154_),
    .B2(_0950_),
    .C1(_1160_),
    .X(_1161_));
 sky130_fd_sc_hd__o32a_1 _4591_ (.A1(_0969_),
    .A2(_1004_),
    .A3(_1038_),
    .B1(_1077_),
    .B2(_1000_),
    .X(_1162_));
 sky130_fd_sc_hd__o221a_1 _4592_ (.A1(_0677_),
    .A2(_0976_),
    .B1(_1046_),
    .B2(_1090_),
    .C1(_1162_),
    .X(_1163_));
 sky130_fd_sc_hd__or2_1 _4593_ (.A(_0683_),
    .B(_0947_),
    .X(_1164_));
 sky130_fd_sc_hd__nor2_2 _4594_ (.A(_0952_),
    .B(_1019_),
    .Y(_1165_));
 sky130_fd_sc_hd__nor2_2 _4595_ (.A(_1107_),
    .B(_0996_),
    .Y(_1166_));
 sky130_fd_sc_hd__or2_1 _4596_ (.A(_0994_),
    .B(_1126_),
    .X(_1167_));
 sky130_fd_sc_hd__o221a_1 _4597_ (.A1(_0990_),
    .A2(_0997_),
    .B1(_0992_),
    .B2(_1166_),
    .C1(_1167_),
    .X(_1168_));
 sky130_fd_sc_hd__o221a_1 _4598_ (.A1(_1003_),
    .A2(_1164_),
    .B1(_1165_),
    .B2(_0943_),
    .C1(_1168_),
    .X(_1169_));
 sky130_fd_sc_hd__and4_2 _4599_ (.A(_1070_),
    .B(_1161_),
    .C(_1163_),
    .D(_1169_),
    .X(_1170_));
 sky130_fd_sc_hd__a2bb2o_1 _4600_ (.A1_N(\sound1.count[10] ),
    .A2_N(_1157_),
    .B1(_1170_),
    .B2(\sound1.count[8] ),
    .X(_1171_));
 sky130_fd_sc_hd__a221o_1 _4601_ (.A1(_1121_),
    .A2(_1122_),
    .B1(_1145_),
    .B2(\sound1.count[4] ),
    .C1(_1171_),
    .X(_1172_));
 sky130_fd_sc_hd__or4_1 _4602_ (.A(_1009_),
    .B(_1051_),
    .C(_1106_),
    .D(_1172_),
    .X(_1173_));
 sky130_fd_sc_hd__a21o_2 _4603_ (.A1(_0695_),
    .A2(net64),
    .B1(net63),
    .X(_1174_));
 sky130_fd_sc_hd__nor2_2 _4604_ (.A(_1001_),
    .B(_1028_),
    .Y(_1175_));
 sky130_fd_sc_hd__or2_2 _4605_ (.A(_0996_),
    .B(_1019_),
    .X(_1176_));
 sky130_fd_sc_hd__o22a_1 _4606_ (.A1(_0950_),
    .A2(_0996_),
    .B1(_1176_),
    .B2(_0981_),
    .X(_1177_));
 sky130_fd_sc_hd__o221a_1 _4607_ (.A1(_0954_),
    .A2(_0994_),
    .B1(_0992_),
    .B2(_1129_),
    .C1(_1177_),
    .X(_1178_));
 sky130_fd_sc_hd__o221a_1 _4608_ (.A1(_0943_),
    .A2(_1028_),
    .B1(_1175_),
    .B2(_0976_),
    .C1(_1178_),
    .X(_1179_));
 sky130_fd_sc_hd__nor2_2 _4609_ (.A(_0983_),
    .B(_0978_),
    .Y(_1180_));
 sky130_fd_sc_hd__or2_1 _4610_ (.A(_0952_),
    .B(_1004_),
    .X(_1181_));
 sky130_fd_sc_hd__nor2_1 _4611_ (.A(_0959_),
    .B(_0944_),
    .Y(_1182_));
 sky130_fd_sc_hd__o22a_1 _4612_ (.A1(_1182_),
    .A2(_1000_),
    .B1(_1003_),
    .B2(_0985_),
    .X(_1183_));
 sky130_fd_sc_hd__o221a_1 _4613_ (.A1(_0969_),
    .A2(_1180_),
    .B1(_1181_),
    .B2(_0967_),
    .C1(_1183_),
    .X(_1184_));
 sky130_fd_sc_hd__o211a_1 _4614_ (.A1(_0958_),
    .A2(_1141_),
    .B1(_1179_),
    .C1(_1184_),
    .X(_1185_));
 sky130_fd_sc_hd__o221ai_4 _4615_ (.A1(_1026_),
    .A2(_0939_),
    .B1(_1174_),
    .B2(_0990_),
    .C1(_1185_),
    .Y(_1186_));
 sky130_fd_sc_hd__xor2_1 _4616_ (.A(\sound1.count[5] ),
    .B(_1186_),
    .X(_1187_));
 sky130_fd_sc_hd__o22a_1 _4617_ (.A1(_0676_),
    .A2(_1003_),
    .B1(_1083_),
    .B2(_1000_),
    .X(_1188_));
 sky130_fd_sc_hd__nor2_4 _4618_ (.A(_1001_),
    .B(net63),
    .Y(_1189_));
 sky130_fd_sc_hd__o22a_1 _4619_ (.A1(_0950_),
    .A2(_1004_),
    .B1(_1189_),
    .B2(_0969_),
    .X(_1190_));
 sky130_fd_sc_hd__o221a_1 _4620_ (.A1(_0677_),
    .A2(_0958_),
    .B1(_1077_),
    .B2(_0981_),
    .C1(_1190_),
    .X(_1191_));
 sky130_fd_sc_hd__o211a_1 _4621_ (.A1(_0939_),
    .A2(_1014_),
    .B1(_1188_),
    .C1(_1191_),
    .X(_1192_));
 sky130_fd_sc_hd__or2_2 _4622_ (.A(_1107_),
    .B(_1100_),
    .X(_1193_));
 sky130_fd_sc_hd__o221a_1 _4623_ (.A1(_0992_),
    .A2(_1028_),
    .B1(_1020_),
    .B2(_0990_),
    .C1(_1130_),
    .X(_1194_));
 sky130_fd_sc_hd__o221a_1 _4624_ (.A1(_1193_),
    .A2(_0967_),
    .B1(_0943_),
    .B2(_1158_),
    .C1(_1194_),
    .X(_1195_));
 sky130_fd_sc_hd__o211a_1 _4625_ (.A1(_0959_),
    .A2(_1082_),
    .B1(_1192_),
    .C1(_1195_),
    .X(_1196_));
 sky130_fd_sc_hd__xnor2_1 _4626_ (.A(\sound1.count[9] ),
    .B(_1196_),
    .Y(_1197_));
 sky130_fd_sc_hd__nand2_2 _4627_ (.A(_0685_),
    .B(_0964_),
    .Y(_1198_));
 sky130_fd_sc_hd__nand2_2 _4628_ (.A(_0970_),
    .B(_1078_),
    .Y(_1199_));
 sky130_fd_sc_hd__inv_2 _4629_ (.A(_1165_),
    .Y(_1200_));
 sky130_fd_sc_hd__o22a_1 _4630_ (.A1(_0686_),
    .A2(_0950_),
    .B1(_0994_),
    .B2(_1146_),
    .X(_1201_));
 sky130_fd_sc_hd__o221a_1 _4631_ (.A1(_0939_),
    .A2(_1200_),
    .B1(_1189_),
    .B2(_0990_),
    .C1(_1201_),
    .X(_1202_));
 sky130_fd_sc_hd__o221a_1 _4632_ (.A1(_1003_),
    .A2(_1134_),
    .B1(_1125_),
    .B2(_0976_),
    .C1(_1202_),
    .X(_1203_));
 sky130_fd_sc_hd__or2_2 _4633_ (.A(_0978_),
    .B(_0996_),
    .X(_1204_));
 sky130_fd_sc_hd__o32a_1 _4634_ (.A1(_0683_),
    .A2(_1107_),
    .A3(_1000_),
    .B1(_0943_),
    .B2(_1014_),
    .X(_1205_));
 sky130_fd_sc_hd__o221a_1 _4635_ (.A1(_0688_),
    .A2(_0967_),
    .B1(_0969_),
    .B2(_1204_),
    .C1(_1205_),
    .X(_1206_));
 sky130_fd_sc_hd__o211a_1 _4636_ (.A1(_0958_),
    .A2(_1027_),
    .B1(_1203_),
    .C1(_1206_),
    .X(_1207_));
 sky130_fd_sc_hd__o221a_2 _4637_ (.A1(_0981_),
    .A2(_1198_),
    .B1(_0992_),
    .B2(_1199_),
    .C1(_1207_),
    .X(_1208_));
 sky130_fd_sc_hd__xnor2_1 _4638_ (.A(\sound1.count[3] ),
    .B(_1208_),
    .Y(_1209_));
 sky130_fd_sc_hd__nand2_1 _4639_ (.A(_0949_),
    .B(_0988_),
    .Y(_1210_));
 sky130_fd_sc_hd__o32a_1 _4640_ (.A1(_0909_),
    .A2(_0937_),
    .A3(_1138_),
    .B1(_0974_),
    .B2(_0688_),
    .X(_1211_));
 sky130_fd_sc_hd__o221a_1 _4641_ (.A1(_1210_),
    .A2(_0869_),
    .B1(_0965_),
    .B2(_1011_),
    .C1(_1211_),
    .X(_1212_));
 sky130_fd_sc_hd__or2_4 _4642_ (.A(_0695_),
    .B(_0977_),
    .X(_1213_));
 sky130_fd_sc_hd__a21o_1 _4643_ (.A1(_0990_),
    .A2(_0941_),
    .B1(_1213_),
    .X(_1214_));
 sky130_fd_sc_hd__o2111a_1 _4644_ (.A1(_0958_),
    .A2(_1058_),
    .B1(_1212_),
    .C1(_1214_),
    .D1(_1070_),
    .X(_1215_));
 sky130_fd_sc_hd__nand2_1 _4645_ (.A(_0988_),
    .B(_0955_),
    .Y(_1216_));
 sky130_fd_sc_hd__a21o_1 _4646_ (.A1(_0990_),
    .A2(_0937_),
    .B1(_1055_),
    .X(_1217_));
 sky130_fd_sc_hd__a21o_1 _4647_ (.A1(_0974_),
    .A2(_1210_),
    .B1(_1010_),
    .X(_1218_));
 sky130_fd_sc_hd__o2111a_1 _4648_ (.A1(_0688_),
    .A2(_1216_),
    .B1(_1070_),
    .C1(_1217_),
    .D1(_1218_),
    .X(_1219_));
 sky130_fd_sc_hd__a22o_1 _4649_ (.A1(\sound1.count[15] ),
    .A2(_1215_),
    .B1(_1219_),
    .B2(\sound1.count[16] ),
    .X(_1220_));
 sky130_fd_sc_hd__o22ai_1 _4650_ (.A1(\sound1.count[15] ),
    .A2(_1215_),
    .B1(_1219_),
    .B2(\sound1.count[16] ),
    .Y(_1221_));
 sky130_fd_sc_hd__nand2_2 _4651_ (.A(_0685_),
    .B(_0684_),
    .Y(_1222_));
 sky130_fd_sc_hd__o21ai_2 _4652_ (.A1(_1222_),
    .A2(_1216_),
    .B1(_1070_),
    .Y(_1223_));
 sky130_fd_sc_hd__xnor2_1 _4653_ (.A(\sound1.count[18] ),
    .B(_1223_),
    .Y(_1224_));
 sky130_fd_sc_hd__a32o_1 _4654_ (.A1(_0988_),
    .A2(_0955_),
    .A3(_0971_),
    .B1(_1069_),
    .B2(_1018_),
    .X(_1225_));
 sky130_fd_sc_hd__xnor2_1 _4655_ (.A(\sound1.count[17] ),
    .B(_1225_),
    .Y(_1226_));
 sky130_fd_sc_hd__o211a_1 _4656_ (.A1(\sound1.count[11] ),
    .A2(_1050_),
    .B1(_1224_),
    .C1(_1226_),
    .X(_1227_));
 sky130_fd_sc_hd__or3b_1 _4657_ (.A(_1220_),
    .B(_1221_),
    .C_N(_1227_),
    .X(_1228_));
 sky130_fd_sc_hd__a21o_1 _4658_ (.A1(_0981_),
    .A2(_0994_),
    .B1(_0687_),
    .X(_1229_));
 sky130_fd_sc_hd__o221a_1 _4659_ (.A1(_0680_),
    .A2(_0950_),
    .B1(_0939_),
    .B2(_0684_),
    .C1(_0992_),
    .X(_1230_));
 sky130_fd_sc_hd__a21o_1 _4660_ (.A1(_1229_),
    .A2(_1230_),
    .B1(_0695_),
    .X(_1231_));
 sky130_fd_sc_hd__a211o_1 _4661_ (.A1(_0685_),
    .A2(_0940_),
    .B1(_0965_),
    .C1(_0964_),
    .X(_1232_));
 sky130_fd_sc_hd__o22a_1 _4662_ (.A1(_0974_),
    .A2(_1058_),
    .B1(_1111_),
    .B2(_0941_),
    .X(_1233_));
 sky130_fd_sc_hd__o211a_1 _4663_ (.A1(_0990_),
    .A2(_1062_),
    .B1(_1232_),
    .C1(_1233_),
    .X(_1234_));
 sky130_fd_sc_hd__o211a_1 _4664_ (.A1(_0958_),
    .A2(_1112_),
    .B1(_1231_),
    .C1(_1234_),
    .X(_1235_));
 sky130_fd_sc_hd__xnor2_1 _4665_ (.A(\sound1.count[14] ),
    .B(_1235_),
    .Y(_1236_));
 sky130_fd_sc_hd__inv_2 _4666_ (.A(\sound1.count[6] ),
    .Y(_1237_));
 sky130_fd_sc_hd__nor2_1 _4667_ (.A(_0681_),
    .B(_0944_),
    .Y(_1238_));
 sky130_fd_sc_hd__o32a_1 _4668_ (.A1(_1004_),
    .A2(_1003_),
    .A3(_1028_),
    .B1(_1238_),
    .B2(_1000_),
    .X(_1239_));
 sky130_fd_sc_hd__or2_2 _4669_ (.A(_0683_),
    .B(_0959_),
    .X(_1240_));
 sky130_fd_sc_hd__o22a_1 _4670_ (.A1(_0969_),
    .A2(_1101_),
    .B1(_1240_),
    .B2(_0943_),
    .X(_1241_));
 sky130_fd_sc_hd__nor2_1 _4671_ (.A(_1012_),
    .B(_1028_),
    .Y(_1242_));
 sky130_fd_sc_hd__o32a_1 _4672_ (.A1(_0958_),
    .A2(_0944_),
    .A3(_1004_),
    .B1(_1025_),
    .B2(_0981_),
    .X(_1243_));
 sky130_fd_sc_hd__o221a_1 _4673_ (.A1(_0985_),
    .A2(_0939_),
    .B1(_1242_),
    .B2(_0950_),
    .C1(_1243_),
    .X(_1244_));
 sky130_fd_sc_hd__or2_2 _4674_ (.A(_1018_),
    .B(_0959_),
    .X(_1245_));
 sky130_fd_sc_hd__o32a_1 _4675_ (.A1(_0994_),
    .A2(_1025_),
    .A3(_1038_),
    .B1(_0954_),
    .B2(_0990_),
    .X(_1246_));
 sky130_fd_sc_hd__o32a_1 _4676_ (.A1(_0967_),
    .A2(_1004_),
    .A3(_1133_),
    .B1(_1110_),
    .B2(_0976_),
    .X(_1247_));
 sky130_fd_sc_hd__o211a_1 _4677_ (.A1(_0992_),
    .A2(_1245_),
    .B1(_1246_),
    .C1(_1247_),
    .X(_1248_));
 sky130_fd_sc_hd__and4_2 _4678_ (.A(_1239_),
    .B(_1241_),
    .C(_1244_),
    .D(_1248_),
    .X(_1249_));
 sky130_fd_sc_hd__o22ai_1 _4679_ (.A1(\sound1.count[4] ),
    .A2(_1145_),
    .B1(_1249_),
    .B2(\sound1.count[12] ),
    .Y(_1250_));
 sky130_fd_sc_hd__a221o_1 _4680_ (.A1(_1237_),
    .A2(_1071_),
    .B1(_1157_),
    .B2(\sound1.count[10] ),
    .C1(_1250_),
    .X(_1251_));
 sky130_fd_sc_hd__o2bb2a_1 _4681_ (.A1_N(\sound1.count[12] ),
    .A2_N(_1249_),
    .B1(_1170_),
    .B2(\sound1.count[8] ),
    .X(_1252_));
 sky130_fd_sc_hd__o221a_1 _4682_ (.A1(_1073_),
    .A2(_1089_),
    .B1(_1104_),
    .B2(\sound1.count[0] ),
    .C1(_1252_),
    .X(_1253_));
 sky130_fd_sc_hd__or4b_1 _4683_ (.A(_1228_),
    .B(_1236_),
    .C(_1251_),
    .D_N(_1253_),
    .X(_1254_));
 sky130_fd_sc_hd__or4_1 _4684_ (.A(_1187_),
    .B(_1197_),
    .C(_1209_),
    .D(_1254_),
    .X(_1255_));
 sky130_fd_sc_hd__o21a_4 _4685_ (.A1(_1173_),
    .A2(_1255_),
    .B1(_1070_),
    .X(_1256_));
 sky130_fd_sc_hd__nand2_1 _4686_ (.A(\sound1.count[0] ),
    .B(_1256_),
    .Y(\sound1.osc.next_count[0] ));
 sky130_fd_sc_hd__or2_1 _4687_ (.A(\sound1.count[0] ),
    .B(\sound1.count[1] ),
    .X(_1257_));
 sky130_fd_sc_hd__nand2_1 _4688_ (.A(\sound1.count[0] ),
    .B(\sound1.count[1] ),
    .Y(_1258_));
 sky130_fd_sc_hd__and3_1 _4689_ (.A(_1256_),
    .B(_1257_),
    .C(_1258_),
    .X(_1259_));
 sky130_fd_sc_hd__clkbuf_1 _4690_ (.A(_1259_),
    .X(\sound1.osc.next_count[1] ));
 sky130_fd_sc_hd__a21o_1 _4691_ (.A1(\sound1.count[0] ),
    .A2(\sound1.count[1] ),
    .B1(\sound1.count[2] ),
    .X(_1260_));
 sky130_fd_sc_hd__nand3_1 _4692_ (.A(\sound1.count[0] ),
    .B(\sound1.count[1] ),
    .C(\sound1.count[2] ),
    .Y(_1261_));
 sky130_fd_sc_hd__and3_1 _4693_ (.A(_1256_),
    .B(_1260_),
    .C(_1261_),
    .X(_1262_));
 sky130_fd_sc_hd__clkbuf_1 _4694_ (.A(_1262_),
    .X(\sound1.osc.next_count[2] ));
 sky130_fd_sc_hd__and4_1 _4695_ (.A(\sound1.count[0] ),
    .B(\sound1.count[1] ),
    .C(\sound1.count[2] ),
    .D(\sound1.count[3] ),
    .X(_1263_));
 sky130_fd_sc_hd__a31o_1 _4696_ (.A1(\sound1.count[0] ),
    .A2(\sound1.count[1] ),
    .A3(\sound1.count[2] ),
    .B1(\sound1.count[3] ),
    .X(_1264_));
 sky130_fd_sc_hd__and3b_1 _4697_ (.A_N(_1263_),
    .B(_1264_),
    .C(_1256_),
    .X(_1265_));
 sky130_fd_sc_hd__clkbuf_1 _4698_ (.A(_1265_),
    .X(\sound1.osc.next_count[3] ));
 sky130_fd_sc_hd__nand2_1 _4699_ (.A(\sound1.count[4] ),
    .B(_1263_),
    .Y(_1266_));
 sky130_fd_sc_hd__or2_1 _4700_ (.A(\sound1.count[4] ),
    .B(_1263_),
    .X(_1267_));
 sky130_fd_sc_hd__and3_1 _4701_ (.A(_1256_),
    .B(_1266_),
    .C(_1267_),
    .X(_1268_));
 sky130_fd_sc_hd__clkbuf_1 _4702_ (.A(_1268_),
    .X(\sound1.osc.next_count[4] ));
 sky130_fd_sc_hd__and3_1 _4703_ (.A(\sound1.count[4] ),
    .B(\sound1.count[5] ),
    .C(_1263_),
    .X(_1269_));
 sky130_fd_sc_hd__a21o_1 _4704_ (.A1(\sound1.count[4] ),
    .A2(_1263_),
    .B1(\sound1.count[5] ),
    .X(_1270_));
 sky130_fd_sc_hd__and3b_1 _4705_ (.A_N(_1269_),
    .B(_1270_),
    .C(_1256_),
    .X(_1271_));
 sky130_fd_sc_hd__clkbuf_1 _4706_ (.A(_1271_),
    .X(\sound1.osc.next_count[5] ));
 sky130_fd_sc_hd__and2_1 _4707_ (.A(\sound1.count[6] ),
    .B(_1269_),
    .X(_1272_));
 sky130_fd_sc_hd__or2_1 _4708_ (.A(\sound1.count[6] ),
    .B(_1269_),
    .X(_1273_));
 sky130_fd_sc_hd__and3b_1 _4709_ (.A_N(_1272_),
    .B(_1273_),
    .C(_1256_),
    .X(_1274_));
 sky130_fd_sc_hd__clkbuf_1 _4710_ (.A(_1274_),
    .X(\sound1.osc.next_count[6] ));
 sky130_fd_sc_hd__nand2_1 _4711_ (.A(\sound1.count[7] ),
    .B(_1272_),
    .Y(_1275_));
 sky130_fd_sc_hd__or2_1 _4712_ (.A(\sound1.count[7] ),
    .B(_1272_),
    .X(_1276_));
 sky130_fd_sc_hd__and3_1 _4713_ (.A(_1256_),
    .B(_1275_),
    .C(_1276_),
    .X(_1277_));
 sky130_fd_sc_hd__clkbuf_1 _4714_ (.A(_1277_),
    .X(\sound1.osc.next_count[7] ));
 sky130_fd_sc_hd__and3_1 _4715_ (.A(\sound1.count[7] ),
    .B(\sound1.count[8] ),
    .C(_1272_),
    .X(_1278_));
 sky130_fd_sc_hd__a31o_1 _4716_ (.A1(\sound1.count[6] ),
    .A2(\sound1.count[7] ),
    .A3(_1269_),
    .B1(\sound1.count[8] ),
    .X(_1279_));
 sky130_fd_sc_hd__and3b_1 _4717_ (.A_N(_1278_),
    .B(_1279_),
    .C(_1256_),
    .X(_1280_));
 sky130_fd_sc_hd__clkbuf_1 _4718_ (.A(_1280_),
    .X(\sound1.osc.next_count[8] ));
 sky130_fd_sc_hd__and2_1 _4719_ (.A(\sound1.count[9] ),
    .B(_1278_),
    .X(_1281_));
 sky130_fd_sc_hd__or2_1 _4720_ (.A(\sound1.count[9] ),
    .B(_1278_),
    .X(_1282_));
 sky130_fd_sc_hd__and3b_1 _4721_ (.A_N(_1281_),
    .B(_1282_),
    .C(_1256_),
    .X(_1283_));
 sky130_fd_sc_hd__clkbuf_1 _4722_ (.A(_1283_),
    .X(\sound1.osc.next_count[9] ));
 sky130_fd_sc_hd__nand2_1 _4723_ (.A(\sound1.count[10] ),
    .B(_1281_),
    .Y(_1284_));
 sky130_fd_sc_hd__or2_1 _4724_ (.A(\sound1.count[10] ),
    .B(_1281_),
    .X(_1285_));
 sky130_fd_sc_hd__and3_1 _4725_ (.A(_1256_),
    .B(_1284_),
    .C(_1285_),
    .X(_1286_));
 sky130_fd_sc_hd__clkbuf_1 _4726_ (.A(_1286_),
    .X(\sound1.osc.next_count[10] ));
 sky130_fd_sc_hd__and3_1 _4727_ (.A(\sound1.count[10] ),
    .B(\sound1.count[11] ),
    .C(_1281_),
    .X(_1287_));
 sky130_fd_sc_hd__a31o_1 _4728_ (.A1(\sound1.count[9] ),
    .A2(\sound1.count[10] ),
    .A3(_1278_),
    .B1(\sound1.count[11] ),
    .X(_1288_));
 sky130_fd_sc_hd__and3b_1 _4729_ (.A_N(_1287_),
    .B(_1288_),
    .C(_1256_),
    .X(_1289_));
 sky130_fd_sc_hd__clkbuf_1 _4730_ (.A(_1289_),
    .X(\sound1.osc.next_count[11] ));
 sky130_fd_sc_hd__and2_1 _4731_ (.A(\sound1.count[12] ),
    .B(_1287_),
    .X(_1290_));
 sky130_fd_sc_hd__or2_1 _4732_ (.A(\sound1.count[12] ),
    .B(_1287_),
    .X(_1291_));
 sky130_fd_sc_hd__and3b_1 _4733_ (.A_N(_1290_),
    .B(_1291_),
    .C(_1256_),
    .X(_1292_));
 sky130_fd_sc_hd__clkbuf_1 _4734_ (.A(_1292_),
    .X(\sound1.osc.next_count[12] ));
 sky130_fd_sc_hd__nand2_1 _4735_ (.A(\sound1.count[13] ),
    .B(_1290_),
    .Y(_1293_));
 sky130_fd_sc_hd__or2_1 _4736_ (.A(\sound1.count[13] ),
    .B(_1290_),
    .X(_1294_));
 sky130_fd_sc_hd__and3_1 _4737_ (.A(_1256_),
    .B(_1293_),
    .C(_1294_),
    .X(_1295_));
 sky130_fd_sc_hd__clkbuf_1 _4738_ (.A(_1295_),
    .X(\sound1.osc.next_count[13] ));
 sky130_fd_sc_hd__and3_1 _4739_ (.A(\sound1.count[13] ),
    .B(\sound1.count[14] ),
    .C(_1290_),
    .X(_1296_));
 sky130_fd_sc_hd__a31o_1 _4740_ (.A1(\sound1.count[12] ),
    .A2(\sound1.count[13] ),
    .A3(_1287_),
    .B1(\sound1.count[14] ),
    .X(_1297_));
 sky130_fd_sc_hd__and3b_1 _4741_ (.A_N(_1296_),
    .B(_1297_),
    .C(_1256_),
    .X(_1298_));
 sky130_fd_sc_hd__clkbuf_1 _4742_ (.A(_1298_),
    .X(\sound1.osc.next_count[14] ));
 sky130_fd_sc_hd__and2_1 _4743_ (.A(\sound1.count[15] ),
    .B(_1296_),
    .X(_1299_));
 sky130_fd_sc_hd__or2_1 _4744_ (.A(\sound1.count[15] ),
    .B(_1296_),
    .X(_1300_));
 sky130_fd_sc_hd__and3b_1 _4745_ (.A_N(_1299_),
    .B(_1300_),
    .C(_1256_),
    .X(_1301_));
 sky130_fd_sc_hd__clkbuf_1 _4746_ (.A(_1301_),
    .X(\sound1.osc.next_count[15] ));
 sky130_fd_sc_hd__nand2_1 _4747_ (.A(\sound1.count[16] ),
    .B(_1299_),
    .Y(_1302_));
 sky130_fd_sc_hd__or2_1 _4748_ (.A(\sound1.count[16] ),
    .B(_1299_),
    .X(_1303_));
 sky130_fd_sc_hd__and3_1 _4749_ (.A(_1256_),
    .B(_1302_),
    .C(_1303_),
    .X(_1304_));
 sky130_fd_sc_hd__clkbuf_1 _4750_ (.A(_1304_),
    .X(\sound1.osc.next_count[16] ));
 sky130_fd_sc_hd__and3_1 _4751_ (.A(\sound1.count[16] ),
    .B(\sound1.count[17] ),
    .C(_1299_),
    .X(_1305_));
 sky130_fd_sc_hd__a31o_1 _4752_ (.A1(\sound1.count[15] ),
    .A2(\sound1.count[16] ),
    .A3(_1296_),
    .B1(\sound1.count[17] ),
    .X(_1306_));
 sky130_fd_sc_hd__and3b_1 _4753_ (.A_N(_1305_),
    .B(_1306_),
    .C(_1256_),
    .X(_1307_));
 sky130_fd_sc_hd__clkbuf_1 _4754_ (.A(_1307_),
    .X(\sound1.osc.next_count[17] ));
 sky130_fd_sc_hd__or2_1 _4755_ (.A(\sound1.count[18] ),
    .B(_1305_),
    .X(_1308_));
 sky130_fd_sc_hd__nand2_1 _4756_ (.A(\sound1.count[18] ),
    .B(_1305_),
    .Y(_1309_));
 sky130_fd_sc_hd__and3_1 _4757_ (.A(_1256_),
    .B(_1308_),
    .C(_1309_),
    .X(_1310_));
 sky130_fd_sc_hd__clkbuf_1 _4758_ (.A(_1310_),
    .X(\sound1.osc.next_count[18] ));
 sky130_fd_sc_hd__nor2_4 _4759_ (.A(_0575_),
    .B(_0560_),
    .Y(_1311_));
 sky130_fd_sc_hd__buf_4 _4760_ (.A(_1311_),
    .X(\sound2.sdiv.next_dived ));
 sky130_fd_sc_hd__and2_1 _4761_ (.A(_0699_),
    .B(net42),
    .X(_1312_));
 sky130_fd_sc_hd__nor2_1 _4762_ (.A(_0698_),
    .B(_0507_),
    .Y(_1313_));
 sky130_fd_sc_hd__or2_2 _4763_ (.A(_1312_),
    .B(_1313_),
    .X(_1314_));
 sky130_fd_sc_hd__or2_2 _4764_ (.A(_0698_),
    .B(_0504_),
    .X(_1315_));
 sky130_fd_sc_hd__nor2_4 _4765_ (.A(_1314_),
    .B(_1315_),
    .Y(_1316_));
 sky130_fd_sc_hd__or2_4 _4766_ (.A(_1314_),
    .B(_1316_),
    .X(_1317_));
 sky130_fd_sc_hd__inv_2 _4767_ (.A(\sound2.count[3] ),
    .Y(_1318_));
 sky130_fd_sc_hd__nand2_1 _4768_ (.A(_0507_),
    .B(_1312_),
    .Y(_1319_));
 sky130_fd_sc_hd__nor2_2 _4769_ (.A(_0499_),
    .B(_1319_),
    .Y(_1320_));
 sky130_fd_sc_hd__nand2_4 _4770_ (.A(net40),
    .B(_1320_),
    .Y(_1321_));
 sky130_fd_sc_hd__nand2_4 _4771_ (.A(_0499_),
    .B(_1316_),
    .Y(_1322_));
 sky130_fd_sc_hd__nand2_8 _4772_ (.A(_0504_),
    .B(_1320_),
    .Y(_1323_));
 sky130_fd_sc_hd__or3_2 _4773_ (.A(_0698_),
    .B(_0507_),
    .C(net42),
    .X(_1324_));
 sky130_fd_sc_hd__or2_2 _4774_ (.A(_0504_),
    .B(_1324_),
    .X(_1325_));
 sky130_fd_sc_hd__or2_1 _4775_ (.A(_0499_),
    .B(_1325_),
    .X(_1326_));
 sky130_fd_sc_hd__buf_4 _4776_ (.A(_1326_),
    .X(_1327_));
 sky130_fd_sc_hd__o22a_1 _4777_ (.A1(_1198_),
    .A2(_1323_),
    .B1(_1327_),
    .B2(_1204_),
    .X(_1328_));
 sky130_fd_sc_hd__o221a_1 _4778_ (.A1(_0686_),
    .A2(_1321_),
    .B1(_1322_),
    .B2(_1134_),
    .C1(_1328_),
    .X(_1329_));
 sky130_fd_sc_hd__or2_1 _4779_ (.A(_0698_),
    .B(_0499_),
    .X(_1330_));
 sky130_fd_sc_hd__nand2_1 _4780_ (.A(_1315_),
    .B(_1330_),
    .Y(_1331_));
 sky130_fd_sc_hd__or2_1 _4781_ (.A(_1319_),
    .B(_1331_),
    .X(_1332_));
 sky130_fd_sc_hd__clkbuf_8 _4782_ (.A(_1332_),
    .X(_1333_));
 sky130_fd_sc_hd__nand2_1 _4783_ (.A(net42),
    .B(_1313_),
    .Y(_1334_));
 sky130_fd_sc_hd__or2_1 _4784_ (.A(_1330_),
    .B(_1334_),
    .X(_1335_));
 sky130_fd_sc_hd__buf_4 _4785_ (.A(_1335_),
    .X(_1336_));
 sky130_fd_sc_hd__or2_1 _4786_ (.A(net39),
    .B(_1325_),
    .X(_1337_));
 sky130_fd_sc_hd__buf_4 _4787_ (.A(_1337_),
    .X(_1338_));
 sky130_fd_sc_hd__nand2_8 _4788_ (.A(net39),
    .B(_1316_),
    .Y(_1339_));
 sky130_fd_sc_hd__or2_1 _4789_ (.A(_1331_),
    .B(_1324_),
    .X(_1340_));
 sky130_fd_sc_hd__buf_4 _4790_ (.A(_1340_),
    .X(_1341_));
 sky130_fd_sc_hd__or3_1 _4791_ (.A(net40),
    .B(_1330_),
    .C(_1324_),
    .X(_1342_));
 sky130_fd_sc_hd__buf_4 _4792_ (.A(_1342_),
    .X(_1343_));
 sky130_fd_sc_hd__or2_1 _4793_ (.A(_1331_),
    .B(_1334_),
    .X(_1344_));
 sky130_fd_sc_hd__buf_4 _4794_ (.A(_1344_),
    .X(_1345_));
 sky130_fd_sc_hd__or3_1 _4795_ (.A(net39),
    .B(_1315_),
    .C(_1319_),
    .X(_1346_));
 sky130_fd_sc_hd__buf_4 _4796_ (.A(_1346_),
    .X(_1347_));
 sky130_fd_sc_hd__o32a_1 _4797_ (.A1(_0683_),
    .A2(_1107_),
    .A3(_1345_),
    .B1(_1347_),
    .B2(_1146_),
    .X(_1348_));
 sky130_fd_sc_hd__o221a_1 _4798_ (.A1(_1199_),
    .A2(_1341_),
    .B1(_1343_),
    .B2(_1200_),
    .C1(_1348_),
    .X(_1349_));
 sky130_fd_sc_hd__o221a_1 _4799_ (.A1(_1014_),
    .A2(_1338_),
    .B1(_1339_),
    .B2(_0688_),
    .C1(_1349_),
    .X(_1350_));
 sky130_fd_sc_hd__o221a_1 _4800_ (.A1(_1189_),
    .A2(_1333_),
    .B1(_1336_),
    .B2(_1125_),
    .C1(_1350_),
    .X(_1351_));
 sky130_fd_sc_hd__nand2_1 _4801_ (.A(_1329_),
    .B(_1351_),
    .Y(_1352_));
 sky130_fd_sc_hd__o32a_1 _4802_ (.A1(_1025_),
    .A2(_1038_),
    .A3(_1347_),
    .B1(_1333_),
    .B2(_0954_),
    .X(_1353_));
 sky130_fd_sc_hd__o221a_1 _4803_ (.A1(_1245_),
    .A2(_1341_),
    .B1(_1343_),
    .B2(_0985_),
    .C1(_1353_),
    .X(_1354_));
 sky130_fd_sc_hd__or3_1 _4804_ (.A(_1004_),
    .B(_1028_),
    .C(_1322_),
    .X(_1355_));
 sky130_fd_sc_hd__o221a_1 _4805_ (.A1(_1025_),
    .A2(_1323_),
    .B1(_1338_),
    .B2(_1240_),
    .C1(_1355_),
    .X(_1356_));
 sky130_fd_sc_hd__or3_1 _4806_ (.A(_1004_),
    .B(_1133_),
    .C(_1339_),
    .X(_1357_));
 sky130_fd_sc_hd__o221a_1 _4807_ (.A1(_1110_),
    .A2(_1336_),
    .B1(_1345_),
    .B2(_1238_),
    .C1(_1357_),
    .X(_1358_));
 sky130_fd_sc_hd__o221a_1 _4808_ (.A1(_1242_),
    .A2(_1321_),
    .B1(_1327_),
    .B2(_1101_),
    .C1(_1358_),
    .X(_1359_));
 sky130_fd_sc_hd__and3_2 _4809_ (.A(_1354_),
    .B(_1356_),
    .C(_1359_),
    .X(_1360_));
 sky130_fd_sc_hd__o32a_1 _4810_ (.A1(_0684_),
    .A2(_1077_),
    .A3(_1343_),
    .B1(_1338_),
    .B2(_0971_),
    .X(_1361_));
 sky130_fd_sc_hd__o221a_1 _4811_ (.A1(_1015_),
    .A2(_1323_),
    .B1(_1327_),
    .B2(_0946_),
    .C1(_1361_),
    .X(_1362_));
 sky130_fd_sc_hd__or2_1 _4812_ (.A(_1039_),
    .B(_1347_),
    .X(_1363_));
 sky130_fd_sc_hd__o221a_1 _4813_ (.A1(_0960_),
    .A2(_1333_),
    .B1(_1345_),
    .B2(_0952_),
    .C1(_1363_),
    .X(_1364_));
 sky130_fd_sc_hd__or2_1 _4814_ (.A(_0680_),
    .B(_1336_),
    .X(_1365_));
 sky130_fd_sc_hd__o221a_1 _4815_ (.A1(_1083_),
    .A2(_1321_),
    .B1(_1341_),
    .B2(_1079_),
    .C1(_1365_),
    .X(_1366_));
 sky130_fd_sc_hd__o221a_1 _4816_ (.A1(_1085_),
    .A2(_1322_),
    .B1(_1339_),
    .B2(_1078_),
    .C1(_1366_),
    .X(_1367_));
 sky130_fd_sc_hd__and3_1 _4817_ (.A(_1362_),
    .B(_1364_),
    .C(_1367_),
    .X(_1368_));
 sky130_fd_sc_hd__a2bb2o_1 _4818_ (.A1_N(\sound2.count[12] ),
    .A2_N(_1360_),
    .B1(_1368_),
    .B2(\sound2.count[7] ),
    .X(_1369_));
 sky130_fd_sc_hd__a221o_1 _4819_ (.A1(_1318_),
    .A2(_1352_),
    .B1(_1360_),
    .B2(\sound2.count[12] ),
    .C1(_1369_),
    .X(_1370_));
 sky130_fd_sc_hd__o32a_1 _4820_ (.A1(_0679_),
    .A2(_1040_),
    .A3(_1321_),
    .B1(_1323_),
    .B2(_1059_),
    .X(_1371_));
 sky130_fd_sc_hd__or2_1 _4821_ (.A(_0944_),
    .B(_1327_),
    .X(_1372_));
 sky130_fd_sc_hd__o221a_1 _4822_ (.A1(_1064_),
    .A2(_1347_),
    .B1(_1322_),
    .B2(_0979_),
    .C1(_1317_),
    .X(_1373_));
 sky130_fd_sc_hd__o22a_1 _4823_ (.A1(_1057_),
    .A2(_1343_),
    .B1(_1333_),
    .B2(_1056_),
    .X(_1374_));
 sky130_fd_sc_hd__o221a_1 _4824_ (.A1(_1053_),
    .A2(_1341_),
    .B1(_1345_),
    .B2(_1063_),
    .C1(_1374_),
    .X(_1375_));
 sky130_fd_sc_hd__o32a_1 _4825_ (.A1(_0677_),
    .A2(_1038_),
    .A3(_1336_),
    .B1(_1339_),
    .B2(_1026_),
    .X(_1376_));
 sky130_fd_sc_hd__o2111a_1 _4826_ (.A1(_0676_),
    .A2(_1372_),
    .B1(_1373_),
    .C1(_1375_),
    .D1(_1376_),
    .X(_1377_));
 sky130_fd_sc_hd__o211ai_4 _4827_ (.A1(_0983_),
    .A2(_1338_),
    .B1(_1371_),
    .C1(_1377_),
    .Y(_1378_));
 sky130_fd_sc_hd__xor2_1 _4828_ (.A(\sound2.count[6] ),
    .B(_1378_),
    .X(_1379_));
 sky130_fd_sc_hd__o22a_1 _4829_ (.A1(_1125_),
    .A2(_1321_),
    .B1(_1327_),
    .B2(_1127_),
    .X(_1380_));
 sky130_fd_sc_hd__o22a_1 _4830_ (.A1(_1042_),
    .A2(_1336_),
    .B1(_1345_),
    .B2(_1154_),
    .X(_1381_));
 sky130_fd_sc_hd__o221a_1 _4831_ (.A1(_1053_),
    .A2(_1347_),
    .B1(_1341_),
    .B2(_0983_),
    .C1(_1381_),
    .X(_1382_));
 sky130_fd_sc_hd__or2_1 _4832_ (.A(_1012_),
    .B(_1338_),
    .X(_1383_));
 sky130_fd_sc_hd__o221a_1 _4833_ (.A1(_1134_),
    .A2(_1343_),
    .B1(_1333_),
    .B2(_1146_),
    .C1(_1383_),
    .X(_1384_));
 sky130_fd_sc_hd__o221a_1 _4834_ (.A1(_1151_),
    .A2(_1323_),
    .B1(_1339_),
    .B2(_1095_),
    .C1(_1384_),
    .X(_1385_));
 sky130_fd_sc_hd__and3_1 _4835_ (.A(_1317_),
    .B(_1382_),
    .C(_1385_),
    .X(_1386_));
 sky130_fd_sc_hd__o311a_2 _4836_ (.A1(_1107_),
    .A2(net63),
    .A3(_1322_),
    .B1(_1380_),
    .C1(_1386_),
    .X(_1387_));
 sky130_fd_sc_hd__xnor2_1 _4837_ (.A(\sound2.count[10] ),
    .B(_1387_),
    .Y(_1388_));
 sky130_fd_sc_hd__o22a_1 _4838_ (.A1(_1129_),
    .A2(_1341_),
    .B1(_1336_),
    .B2(_1175_),
    .X(_1389_));
 sky130_fd_sc_hd__o221a_1 _4839_ (.A1(_0954_),
    .A2(_1347_),
    .B1(_1345_),
    .B2(_1182_),
    .C1(_1389_),
    .X(_1390_));
 sky130_fd_sc_hd__or2_1 _4840_ (.A(_1180_),
    .B(_1327_),
    .X(_1391_));
 sky130_fd_sc_hd__o221a_1 _4841_ (.A1(_1176_),
    .A2(_1323_),
    .B1(_1338_),
    .B2(_1028_),
    .C1(_1391_),
    .X(_1392_));
 sky130_fd_sc_hd__or2_1 _4842_ (.A(_0996_),
    .B(_1321_),
    .X(_1393_));
 sky130_fd_sc_hd__o221a_1 _4843_ (.A1(_1026_),
    .A2(_1343_),
    .B1(_1333_),
    .B2(_1174_),
    .C1(_1393_),
    .X(_1394_));
 sky130_fd_sc_hd__o221a_1 _4844_ (.A1(_0985_),
    .A2(_1322_),
    .B1(_1339_),
    .B2(_1181_),
    .C1(_1394_),
    .X(_1395_));
 sky130_fd_sc_hd__and3_2 _4845_ (.A(_1390_),
    .B(_1392_),
    .C(_1395_),
    .X(_1396_));
 sky130_fd_sc_hd__a2bb2o_1 _4846_ (.A1_N(\sound2.count[7] ),
    .A2_N(_1368_),
    .B1(_1396_),
    .B2(\sound2.count[5] ),
    .X(_1397_));
 sky130_fd_sc_hd__o32a_1 _4847_ (.A1(_0959_),
    .A2(_0993_),
    .A3(_1341_),
    .B1(_1336_),
    .B2(_0979_),
    .X(_1398_));
 sky130_fd_sc_hd__o22a_1 _4848_ (.A1(_0954_),
    .A2(_1321_),
    .B1(_1327_),
    .B2(_0973_),
    .X(_1399_));
 sky130_fd_sc_hd__o221a_1 _4849_ (.A1(_0985_),
    .A2(_1323_),
    .B1(_1338_),
    .B2(_0948_),
    .C1(_1399_),
    .X(_1400_));
 sky130_fd_sc_hd__o32a_1 _4850_ (.A1(_0978_),
    .A2(_0944_),
    .A3(_1333_),
    .B1(_1347_),
    .B2(_0997_),
    .X(_1401_));
 sky130_fd_sc_hd__o221a_1 _4851_ (.A1(_0869_),
    .A2(_1343_),
    .B1(_1345_),
    .B2(_1001_),
    .C1(_1401_),
    .X(_1402_));
 sky130_fd_sc_hd__o221a_1 _4852_ (.A1(_1005_),
    .A2(_1322_),
    .B1(_1339_),
    .B2(_0964_),
    .C1(_1402_),
    .X(_1403_));
 sky130_fd_sc_hd__and3_1 _4853_ (.A(_1398_),
    .B(_1400_),
    .C(_1403_),
    .X(_1404_));
 sky130_fd_sc_hd__o22a_1 _4854_ (.A1(_0677_),
    .A2(_1336_),
    .B1(_1345_),
    .B2(_1077_),
    .X(_1405_));
 sky130_fd_sc_hd__o22a_1 _4855_ (.A1(_1159_),
    .A2(_1343_),
    .B1(_1333_),
    .B2(_0997_),
    .X(_1406_));
 sky130_fd_sc_hd__o221a_1 _4856_ (.A1(_1126_),
    .A2(_1347_),
    .B1(_1341_),
    .B2(_1166_),
    .C1(_1406_),
    .X(_1407_));
 sky130_fd_sc_hd__o221a_1 _4857_ (.A1(_0685_),
    .A2(_1323_),
    .B1(_1338_),
    .B2(_1165_),
    .C1(_1407_),
    .X(_1408_));
 sky130_fd_sc_hd__o32a_1 _4858_ (.A1(_1025_),
    .A2(_1046_),
    .A3(_1339_),
    .B1(_1322_),
    .B2(_1164_),
    .X(_1409_));
 sky130_fd_sc_hd__o32a_1 _4859_ (.A1(_1004_),
    .A2(_1038_),
    .A3(_1327_),
    .B1(_1321_),
    .B2(_1154_),
    .X(_1410_));
 sky130_fd_sc_hd__and3_1 _4860_ (.A(_1317_),
    .B(_1409_),
    .C(_1410_),
    .X(_1411_));
 sky130_fd_sc_hd__and3_1 _4861_ (.A(_1405_),
    .B(_1408_),
    .C(_1411_),
    .X(_1412_));
 sky130_fd_sc_hd__a2bb2o_1 _4862_ (.A1_N(\sound2.count[1] ),
    .A2_N(_1404_),
    .B1(_1412_),
    .B2(\sound2.count[8] ),
    .X(_1413_));
 sky130_fd_sc_hd__or4_1 _4863_ (.A(_1379_),
    .B(_1388_),
    .C(_1397_),
    .D(_1413_),
    .X(_1414_));
 sky130_fd_sc_hd__o221a_1 _4864_ (.A1(_0684_),
    .A2(_1343_),
    .B1(_1333_),
    .B2(_0686_),
    .C1(_1341_),
    .X(_1415_));
 sky130_fd_sc_hd__a21o_1 _4865_ (.A1(_1347_),
    .A2(_1323_),
    .B1(_0687_),
    .X(_1416_));
 sky130_fd_sc_hd__o211a_1 _4866_ (.A1(_0680_),
    .A2(_1321_),
    .B1(_1415_),
    .C1(_1416_),
    .X(_1417_));
 sky130_fd_sc_hd__or2_1 _4867_ (.A(_1314_),
    .B(_1315_),
    .X(_1418_));
 sky130_fd_sc_hd__or2_1 _4868_ (.A(_0695_),
    .B(_0499_),
    .X(_1419_));
 sky130_fd_sc_hd__or3b_1 _4869_ (.A(_0964_),
    .B(_1418_),
    .C_N(_1419_),
    .X(_1420_));
 sky130_fd_sc_hd__o221a_1 _4870_ (.A1(_1111_),
    .A2(_1325_),
    .B1(_1334_),
    .B2(_1058_),
    .C1(_1420_),
    .X(_1421_));
 sky130_fd_sc_hd__o21ai_2 _4871_ (.A1(_0695_),
    .A2(_1417_),
    .B1(_1421_),
    .Y(_1422_));
 sky130_fd_sc_hd__nand2_1 _4872_ (.A(\sound2.count[14] ),
    .B(_1422_),
    .Y(_1423_));
 sky130_fd_sc_hd__or2_1 _4873_ (.A(\sound2.count[14] ),
    .B(_1422_),
    .X(_1424_));
 sky130_fd_sc_hd__or2_1 _4874_ (.A(_0683_),
    .B(_1323_),
    .X(_1425_));
 sky130_fd_sc_hd__a31o_1 _4875_ (.A1(_1341_),
    .A2(_1372_),
    .A3(_1425_),
    .B1(_1107_),
    .X(_1426_));
 sky130_fd_sc_hd__or2_1 _4876_ (.A(_0676_),
    .B(_1322_),
    .X(_1427_));
 sky130_fd_sc_hd__or3_1 _4877_ (.A(_0677_),
    .B(_1083_),
    .C(_1321_),
    .X(_1428_));
 sky130_fd_sc_hd__o22a_1 _4878_ (.A1(_1116_),
    .A2(_1347_),
    .B1(_1345_),
    .B2(_1113_),
    .X(_1429_));
 sky130_fd_sc_hd__o221a_1 _4879_ (.A1(_0997_),
    .A2(_1343_),
    .B1(_1333_),
    .B2(_1064_),
    .C1(_1429_),
    .X(_1430_));
 sky130_fd_sc_hd__o211a_1 _4880_ (.A1(_1034_),
    .A2(_1427_),
    .B1(_1428_),
    .C1(_1430_),
    .X(_1431_));
 sky130_fd_sc_hd__o32a_1 _4881_ (.A1(_0687_),
    .A2(_1001_),
    .A3(_1338_),
    .B1(_1336_),
    .B2(_1112_),
    .X(_1432_));
 sky130_fd_sc_hd__o31a_1 _4882_ (.A1(_0952_),
    .A2(_1025_),
    .A3(_1339_),
    .B1(_1432_),
    .X(_1433_));
 sky130_fd_sc_hd__and4_2 _4883_ (.A(_1317_),
    .B(_1426_),
    .C(_1431_),
    .D(_1433_),
    .X(_1434_));
 sky130_fd_sc_hd__o22a_1 _4884_ (.A1(_1134_),
    .A2(_1338_),
    .B1(_1322_),
    .B2(_1041_),
    .X(_1435_));
 sky130_fd_sc_hd__o22a_1 _4885_ (.A1(_1135_),
    .A2(_1321_),
    .B1(_1333_),
    .B2(_1127_),
    .X(_1436_));
 sky130_fd_sc_hd__o22a_1 _4886_ (.A1(_1129_),
    .A2(_1347_),
    .B1(_1345_),
    .B2(_1140_),
    .X(_1437_));
 sky130_fd_sc_hd__o221a_1 _4887_ (.A1(_1138_),
    .A2(_1323_),
    .B1(_1341_),
    .B2(_1126_),
    .C1(_1437_),
    .X(_1438_));
 sky130_fd_sc_hd__o221a_1 _4888_ (.A1(_1123_),
    .A2(_1339_),
    .B1(_1336_),
    .B2(_1141_),
    .C1(_1438_),
    .X(_1439_));
 sky130_fd_sc_hd__o211a_1 _4889_ (.A1(_0696_),
    .A2(_1343_),
    .B1(_1436_),
    .C1(_1439_),
    .X(_1440_));
 sky130_fd_sc_hd__o2111ai_4 _4890_ (.A1(_1139_),
    .A2(_1327_),
    .B1(_1435_),
    .C1(_1440_),
    .D1(_1317_),
    .Y(_1441_));
 sky130_fd_sc_hd__xor2_1 _4891_ (.A(\sound2.count[4] ),
    .B(_1441_),
    .X(_1442_));
 sky130_fd_sc_hd__a221o_1 _4892_ (.A1(_1423_),
    .A2(_1424_),
    .B1(_1434_),
    .B2(\sound2.count[13] ),
    .C1(_1442_),
    .X(_1443_));
 sky130_fd_sc_hd__nor2_1 _4893_ (.A(\sound2.count[13] ),
    .B(_1434_),
    .Y(_1444_));
 sky130_fd_sc_hd__o31a_1 _4894_ (.A1(_0695_),
    .A2(_0964_),
    .A3(_1418_),
    .B1(_1317_),
    .X(_1445_));
 sky130_fd_sc_hd__a22o_1 _4895_ (.A1(_1018_),
    .A2(_1314_),
    .B1(_1316_),
    .B2(_0971_),
    .X(_1446_));
 sky130_fd_sc_hd__xnor2_1 _4896_ (.A(\sound2.count[17] ),
    .B(_1446_),
    .Y(_1447_));
 sky130_fd_sc_hd__o21ai_1 _4897_ (.A1(\sound2.count[18] ),
    .A2(_1445_),
    .B1(_1447_),
    .Y(_1448_));
 sky130_fd_sc_hd__nand2_1 _4898_ (.A(_1333_),
    .B(_1325_),
    .Y(_1449_));
 sky130_fd_sc_hd__a21oi_1 _4899_ (.A1(_0499_),
    .A2(_1315_),
    .B1(_1319_),
    .Y(_1450_));
 sky130_fd_sc_hd__a22o_1 _4900_ (.A1(net63),
    .A2(_1449_),
    .B1(_1450_),
    .B2(_0944_),
    .X(_1451_));
 sky130_fd_sc_hd__or3b_1 _4901_ (.A(_1138_),
    .B(_1324_),
    .C_N(_1315_),
    .X(_1452_));
 sky130_fd_sc_hd__o211ai_1 _4902_ (.A1(_0688_),
    .A2(_1334_),
    .B1(_1452_),
    .C1(_1317_),
    .Y(_1453_));
 sky130_fd_sc_hd__a211o_2 _4903_ (.A1(_0683_),
    .A2(_1316_),
    .B1(_1451_),
    .C1(_1453_),
    .X(_1454_));
 sky130_fd_sc_hd__xor2_1 _4904_ (.A(\sound2.count[15] ),
    .B(_1454_),
    .X(_1455_));
 sky130_fd_sc_hd__and2b_1 _4905_ (.A_N(_1450_),
    .B(_1334_),
    .X(_1456_));
 sky130_fd_sc_hd__a21o_1 _4906_ (.A1(_1324_),
    .A2(_1333_),
    .B1(_1055_),
    .X(_1457_));
 sky130_fd_sc_hd__o211a_1 _4907_ (.A1(_0688_),
    .A2(_1418_),
    .B1(_1317_),
    .C1(_1457_),
    .X(_1458_));
 sky130_fd_sc_hd__o21ai_4 _4908_ (.A1(_1010_),
    .A2(_1456_),
    .B1(_1458_),
    .Y(_1459_));
 sky130_fd_sc_hd__xor2_1 _4909_ (.A(\sound2.count[16] ),
    .B(_1459_),
    .X(_1460_));
 sky130_fd_sc_hd__a2111o_1 _4910_ (.A1(\sound2.count[18] ),
    .A2(_1445_),
    .B1(_1448_),
    .C1(_1455_),
    .D1(_1460_),
    .X(_1461_));
 sky130_fd_sc_hd__o22a_1 _4911_ (.A1(_1017_),
    .A2(_1321_),
    .B1(_1341_),
    .B2(_1016_),
    .X(_1462_));
 sky130_fd_sc_hd__o22a_1 _4912_ (.A1(_1020_),
    .A2(_1347_),
    .B1(_1333_),
    .B2(_0973_),
    .X(_1463_));
 sky130_fd_sc_hd__o221a_1 _4913_ (.A1(_0997_),
    .A2(_1323_),
    .B1(_1343_),
    .B2(_1010_),
    .C1(_1463_),
    .X(_1464_));
 sky130_fd_sc_hd__o221a_1 _4914_ (.A1(_1005_),
    .A2(_1338_),
    .B1(_1336_),
    .B2(_1027_),
    .C1(_1464_),
    .X(_1465_));
 sky130_fd_sc_hd__o211a_1 _4915_ (.A1(_1025_),
    .A2(_1345_),
    .B1(_1462_),
    .C1(_1465_),
    .X(_1466_));
 sky130_fd_sc_hd__o32a_1 _4916_ (.A1(_1025_),
    .A2(_1028_),
    .A3(_1325_),
    .B1(_1418_),
    .B2(_1011_),
    .X(_1467_));
 sky130_fd_sc_hd__o22a_1 _4917_ (.A1(_1014_),
    .A2(_1322_),
    .B1(_1467_),
    .B2(_0499_),
    .X(_1468_));
 sky130_fd_sc_hd__nand2_1 _4918_ (.A(_1466_),
    .B(_1468_),
    .Y(_1469_));
 sky130_fd_sc_hd__inv_2 _4919_ (.A(\sound2.count[2] ),
    .Y(_1470_));
 sky130_fd_sc_hd__o32a_1 _4920_ (.A1(_0996_),
    .A2(_1025_),
    .A3(_1339_),
    .B1(_1393_),
    .B2(_0977_),
    .X(_1471_));
 sky130_fd_sc_hd__a21o_1 _4921_ (.A1(_1341_),
    .A2(_1322_),
    .B1(_0948_),
    .X(_1472_));
 sky130_fd_sc_hd__o22a_1 _4922_ (.A1(_1101_),
    .A2(_1333_),
    .B1(_1345_),
    .B2(_1097_),
    .X(_1473_));
 sky130_fd_sc_hd__a21o_1 _4923_ (.A1(_1347_),
    .A2(_1336_),
    .B1(_0960_),
    .X(_1474_));
 sky130_fd_sc_hd__o221a_1 _4924_ (.A1(_1041_),
    .A2(_1323_),
    .B1(_1327_),
    .B2(_1096_),
    .C1(_1474_),
    .X(_1475_));
 sky130_fd_sc_hd__o2111a_1 _4925_ (.A1(_1095_),
    .A2(_1343_),
    .B1(_1472_),
    .C1(_1473_),
    .D1(_1475_),
    .X(_1476_));
 sky130_fd_sc_hd__o211ai_2 _4926_ (.A1(_0993_),
    .A2(_1383_),
    .B1(_1471_),
    .C1(_1476_),
    .Y(_1477_));
 sky130_fd_sc_hd__xor2_1 _4927_ (.A(\sound2.count[0] ),
    .B(_1477_),
    .X(_1478_));
 sky130_fd_sc_hd__a221o_1 _4928_ (.A1(\sound2.count[1] ),
    .A2(_1404_),
    .B1(_1469_),
    .B2(_1470_),
    .C1(_1478_),
    .X(_1479_));
 sky130_fd_sc_hd__o21a_1 _4929_ (.A1(_1046_),
    .A2(_1347_),
    .B1(_1393_),
    .X(_1480_));
 sky130_fd_sc_hd__or2_1 _4930_ (.A(_1043_),
    .B(_1339_),
    .X(_1481_));
 sky130_fd_sc_hd__o221a_1 _4931_ (.A1(_1035_),
    .A2(_1323_),
    .B1(_1322_),
    .B2(_1039_),
    .C1(_1481_),
    .X(_1482_));
 sky130_fd_sc_hd__o21a_1 _4932_ (.A1(_0944_),
    .A2(_1336_),
    .B1(_1345_),
    .X(_1483_));
 sky130_fd_sc_hd__o22a_1 _4933_ (.A1(_1041_),
    .A2(_1343_),
    .B1(_1333_),
    .B2(_1129_),
    .X(_1484_));
 sky130_fd_sc_hd__nor2_1 _4934_ (.A(_0977_),
    .B(_1419_),
    .Y(_1485_));
 sky130_fd_sc_hd__o32a_1 _4935_ (.A1(_0947_),
    .A2(_1325_),
    .A3(_1485_),
    .B1(_1033_),
    .B2(_1341_),
    .X(_1486_));
 sky130_fd_sc_hd__o211a_1 _4936_ (.A1(_1004_),
    .A2(_1483_),
    .B1(_1484_),
    .C1(_1486_),
    .X(_1487_));
 sky130_fd_sc_hd__o211a_2 _4937_ (.A1(_1001_),
    .A2(_1480_),
    .B1(_1482_),
    .C1(_1487_),
    .X(_1488_));
 sky130_fd_sc_hd__o22a_1 _4938_ (.A1(_1077_),
    .A2(_1323_),
    .B1(_1339_),
    .B2(_1193_),
    .X(_1489_));
 sky130_fd_sc_hd__o221a_1 _4939_ (.A1(_1189_),
    .A2(_1327_),
    .B1(_1365_),
    .B2(_0959_),
    .C1(_1489_),
    .X(_1490_));
 sky130_fd_sc_hd__or2_1 _4940_ (.A(_1028_),
    .B(_1341_),
    .X(_1491_));
 sky130_fd_sc_hd__o221a_1 _4941_ (.A1(_1020_),
    .A2(_1333_),
    .B1(_1345_),
    .B2(_1083_),
    .C1(_1491_),
    .X(_1492_));
 sky130_fd_sc_hd__o221a_1 _4942_ (.A1(_1129_),
    .A2(_1347_),
    .B1(_1343_),
    .B2(_1014_),
    .C1(_1427_),
    .X(_1493_));
 sky130_fd_sc_hd__o221a_1 _4943_ (.A1(_1004_),
    .A2(_1321_),
    .B1(_1338_),
    .B2(_1158_),
    .C1(_1493_),
    .X(_1494_));
 sky130_fd_sc_hd__and3_1 _4944_ (.A(_1490_),
    .B(_1492_),
    .C(_1494_),
    .X(_1495_));
 sky130_fd_sc_hd__o22a_1 _4945_ (.A1(\sound2.count[11] ),
    .A2(_1488_),
    .B1(_1495_),
    .B2(\sound2.count[9] ),
    .X(_1496_));
 sky130_fd_sc_hd__o221a_1 _4946_ (.A1(_1318_),
    .A2(_1352_),
    .B1(_1396_),
    .B2(\sound2.count[5] ),
    .C1(_1496_),
    .X(_1497_));
 sky130_fd_sc_hd__a22oi_1 _4947_ (.A1(\sound2.count[11] ),
    .A2(_1488_),
    .B1(_1495_),
    .B2(\sound2.count[9] ),
    .Y(_1498_));
 sky130_fd_sc_hd__o221a_1 _4948_ (.A1(\sound2.count[8] ),
    .A2(_1412_),
    .B1(_1469_),
    .B2(_1470_),
    .C1(_1498_),
    .X(_1499_));
 sky130_fd_sc_hd__nand2_1 _4949_ (.A(_1497_),
    .B(_1499_),
    .Y(_1500_));
 sky130_fd_sc_hd__or4_1 _4950_ (.A(_1444_),
    .B(_1461_),
    .C(_1479_),
    .D(_1500_),
    .X(_1501_));
 sky130_fd_sc_hd__or4_1 _4951_ (.A(_1370_),
    .B(_1414_),
    .C(_1443_),
    .D(_1501_),
    .X(_1502_));
 sky130_fd_sc_hd__and2_1 _4952_ (.A(_1317_),
    .B(_1502_),
    .X(_1503_));
 sky130_fd_sc_hd__buf_4 _4953_ (.A(_1503_),
    .X(_1504_));
 sky130_fd_sc_hd__nand2_1 _4954_ (.A(\sound2.count[0] ),
    .B(_1504_),
    .Y(\sound2.osc.next_count[0] ));
 sky130_fd_sc_hd__or2_1 _4955_ (.A(\sound2.count[0] ),
    .B(\sound2.count[1] ),
    .X(_1505_));
 sky130_fd_sc_hd__nand2_1 _4956_ (.A(\sound2.count[0] ),
    .B(\sound2.count[1] ),
    .Y(_1506_));
 sky130_fd_sc_hd__and3_1 _4957_ (.A(_1504_),
    .B(_1505_),
    .C(_1506_),
    .X(_1507_));
 sky130_fd_sc_hd__clkbuf_1 _4958_ (.A(_1507_),
    .X(\sound2.osc.next_count[1] ));
 sky130_fd_sc_hd__nor2_1 _4959_ (.A(_1470_),
    .B(_1506_),
    .Y(_1508_));
 sky130_fd_sc_hd__nand2_1 _4960_ (.A(_1470_),
    .B(_1506_),
    .Y(_1509_));
 sky130_fd_sc_hd__and3b_1 _4961_ (.A_N(_1508_),
    .B(_1504_),
    .C(_1509_),
    .X(_1510_));
 sky130_fd_sc_hd__clkbuf_1 _4962_ (.A(_1510_),
    .X(\sound2.osc.next_count[2] ));
 sky130_fd_sc_hd__and2_1 _4963_ (.A(\sound2.count[3] ),
    .B(_1508_),
    .X(_1511_));
 sky130_fd_sc_hd__or2_1 _4964_ (.A(\sound2.count[3] ),
    .B(_1508_),
    .X(_1512_));
 sky130_fd_sc_hd__and3b_1 _4965_ (.A_N(_1511_),
    .B(_1512_),
    .C(_1504_),
    .X(_1513_));
 sky130_fd_sc_hd__clkbuf_1 _4966_ (.A(_1513_),
    .X(\sound2.osc.next_count[3] ));
 sky130_fd_sc_hd__o21ai_1 _4967_ (.A1(\sound2.count[4] ),
    .A2(_1511_),
    .B1(_1504_),
    .Y(_1514_));
 sky130_fd_sc_hd__a21oi_1 _4968_ (.A1(\sound2.count[4] ),
    .A2(_1511_),
    .B1(_1514_),
    .Y(\sound2.osc.next_count[4] ));
 sky130_fd_sc_hd__and3_1 _4969_ (.A(\sound2.count[4] ),
    .B(\sound2.count[5] ),
    .C(_1511_),
    .X(_1515_));
 sky130_fd_sc_hd__a31o_1 _4970_ (.A1(\sound2.count[3] ),
    .A2(\sound2.count[4] ),
    .A3(_1508_),
    .B1(\sound2.count[5] ),
    .X(_1516_));
 sky130_fd_sc_hd__and3b_1 _4971_ (.A_N(_1515_),
    .B(_1516_),
    .C(_1504_),
    .X(_1517_));
 sky130_fd_sc_hd__clkbuf_1 _4972_ (.A(_1517_),
    .X(\sound2.osc.next_count[5] ));
 sky130_fd_sc_hd__and2_1 _4973_ (.A(\sound2.count[6] ),
    .B(_1515_),
    .X(_1518_));
 sky130_fd_sc_hd__o21ai_1 _4974_ (.A1(\sound2.count[6] ),
    .A2(_1515_),
    .B1(_1504_),
    .Y(_1519_));
 sky130_fd_sc_hd__nor2_1 _4975_ (.A(_1518_),
    .B(_1519_),
    .Y(\sound2.osc.next_count[6] ));
 sky130_fd_sc_hd__and3_1 _4976_ (.A(\sound2.count[6] ),
    .B(\sound2.count[7] ),
    .C(_1515_),
    .X(_1520_));
 sky130_fd_sc_hd__o21ai_1 _4977_ (.A1(\sound2.count[7] ),
    .A2(_1518_),
    .B1(_1504_),
    .Y(_1521_));
 sky130_fd_sc_hd__nor2_1 _4978_ (.A(_1520_),
    .B(_1521_),
    .Y(\sound2.osc.next_count[7] ));
 sky130_fd_sc_hd__and2_1 _4979_ (.A(\sound2.count[8] ),
    .B(_1520_),
    .X(_1522_));
 sky130_fd_sc_hd__o21ai_1 _4980_ (.A1(\sound2.count[8] ),
    .A2(_1520_),
    .B1(_1504_),
    .Y(_1523_));
 sky130_fd_sc_hd__nor2_1 _4981_ (.A(_1522_),
    .B(_1523_),
    .Y(\sound2.osc.next_count[8] ));
 sky130_fd_sc_hd__and3_1 _4982_ (.A(\sound2.count[8] ),
    .B(\sound2.count[9] ),
    .C(_1520_),
    .X(_1524_));
 sky130_fd_sc_hd__o21ai_1 _4983_ (.A1(\sound2.count[9] ),
    .A2(_1522_),
    .B1(_1504_),
    .Y(_1525_));
 sky130_fd_sc_hd__nor2_1 _4984_ (.A(_1524_),
    .B(_1525_),
    .Y(\sound2.osc.next_count[9] ));
 sky130_fd_sc_hd__o21ai_1 _4985_ (.A1(\sound2.count[10] ),
    .A2(_1524_),
    .B1(_1504_),
    .Y(_1526_));
 sky130_fd_sc_hd__a21oi_1 _4986_ (.A1(\sound2.count[10] ),
    .A2(_1524_),
    .B1(_1526_),
    .Y(\sound2.osc.next_count[10] ));
 sky130_fd_sc_hd__and3_1 _4987_ (.A(\sound2.count[10] ),
    .B(\sound2.count[11] ),
    .C(_1524_),
    .X(_1527_));
 sky130_fd_sc_hd__a21o_1 _4988_ (.A1(\sound2.count[10] ),
    .A2(_1524_),
    .B1(\sound2.count[11] ),
    .X(_1528_));
 sky130_fd_sc_hd__and3b_1 _4989_ (.A_N(_1527_),
    .B(_1528_),
    .C(_1504_),
    .X(_1529_));
 sky130_fd_sc_hd__clkbuf_1 _4990_ (.A(_1529_),
    .X(\sound2.osc.next_count[11] ));
 sky130_fd_sc_hd__and2_1 _4991_ (.A(\sound2.count[12] ),
    .B(_1527_),
    .X(_1530_));
 sky130_fd_sc_hd__o21ai_1 _4992_ (.A1(\sound2.count[12] ),
    .A2(_1527_),
    .B1(_1504_),
    .Y(_1531_));
 sky130_fd_sc_hd__nor2_1 _4993_ (.A(_1530_),
    .B(_1531_),
    .Y(\sound2.osc.next_count[12] ));
 sky130_fd_sc_hd__o21ai_1 _4994_ (.A1(\sound2.count[13] ),
    .A2(_1530_),
    .B1(_1504_),
    .Y(_1532_));
 sky130_fd_sc_hd__a21oi_1 _4995_ (.A1(\sound2.count[13] ),
    .A2(_1530_),
    .B1(_1532_),
    .Y(\sound2.osc.next_count[13] ));
 sky130_fd_sc_hd__and3_1 _4996_ (.A(\sound2.count[13] ),
    .B(\sound2.count[14] ),
    .C(_1530_),
    .X(_1533_));
 sky130_fd_sc_hd__a31o_1 _4997_ (.A1(\sound2.count[12] ),
    .A2(\sound2.count[13] ),
    .A3(_1527_),
    .B1(\sound2.count[14] ),
    .X(_1534_));
 sky130_fd_sc_hd__and3b_1 _4998_ (.A_N(_1533_),
    .B(_1534_),
    .C(_1504_),
    .X(_1535_));
 sky130_fd_sc_hd__clkbuf_1 _4999_ (.A(_1535_),
    .X(\sound2.osc.next_count[14] ));
 sky130_fd_sc_hd__and2_1 _5000_ (.A(\sound2.count[15] ),
    .B(_1533_),
    .X(_1536_));
 sky130_fd_sc_hd__o21ai_1 _5001_ (.A1(\sound2.count[15] ),
    .A2(_1533_),
    .B1(_1504_),
    .Y(_1537_));
 sky130_fd_sc_hd__nor2_1 _5002_ (.A(_1536_),
    .B(_1537_),
    .Y(\sound2.osc.next_count[15] ));
 sky130_fd_sc_hd__o21ai_1 _5003_ (.A1(\sound2.count[16] ),
    .A2(_1536_),
    .B1(_1504_),
    .Y(_1538_));
 sky130_fd_sc_hd__a21oi_1 _5004_ (.A1(\sound2.count[16] ),
    .A2(_1536_),
    .B1(_1538_),
    .Y(\sound2.osc.next_count[16] ));
 sky130_fd_sc_hd__and3_1 _5005_ (.A(\sound2.count[16] ),
    .B(\sound2.count[17] ),
    .C(_1536_),
    .X(_1539_));
 sky130_fd_sc_hd__a31o_1 _5006_ (.A1(\sound2.count[15] ),
    .A2(\sound2.count[16] ),
    .A3(_1533_),
    .B1(\sound2.count[17] ),
    .X(_1540_));
 sky130_fd_sc_hd__and3b_1 _5007_ (.A_N(_1539_),
    .B(_1540_),
    .C(_1504_),
    .X(_1541_));
 sky130_fd_sc_hd__clkbuf_1 _5008_ (.A(_1541_),
    .X(\sound2.osc.next_count[17] ));
 sky130_fd_sc_hd__or2_1 _5009_ (.A(\sound2.count[18] ),
    .B(_1539_),
    .X(_1542_));
 sky130_fd_sc_hd__nand2_1 _5010_ (.A(\sound2.count[18] ),
    .B(_1539_),
    .Y(_1543_));
 sky130_fd_sc_hd__and3_1 _5011_ (.A(_1504_),
    .B(_1542_),
    .C(_1543_),
    .X(_1544_));
 sky130_fd_sc_hd__clkbuf_1 _5012_ (.A(_1544_),
    .X(\sound2.osc.next_count[18] ));
 sky130_fd_sc_hd__nor2_2 _5013_ (.A(_0575_),
    .B(_0563_),
    .Y(_1545_));
 sky130_fd_sc_hd__buf_4 _5014_ (.A(_1545_),
    .X(\sound3.sdiv.next_dived ));
 sky130_fd_sc_hd__and2_1 _5015_ (.A(_0699_),
    .B(net46),
    .X(_1546_));
 sky130_fd_sc_hd__nand2_1 _5016_ (.A(_0546_),
    .B(_1546_),
    .Y(_1547_));
 sky130_fd_sc_hd__or2_1 _5017_ (.A(net56),
    .B(_1547_),
    .X(_1548_));
 sky130_fd_sc_hd__or2_1 _5018_ (.A(_0540_),
    .B(_1548_),
    .X(_1549_));
 sky130_fd_sc_hd__buf_4 _5019_ (.A(_1549_),
    .X(_1550_));
 sky130_fd_sc_hd__or3_4 _5020_ (.A(_0698_),
    .B(_0546_),
    .C(net46),
    .X(_1551_));
 sky130_fd_sc_hd__nor2_4 _5021_ (.A(net56),
    .B(_1551_),
    .Y(_1552_));
 sky130_fd_sc_hd__nand2_8 _5022_ (.A(net43),
    .B(_1552_),
    .Y(_1553_));
 sky130_fd_sc_hd__o32a_1 _5023_ (.A1(_0977_),
    .A2(_0996_),
    .A3(_1550_),
    .B1(_1553_),
    .B2(_1096_),
    .X(_1554_));
 sky130_fd_sc_hd__nor2_1 _5024_ (.A(_0698_),
    .B(_0546_),
    .Y(_1555_));
 sky130_fd_sc_hd__or2_1 _5025_ (.A(_1555_),
    .B(_1546_),
    .X(_1556_));
 sky130_fd_sc_hd__or2_1 _5026_ (.A(_0698_),
    .B(net56),
    .X(_1557_));
 sky130_fd_sc_hd__or2_1 _5027_ (.A(_1556_),
    .B(_1557_),
    .X(_1558_));
 sky130_fd_sc_hd__buf_4 _5028_ (.A(_1558_),
    .X(_1559_));
 sky130_fd_sc_hd__or3_2 _5029_ (.A(_0698_),
    .B(_0540_),
    .C(net44),
    .X(_1560_));
 sky130_fd_sc_hd__or2_1 _5030_ (.A(_1547_),
    .B(_1560_),
    .X(_1561_));
 sky130_fd_sc_hd__clkbuf_8 _5031_ (.A(_1561_),
    .X(_1562_));
 sky130_fd_sc_hd__o21ai_1 _5032_ (.A1(_0698_),
    .A2(_0540_),
    .B1(_1557_),
    .Y(_1563_));
 sky130_fd_sc_hd__or2_1 _5033_ (.A(_1547_),
    .B(_1563_),
    .X(_1564_));
 sky130_fd_sc_hd__buf_4 _5034_ (.A(_1564_),
    .X(_1565_));
 sky130_fd_sc_hd__or2_1 _5035_ (.A(_1560_),
    .B(_1551_),
    .X(_1566_));
 sky130_fd_sc_hd__buf_4 _5036_ (.A(_1566_),
    .X(_1567_));
 sky130_fd_sc_hd__nand2_2 _5037_ (.A(net46),
    .B(_1555_),
    .Y(_1568_));
 sky130_fd_sc_hd__or2_1 _5038_ (.A(_1563_),
    .B(_1568_),
    .X(_1569_));
 sky130_fd_sc_hd__buf_4 _5039_ (.A(_1569_),
    .X(_1570_));
 sky130_fd_sc_hd__or2_1 _5040_ (.A(net43),
    .B(_1548_),
    .X(_1571_));
 sky130_fd_sc_hd__buf_4 _5041_ (.A(_1571_),
    .X(_1572_));
 sky130_fd_sc_hd__or2_1 _5042_ (.A(_1560_),
    .B(_1568_),
    .X(_1573_));
 sky130_fd_sc_hd__buf_4 _5043_ (.A(_1573_),
    .X(_1574_));
 sky130_fd_sc_hd__a21o_1 _5044_ (.A1(_1572_),
    .A2(_1574_),
    .B1(_0960_),
    .X(_1575_));
 sky130_fd_sc_hd__o221a_1 _5045_ (.A1(_1095_),
    .A2(_1567_),
    .B1(_1570_),
    .B2(_1097_),
    .C1(_1575_),
    .X(_1576_));
 sky130_fd_sc_hd__o221a_1 _5046_ (.A1(_1041_),
    .A2(_1562_),
    .B1(_1565_),
    .B2(_1101_),
    .C1(_1576_),
    .X(_1577_));
 sky130_fd_sc_hd__nand2_8 _5047_ (.A(_0540_),
    .B(_1552_),
    .Y(_1578_));
 sky130_fd_sc_hd__or2_1 _5048_ (.A(_1551_),
    .B(_1563_),
    .X(_1579_));
 sky130_fd_sc_hd__buf_4 _5049_ (.A(_1579_),
    .X(_1580_));
 sky130_fd_sc_hd__o32a_1 _5050_ (.A1(_0993_),
    .A2(_1012_),
    .A3(_1578_),
    .B1(_1580_),
    .B2(_0948_),
    .X(_1581_));
 sky130_fd_sc_hd__o311a_1 _5051_ (.A1(_0996_),
    .A2(_1025_),
    .A3(_1559_),
    .B1(_1577_),
    .C1(_1581_),
    .X(_1582_));
 sky130_fd_sc_hd__nand2_1 _5052_ (.A(_1554_),
    .B(_1582_),
    .Y(_1583_));
 sky130_fd_sc_hd__xor2_1 _5053_ (.A(\sound3.count[0] ),
    .B(_1583_),
    .X(_1584_));
 sky130_fd_sc_hd__o32a_1 _5054_ (.A1(_0959_),
    .A2(_1133_),
    .A3(_1553_),
    .B1(_1578_),
    .B2(_0983_),
    .X(_1585_));
 sky130_fd_sc_hd__o221a_1 _5055_ (.A1(_1057_),
    .A2(_1567_),
    .B1(_1565_),
    .B2(_1056_),
    .C1(_1585_),
    .X(_1586_));
 sky130_fd_sc_hd__or2_1 _5056_ (.A(_0677_),
    .B(_1574_),
    .X(_1587_));
 sky130_fd_sc_hd__o32a_1 _5057_ (.A1(_0679_),
    .A2(net63),
    .A3(_1550_),
    .B1(_1580_),
    .B2(_1053_),
    .X(_1588_));
 sky130_fd_sc_hd__o221a_1 _5058_ (.A1(_1059_),
    .A2(_1562_),
    .B1(_1570_),
    .B2(_1063_),
    .C1(_1588_),
    .X(_1589_));
 sky130_fd_sc_hd__inv_2 _5059_ (.A(_1557_),
    .Y(_1590_));
 sky130_fd_sc_hd__or2_4 _5060_ (.A(_1556_),
    .B(_1590_),
    .X(_1591_));
 sky130_fd_sc_hd__o221a_1 _5061_ (.A1(_1026_),
    .A2(_1559_),
    .B1(_1572_),
    .B2(_1064_),
    .C1(_1591_),
    .X(_1592_));
 sky130_fd_sc_hd__o211a_1 _5062_ (.A1(_1038_),
    .A2(_1587_),
    .B1(_1589_),
    .C1(_1592_),
    .X(_1593_));
 sky130_fd_sc_hd__nand2_1 _5063_ (.A(_1586_),
    .B(_1593_),
    .Y(_1594_));
 sky130_fd_sc_hd__xor2_1 _5064_ (.A(\sound3.count[6] ),
    .B(_1594_),
    .X(_1595_));
 sky130_fd_sc_hd__o22a_1 _5065_ (.A1(_1138_),
    .A2(_1562_),
    .B1(_1567_),
    .B2(_0696_),
    .X(_1596_));
 sky130_fd_sc_hd__o221a_1 _5066_ (.A1(_1129_),
    .A2(_1572_),
    .B1(_1574_),
    .B2(_1141_),
    .C1(_1596_),
    .X(_1597_));
 sky130_fd_sc_hd__o221a_1 _5067_ (.A1(_1134_),
    .A2(_1578_),
    .B1(_1553_),
    .B2(_1139_),
    .C1(_1597_),
    .X(_1598_));
 sky130_fd_sc_hd__o221a_1 _5068_ (.A1(_1123_),
    .A2(_1559_),
    .B1(_1565_),
    .B2(_1127_),
    .C1(_1591_),
    .X(_1599_));
 sky130_fd_sc_hd__o211a_1 _5069_ (.A1(_1126_),
    .A2(_1580_),
    .B1(_1598_),
    .C1(_1599_),
    .X(_1600_));
 sky130_fd_sc_hd__o221a_1 _5070_ (.A1(_1135_),
    .A2(_1550_),
    .B1(_1570_),
    .B2(_1140_),
    .C1(_1600_),
    .X(_1601_));
 sky130_fd_sc_hd__xnor2_1 _5071_ (.A(\sound3.count[4] ),
    .B(_1601_),
    .Y(_1602_));
 sky130_fd_sc_hd__nor2_1 _5072_ (.A(_1556_),
    .B(_1557_),
    .Y(_1603_));
 sky130_fd_sc_hd__a22o_1 _5073_ (.A1(_1018_),
    .A2(_1556_),
    .B1(_1603_),
    .B2(_0971_),
    .X(_1604_));
 sky130_fd_sc_hd__xor2_1 _5074_ (.A(\sound3.count[17] ),
    .B(_1604_),
    .X(_1605_));
 sky130_fd_sc_hd__a31o_1 _5075_ (.A1(_1562_),
    .A2(_1548_),
    .A3(_1568_),
    .B1(_1010_),
    .X(_1606_));
 sky130_fd_sc_hd__a21o_1 _5076_ (.A1(_1551_),
    .A2(_1565_),
    .B1(_1055_),
    .X(_1607_));
 sky130_fd_sc_hd__o2111a_1 _5077_ (.A1(_0688_),
    .A2(_1559_),
    .B1(_1591_),
    .C1(_1606_),
    .D1(_1607_),
    .X(_1608_));
 sky130_fd_sc_hd__xnor2_1 _5078_ (.A(\sound3.count[16] ),
    .B(_1608_),
    .Y(_1609_));
 sky130_fd_sc_hd__a21o_1 _5079_ (.A1(_1562_),
    .A2(_1548_),
    .B1(_0869_),
    .X(_1610_));
 sky130_fd_sc_hd__or2_1 _5080_ (.A(net56),
    .B(_1551_),
    .X(_1611_));
 sky130_fd_sc_hd__a21o_1 _5081_ (.A1(_1611_),
    .A2(_1565_),
    .B1(_1213_),
    .X(_1612_));
 sky130_fd_sc_hd__o22a_1 _5082_ (.A1(_1138_),
    .A2(_1551_),
    .B1(_1568_),
    .B2(_0688_),
    .X(_1613_));
 sky130_fd_sc_hd__o221a_1 _5083_ (.A1(_1011_),
    .A2(_1559_),
    .B1(_1613_),
    .B2(_1590_),
    .C1(_1591_),
    .X(_1614_));
 sky130_fd_sc_hd__and3_1 _5084_ (.A(_1610_),
    .B(_1612_),
    .C(_1614_),
    .X(_1615_));
 sky130_fd_sc_hd__xnor2_1 _5085_ (.A(\sound3.count[15] ),
    .B(_1615_),
    .Y(_1616_));
 sky130_fd_sc_hd__nand2_1 _5086_ (.A(net64),
    .B(_1603_),
    .Y(_1617_));
 sky130_fd_sc_hd__o21a_1 _5087_ (.A1(_0695_),
    .A2(_1617_),
    .B1(_1591_),
    .X(_1618_));
 sky130_fd_sc_hd__xnor2_1 _5088_ (.A(\sound3.count[18] ),
    .B(_1618_),
    .Y(_1619_));
 sky130_fd_sc_hd__or4_1 _5089_ (.A(_1605_),
    .B(_1609_),
    .C(_1616_),
    .D(_1619_),
    .X(_1620_));
 sky130_fd_sc_hd__or4_1 _5090_ (.A(_1584_),
    .B(_1595_),
    .C(_1602_),
    .D(_1620_),
    .X(_1621_));
 sky130_fd_sc_hd__nor2_1 _5091_ (.A(_0695_),
    .B(_0540_),
    .Y(_1622_));
 sky130_fd_sc_hd__o22a_1 _5092_ (.A1(_1111_),
    .A2(_1611_),
    .B1(_1568_),
    .B2(_1058_),
    .X(_1623_));
 sky130_fd_sc_hd__o221a_1 _5093_ (.A1(_1062_),
    .A2(_1565_),
    .B1(_1617_),
    .B2(_1622_),
    .C1(_1623_),
    .X(_1624_));
 sky130_fd_sc_hd__and2_1 _5094_ (.A(_1562_),
    .B(_1572_),
    .X(_1625_));
 sky130_fd_sc_hd__o221a_1 _5095_ (.A1(net64),
    .A2(_1567_),
    .B1(_1625_),
    .B2(_0687_),
    .C1(_1580_),
    .X(_1626_));
 sky130_fd_sc_hd__o22a_1 _5096_ (.A1(_1095_),
    .A2(_1550_),
    .B1(_1626_),
    .B2(_0695_),
    .X(_1627_));
 sky130_fd_sc_hd__nand2_1 _5097_ (.A(_1624_),
    .B(_1627_),
    .Y(_1628_));
 sky130_fd_sc_hd__xor2_1 _5098_ (.A(\sound3.count[14] ),
    .B(_1628_),
    .X(_1629_));
 sky130_fd_sc_hd__o22a_1 _5099_ (.A1(_1180_),
    .A2(_1553_),
    .B1(_1565_),
    .B2(_1174_),
    .X(_1630_));
 sky130_fd_sc_hd__o22a_1 _5100_ (.A1(_1026_),
    .A2(_1567_),
    .B1(_1574_),
    .B2(_1175_),
    .X(_1631_));
 sky130_fd_sc_hd__o221a_1 _5101_ (.A1(_1129_),
    .A2(_1580_),
    .B1(_1570_),
    .B2(_1182_),
    .C1(_1631_),
    .X(_1632_));
 sky130_fd_sc_hd__o211a_1 _5102_ (.A1(_0996_),
    .A2(_1550_),
    .B1(_1630_),
    .C1(_1632_),
    .X(_1633_));
 sky130_fd_sc_hd__o221a_1 _5103_ (.A1(_1176_),
    .A2(_1562_),
    .B1(_1572_),
    .B2(_0954_),
    .C1(_1633_),
    .X(_1634_));
 sky130_fd_sc_hd__o221a_2 _5104_ (.A1(_1181_),
    .A2(_1559_),
    .B1(_1578_),
    .B2(_1028_),
    .C1(_1634_),
    .X(_1635_));
 sky130_fd_sc_hd__o32a_1 _5105_ (.A1(_0683_),
    .A2(_1107_),
    .A3(_1570_),
    .B1(_1562_),
    .B2(_1198_),
    .X(_1636_));
 sky130_fd_sc_hd__o221a_1 _5106_ (.A1(_1200_),
    .A2(_1567_),
    .B1(_1550_),
    .B2(_0686_),
    .C1(_1636_),
    .X(_1637_));
 sky130_fd_sc_hd__o22a_1 _5107_ (.A1(_1204_),
    .A2(_1553_),
    .B1(_1580_),
    .B2(_1199_),
    .X(_1638_));
 sky130_fd_sc_hd__o211a_1 _5108_ (.A1(_1189_),
    .A2(_1565_),
    .B1(_1637_),
    .C1(_1638_),
    .X(_1639_));
 sky130_fd_sc_hd__o221a_1 _5109_ (.A1(_1146_),
    .A2(_1572_),
    .B1(_1574_),
    .B2(_1125_),
    .C1(_1639_),
    .X(_1640_));
 sky130_fd_sc_hd__o221a_2 _5110_ (.A1(_0688_),
    .A2(_1559_),
    .B1(_1578_),
    .B2(_1014_),
    .C1(_1640_),
    .X(_1641_));
 sky130_fd_sc_hd__inv_2 _5111_ (.A(\sound3.count[7] ),
    .Y(_1642_));
 sky130_fd_sc_hd__o32a_1 _5112_ (.A1(net64),
    .A2(_1077_),
    .A3(_1567_),
    .B1(_1553_),
    .B2(_0946_),
    .X(_1643_));
 sky130_fd_sc_hd__o22a_1 _5113_ (.A1(_1079_),
    .A2(_1580_),
    .B1(_1574_),
    .B2(_0680_),
    .X(_1644_));
 sky130_fd_sc_hd__o221a_1 _5114_ (.A1(_1015_),
    .A2(_1562_),
    .B1(_1570_),
    .B2(_0952_),
    .C1(_1644_),
    .X(_1645_));
 sky130_fd_sc_hd__o22a_1 _5115_ (.A1(_1078_),
    .A2(_1559_),
    .B1(_1572_),
    .B2(_1039_),
    .X(_1646_));
 sky130_fd_sc_hd__o221a_1 _5116_ (.A1(_1083_),
    .A2(_1550_),
    .B1(_1565_),
    .B2(_0960_),
    .C1(_1646_),
    .X(_1647_));
 sky130_fd_sc_hd__o211a_1 _5117_ (.A1(_0971_),
    .A2(_1578_),
    .B1(_1645_),
    .C1(_1647_),
    .X(_1648_));
 sky130_fd_sc_hd__nand2_1 _5118_ (.A(_1643_),
    .B(_1648_),
    .Y(_1649_));
 sky130_fd_sc_hd__o22a_1 _5119_ (.A1(_1010_),
    .A2(_1567_),
    .B1(_1574_),
    .B2(_1027_),
    .X(_1650_));
 sky130_fd_sc_hd__o22a_1 _5120_ (.A1(_1016_),
    .A2(_1580_),
    .B1(_1570_),
    .B2(_1024_),
    .X(_1651_));
 sky130_fd_sc_hd__o221a_1 _5121_ (.A1(_0997_),
    .A2(_1562_),
    .B1(_1565_),
    .B2(_0973_),
    .C1(_1651_),
    .X(_1652_));
 sky130_fd_sc_hd__o221a_1 _5122_ (.A1(_1011_),
    .A2(_1559_),
    .B1(_1572_),
    .B2(_1020_),
    .C1(_1652_),
    .X(_1653_));
 sky130_fd_sc_hd__o311a_1 _5123_ (.A1(_1025_),
    .A2(_1028_),
    .A3(_1553_),
    .B1(_1650_),
    .C1(_1653_),
    .X(_1654_));
 sky130_fd_sc_hd__o221a_2 _5124_ (.A1(_1005_),
    .A2(_1578_),
    .B1(_1550_),
    .B2(_1017_),
    .C1(_1654_),
    .X(_1655_));
 sky130_fd_sc_hd__a22o_1 _5125_ (.A1(_1642_),
    .A2(_1649_),
    .B1(_1655_),
    .B2(\sound3.count[2] ),
    .X(_1656_));
 sky130_fd_sc_hd__a221o_1 _5126_ (.A1(\sound3.count[5] ),
    .A2(_1635_),
    .B1(_1641_),
    .B2(\sound3.count[3] ),
    .C1(_1656_),
    .X(_1657_));
 sky130_fd_sc_hd__inv_2 _5127_ (.A(\sound3.count[13] ),
    .Y(_1658_));
 sky130_fd_sc_hd__o21a_1 _5128_ (.A1(_0683_),
    .A2(_1562_),
    .B1(_1580_),
    .X(_1659_));
 sky130_fd_sc_hd__o32a_1 _5129_ (.A1(_0677_),
    .A2(_1083_),
    .A3(_1550_),
    .B1(_1659_),
    .B2(_1107_),
    .X(_1660_));
 sky130_fd_sc_hd__o32a_1 _5130_ (.A1(_0687_),
    .A2(_1001_),
    .A3(_1578_),
    .B1(_1572_),
    .B2(_1116_),
    .X(_1661_));
 sky130_fd_sc_hd__or2_1 _5131_ (.A(_1064_),
    .B(_1565_),
    .X(_1662_));
 sky130_fd_sc_hd__o221a_1 _5132_ (.A1(_1113_),
    .A2(_1570_),
    .B1(_1574_),
    .B2(_1112_),
    .C1(_1662_),
    .X(_1663_));
 sky130_fd_sc_hd__o221a_1 _5133_ (.A1(_1016_),
    .A2(_1553_),
    .B1(_1567_),
    .B2(_0997_),
    .C1(_1663_),
    .X(_1664_));
 sky130_fd_sc_hd__o311a_1 _5134_ (.A1(_0952_),
    .A2(_1025_),
    .A3(_1559_),
    .B1(_1661_),
    .C1(_1664_),
    .X(_1665_));
 sky130_fd_sc_hd__and3_1 _5135_ (.A(_1591_),
    .B(_1660_),
    .C(_1665_),
    .X(_1666_));
 sky130_fd_sc_hd__inv_2 _5136_ (.A(_1666_),
    .Y(_1667_));
 sky130_fd_sc_hd__o32a_1 _5137_ (.A1(_0978_),
    .A2(_0944_),
    .A3(_1565_),
    .B1(_1572_),
    .B2(_0997_),
    .X(_1668_));
 sky130_fd_sc_hd__o32a_1 _5138_ (.A1(_0959_),
    .A2(_0993_),
    .A3(_1580_),
    .B1(_1562_),
    .B2(_0985_),
    .X(_1669_));
 sky130_fd_sc_hd__o221a_1 _5139_ (.A1(_0869_),
    .A2(_1567_),
    .B1(_1550_),
    .B2(_0954_),
    .C1(_1669_),
    .X(_1670_));
 sky130_fd_sc_hd__o221a_1 _5140_ (.A1(_0973_),
    .A2(_1553_),
    .B1(_1574_),
    .B2(_0979_),
    .C1(_1670_),
    .X(_1671_));
 sky130_fd_sc_hd__o211a_1 _5141_ (.A1(_1001_),
    .A2(_1570_),
    .B1(_1668_),
    .C1(_1671_),
    .X(_1672_));
 sky130_fd_sc_hd__o211a_2 _5142_ (.A1(_0948_),
    .A2(_1578_),
    .B1(_1617_),
    .C1(_1672_),
    .X(_1673_));
 sky130_fd_sc_hd__o22a_1 _5143_ (.A1(\sound3.count[1] ),
    .A2(_1673_),
    .B1(_1635_),
    .B2(\sound3.count[5] ),
    .X(_1674_));
 sky130_fd_sc_hd__o32a_1 _5144_ (.A1(_1004_),
    .A2(_1133_),
    .A3(_1559_),
    .B1(_1565_),
    .B2(_0954_),
    .X(_1675_));
 sky130_fd_sc_hd__o22a_1 _5145_ (.A1(_0985_),
    .A2(_1567_),
    .B1(_1570_),
    .B2(_1238_),
    .X(_1676_));
 sky130_fd_sc_hd__o221a_1 _5146_ (.A1(_1245_),
    .A2(_1580_),
    .B1(_1574_),
    .B2(_1110_),
    .C1(_1676_),
    .X(_1677_));
 sky130_fd_sc_hd__a211o_1 _5147_ (.A1(_1038_),
    .A2(_1562_),
    .B1(_1625_),
    .C1(_1025_),
    .X(_1678_));
 sky130_fd_sc_hd__o22a_1 _5148_ (.A1(_1240_),
    .A2(_1578_),
    .B1(_1550_),
    .B2(_1242_),
    .X(_1679_));
 sky130_fd_sc_hd__o211a_1 _5149_ (.A1(_1101_),
    .A2(_1553_),
    .B1(_1678_),
    .C1(_1679_),
    .X(_1680_));
 sky130_fd_sc_hd__and3_2 _5150_ (.A(_1675_),
    .B(_1677_),
    .C(_1680_),
    .X(_1681_));
 sky130_fd_sc_hd__o2bb2a_1 _5151_ (.A1_N(\sound3.count[1] ),
    .A2_N(_1673_),
    .B1(_1666_),
    .B2(\sound3.count[13] ),
    .X(_1682_));
 sky130_fd_sc_hd__o221a_1 _5152_ (.A1(\sound3.count[12] ),
    .A2(_1681_),
    .B1(_1655_),
    .B2(\sound3.count[2] ),
    .C1(_1682_),
    .X(_1683_));
 sky130_fd_sc_hd__o221a_1 _5153_ (.A1(_1095_),
    .A2(_1559_),
    .B1(_1553_),
    .B2(_1127_),
    .C1(_1591_),
    .X(_1684_));
 sky130_fd_sc_hd__o22a_1 _5154_ (.A1(_1151_),
    .A2(_1562_),
    .B1(_1574_),
    .B2(_1042_),
    .X(_1685_));
 sky130_fd_sc_hd__o221a_1 _5155_ (.A1(_1134_),
    .A2(_1567_),
    .B1(_1570_),
    .B2(_1154_),
    .C1(_1685_),
    .X(_1686_));
 sky130_fd_sc_hd__o22a_1 _5156_ (.A1(_0983_),
    .A2(_1580_),
    .B1(_1565_),
    .B2(_1146_),
    .X(_1687_));
 sky130_fd_sc_hd__o221a_1 _5157_ (.A1(_1053_),
    .A2(_1572_),
    .B1(_1550_),
    .B2(_1125_),
    .C1(_1687_),
    .X(_1688_));
 sky130_fd_sc_hd__o211a_1 _5158_ (.A1(_1012_),
    .A2(_1578_),
    .B1(_1686_),
    .C1(_1688_),
    .X(_1689_));
 sky130_fd_sc_hd__nand2_2 _5159_ (.A(_1684_),
    .B(_1689_),
    .Y(_1690_));
 sky130_fd_sc_hd__xnor2_1 _5160_ (.A(\sound3.count[10] ),
    .B(_1690_),
    .Y(_1691_));
 sky130_fd_sc_hd__o2111ai_1 _5161_ (.A1(_1658_),
    .A2(_1667_),
    .B1(_1674_),
    .C1(_1683_),
    .D1(_1691_),
    .Y(_1692_));
 sky130_fd_sc_hd__o21a_1 _5162_ (.A1(_0944_),
    .A2(_1574_),
    .B1(_1570_),
    .X(_1693_));
 sky130_fd_sc_hd__o22a_1 _5163_ (.A1(_1046_),
    .A2(_1572_),
    .B1(_1550_),
    .B2(_0996_),
    .X(_1694_));
 sky130_fd_sc_hd__nor2_1 _5164_ (.A(_0540_),
    .B(_1213_),
    .Y(_1695_));
 sky130_fd_sc_hd__o32a_1 _5165_ (.A1(_0947_),
    .A2(_1611_),
    .A3(_1695_),
    .B1(_1035_),
    .B2(_1562_),
    .X(_1696_));
 sky130_fd_sc_hd__o221a_1 _5166_ (.A1(_1041_),
    .A2(_1567_),
    .B1(_1565_),
    .B2(_1129_),
    .C1(_1696_),
    .X(_1697_));
 sky130_fd_sc_hd__o221a_1 _5167_ (.A1(_1004_),
    .A2(_1693_),
    .B1(_1694_),
    .B2(_1001_),
    .C1(_1697_),
    .X(_1698_));
 sky130_fd_sc_hd__o221a_2 _5168_ (.A1(_1043_),
    .A2(_1559_),
    .B1(_1580_),
    .B2(_1033_),
    .C1(_1698_),
    .X(_1699_));
 sky130_fd_sc_hd__o22a_1 _5169_ (.A1(_1154_),
    .A2(_1550_),
    .B1(_1570_),
    .B2(_1077_),
    .X(_1700_));
 sky130_fd_sc_hd__o221a_1 _5170_ (.A1(_0685_),
    .A2(_1562_),
    .B1(_1572_),
    .B2(_1126_),
    .C1(_1700_),
    .X(_1701_));
 sky130_fd_sc_hd__o32a_1 _5171_ (.A1(_1004_),
    .A2(_1038_),
    .A3(_1553_),
    .B1(_1580_),
    .B2(_1166_),
    .X(_1702_));
 sky130_fd_sc_hd__o221a_1 _5172_ (.A1(_1159_),
    .A2(_1567_),
    .B1(_1565_),
    .B2(_0997_),
    .C1(_1702_),
    .X(_1703_));
 sky130_fd_sc_hd__o32a_1 _5173_ (.A1(_1025_),
    .A2(_1046_),
    .A3(_1559_),
    .B1(_1578_),
    .B2(_1165_),
    .X(_1704_));
 sky130_fd_sc_hd__and4_1 _5174_ (.A(_1591_),
    .B(_1703_),
    .C(_1587_),
    .D(_1704_),
    .X(_1705_));
 sky130_fd_sc_hd__and2_1 _5175_ (.A(_1701_),
    .B(_1705_),
    .X(_1706_));
 sky130_fd_sc_hd__xnor2_1 _5176_ (.A(\sound3.count[8] ),
    .B(_1706_),
    .Y(_1707_));
 sky130_fd_sc_hd__o22a_1 _5177_ (.A1(_1014_),
    .A2(_1567_),
    .B1(_1570_),
    .B2(_1083_),
    .X(_1708_));
 sky130_fd_sc_hd__o221a_1 _5178_ (.A1(_1158_),
    .A2(_1578_),
    .B1(_1550_),
    .B2(_1004_),
    .C1(_1708_),
    .X(_1709_));
 sky130_fd_sc_hd__or3_1 _5179_ (.A(_0680_),
    .B(_0959_),
    .C(_1574_),
    .X(_1710_));
 sky130_fd_sc_hd__o221a_1 _5180_ (.A1(_1193_),
    .A2(_1559_),
    .B1(_1572_),
    .B2(_1129_),
    .C1(_1710_),
    .X(_1711_));
 sky130_fd_sc_hd__o22a_1 _5181_ (.A1(_1077_),
    .A2(_1562_),
    .B1(_1565_),
    .B2(_1020_),
    .X(_1712_));
 sky130_fd_sc_hd__o221a_1 _5182_ (.A1(_1189_),
    .A2(_1553_),
    .B1(_1580_),
    .B2(_1028_),
    .C1(_1712_),
    .X(_1713_));
 sky130_fd_sc_hd__and3_1 _5183_ (.A(_1709_),
    .B(_1711_),
    .C(_1713_),
    .X(_1714_));
 sky130_fd_sc_hd__o2bb2a_1 _5184_ (.A1_N(\sound3.count[9] ),
    .A2_N(_1714_),
    .B1(_1699_),
    .B2(\sound3.count[11] ),
    .X(_1715_));
 sky130_fd_sc_hd__o221ai_1 _5185_ (.A1(_1642_),
    .A2(_1649_),
    .B1(_1714_),
    .B2(\sound3.count[9] ),
    .C1(_1715_),
    .Y(_1716_));
 sky130_fd_sc_hd__a2bb2o_1 _5186_ (.A1_N(\sound3.count[3] ),
    .A2_N(_1641_),
    .B1(_1681_),
    .B2(\sound3.count[12] ),
    .X(_1717_));
 sky130_fd_sc_hd__a2111o_1 _5187_ (.A1(\sound3.count[11] ),
    .A2(_1699_),
    .B1(_1707_),
    .C1(_1716_),
    .D1(_1717_),
    .X(_1718_));
 sky130_fd_sc_hd__or4_1 _5188_ (.A(_1629_),
    .B(_1657_),
    .C(_1692_),
    .D(_1718_),
    .X(_1719_));
 sky130_fd_sc_hd__o21a_1 _5189_ (.A1(_1621_),
    .A2(_1719_),
    .B1(_1591_),
    .X(_1720_));
 sky130_fd_sc_hd__buf_4 _5190_ (.A(_1720_),
    .X(_1721_));
 sky130_fd_sc_hd__nand2_1 _5191_ (.A(\sound3.count[0] ),
    .B(_1721_),
    .Y(\sound3.osc.next_count[0] ));
 sky130_fd_sc_hd__or2_1 _5192_ (.A(\sound3.count[0] ),
    .B(\sound3.count[1] ),
    .X(_1722_));
 sky130_fd_sc_hd__nand2_1 _5193_ (.A(\sound3.count[0] ),
    .B(\sound3.count[1] ),
    .Y(_1723_));
 sky130_fd_sc_hd__and3_1 _5194_ (.A(_1721_),
    .B(_1722_),
    .C(_1723_),
    .X(_1724_));
 sky130_fd_sc_hd__clkbuf_1 _5195_ (.A(_1724_),
    .X(\sound3.osc.next_count[1] ));
 sky130_fd_sc_hd__a21o_1 _5196_ (.A1(\sound3.count[0] ),
    .A2(\sound3.count[1] ),
    .B1(\sound3.count[2] ),
    .X(_1725_));
 sky130_fd_sc_hd__nand3_1 _5197_ (.A(\sound3.count[0] ),
    .B(\sound3.count[1] ),
    .C(\sound3.count[2] ),
    .Y(_1726_));
 sky130_fd_sc_hd__and3_1 _5198_ (.A(_1721_),
    .B(_1725_),
    .C(_1726_),
    .X(_1727_));
 sky130_fd_sc_hd__clkbuf_1 _5199_ (.A(_1727_),
    .X(\sound3.osc.next_count[2] ));
 sky130_fd_sc_hd__and4_1 _5200_ (.A(\sound3.count[0] ),
    .B(\sound3.count[1] ),
    .C(\sound3.count[2] ),
    .D(\sound3.count[3] ),
    .X(_1728_));
 sky130_fd_sc_hd__a31o_1 _5201_ (.A1(\sound3.count[0] ),
    .A2(\sound3.count[1] ),
    .A3(\sound3.count[2] ),
    .B1(\sound3.count[3] ),
    .X(_1729_));
 sky130_fd_sc_hd__and3b_1 _5202_ (.A_N(_1728_),
    .B(_1729_),
    .C(_1721_),
    .X(_1730_));
 sky130_fd_sc_hd__clkbuf_1 _5203_ (.A(_1730_),
    .X(\sound3.osc.next_count[3] ));
 sky130_fd_sc_hd__o21ai_1 _5204_ (.A1(\sound3.count[4] ),
    .A2(_1728_),
    .B1(_1721_),
    .Y(_1731_));
 sky130_fd_sc_hd__a21oi_1 _5205_ (.A1(\sound3.count[4] ),
    .A2(_1728_),
    .B1(_1731_),
    .Y(\sound3.osc.next_count[4] ));
 sky130_fd_sc_hd__and3_1 _5206_ (.A(\sound3.count[4] ),
    .B(\sound3.count[5] ),
    .C(_1728_),
    .X(_1732_));
 sky130_fd_sc_hd__a21o_1 _5207_ (.A1(\sound3.count[4] ),
    .A2(_1728_),
    .B1(\sound3.count[5] ),
    .X(_1733_));
 sky130_fd_sc_hd__and3b_1 _5208_ (.A_N(_1732_),
    .B(_1733_),
    .C(_1721_),
    .X(_1734_));
 sky130_fd_sc_hd__clkbuf_1 _5209_ (.A(_1734_),
    .X(\sound3.osc.next_count[5] ));
 sky130_fd_sc_hd__and2_1 _5210_ (.A(\sound3.count[6] ),
    .B(_1732_),
    .X(_1735_));
 sky130_fd_sc_hd__o21ai_1 _5211_ (.A1(\sound3.count[6] ),
    .A2(_1732_),
    .B1(_1721_),
    .Y(_1736_));
 sky130_fd_sc_hd__nor2_1 _5212_ (.A(_1735_),
    .B(_1736_),
    .Y(\sound3.osc.next_count[6] ));
 sky130_fd_sc_hd__o21ai_1 _5213_ (.A1(\sound3.count[7] ),
    .A2(_1735_),
    .B1(_1721_),
    .Y(_1737_));
 sky130_fd_sc_hd__a21oi_1 _5214_ (.A1(\sound3.count[7] ),
    .A2(_1735_),
    .B1(_1737_),
    .Y(\sound3.osc.next_count[7] ));
 sky130_fd_sc_hd__and3_1 _5215_ (.A(\sound3.count[7] ),
    .B(\sound3.count[8] ),
    .C(_1735_),
    .X(_1738_));
 sky130_fd_sc_hd__a31o_1 _5216_ (.A1(\sound3.count[6] ),
    .A2(\sound3.count[7] ),
    .A3(_1732_),
    .B1(\sound3.count[8] ),
    .X(_1739_));
 sky130_fd_sc_hd__and3b_1 _5217_ (.A_N(_1738_),
    .B(_1739_),
    .C(_1721_),
    .X(_1740_));
 sky130_fd_sc_hd__clkbuf_1 _5218_ (.A(_1740_),
    .X(\sound3.osc.next_count[8] ));
 sky130_fd_sc_hd__and2_1 _5219_ (.A(\sound3.count[9] ),
    .B(_1738_),
    .X(_1741_));
 sky130_fd_sc_hd__o21ai_1 _5220_ (.A1(\sound3.count[9] ),
    .A2(_1738_),
    .B1(_1721_),
    .Y(_1742_));
 sky130_fd_sc_hd__nor2_1 _5221_ (.A(_1741_),
    .B(_1742_),
    .Y(\sound3.osc.next_count[9] ));
 sky130_fd_sc_hd__o21ai_1 _5222_ (.A1(\sound3.count[10] ),
    .A2(_1741_),
    .B1(_1721_),
    .Y(_1743_));
 sky130_fd_sc_hd__a21oi_1 _5223_ (.A1(\sound3.count[10] ),
    .A2(_1741_),
    .B1(_1743_),
    .Y(\sound3.osc.next_count[10] ));
 sky130_fd_sc_hd__and3_1 _5224_ (.A(\sound3.count[10] ),
    .B(\sound3.count[11] ),
    .C(_1741_),
    .X(_1744_));
 sky130_fd_sc_hd__a31o_1 _5225_ (.A1(\sound3.count[9] ),
    .A2(\sound3.count[10] ),
    .A3(_1738_),
    .B1(\sound3.count[11] ),
    .X(_1745_));
 sky130_fd_sc_hd__and3b_1 _5226_ (.A_N(_1744_),
    .B(_1745_),
    .C(_1721_),
    .X(_1746_));
 sky130_fd_sc_hd__clkbuf_1 _5227_ (.A(_1746_),
    .X(\sound3.osc.next_count[11] ));
 sky130_fd_sc_hd__and2_1 _5228_ (.A(\sound3.count[12] ),
    .B(_1744_),
    .X(_1747_));
 sky130_fd_sc_hd__o21ai_1 _5229_ (.A1(\sound3.count[12] ),
    .A2(_1744_),
    .B1(_1721_),
    .Y(_1748_));
 sky130_fd_sc_hd__nor2_1 _5230_ (.A(_1747_),
    .B(_1748_),
    .Y(\sound3.osc.next_count[12] ));
 sky130_fd_sc_hd__o21ai_1 _5231_ (.A1(\sound3.count[13] ),
    .A2(_1747_),
    .B1(_1721_),
    .Y(_1749_));
 sky130_fd_sc_hd__a21oi_1 _5232_ (.A1(\sound3.count[13] ),
    .A2(_1747_),
    .B1(_1749_),
    .Y(\sound3.osc.next_count[13] ));
 sky130_fd_sc_hd__and3_1 _5233_ (.A(\sound3.count[13] ),
    .B(\sound3.count[14] ),
    .C(_1747_),
    .X(_1750_));
 sky130_fd_sc_hd__a31o_1 _5234_ (.A1(\sound3.count[12] ),
    .A2(\sound3.count[13] ),
    .A3(_1744_),
    .B1(\sound3.count[14] ),
    .X(_1751_));
 sky130_fd_sc_hd__and3b_1 _5235_ (.A_N(_1750_),
    .B(_1751_),
    .C(_1721_),
    .X(_1752_));
 sky130_fd_sc_hd__clkbuf_1 _5236_ (.A(_1752_),
    .X(\sound3.osc.next_count[14] ));
 sky130_fd_sc_hd__and2_1 _5237_ (.A(\sound3.count[15] ),
    .B(_1750_),
    .X(_1753_));
 sky130_fd_sc_hd__o21ai_1 _5238_ (.A1(\sound3.count[15] ),
    .A2(_1750_),
    .B1(_1721_),
    .Y(_1754_));
 sky130_fd_sc_hd__nor2_1 _5239_ (.A(_1753_),
    .B(_1754_),
    .Y(\sound3.osc.next_count[15] ));
 sky130_fd_sc_hd__o21ai_1 _5240_ (.A1(\sound3.count[16] ),
    .A2(_1753_),
    .B1(_1721_),
    .Y(_1755_));
 sky130_fd_sc_hd__a21oi_1 _5241_ (.A1(\sound3.count[16] ),
    .A2(_1753_),
    .B1(_1755_),
    .Y(\sound3.osc.next_count[16] ));
 sky130_fd_sc_hd__and3_1 _5242_ (.A(\sound3.count[16] ),
    .B(\sound3.count[17] ),
    .C(_1753_),
    .X(_1756_));
 sky130_fd_sc_hd__a31o_1 _5243_ (.A1(\sound3.count[15] ),
    .A2(\sound3.count[16] ),
    .A3(_1750_),
    .B1(\sound3.count[17] ),
    .X(_1757_));
 sky130_fd_sc_hd__and3b_1 _5244_ (.A_N(_1756_),
    .B(_1757_),
    .C(_1721_),
    .X(_1758_));
 sky130_fd_sc_hd__clkbuf_1 _5245_ (.A(_1758_),
    .X(\sound3.osc.next_count[17] ));
 sky130_fd_sc_hd__or2_1 _5246_ (.A(\sound3.count[18] ),
    .B(_1756_),
    .X(_1759_));
 sky130_fd_sc_hd__nand2_1 _5247_ (.A(\sound3.count[18] ),
    .B(_1756_),
    .Y(_1760_));
 sky130_fd_sc_hd__and3_1 _5248_ (.A(_1721_),
    .B(_1759_),
    .C(_1760_),
    .X(_1761_));
 sky130_fd_sc_hd__clkbuf_1 _5249_ (.A(_1761_),
    .X(\sound3.osc.next_count[18] ));
 sky130_fd_sc_hd__or2_1 _5250_ (.A(_0575_),
    .B(_0557_),
    .X(_1762_));
 sky130_fd_sc_hd__buf_2 _5251_ (.A(_1762_),
    .X(_1763_));
 sky130_fd_sc_hd__inv_2 _5252_ (.A(_1763_),
    .Y(_1764_));
 sky130_fd_sc_hd__buf_4 _5253_ (.A(_1764_),
    .X(\sound4.sdiv.next_dived ));
 sky130_fd_sc_hd__or3_4 _5254_ (.A(_0698_),
    .B(_0606_),
    .C(net49),
    .X(_1765_));
 sky130_fd_sc_hd__and2_1 _5255_ (.A(_0699_),
    .B(net47),
    .X(_1766_));
 sky130_fd_sc_hd__nand2_1 _5256_ (.A(_0673_),
    .B(_1766_),
    .Y(_1767_));
 sky130_fd_sc_hd__or2_1 _5257_ (.A(_1765_),
    .B(_1767_),
    .X(_1768_));
 sky130_fd_sc_hd__clkbuf_8 _5258_ (.A(_1768_),
    .X(_1769_));
 sky130_fd_sc_hd__or2_1 _5259_ (.A(_0673_),
    .B(_1765_),
    .X(_1770_));
 sky130_fd_sc_hd__or2_4 _5260_ (.A(_0698_),
    .B(_0605_),
    .X(_1771_));
 sky130_fd_sc_hd__and3_1 _5261_ (.A(_1769_),
    .B(_1770_),
    .C(_1771_),
    .X(_1772_));
 sky130_fd_sc_hd__or2_4 _5262_ (.A(_0698_),
    .B(_0587_),
    .X(_1773_));
 sky130_fd_sc_hd__nor2_1 _5263_ (.A(_0698_),
    .B(_0673_),
    .Y(_1774_));
 sky130_fd_sc_hd__or2_1 _5264_ (.A(_1766_),
    .B(_1774_),
    .X(_1775_));
 sky130_fd_sc_hd__or2_1 _5265_ (.A(_1765_),
    .B(_1775_),
    .X(_1776_));
 sky130_fd_sc_hd__buf_6 _5266_ (.A(_1776_),
    .X(_1777_));
 sky130_fd_sc_hd__nand3_4 _5267_ (.A(_1772_),
    .B(_1773_),
    .C(_1777_),
    .Y(_1778_));
 sky130_fd_sc_hd__buf_4 _5268_ (.A(_1778_),
    .X(_1779_));
 sky130_fd_sc_hd__nor2_2 _5269_ (.A(net47),
    .B(_1770_),
    .Y(_1780_));
 sky130_fd_sc_hd__clkinv_4 _5270_ (.A(_1780_),
    .Y(_1781_));
 sky130_fd_sc_hd__inv_2 _5271_ (.A(_1766_),
    .Y(_1782_));
 sky130_fd_sc_hd__or2_1 _5272_ (.A(_1782_),
    .B(_1770_),
    .X(_1783_));
 sky130_fd_sc_hd__buf_4 _5273_ (.A(_1783_),
    .X(_1784_));
 sky130_fd_sc_hd__or4_2 _5274_ (.A(_0719_),
    .B(_0587_),
    .C(_0672_),
    .D(_0673_),
    .X(_1785_));
 sky130_fd_sc_hd__buf_4 _5275_ (.A(_1785_),
    .X(_1786_));
 sky130_fd_sc_hd__o22a_1 _5276_ (.A1(_1125_),
    .A2(_1784_),
    .B1(_1786_),
    .B2(_1127_),
    .X(_1787_));
 sky130_fd_sc_hd__or2_1 _5277_ (.A(_0673_),
    .B(_1773_),
    .X(_1788_));
 sky130_fd_sc_hd__or2_1 _5278_ (.A(net47),
    .B(_1788_),
    .X(_1789_));
 sky130_fd_sc_hd__clkbuf_4 _5279_ (.A(_1789_),
    .X(_1790_));
 sky130_fd_sc_hd__or2_1 _5280_ (.A(_1767_),
    .B(_1773_),
    .X(_1791_));
 sky130_fd_sc_hd__clkbuf_8 _5281_ (.A(_1791_),
    .X(_1792_));
 sky130_fd_sc_hd__or2_1 _5282_ (.A(_1771_),
    .B(_1775_),
    .X(_1793_));
 sky130_fd_sc_hd__buf_4 _5283_ (.A(_1793_),
    .X(_1794_));
 sky130_fd_sc_hd__or2_1 _5284_ (.A(_1782_),
    .B(_1771_),
    .X(_1795_));
 sky130_fd_sc_hd__clkbuf_4 _5285_ (.A(_1795_),
    .X(_1796_));
 sky130_fd_sc_hd__o22a_1 _5286_ (.A1(_1154_),
    .A2(_1794_),
    .B1(_1796_),
    .B2(_1042_),
    .X(_1797_));
 sky130_fd_sc_hd__o221a_1 _5287_ (.A1(_1146_),
    .A2(_1777_),
    .B1(_1792_),
    .B2(_1134_),
    .C1(_1797_),
    .X(_1798_));
 sky130_fd_sc_hd__or2_1 _5288_ (.A(_1773_),
    .B(_1775_),
    .X(_1799_));
 sky130_fd_sc_hd__buf_4 _5289_ (.A(_1799_),
    .X(_1800_));
 sky130_fd_sc_hd__o22a_1 _5290_ (.A1(_1151_),
    .A2(_1769_),
    .B1(_1800_),
    .B2(_0983_),
    .X(_1801_));
 sky130_fd_sc_hd__o2111a_1 _5291_ (.A1(_1012_),
    .A2(_1790_),
    .B1(_1798_),
    .C1(_1801_),
    .D1(_1778_),
    .X(_1802_));
 sky130_fd_sc_hd__o211ai_4 _5292_ (.A1(_1053_),
    .A2(_1781_),
    .B1(_1787_),
    .C1(_1802_),
    .Y(_1803_));
 sky130_fd_sc_hd__xor2_1 _5293_ (.A(\sound4.count[10] ),
    .B(_1803_),
    .X(_1804_));
 sky130_fd_sc_hd__o22a_1 _5294_ (.A1(_1180_),
    .A2(_1786_),
    .B1(_1790_),
    .B2(_1028_),
    .X(_1805_));
 sky130_fd_sc_hd__o22a_1 _5295_ (.A1(_1176_),
    .A2(_1769_),
    .B1(_1777_),
    .B2(_1174_),
    .X(_1806_));
 sky130_fd_sc_hd__o22a_1 _5296_ (.A1(_1129_),
    .A2(_1800_),
    .B1(_1792_),
    .B2(_1026_),
    .X(_1807_));
 sky130_fd_sc_hd__o221a_1 _5297_ (.A1(_1182_),
    .A2(_1794_),
    .B1(_1796_),
    .B2(_1175_),
    .C1(_1807_),
    .X(_1808_));
 sky130_fd_sc_hd__o211a_1 _5298_ (.A1(_0996_),
    .A2(_1784_),
    .B1(_1806_),
    .C1(_1808_),
    .X(_1809_));
 sky130_fd_sc_hd__o211ai_4 _5299_ (.A1(_0954_),
    .A2(_1781_),
    .B1(_1805_),
    .C1(_1809_),
    .Y(_1810_));
 sky130_fd_sc_hd__nand2_1 _5300_ (.A(\sound4.count[5] ),
    .B(_1810_),
    .Y(_1811_));
 sky130_fd_sc_hd__or2_1 _5301_ (.A(\sound4.count[5] ),
    .B(_1810_),
    .X(_1812_));
 sky130_fd_sc_hd__o22a_1 _5302_ (.A1(_1058_),
    .A2(_1771_),
    .B1(_1788_),
    .B2(_1111_),
    .X(_1813_));
 sky130_fd_sc_hd__a21o_1 _5303_ (.A1(_1769_),
    .A2(_1781_),
    .B1(_0687_),
    .X(_1814_));
 sky130_fd_sc_hd__o221a_1 _5304_ (.A1(_0680_),
    .A2(_1784_),
    .B1(_1792_),
    .B2(_0684_),
    .C1(_1800_),
    .X(_1815_));
 sky130_fd_sc_hd__a21o_1 _5305_ (.A1(_1814_),
    .A2(_1815_),
    .B1(_0695_),
    .X(_1816_));
 sky130_fd_sc_hd__o211a_2 _5306_ (.A1(_1062_),
    .A2(_1777_),
    .B1(_1813_),
    .C1(_1816_),
    .X(_1817_));
 sky130_fd_sc_hd__xnor2_1 _5307_ (.A(\sound4.count[14] ),
    .B(_1817_),
    .Y(_1818_));
 sky130_fd_sc_hd__a21o_1 _5308_ (.A1(_1773_),
    .A2(_1777_),
    .B1(_1055_),
    .X(_1819_));
 sky130_fd_sc_hd__o211a_1 _5309_ (.A1(_1010_),
    .A2(_1772_),
    .B1(_1778_),
    .C1(_1819_),
    .X(_1820_));
 sky130_fd_sc_hd__xnor2_1 _5310_ (.A(\sound4.count[16] ),
    .B(_1820_),
    .Y(_1821_));
 sky130_fd_sc_hd__a211o_1 _5311_ (.A1(_1811_),
    .A2(_1812_),
    .B1(_1818_),
    .C1(_1821_),
    .X(_1822_));
 sky130_fd_sc_hd__or3_1 _5312_ (.A(_1004_),
    .B(_1038_),
    .C(_1786_),
    .X(_1823_));
 sky130_fd_sc_hd__o221a_1 _5313_ (.A1(_1126_),
    .A2(_1781_),
    .B1(_1790_),
    .B2(_1165_),
    .C1(_1823_),
    .X(_1824_));
 sky130_fd_sc_hd__o22a_1 _5314_ (.A1(_0997_),
    .A2(_1777_),
    .B1(_1792_),
    .B2(_1159_),
    .X(_1825_));
 sky130_fd_sc_hd__o221a_1 _5315_ (.A1(_0685_),
    .A2(_1769_),
    .B1(_1794_),
    .B2(_1077_),
    .C1(_1825_),
    .X(_1826_));
 sky130_fd_sc_hd__o22a_1 _5316_ (.A1(_1166_),
    .A2(_1800_),
    .B1(_1796_),
    .B2(_0677_),
    .X(_1827_));
 sky130_fd_sc_hd__o211a_1 _5317_ (.A1(_1154_),
    .A2(_1784_),
    .B1(_1826_),
    .C1(_1827_),
    .X(_1828_));
 sky130_fd_sc_hd__and3_1 _5318_ (.A(_1778_),
    .B(_1824_),
    .C(_1828_),
    .X(_1829_));
 sky130_fd_sc_hd__and2_1 _5319_ (.A(\sound4.count[8] ),
    .B(_1829_),
    .X(_1830_));
 sky130_fd_sc_hd__nor2_1 _5320_ (.A(\sound4.count[8] ),
    .B(_1829_),
    .Y(_1831_));
 sky130_fd_sc_hd__nor2_1 _5321_ (.A(_1782_),
    .B(_1771_),
    .Y(_1832_));
 sky130_fd_sc_hd__nand2_1 _5322_ (.A(_0677_),
    .B(_1832_),
    .Y(_1833_));
 sky130_fd_sc_hd__or3_1 _5323_ (.A(net47),
    .B(_1129_),
    .C(_1770_),
    .X(_1834_));
 sky130_fd_sc_hd__o22a_1 _5324_ (.A1(_1004_),
    .A2(_1784_),
    .B1(_1786_),
    .B2(_1189_),
    .X(_1835_));
 sky130_fd_sc_hd__o22a_1 _5325_ (.A1(_1028_),
    .A2(_1800_),
    .B1(_1794_),
    .B2(_1083_),
    .X(_1836_));
 sky130_fd_sc_hd__or2_1 _5326_ (.A(_1158_),
    .B(_1790_),
    .X(_1837_));
 sky130_fd_sc_hd__o221a_1 _5327_ (.A1(_1020_),
    .A2(_1777_),
    .B1(_1792_),
    .B2(_1014_),
    .C1(_1837_),
    .X(_1838_));
 sky130_fd_sc_hd__o211a_1 _5328_ (.A1(_1077_),
    .A2(_1769_),
    .B1(_1836_),
    .C1(_1838_),
    .X(_1839_));
 sky130_fd_sc_hd__o2111a_1 _5329_ (.A1(_0959_),
    .A2(_1833_),
    .B1(_1834_),
    .C1(_1835_),
    .D1(_1839_),
    .X(_1840_));
 sky130_fd_sc_hd__xnor2_1 _5330_ (.A(\sound4.count[9] ),
    .B(_1840_),
    .Y(_1841_));
 sky130_fd_sc_hd__nor2_1 _5331_ (.A(_1771_),
    .B(_1775_),
    .Y(_1842_));
 sky130_fd_sc_hd__nor2_1 _5332_ (.A(_1200_),
    .B(_1792_),
    .Y(_1843_));
 sky130_fd_sc_hd__a31o_1 _5333_ (.A1(_1011_),
    .A2(_1015_),
    .A3(_1842_),
    .B1(_1843_),
    .X(_1844_));
 sky130_fd_sc_hd__o22ai_1 _5334_ (.A1(_0686_),
    .A2(_1784_),
    .B1(_1781_),
    .B2(_1146_),
    .Y(_1845_));
 sky130_fd_sc_hd__o22a_1 _5335_ (.A1(_1204_),
    .A2(_1786_),
    .B1(_1790_),
    .B2(_1014_),
    .X(_1846_));
 sky130_fd_sc_hd__o22a_1 _5336_ (.A1(_1198_),
    .A2(_1769_),
    .B1(_1777_),
    .B2(_1189_),
    .X(_1847_));
 sky130_fd_sc_hd__o211a_1 _5337_ (.A1(_1199_),
    .A2(_1800_),
    .B1(_1846_),
    .C1(_1847_),
    .X(_1848_));
 sky130_fd_sc_hd__o21ai_1 _5338_ (.A1(_1125_),
    .A2(_1796_),
    .B1(_1848_),
    .Y(_1849_));
 sky130_fd_sc_hd__or3_2 _5339_ (.A(_1844_),
    .B(_1845_),
    .C(_1849_),
    .X(_1850_));
 sky130_fd_sc_hd__xor2_1 _5340_ (.A(\sound4.count[3] ),
    .B(_1850_),
    .X(_1851_));
 sky130_fd_sc_hd__or4_1 _5341_ (.A(_1830_),
    .B(_1831_),
    .C(_1841_),
    .D(_1851_),
    .X(_1852_));
 sky130_fd_sc_hd__o22a_1 _5342_ (.A1(_1096_),
    .A2(_1786_),
    .B1(_1794_),
    .B2(_1097_),
    .X(_1853_));
 sky130_fd_sc_hd__nor2_1 _5343_ (.A(_1780_),
    .B(_1832_),
    .Y(_1854_));
 sky130_fd_sc_hd__o32a_1 _5344_ (.A1(_0977_),
    .A2(_0996_),
    .A3(_1784_),
    .B1(_1854_),
    .B2(_0960_),
    .X(_1855_));
 sky130_fd_sc_hd__or3_1 _5345_ (.A(_0993_),
    .B(_1012_),
    .C(_1790_),
    .X(_1856_));
 sky130_fd_sc_hd__o211a_1 _5346_ (.A1(_1095_),
    .A2(_1792_),
    .B1(_1855_),
    .C1(_1856_),
    .X(_1857_));
 sky130_fd_sc_hd__o211a_1 _5347_ (.A1(_0948_),
    .A2(_1800_),
    .B1(_1853_),
    .C1(_1857_),
    .X(_1858_));
 sky130_fd_sc_hd__o221ai_4 _5348_ (.A1(_1041_),
    .A2(_1769_),
    .B1(_1777_),
    .B2(_1101_),
    .C1(_1858_),
    .Y(_1859_));
 sky130_fd_sc_hd__xor2_1 _5349_ (.A(\sound4.count[0] ),
    .B(_1859_),
    .X(_1860_));
 sky130_fd_sc_hd__or4_1 _5350_ (.A(_1804_),
    .B(_1822_),
    .C(_1852_),
    .D(_1860_),
    .X(_1861_));
 sky130_fd_sc_hd__o221a_1 _5351_ (.A1(_1139_),
    .A2(_1786_),
    .B1(_1790_),
    .B2(_1134_),
    .C1(_1834_),
    .X(_1862_));
 sky130_fd_sc_hd__o221a_1 _5352_ (.A1(_1127_),
    .A2(_1777_),
    .B1(_1800_),
    .B2(_1126_),
    .C1(_1862_),
    .X(_1863_));
 sky130_fd_sc_hd__o221a_1 _5353_ (.A1(_1135_),
    .A2(_1784_),
    .B1(_1796_),
    .B2(_1141_),
    .C1(_1863_),
    .X(_1864_));
 sky130_fd_sc_hd__o211a_1 _5354_ (.A1(_1138_),
    .A2(_1769_),
    .B1(_1778_),
    .C1(_1864_),
    .X(_1865_));
 sky130_fd_sc_hd__o221ai_4 _5355_ (.A1(_0696_),
    .A2(_1792_),
    .B1(_1794_),
    .B2(_1140_),
    .C1(_1865_),
    .Y(_1866_));
 sky130_fd_sc_hd__nand2_1 _5356_ (.A(\sound4.count[4] ),
    .B(_1866_),
    .Y(_1867_));
 sky130_fd_sc_hd__or2_1 _5357_ (.A(\sound4.count[4] ),
    .B(_1866_),
    .X(_1868_));
 sky130_fd_sc_hd__o221a_1 _5358_ (.A1(_0683_),
    .A2(_1769_),
    .B1(_1794_),
    .B2(_0996_),
    .C1(_1800_),
    .X(_1869_));
 sky130_fd_sc_hd__or3_1 _5359_ (.A(_0687_),
    .B(_1001_),
    .C(_1790_),
    .X(_1870_));
 sky130_fd_sc_hd__o221a_1 _5360_ (.A1(_1016_),
    .A2(_1786_),
    .B1(_1781_),
    .B2(_1116_),
    .C1(_1870_),
    .X(_1871_));
 sky130_fd_sc_hd__o221a_1 _5361_ (.A1(_0997_),
    .A2(_1792_),
    .B1(_1796_),
    .B2(_1112_),
    .C1(_1871_),
    .X(_1872_));
 sky130_fd_sc_hd__o32a_1 _5362_ (.A1(_0677_),
    .A2(_1083_),
    .A3(_1784_),
    .B1(_1777_),
    .B2(_1064_),
    .X(_1873_));
 sky130_fd_sc_hd__o211a_1 _5363_ (.A1(_1107_),
    .A2(_1869_),
    .B1(_1872_),
    .C1(_1873_),
    .X(_1874_));
 sky130_fd_sc_hd__nand2_2 _5364_ (.A(_1778_),
    .B(_1874_),
    .Y(_1875_));
 sky130_fd_sc_hd__nand2_1 _5365_ (.A(\sound4.count[13] ),
    .B(_1875_),
    .Y(_1876_));
 sky130_fd_sc_hd__or2_1 _5366_ (.A(\sound4.count[13] ),
    .B(_1875_),
    .X(_1877_));
 sky130_fd_sc_hd__o32a_1 _5367_ (.A1(_0959_),
    .A2(_1133_),
    .A3(_1786_),
    .B1(_1790_),
    .B2(_0983_),
    .X(_1878_));
 sky130_fd_sc_hd__o32a_1 _5368_ (.A1(_0677_),
    .A2(_1038_),
    .A3(_1796_),
    .B1(_1769_),
    .B2(_1059_),
    .X(_1879_));
 sky130_fd_sc_hd__o211a_1 _5369_ (.A1(_1064_),
    .A2(_1781_),
    .B1(_1878_),
    .C1(_1879_),
    .X(_1880_));
 sky130_fd_sc_hd__o22a_1 _5370_ (.A1(_1056_),
    .A2(_1777_),
    .B1(_1800_),
    .B2(_1053_),
    .X(_1881_));
 sky130_fd_sc_hd__o221a_1 _5371_ (.A1(_1057_),
    .A2(_1792_),
    .B1(_1794_),
    .B2(_1063_),
    .C1(_1881_),
    .X(_1882_));
 sky130_fd_sc_hd__o311a_1 _5372_ (.A1(_0679_),
    .A2(net63),
    .A3(_1784_),
    .B1(_1882_),
    .C1(_1778_),
    .X(_1883_));
 sky130_fd_sc_hd__nand2_1 _5373_ (.A(_1880_),
    .B(_1883_),
    .Y(_1884_));
 sky130_fd_sc_hd__xor2_1 _5374_ (.A(\sound4.count[6] ),
    .B(_1884_),
    .X(_1885_));
 sky130_fd_sc_hd__a221o_1 _5375_ (.A1(_1867_),
    .A2(_1868_),
    .B1(_1876_),
    .B2(_1877_),
    .C1(_1885_),
    .X(_1886_));
 sky130_fd_sc_hd__a21o_1 _5376_ (.A1(_1777_),
    .A2(_1788_),
    .B1(_1213_),
    .X(_1887_));
 sky130_fd_sc_hd__nor2_1 _5377_ (.A(_0869_),
    .B(_1765_),
    .Y(_1888_));
 sky130_fd_sc_hd__o22a_1 _5378_ (.A1(_0688_),
    .A2(_1771_),
    .B1(_1773_),
    .B2(_1138_),
    .X(_1889_));
 sky130_fd_sc_hd__o2bb2a_1 _5379_ (.A1_N(_1775_),
    .A2_N(_1888_),
    .B1(_1889_),
    .B2(_1774_),
    .X(_1890_));
 sky130_fd_sc_hd__and3_2 _5380_ (.A(_1778_),
    .B(_1887_),
    .C(_1890_),
    .X(_1891_));
 sky130_fd_sc_hd__o22a_1 _5381_ (.A1(_0946_),
    .A2(_1786_),
    .B1(_1790_),
    .B2(_0971_),
    .X(_1892_));
 sky130_fd_sc_hd__o32a_1 _5382_ (.A1(_0684_),
    .A2(_1077_),
    .A3(_1792_),
    .B1(_1781_),
    .B2(_1039_),
    .X(_1893_));
 sky130_fd_sc_hd__o22a_1 _5383_ (.A1(_1079_),
    .A2(_1800_),
    .B1(_1794_),
    .B2(_0952_),
    .X(_1894_));
 sky130_fd_sc_hd__o221a_1 _5384_ (.A1(_1015_),
    .A2(_1769_),
    .B1(_1784_),
    .B2(_1083_),
    .C1(_1833_),
    .X(_1895_));
 sky130_fd_sc_hd__o211a_1 _5385_ (.A1(_0960_),
    .A2(_1777_),
    .B1(_1894_),
    .C1(_1895_),
    .X(_1896_));
 sky130_fd_sc_hd__and3_2 _5386_ (.A(_1892_),
    .B(_1893_),
    .C(_1896_),
    .X(_1897_));
 sky130_fd_sc_hd__or3_1 _5387_ (.A(_1024_),
    .B(_1028_),
    .C(_1786_),
    .X(_1898_));
 sky130_fd_sc_hd__o221a_1 _5388_ (.A1(_1025_),
    .A2(_1794_),
    .B1(_1796_),
    .B2(_1027_),
    .C1(_1898_),
    .X(_1899_));
 sky130_fd_sc_hd__o221a_1 _5389_ (.A1(_1017_),
    .A2(_1784_),
    .B1(_1781_),
    .B2(_1020_),
    .C1(_1899_),
    .X(_1900_));
 sky130_fd_sc_hd__o22a_1 _5390_ (.A1(_0973_),
    .A2(_1777_),
    .B1(_1800_),
    .B2(_1016_),
    .X(_1901_));
 sky130_fd_sc_hd__o221a_1 _5391_ (.A1(_0997_),
    .A2(_1769_),
    .B1(_1792_),
    .B2(_1010_),
    .C1(_1901_),
    .X(_1902_));
 sky130_fd_sc_hd__o211a_1 _5392_ (.A1(_0993_),
    .A2(_1837_),
    .B1(_1900_),
    .C1(_1902_),
    .X(_1903_));
 sky130_fd_sc_hd__a21oi_1 _5393_ (.A1(_0869_),
    .A2(_1832_),
    .B1(_1842_),
    .Y(_1904_));
 sky130_fd_sc_hd__o32a_1 _5394_ (.A1(_1001_),
    .A2(_0996_),
    .A3(_1784_),
    .B1(_1904_),
    .B2(_1004_),
    .X(_1905_));
 sky130_fd_sc_hd__a211o_1 _5395_ (.A1(net47),
    .A2(net63),
    .B1(_1788_),
    .C1(_0947_),
    .X(_1906_));
 sky130_fd_sc_hd__o2bb2a_1 _5396_ (.A1_N(_1125_),
    .A2_N(_1780_),
    .B1(_1800_),
    .B2(_1033_),
    .X(_1907_));
 sky130_fd_sc_hd__o2111a_1 _5397_ (.A1(_1129_),
    .A2(_1777_),
    .B1(_1905_),
    .C1(_1906_),
    .D1(_1907_),
    .X(_1908_));
 sky130_fd_sc_hd__o221a_2 _5398_ (.A1(_1035_),
    .A2(_1769_),
    .B1(_1792_),
    .B2(_1041_),
    .C1(_1908_),
    .X(_1909_));
 sky130_fd_sc_hd__a2bb2o_1 _5399_ (.A1_N(\sound4.count[2] ),
    .A2_N(_1903_),
    .B1(_1909_),
    .B2(\sound4.count[11] ),
    .X(_1910_));
 sky130_fd_sc_hd__a221o_1 _5400_ (.A1(\sound4.count[15] ),
    .A2(_1891_),
    .B1(_1897_),
    .B2(\sound4.count[7] ),
    .C1(_1910_),
    .X(_1911_));
 sky130_fd_sc_hd__a2bb2o_1 _5401_ (.A1_N(\sound4.count[7] ),
    .A2_N(_1897_),
    .B1(_1903_),
    .B2(\sound4.count[2] ),
    .X(_1912_));
 sky130_fd_sc_hd__and3_1 _5402_ (.A(_1772_),
    .B(_1773_),
    .C(_1777_),
    .X(_1913_));
 sky130_fd_sc_hd__o21a_1 _5403_ (.A1(_1222_),
    .A2(_1913_),
    .B1(\sound4.count[17] ),
    .X(_1914_));
 sky130_fd_sc_hd__nand2_1 _5404_ (.A(\sound4.count[18] ),
    .B(_1778_),
    .Y(_1915_));
 sky130_fd_sc_hd__or2_1 _5405_ (.A(\sound4.count[18] ),
    .B(_1778_),
    .X(_1916_));
 sky130_fd_sc_hd__o311a_1 _5406_ (.A1(\sound4.count[17] ),
    .A2(_1222_),
    .A3(_1913_),
    .B1(_1915_),
    .C1(_1916_),
    .X(_1917_));
 sky130_fd_sc_hd__or3b_1 _5407_ (.A(_1912_),
    .B(_1914_),
    .C_N(_1917_),
    .X(_1918_));
 sky130_fd_sc_hd__o22ai_1 _5408_ (.A1(_0954_),
    .A2(_1777_),
    .B1(_1792_),
    .B2(_0985_),
    .Y(_1919_));
 sky130_fd_sc_hd__o221a_1 _5409_ (.A1(net63),
    .A2(_1784_),
    .B1(_1781_),
    .B2(_1038_),
    .C1(_1769_),
    .X(_1920_));
 sky130_fd_sc_hd__o22a_1 _5410_ (.A1(_1101_),
    .A2(_1786_),
    .B1(_1790_),
    .B2(_1240_),
    .X(_1921_));
 sky130_fd_sc_hd__o221a_1 _5411_ (.A1(_1245_),
    .A2(_1800_),
    .B1(_1796_),
    .B2(_1110_),
    .C1(_1921_),
    .X(_1922_));
 sky130_fd_sc_hd__o21ai_1 _5412_ (.A1(_1025_),
    .A2(_1920_),
    .B1(_1922_),
    .Y(_1923_));
 sky130_fd_sc_hd__a211o_2 _5413_ (.A1(_1079_),
    .A2(_1842_),
    .B1(_1919_),
    .C1(_1923_),
    .X(_1924_));
 sky130_fd_sc_hd__xor2_1 _5414_ (.A(\sound4.count[12] ),
    .B(_1924_),
    .X(_1925_));
 sky130_fd_sc_hd__o22a_1 _5415_ (.A1(_0954_),
    .A2(_1784_),
    .B1(_1790_),
    .B2(_0948_),
    .X(_1926_));
 sky130_fd_sc_hd__o32a_1 _5416_ (.A1(_0978_),
    .A2(_0944_),
    .A3(_1777_),
    .B1(_1794_),
    .B2(_1001_),
    .X(_1927_));
 sky130_fd_sc_hd__o221a_1 _5417_ (.A1(_0985_),
    .A2(_1769_),
    .B1(_1796_),
    .B2(_0979_),
    .C1(_1927_),
    .X(_1928_));
 sky130_fd_sc_hd__o32a_1 _5418_ (.A1(_0959_),
    .A2(_0993_),
    .A3(_1800_),
    .B1(_1792_),
    .B2(_0869_),
    .X(_1929_));
 sky130_fd_sc_hd__o211a_1 _5419_ (.A1(_0973_),
    .A2(_1786_),
    .B1(_1928_),
    .C1(_1929_),
    .X(_1930_));
 sky130_fd_sc_hd__o211a_2 _5420_ (.A1(_0997_),
    .A2(_1781_),
    .B1(_1926_),
    .C1(_1930_),
    .X(_1931_));
 sky130_fd_sc_hd__o2bb2a_1 _5421_ (.A1_N(\sound4.count[1] ),
    .A2_N(_1931_),
    .B1(_1891_),
    .B2(\sound4.count[15] ),
    .X(_1932_));
 sky130_fd_sc_hd__o221a_1 _5422_ (.A1(\sound4.count[1] ),
    .A2(_1931_),
    .B1(_1909_),
    .B2(\sound4.count[11] ),
    .C1(_1932_),
    .X(_1933_));
 sky130_fd_sc_hd__or4b_1 _5423_ (.A(_1911_),
    .B(_1918_),
    .C(_1925_),
    .D_N(_1933_),
    .X(_1934_));
 sky130_fd_sc_hd__or3_1 _5424_ (.A(_1861_),
    .B(_1886_),
    .C(_1934_),
    .X(_1935_));
 sky130_fd_sc_hd__buf_4 _5425_ (.A(_1935_),
    .X(_1936_));
 sky130_fd_sc_hd__nand3_1 _5426_ (.A(\sound4.count[0] ),
    .B(_1779_),
    .C(_1936_),
    .Y(\sound4.osc.next_count[0] ));
 sky130_fd_sc_hd__nand2_1 _5427_ (.A(\sound4.count[0] ),
    .B(\sound4.count[1] ),
    .Y(_1937_));
 sky130_fd_sc_hd__or2_1 _5428_ (.A(\sound4.count[0] ),
    .B(\sound4.count[1] ),
    .X(_1938_));
 sky130_fd_sc_hd__and4_1 _5429_ (.A(_1779_),
    .B(_1936_),
    .C(_1937_),
    .D(_1938_),
    .X(_1939_));
 sky130_fd_sc_hd__clkbuf_1 _5430_ (.A(_1939_),
    .X(\sound4.osc.next_count[1] ));
 sky130_fd_sc_hd__and3_1 _5431_ (.A(\sound4.count[0] ),
    .B(\sound4.count[1] ),
    .C(\sound4.count[2] ),
    .X(_1940_));
 sky130_fd_sc_hd__inv_2 _5432_ (.A(_1940_),
    .Y(_1941_));
 sky130_fd_sc_hd__a21o_1 _5433_ (.A1(\sound4.count[0] ),
    .A2(\sound4.count[1] ),
    .B1(\sound4.count[2] ),
    .X(_1942_));
 sky130_fd_sc_hd__and4_1 _5434_ (.A(_1779_),
    .B(_1936_),
    .C(_1941_),
    .D(_1942_),
    .X(_1943_));
 sky130_fd_sc_hd__clkbuf_1 _5435_ (.A(_1943_),
    .X(\sound4.osc.next_count[2] ));
 sky130_fd_sc_hd__and2_1 _5436_ (.A(\sound4.count[3] ),
    .B(_1940_),
    .X(_1944_));
 sky130_fd_sc_hd__inv_2 _5437_ (.A(_1944_),
    .Y(_1945_));
 sky130_fd_sc_hd__or2_1 _5438_ (.A(\sound4.count[3] ),
    .B(_1940_),
    .X(_1946_));
 sky130_fd_sc_hd__and4_1 _5439_ (.A(_1779_),
    .B(_1936_),
    .C(_1945_),
    .D(_1946_),
    .X(_1947_));
 sky130_fd_sc_hd__clkbuf_1 _5440_ (.A(_1947_),
    .X(\sound4.osc.next_count[3] ));
 sky130_fd_sc_hd__nand2_1 _5441_ (.A(\sound4.count[4] ),
    .B(_1944_),
    .Y(_1948_));
 sky130_fd_sc_hd__or2_1 _5442_ (.A(\sound4.count[4] ),
    .B(_1944_),
    .X(_1949_));
 sky130_fd_sc_hd__and4_1 _5443_ (.A(_1779_),
    .B(_1936_),
    .C(_1948_),
    .D(_1949_),
    .X(_1950_));
 sky130_fd_sc_hd__clkbuf_1 _5444_ (.A(_1950_),
    .X(\sound4.osc.next_count[4] ));
 sky130_fd_sc_hd__and3_1 _5445_ (.A(\sound4.count[4] ),
    .B(\sound4.count[5] ),
    .C(_1944_),
    .X(_1951_));
 sky130_fd_sc_hd__inv_2 _5446_ (.A(_1951_),
    .Y(_1952_));
 sky130_fd_sc_hd__a31o_1 _5447_ (.A1(\sound4.count[3] ),
    .A2(\sound4.count[4] ),
    .A3(_1940_),
    .B1(\sound4.count[5] ),
    .X(_1953_));
 sky130_fd_sc_hd__and4_1 _5448_ (.A(_1779_),
    .B(_1936_),
    .C(_1952_),
    .D(_1953_),
    .X(_1954_));
 sky130_fd_sc_hd__clkbuf_1 _5449_ (.A(_1954_),
    .X(\sound4.osc.next_count[5] ));
 sky130_fd_sc_hd__and2_1 _5450_ (.A(\sound4.count[6] ),
    .B(_1951_),
    .X(_1955_));
 sky130_fd_sc_hd__inv_2 _5451_ (.A(_1955_),
    .Y(_1956_));
 sky130_fd_sc_hd__or2_1 _5452_ (.A(\sound4.count[6] ),
    .B(_1951_),
    .X(_1957_));
 sky130_fd_sc_hd__and4_1 _5453_ (.A(_1779_),
    .B(_1936_),
    .C(_1956_),
    .D(_1957_),
    .X(_1958_));
 sky130_fd_sc_hd__clkbuf_1 _5454_ (.A(_1958_),
    .X(\sound4.osc.next_count[6] ));
 sky130_fd_sc_hd__nand2_1 _5455_ (.A(\sound4.count[7] ),
    .B(_1955_),
    .Y(_1959_));
 sky130_fd_sc_hd__or2_1 _5456_ (.A(\sound4.count[7] ),
    .B(_1955_),
    .X(_1960_));
 sky130_fd_sc_hd__and4_1 _5457_ (.A(_1779_),
    .B(_1936_),
    .C(_1959_),
    .D(_1960_),
    .X(_1961_));
 sky130_fd_sc_hd__clkbuf_1 _5458_ (.A(_1961_),
    .X(\sound4.osc.next_count[7] ));
 sky130_fd_sc_hd__and3_1 _5459_ (.A(\sound4.count[7] ),
    .B(\sound4.count[8] ),
    .C(_1955_),
    .X(_1962_));
 sky130_fd_sc_hd__inv_2 _5460_ (.A(_1962_),
    .Y(_1963_));
 sky130_fd_sc_hd__a31o_1 _5461_ (.A1(\sound4.count[6] ),
    .A2(\sound4.count[7] ),
    .A3(_1951_),
    .B1(\sound4.count[8] ),
    .X(_1964_));
 sky130_fd_sc_hd__and4_1 _5462_ (.A(_1779_),
    .B(_1936_),
    .C(_1963_),
    .D(_1964_),
    .X(_1965_));
 sky130_fd_sc_hd__clkbuf_1 _5463_ (.A(_1965_),
    .X(\sound4.osc.next_count[8] ));
 sky130_fd_sc_hd__and2_1 _5464_ (.A(\sound4.count[9] ),
    .B(_1962_),
    .X(_1966_));
 sky130_fd_sc_hd__inv_2 _5465_ (.A(_1966_),
    .Y(_1967_));
 sky130_fd_sc_hd__or2_1 _5466_ (.A(\sound4.count[9] ),
    .B(_1962_),
    .X(_1968_));
 sky130_fd_sc_hd__and4_1 _5467_ (.A(_1779_),
    .B(_1936_),
    .C(_1967_),
    .D(_1968_),
    .X(_1969_));
 sky130_fd_sc_hd__clkbuf_1 _5468_ (.A(_1969_),
    .X(\sound4.osc.next_count[9] ));
 sky130_fd_sc_hd__nand2_1 _5469_ (.A(\sound4.count[10] ),
    .B(_1966_),
    .Y(_1970_));
 sky130_fd_sc_hd__or2_1 _5470_ (.A(\sound4.count[10] ),
    .B(_1966_),
    .X(_1971_));
 sky130_fd_sc_hd__and4_1 _5471_ (.A(_1779_),
    .B(_1936_),
    .C(_1970_),
    .D(_1971_),
    .X(_1972_));
 sky130_fd_sc_hd__clkbuf_1 _5472_ (.A(_1972_),
    .X(\sound4.osc.next_count[10] ));
 sky130_fd_sc_hd__and3_1 _5473_ (.A(\sound4.count[10] ),
    .B(\sound4.count[11] ),
    .C(_1966_),
    .X(_1973_));
 sky130_fd_sc_hd__inv_2 _5474_ (.A(_1973_),
    .Y(_1974_));
 sky130_fd_sc_hd__a31o_1 _5475_ (.A1(\sound4.count[9] ),
    .A2(\sound4.count[10] ),
    .A3(_1962_),
    .B1(\sound4.count[11] ),
    .X(_1975_));
 sky130_fd_sc_hd__and4_1 _5476_ (.A(_1779_),
    .B(_1936_),
    .C(_1974_),
    .D(_1975_),
    .X(_1976_));
 sky130_fd_sc_hd__clkbuf_1 _5477_ (.A(_1976_),
    .X(\sound4.osc.next_count[11] ));
 sky130_fd_sc_hd__and2_1 _5478_ (.A(\sound4.count[12] ),
    .B(_1973_),
    .X(_1977_));
 sky130_fd_sc_hd__inv_2 _5479_ (.A(_1977_),
    .Y(_1978_));
 sky130_fd_sc_hd__or2_1 _5480_ (.A(\sound4.count[12] ),
    .B(_1973_),
    .X(_1979_));
 sky130_fd_sc_hd__and4_1 _5481_ (.A(_1779_),
    .B(_1936_),
    .C(_1978_),
    .D(_1979_),
    .X(_1980_));
 sky130_fd_sc_hd__clkbuf_1 _5482_ (.A(_1980_),
    .X(\sound4.osc.next_count[12] ));
 sky130_fd_sc_hd__nand2_1 _5483_ (.A(\sound4.count[13] ),
    .B(_1977_),
    .Y(_1981_));
 sky130_fd_sc_hd__or2_1 _5484_ (.A(\sound4.count[13] ),
    .B(_1977_),
    .X(_1982_));
 sky130_fd_sc_hd__and4_1 _5485_ (.A(_1779_),
    .B(_1936_),
    .C(_1981_),
    .D(_1982_),
    .X(_1983_));
 sky130_fd_sc_hd__clkbuf_1 _5486_ (.A(_1983_),
    .X(\sound4.osc.next_count[13] ));
 sky130_fd_sc_hd__and3_2 _5487_ (.A(\sound4.count[13] ),
    .B(\sound4.count[14] ),
    .C(_1977_),
    .X(_1984_));
 sky130_fd_sc_hd__inv_2 _5488_ (.A(_1984_),
    .Y(_1985_));
 sky130_fd_sc_hd__a31o_1 _5489_ (.A1(\sound4.count[12] ),
    .A2(\sound4.count[13] ),
    .A3(_1973_),
    .B1(\sound4.count[14] ),
    .X(_1986_));
 sky130_fd_sc_hd__and4_1 _5490_ (.A(_1779_),
    .B(_1936_),
    .C(_1985_),
    .D(_1986_),
    .X(_1987_));
 sky130_fd_sc_hd__clkbuf_1 _5491_ (.A(_1987_),
    .X(\sound4.osc.next_count[14] ));
 sky130_fd_sc_hd__and2_2 _5492_ (.A(\sound4.count[15] ),
    .B(_1984_),
    .X(_1988_));
 sky130_fd_sc_hd__inv_2 _5493_ (.A(_1988_),
    .Y(_1989_));
 sky130_fd_sc_hd__or2_1 _5494_ (.A(\sound4.count[15] ),
    .B(_1984_),
    .X(_1990_));
 sky130_fd_sc_hd__and4_1 _5495_ (.A(_1779_),
    .B(_1936_),
    .C(_1989_),
    .D(_1990_),
    .X(_1991_));
 sky130_fd_sc_hd__clkbuf_1 _5496_ (.A(_1991_),
    .X(\sound4.osc.next_count[15] ));
 sky130_fd_sc_hd__nand2_1 _5497_ (.A(\sound4.count[16] ),
    .B(_1988_),
    .Y(_1992_));
 sky130_fd_sc_hd__or2_1 _5498_ (.A(\sound4.count[16] ),
    .B(_1988_),
    .X(_1993_));
 sky130_fd_sc_hd__and4_1 _5499_ (.A(_1779_),
    .B(_1936_),
    .C(_1992_),
    .D(_1993_),
    .X(_1994_));
 sky130_fd_sc_hd__clkbuf_1 _5500_ (.A(_1994_),
    .X(\sound4.osc.next_count[16] ));
 sky130_fd_sc_hd__nand3_1 _5501_ (.A(\sound4.count[16] ),
    .B(\sound4.count[17] ),
    .C(_1988_),
    .Y(_1995_));
 sky130_fd_sc_hd__a31o_1 _5502_ (.A1(\sound4.count[15] ),
    .A2(\sound4.count[16] ),
    .A3(_1984_),
    .B1(\sound4.count[17] ),
    .X(_1996_));
 sky130_fd_sc_hd__and4_1 _5503_ (.A(_1779_),
    .B(_1936_),
    .C(_1995_),
    .D(_1996_),
    .X(_1997_));
 sky130_fd_sc_hd__clkbuf_1 _5504_ (.A(_1997_),
    .X(\sound4.osc.next_count[17] ));
 sky130_fd_sc_hd__a31o_1 _5505_ (.A1(\sound4.count[16] ),
    .A2(\sound4.count[17] ),
    .A3(_1988_),
    .B1(\sound4.count[18] ),
    .X(_1998_));
 sky130_fd_sc_hd__nand4_1 _5506_ (.A(\sound4.count[16] ),
    .B(\sound4.count[17] ),
    .C(\sound4.count[18] ),
    .D(_1988_),
    .Y(_1999_));
 sky130_fd_sc_hd__and3_1 _5507_ (.A(_1779_),
    .B(_1998_),
    .C(_1999_),
    .X(_2000_));
 sky130_fd_sc_hd__clkbuf_1 _5508_ (.A(_2000_),
    .X(\sound4.osc.next_count[18] ));
 sky130_fd_sc_hd__inv_2 _5509_ (.A(\rate_clk.count[0] ),
    .Y(\rate_clk.next_count[0] ));
 sky130_fd_sc_hd__xor2_1 _5510_ (.A(\rate_clk.count[1] ),
    .B(\rate_clk.count[0] ),
    .X(\rate_clk.next_count[1] ));
 sky130_fd_sc_hd__a21oi_1 _5511_ (.A1(\rate_clk.count[1] ),
    .A2(\rate_clk.count[0] ),
    .B1(\rate_clk.count[2] ),
    .Y(_2001_));
 sky130_fd_sc_hd__nor2_1 _5512_ (.A(_0550_),
    .B(_2001_),
    .Y(\rate_clk.next_count[2] ));
 sky130_fd_sc_hd__nor2_1 _5513_ (.A(\rate_clk.count[3] ),
    .B(_0550_),
    .Y(_2002_));
 sky130_fd_sc_hd__nor2_1 _5514_ (.A(_0551_),
    .B(_2002_),
    .Y(\rate_clk.next_count[3] ));
 sky130_fd_sc_hd__xor2_1 _5515_ (.A(\rate_clk.count[4] ),
    .B(_0551_),
    .X(\rate_clk.next_count[4] ));
 sky130_fd_sc_hd__a21oi_1 _5516_ (.A1(\rate_clk.count[4] ),
    .A2(_0551_),
    .B1(\rate_clk.count[5] ),
    .Y(_2003_));
 sky130_fd_sc_hd__nor2_1 _5517_ (.A(_0552_),
    .B(_2003_),
    .Y(\rate_clk.next_count[5] ));
 sky130_fd_sc_hd__nor2_1 _5518_ (.A(\rate_clk.count[6] ),
    .B(_0552_),
    .Y(_2004_));
 sky130_fd_sc_hd__nor2_1 _5519_ (.A(_0553_),
    .B(_2004_),
    .Y(\rate_clk.next_count[6] ));
 sky130_fd_sc_hd__clkbuf_16 _5520_ (.A(_0575_),
    .X(_2005_));
 sky130_fd_sc_hd__nor2_1 _5521_ (.A(\rate_clk.count[7] ),
    .B(_0553_),
    .Y(_2006_));
 sky130_fd_sc_hd__nor2_1 _5522_ (.A(_2005_),
    .B(_2006_),
    .Y(\rate_clk.next_count[7] ));
 sky130_fd_sc_hd__inv_2 _5523_ (.A(\pm.count[6] ),
    .Y(_2007_));
 sky130_fd_sc_hd__and2_1 _5524_ (.A(_2007_),
    .B(\pm.current_waveform[6] ),
    .X(_2008_));
 sky130_fd_sc_hd__inv_2 _5525_ (.A(\pm.count[5] ),
    .Y(_2009_));
 sky130_fd_sc_hd__and2_1 _5526_ (.A(_2009_),
    .B(\pm.current_waveform[5] ),
    .X(_2010_));
 sky130_fd_sc_hd__and2_1 _5527_ (.A(_0651_),
    .B(\pm.current_waveform[4] ),
    .X(_2011_));
 sky130_fd_sc_hd__inv_2 _5528_ (.A(\pm.count[3] ),
    .Y(_2012_));
 sky130_fd_sc_hd__and2_1 _5529_ (.A(_2012_),
    .B(\pm.current_waveform[3] ),
    .X(_2013_));
 sky130_fd_sc_hd__inv_2 _5530_ (.A(\pm.count[2] ),
    .Y(_2014_));
 sky130_fd_sc_hd__inv_2 _5531_ (.A(\pm.count[1] ),
    .Y(_2015_));
 sky130_fd_sc_hd__or2_1 _5532_ (.A(_2015_),
    .B(\pm.current_waveform[1] ),
    .X(_2016_));
 sky130_fd_sc_hd__a22o_1 _5533_ (.A1(_2014_),
    .A2(\pm.current_waveform[2] ),
    .B1(\pm.current_waveform[1] ),
    .B2(_2015_),
    .X(_2017_));
 sky130_fd_sc_hd__a31o_1 _5534_ (.A1(\pm.next_count[0] ),
    .A2(\pm.current_waveform[0] ),
    .A3(_2016_),
    .B1(_2017_),
    .X(_2018_));
 sky130_fd_sc_hd__o221a_1 _5535_ (.A1(_2012_),
    .A2(\pm.current_waveform[3] ),
    .B1(\pm.current_waveform[2] ),
    .B2(_2014_),
    .C1(_2018_),
    .X(_2019_));
 sky130_fd_sc_hd__o22a_1 _5536_ (.A1(_0651_),
    .A2(\pm.current_waveform[4] ),
    .B1(_2013_),
    .B2(_2019_),
    .X(_2020_));
 sky130_fd_sc_hd__o22a_1 _5537_ (.A1(_2009_),
    .A2(\pm.current_waveform[5] ),
    .B1(_2011_),
    .B2(_2020_),
    .X(_2021_));
 sky130_fd_sc_hd__o22a_1 _5538_ (.A1(_2007_),
    .A2(\pm.current_waveform[6] ),
    .B1(_2010_),
    .B2(_2021_),
    .X(_2022_));
 sky130_fd_sc_hd__o22a_1 _5539_ (.A1(_0657_),
    .A2(\pm.current_waveform[7] ),
    .B1(_2008_),
    .B2(_2022_),
    .X(_2023_));
 sky130_fd_sc_hd__a21o_1 _5540_ (.A1(_0657_),
    .A2(\pm.current_waveform[7] ),
    .B1(_2023_),
    .X(_2024_));
 sky130_fd_sc_hd__a21bo_1 _5541_ (.A1(\pm.current_waveform[8] ),
    .A2(_2024_),
    .B1_N(\pm.count[8] ),
    .X(_2025_));
 sky130_fd_sc_hd__o21a_1 _5542_ (.A1(\pm.current_waveform[8] ),
    .A2(_2024_),
    .B1(_2025_),
    .X(\pm.next_pwm_o ));
 sky130_fd_sc_hd__or4_1 _5543_ (.A(\sound4.divisor_m[3] ),
    .B(\sound4.divisor_m[2] ),
    .C(\sound4.divisor_m[1] ),
    .D(\sound4.divisor_m[0] ),
    .X(_2026_));
 sky130_fd_sc_hd__or3_1 _5544_ (.A(\sound4.divisor_m[5] ),
    .B(\sound4.divisor_m[4] ),
    .C(_2026_),
    .X(_2027_));
 sky130_fd_sc_hd__or2_1 _5545_ (.A(\sound4.divisor_m[6] ),
    .B(_2027_),
    .X(_2028_));
 sky130_fd_sc_hd__or3_1 _5546_ (.A(\sound4.divisor_m[8] ),
    .B(\sound4.divisor_m[7] ),
    .C(_2028_),
    .X(_2029_));
 sky130_fd_sc_hd__or2_1 _5547_ (.A(\sound4.divisor_m[9] ),
    .B(_2029_),
    .X(_2030_));
 sky130_fd_sc_hd__or3_1 _5548_ (.A(\sound4.divisor_m[11] ),
    .B(\sound4.divisor_m[10] ),
    .C(_2030_),
    .X(_2031_));
 sky130_fd_sc_hd__or2_1 _5549_ (.A(\sound4.divisor_m[12] ),
    .B(_2031_),
    .X(_2032_));
 sky130_fd_sc_hd__or4_1 _5550_ (.A(\sound4.divisor_m[15] ),
    .B(\sound4.divisor_m[14] ),
    .C(\sound4.divisor_m[13] ),
    .D(_2032_),
    .X(_2033_));
 sky130_fd_sc_hd__or2_1 _5551_ (.A(\sound4.divisor_m[16] ),
    .B(_2033_),
    .X(_2034_));
 sky130_fd_sc_hd__or2_1 _5552_ (.A(\sound4.divisor_m[17] ),
    .B(_2034_),
    .X(_2035_));
 sky130_fd_sc_hd__clkinv_4 _5553_ (.A(\sound4.sdiv.A[26] ),
    .Y(_2036_));
 sky130_fd_sc_hd__o21a_1 _5554_ (.A1(\sound4.divisor_m[18] ),
    .A2(_2035_),
    .B1(_2036_),
    .X(_2037_));
 sky130_fd_sc_hd__clkbuf_8 _5555_ (.A(_2037_),
    .X(_2038_));
 sky130_fd_sc_hd__nand2_1 _5556_ (.A(\sound4.sdiv.A[25] ),
    .B(_2038_),
    .Y(_2039_));
 sky130_fd_sc_hd__xnor2_1 _5557_ (.A(\sound4.sdiv.A[20] ),
    .B(_2038_),
    .Y(_2040_));
 sky130_fd_sc_hd__xnor2_1 _5558_ (.A(\sound4.sdiv.A[19] ),
    .B(_2038_),
    .Y(_2041_));
 sky130_fd_sc_hd__or2_1 _5559_ (.A(_2040_),
    .B(_2041_),
    .X(_2042_));
 sky130_fd_sc_hd__xor2_2 _5560_ (.A(\sound4.sdiv.A[22] ),
    .B(_2038_),
    .X(_2043_));
 sky130_fd_sc_hd__inv_2 _5561_ (.A(_2043_),
    .Y(_2044_));
 sky130_fd_sc_hd__xnor2_1 _5562_ (.A(\sound4.sdiv.A[21] ),
    .B(_2038_),
    .Y(_2045_));
 sky130_fd_sc_hd__inv_2 _5563_ (.A(\sound4.sdiv.A[16] ),
    .Y(_2046_));
 sky130_fd_sc_hd__nand2_1 _5564_ (.A(_2036_),
    .B(_2034_),
    .Y(_2047_));
 sky130_fd_sc_hd__xor2_1 _5565_ (.A(\sound4.divisor_m[17] ),
    .B(_2047_),
    .X(_2048_));
 sky130_fd_sc_hd__nand2_1 _5566_ (.A(_2046_),
    .B(_2048_),
    .Y(_2049_));
 sky130_fd_sc_hd__inv_2 _5567_ (.A(\sound4.sdiv.A[15] ),
    .Y(_2050_));
 sky130_fd_sc_hd__and2_1 _5568_ (.A(_2036_),
    .B(_2033_),
    .X(_2051_));
 sky130_fd_sc_hd__xnor2_1 _5569_ (.A(\sound4.divisor_m[16] ),
    .B(_2051_),
    .Y(_2052_));
 sky130_fd_sc_hd__nor2_1 _5570_ (.A(_2050_),
    .B(_2052_),
    .Y(_2053_));
 sky130_fd_sc_hd__nor2_1 _5571_ (.A(\sound4.divisor_m[13] ),
    .B(_2032_),
    .Y(_2054_));
 sky130_fd_sc_hd__nor2_1 _5572_ (.A(\sound4.sdiv.A[26] ),
    .B(_2054_),
    .Y(_2055_));
 sky130_fd_sc_hd__xnor2_1 _5573_ (.A(\sound4.divisor_m[14] ),
    .B(_2055_),
    .Y(_2056_));
 sky130_fd_sc_hd__xnor2_1 _5574_ (.A(\sound4.sdiv.A[13] ),
    .B(_2056_),
    .Y(_2057_));
 sky130_fd_sc_hd__inv_2 _5575_ (.A(\sound4.sdiv.A[12] ),
    .Y(_2058_));
 sky130_fd_sc_hd__and2_1 _5576_ (.A(_2036_),
    .B(_2032_),
    .X(_2059_));
 sky130_fd_sc_hd__xnor2_2 _5577_ (.A(\sound4.divisor_m[13] ),
    .B(_2059_),
    .Y(_2060_));
 sky130_fd_sc_hd__nand2_1 _5578_ (.A(_2058_),
    .B(_2060_),
    .Y(_2061_));
 sky130_fd_sc_hd__inv_2 _5579_ (.A(_2060_),
    .Y(_2062_));
 sky130_fd_sc_hd__inv_2 _5580_ (.A(\sound4.sdiv.A[11] ),
    .Y(_2063_));
 sky130_fd_sc_hd__nand2_1 _5581_ (.A(_2036_),
    .B(_2031_),
    .Y(_2064_));
 sky130_fd_sc_hd__xor2_1 _5582_ (.A(\sound4.divisor_m[12] ),
    .B(_2064_),
    .X(_2065_));
 sky130_fd_sc_hd__or2_1 _5583_ (.A(_2063_),
    .B(_2065_),
    .X(_2066_));
 sky130_fd_sc_hd__inv_2 _5584_ (.A(_2066_),
    .Y(_2067_));
 sky130_fd_sc_hd__and2_1 _5585_ (.A(_2063_),
    .B(_2065_),
    .X(_2068_));
 sky130_fd_sc_hd__nor2_1 _5586_ (.A(_2067_),
    .B(_2068_),
    .Y(_2069_));
 sky130_fd_sc_hd__inv_2 _5587_ (.A(\sound4.sdiv.A[10] ),
    .Y(_2070_));
 sky130_fd_sc_hd__o21a_1 _5588_ (.A1(\sound4.divisor_m[10] ),
    .A2(_2030_),
    .B1(_2036_),
    .X(_2071_));
 sky130_fd_sc_hd__xnor2_1 _5589_ (.A(\sound4.divisor_m[11] ),
    .B(_2071_),
    .Y(_2072_));
 sky130_fd_sc_hd__nand2_1 _5590_ (.A(_2070_),
    .B(_2072_),
    .Y(_2073_));
 sky130_fd_sc_hd__and2_1 _5591_ (.A(_2036_),
    .B(_2030_),
    .X(_2074_));
 sky130_fd_sc_hd__xnor2_1 _5592_ (.A(\sound4.divisor_m[10] ),
    .B(_2074_),
    .Y(_2075_));
 sky130_fd_sc_hd__inv_2 _5593_ (.A(_2075_),
    .Y(_2076_));
 sky130_fd_sc_hd__nand2_1 _5594_ (.A(\sound4.sdiv.A[9] ),
    .B(_2076_),
    .Y(_2077_));
 sky130_fd_sc_hd__or2_1 _5595_ (.A(\sound4.sdiv.A[9] ),
    .B(_2076_),
    .X(_2078_));
 sky130_fd_sc_hd__nand2_1 _5596_ (.A(_2077_),
    .B(_2078_),
    .Y(_2079_));
 sky130_fd_sc_hd__and2_1 _5597_ (.A(_2036_),
    .B(_2029_),
    .X(_2080_));
 sky130_fd_sc_hd__xnor2_1 _5598_ (.A(\sound4.divisor_m[9] ),
    .B(_2080_),
    .Y(_2081_));
 sky130_fd_sc_hd__inv_2 _5599_ (.A(_2081_),
    .Y(_2082_));
 sky130_fd_sc_hd__or2_1 _5600_ (.A(\sound4.sdiv.A[8] ),
    .B(_2082_),
    .X(_2083_));
 sky130_fd_sc_hd__o21a_1 _5601_ (.A1(\sound4.divisor_m[7] ),
    .A2(_2028_),
    .B1(_2036_),
    .X(_2084_));
 sky130_fd_sc_hd__xnor2_1 _5602_ (.A(\sound4.divisor_m[8] ),
    .B(_2084_),
    .Y(_2085_));
 sky130_fd_sc_hd__inv_2 _5603_ (.A(_2085_),
    .Y(_2086_));
 sky130_fd_sc_hd__nand2_1 _5604_ (.A(\sound4.sdiv.A[7] ),
    .B(_2086_),
    .Y(_2087_));
 sky130_fd_sc_hd__or2_1 _5605_ (.A(\sound4.sdiv.A[7] ),
    .B(_2086_),
    .X(_2088_));
 sky130_fd_sc_hd__nand2_1 _5606_ (.A(_2087_),
    .B(_2088_),
    .Y(_2089_));
 sky130_fd_sc_hd__and2_1 _5607_ (.A(_2036_),
    .B(_2028_),
    .X(_2090_));
 sky130_fd_sc_hd__xnor2_1 _5608_ (.A(\sound4.divisor_m[7] ),
    .B(_2090_),
    .Y(_2091_));
 sky130_fd_sc_hd__inv_2 _5609_ (.A(_2091_),
    .Y(_2092_));
 sky130_fd_sc_hd__or2_1 _5610_ (.A(\sound4.sdiv.A[6] ),
    .B(_2092_),
    .X(_2093_));
 sky130_fd_sc_hd__and2_1 _5611_ (.A(_2036_),
    .B(_2027_),
    .X(_2094_));
 sky130_fd_sc_hd__xnor2_1 _5612_ (.A(\sound4.divisor_m[6] ),
    .B(_2094_),
    .Y(_2095_));
 sky130_fd_sc_hd__inv_2 _5613_ (.A(_2095_),
    .Y(_2096_));
 sky130_fd_sc_hd__nand2_1 _5614_ (.A(\sound4.sdiv.A[5] ),
    .B(_2096_),
    .Y(_2097_));
 sky130_fd_sc_hd__or2_1 _5615_ (.A(\sound4.sdiv.A[5] ),
    .B(_2096_),
    .X(_2098_));
 sky130_fd_sc_hd__nand2_1 _5616_ (.A(_2097_),
    .B(_2098_),
    .Y(_2099_));
 sky130_fd_sc_hd__o21a_1 _5617_ (.A1(\sound4.divisor_m[4] ),
    .A2(_2026_),
    .B1(_2036_),
    .X(_2100_));
 sky130_fd_sc_hd__xnor2_1 _5618_ (.A(\sound4.divisor_m[5] ),
    .B(_2100_),
    .Y(_2101_));
 sky130_fd_sc_hd__inv_2 _5619_ (.A(_2101_),
    .Y(_2102_));
 sky130_fd_sc_hd__or2_1 _5620_ (.A(\sound4.sdiv.A[4] ),
    .B(_2102_),
    .X(_2103_));
 sky130_fd_sc_hd__inv_2 _5621_ (.A(\sound4.sdiv.A[3] ),
    .Y(_2104_));
 sky130_fd_sc_hd__nand2_1 _5622_ (.A(_2036_),
    .B(_2026_),
    .Y(_2105_));
 sky130_fd_sc_hd__xor2_1 _5623_ (.A(\sound4.divisor_m[4] ),
    .B(_2105_),
    .X(_2106_));
 sky130_fd_sc_hd__nor2_1 _5624_ (.A(_2104_),
    .B(_2106_),
    .Y(_2107_));
 sky130_fd_sc_hd__and2_1 _5625_ (.A(_2104_),
    .B(_2106_),
    .X(_2108_));
 sky130_fd_sc_hd__or2_1 _5626_ (.A(_2107_),
    .B(_2108_),
    .X(_2109_));
 sky130_fd_sc_hd__inv_2 _5627_ (.A(_2109_),
    .Y(_2110_));
 sky130_fd_sc_hd__inv_2 _5628_ (.A(\sound4.sdiv.A[2] ),
    .Y(_2111_));
 sky130_fd_sc_hd__o31a_1 _5629_ (.A1(\sound4.divisor_m[2] ),
    .A2(\sound4.divisor_m[1] ),
    .A3(\sound4.divisor_m[0] ),
    .B1(_2036_),
    .X(_2112_));
 sky130_fd_sc_hd__xnor2_1 _5630_ (.A(\sound4.divisor_m[3] ),
    .B(_2112_),
    .Y(_2113_));
 sky130_fd_sc_hd__or2_1 _5631_ (.A(_2111_),
    .B(_2113_),
    .X(_2114_));
 sky130_fd_sc_hd__nand2_1 _5632_ (.A(_2111_),
    .B(_2113_),
    .Y(_2115_));
 sky130_fd_sc_hd__nand2_1 _5633_ (.A(_2114_),
    .B(_2115_),
    .Y(_2116_));
 sky130_fd_sc_hd__inv_2 _5634_ (.A(\sound4.sdiv.A[1] ),
    .Y(_2117_));
 sky130_fd_sc_hd__o21a_1 _5635_ (.A1(\sound4.divisor_m[1] ),
    .A2(\sound4.divisor_m[0] ),
    .B1(_2036_),
    .X(_2118_));
 sky130_fd_sc_hd__xnor2_1 _5636_ (.A(\sound4.divisor_m[2] ),
    .B(_2118_),
    .Y(_2119_));
 sky130_fd_sc_hd__xnor2_1 _5637_ (.A(_2117_),
    .B(_2119_),
    .Y(_2120_));
 sky130_fd_sc_hd__and2b_1 _5638_ (.A_N(\sound4.sdiv.A[26] ),
    .B(\sound4.divisor_m[0] ),
    .X(_2121_));
 sky130_fd_sc_hd__xnor2_2 _5639_ (.A(\sound4.divisor_m[1] ),
    .B(_2121_),
    .Y(_2122_));
 sky130_fd_sc_hd__xnor2_2 _5640_ (.A(\sound4.sdiv.A[0] ),
    .B(_2122_),
    .Y(_2123_));
 sky130_fd_sc_hd__and2b_1 _5641_ (.A_N(_2122_),
    .B(\sound4.sdiv.A[0] ),
    .X(_2124_));
 sky130_fd_sc_hd__a31oi_2 _5642_ (.A1(\sound4.divisor_m[0] ),
    .A2(\sound4.sdiv.Q[27] ),
    .A3(_2123_),
    .B1(_2124_),
    .Y(_2125_));
 sky130_fd_sc_hd__or2_1 _5643_ (.A(_2117_),
    .B(_2119_),
    .X(_2126_));
 sky130_fd_sc_hd__o21a_1 _5644_ (.A1(_2120_),
    .A2(_2125_),
    .B1(_2126_),
    .X(_2127_));
 sky130_fd_sc_hd__o21ai_1 _5645_ (.A1(_2116_),
    .A2(_2127_),
    .B1(_2114_),
    .Y(_2128_));
 sky130_fd_sc_hd__a21o_1 _5646_ (.A1(_2110_),
    .A2(_2128_),
    .B1(_2107_),
    .X(_2129_));
 sky130_fd_sc_hd__nand2_1 _5647_ (.A(\sound4.sdiv.A[4] ),
    .B(_2102_),
    .Y(_2130_));
 sky130_fd_sc_hd__a21boi_1 _5648_ (.A1(_2103_),
    .A2(_2129_),
    .B1_N(_2130_),
    .Y(_2131_));
 sky130_fd_sc_hd__o21ai_1 _5649_ (.A1(_2099_),
    .A2(_2131_),
    .B1(_2097_),
    .Y(_2132_));
 sky130_fd_sc_hd__nand2_1 _5650_ (.A(\sound4.sdiv.A[6] ),
    .B(_2092_),
    .Y(_2133_));
 sky130_fd_sc_hd__a21boi_1 _5651_ (.A1(_2093_),
    .A2(_2132_),
    .B1_N(_2133_),
    .Y(_2134_));
 sky130_fd_sc_hd__o21ai_1 _5652_ (.A1(_2089_),
    .A2(_2134_),
    .B1(_2087_),
    .Y(_2135_));
 sky130_fd_sc_hd__nand2_1 _5653_ (.A(\sound4.sdiv.A[8] ),
    .B(_2082_),
    .Y(_2136_));
 sky130_fd_sc_hd__a21boi_1 _5654_ (.A1(_2083_),
    .A2(_2135_),
    .B1_N(_2136_),
    .Y(_2137_));
 sky130_fd_sc_hd__o21ai_1 _5655_ (.A1(_2079_),
    .A2(_2137_),
    .B1(_2077_),
    .Y(_2138_));
 sky130_fd_sc_hd__nor2_1 _5656_ (.A(_2070_),
    .B(_2072_),
    .Y(_2139_));
 sky130_fd_sc_hd__a21o_1 _5657_ (.A1(_2073_),
    .A2(_2138_),
    .B1(_2139_),
    .X(_2140_));
 sky130_fd_sc_hd__a221o_1 _5658_ (.A1(\sound4.sdiv.A[12] ),
    .A2(_2062_),
    .B1(_2069_),
    .B2(_2140_),
    .C1(_2067_),
    .X(_2141_));
 sky130_fd_sc_hd__inv_2 _5659_ (.A(\sound4.divisor_m[14] ),
    .Y(_2142_));
 sky130_fd_sc_hd__a21o_1 _5660_ (.A1(_2142_),
    .A2(_2054_),
    .B1(\sound4.sdiv.A[26] ),
    .X(_2143_));
 sky130_fd_sc_hd__xnor2_1 _5661_ (.A(\sound4.divisor_m[15] ),
    .B(_2143_),
    .Y(_2144_));
 sky130_fd_sc_hd__nand2_1 _5662_ (.A(\sound4.sdiv.A[14] ),
    .B(_2144_),
    .Y(_2145_));
 sky130_fd_sc_hd__inv_2 _5663_ (.A(_2145_),
    .Y(_2146_));
 sky130_fd_sc_hd__nor2_1 _5664_ (.A(\sound4.sdiv.A[14] ),
    .B(_2144_),
    .Y(_2147_));
 sky130_fd_sc_hd__nor2_1 _5665_ (.A(_2146_),
    .B(_2147_),
    .Y(_2148_));
 sky130_fd_sc_hd__inv_2 _5666_ (.A(\sound4.sdiv.A[13] ),
    .Y(_2149_));
 sky130_fd_sc_hd__or2_1 _5667_ (.A(_2149_),
    .B(_2056_),
    .X(_2150_));
 sky130_fd_sc_hd__a21oi_1 _5668_ (.A1(_2145_),
    .A2(_2150_),
    .B1(_2147_),
    .Y(_2151_));
 sky130_fd_sc_hd__a41o_1 _5669_ (.A1(_2057_),
    .A2(_2061_),
    .A3(_2141_),
    .A4(_2148_),
    .B1(_2151_),
    .X(_2152_));
 sky130_fd_sc_hd__and2_1 _5670_ (.A(_2050_),
    .B(_2052_),
    .X(_2153_));
 sky130_fd_sc_hd__or2_1 _5671_ (.A(_2053_),
    .B(_2153_),
    .X(_2154_));
 sky130_fd_sc_hd__nor2_1 _5672_ (.A(_2046_),
    .B(_2048_),
    .Y(_2155_));
 sky130_fd_sc_hd__or2b_1 _5673_ (.A(_2155_),
    .B_N(_2049_),
    .X(_2156_));
 sky130_fd_sc_hd__nor2_1 _5674_ (.A(_2154_),
    .B(_2156_),
    .Y(_2157_));
 sky130_fd_sc_hd__a221o_1 _5675_ (.A1(_2049_),
    .A2(_2053_),
    .B1(_2152_),
    .B2(_2157_),
    .C1(_2155_),
    .X(_2158_));
 sky130_fd_sc_hd__inv_2 _5676_ (.A(\sound4.sdiv.A[17] ),
    .Y(_2159_));
 sky130_fd_sc_hd__and2_1 _5677_ (.A(_2036_),
    .B(_2035_),
    .X(_2160_));
 sky130_fd_sc_hd__xnor2_1 _5678_ (.A(\sound4.divisor_m[18] ),
    .B(_2160_),
    .Y(_2161_));
 sky130_fd_sc_hd__nor2_1 _5679_ (.A(_2159_),
    .B(_2161_),
    .Y(_2162_));
 sky130_fd_sc_hd__nand2_1 _5680_ (.A(_2159_),
    .B(_2161_),
    .Y(_2163_));
 sky130_fd_sc_hd__or2b_1 _5681_ (.A(_2162_),
    .B_N(_2163_),
    .X(_2164_));
 sky130_fd_sc_hd__xnor2_1 _5682_ (.A(\sound4.sdiv.A[18] ),
    .B(_2037_),
    .Y(_2165_));
 sky130_fd_sc_hd__nor2_1 _5683_ (.A(_2164_),
    .B(_2165_),
    .Y(_2166_));
 sky130_fd_sc_hd__o21a_1 _5684_ (.A1(\sound4.sdiv.A[18] ),
    .A2(_2038_),
    .B1(_2162_),
    .X(_2167_));
 sky130_fd_sc_hd__a221o_1 _5685_ (.A1(\sound4.sdiv.A[18] ),
    .A2(_2038_),
    .B1(_2158_),
    .B2(_2166_),
    .C1(_2167_),
    .X(_2168_));
 sky130_fd_sc_hd__or4b_2 _5686_ (.A(_2042_),
    .B(_2044_),
    .C(_2045_),
    .D_N(_2168_),
    .X(_2169_));
 sky130_fd_sc_hd__o21ai_2 _5687_ (.A1(\sound4.sdiv.A[22] ),
    .A2(\sound4.sdiv.A[21] ),
    .B1(_2038_),
    .Y(_2170_));
 sky130_fd_sc_hd__o21ai_4 _5688_ (.A1(\sound4.sdiv.A[20] ),
    .A2(\sound4.sdiv.A[19] ),
    .B1(_2038_),
    .Y(_2171_));
 sky130_fd_sc_hd__nor2_1 _5689_ (.A(\sound4.sdiv.A[23] ),
    .B(_2038_),
    .Y(_2172_));
 sky130_fd_sc_hd__and2_2 _5690_ (.A(\sound4.sdiv.A[23] ),
    .B(_2038_),
    .X(_2173_));
 sky130_fd_sc_hd__a311oi_4 _5691_ (.A1(_2169_),
    .A2(_2170_),
    .A3(_2171_),
    .B1(_2172_),
    .C1(_2173_),
    .Y(_2174_));
 sky130_fd_sc_hd__o21ai_1 _5692_ (.A1(\sound4.sdiv.A[24] ),
    .A2(_2038_),
    .B1(_2174_),
    .Y(_2175_));
 sky130_fd_sc_hd__o21ai_1 _5693_ (.A1(\sound4.sdiv.A[24] ),
    .A2(\sound4.sdiv.A[23] ),
    .B1(_2038_),
    .Y(_2176_));
 sky130_fd_sc_hd__or2_1 _5694_ (.A(\sound4.sdiv.A[25] ),
    .B(_2038_),
    .X(_2177_));
 sky130_fd_sc_hd__nand2_1 _5695_ (.A(_2039_),
    .B(_2177_),
    .Y(_2178_));
 sky130_fd_sc_hd__a21o_1 _5696_ (.A1(_2175_),
    .A2(_2176_),
    .B1(_2178_),
    .X(_2179_));
 sky130_fd_sc_hd__o311a_1 _5697_ (.A1(\sound4.divisor_m[18] ),
    .A2(\sound4.sdiv.A[26] ),
    .A3(_2035_),
    .B1(_2039_),
    .C1(_2179_),
    .X(_2180_));
 sky130_fd_sc_hd__and2_2 _5698_ (.A(\sound4.sdiv.Q[0] ),
    .B(_0576_),
    .X(_2181_));
 sky130_fd_sc_hd__o21bai_1 _5699_ (.A1(_1763_),
    .A2(_2180_),
    .B1_N(_2181_),
    .Y(_0000_));
 sky130_fd_sc_hd__clkbuf_8 _5700_ (.A(_0576_),
    .X(_2182_));
 sky130_fd_sc_hd__clkbuf_8 _5701_ (.A(_2182_),
    .X(_2183_));
 sky130_fd_sc_hd__a22o_1 _5702_ (.A1(\sound4.sdiv.Q[1] ),
    .A2(_2183_),
    .B1(\sound4.sdiv.next_dived ),
    .B2(\sound4.sdiv.Q[0] ),
    .X(_0001_));
 sky130_fd_sc_hd__a22o_1 _5703_ (.A1(\sound4.sdiv.Q[2] ),
    .A2(_2183_),
    .B1(\sound4.sdiv.next_dived ),
    .B2(\sound4.sdiv.Q[1] ),
    .X(_0002_));
 sky130_fd_sc_hd__a22o_1 _5704_ (.A1(\sound4.sdiv.Q[3] ),
    .A2(_2183_),
    .B1(\sound4.sdiv.next_dived ),
    .B2(\sound4.sdiv.Q[2] ),
    .X(_0003_));
 sky130_fd_sc_hd__a22o_1 _5705_ (.A1(\sound4.sdiv.Q[4] ),
    .A2(_2183_),
    .B1(\sound4.sdiv.next_dived ),
    .B2(\sound4.sdiv.Q[3] ),
    .X(_0004_));
 sky130_fd_sc_hd__a22o_1 _5706_ (.A1(\sound4.sdiv.Q[5] ),
    .A2(_2183_),
    .B1(\sound4.sdiv.next_dived ),
    .B2(\sound4.sdiv.Q[4] ),
    .X(_0005_));
 sky130_fd_sc_hd__a22o_1 _5707_ (.A1(\sound4.sdiv.Q[6] ),
    .A2(_2183_),
    .B1(\sound4.sdiv.next_dived ),
    .B2(\sound4.sdiv.Q[5] ),
    .X(_0006_));
 sky130_fd_sc_hd__a22o_1 _5708_ (.A1(\sound4.sdiv.Q[7] ),
    .A2(_2183_),
    .B1(\sound4.sdiv.next_dived ),
    .B2(\sound4.sdiv.Q[6] ),
    .X(_0007_));
 sky130_fd_sc_hd__buf_6 _5709_ (.A(_0576_),
    .X(_2184_));
 sky130_fd_sc_hd__clkbuf_8 _5710_ (.A(_1764_),
    .X(_2185_));
 sky130_fd_sc_hd__buf_4 _5711_ (.A(_0575_),
    .X(_2186_));
 sky130_fd_sc_hd__and2_1 _5712_ (.A(\sound4.count[0] ),
    .B(_2186_),
    .X(_2187_));
 sky130_fd_sc_hd__a221o_1 _5713_ (.A1(\sound4.sdiv.Q[8] ),
    .A2(_2184_),
    .B1(_2185_),
    .B2(\sound4.sdiv.Q[7] ),
    .C1(_2187_),
    .X(_0008_));
 sky130_fd_sc_hd__and2_1 _5714_ (.A(\sound4.count[1] ),
    .B(_2186_),
    .X(_2188_));
 sky130_fd_sc_hd__a221o_1 _5715_ (.A1(\sound4.sdiv.Q[9] ),
    .A2(_2184_),
    .B1(_2185_),
    .B2(\sound4.sdiv.Q[8] ),
    .C1(_2188_),
    .X(_0009_));
 sky130_fd_sc_hd__and2_1 _5716_ (.A(\sound4.count[2] ),
    .B(_2186_),
    .X(_2189_));
 sky130_fd_sc_hd__a221o_1 _5717_ (.A1(\sound4.sdiv.Q[10] ),
    .A2(_2182_),
    .B1(_2185_),
    .B2(\sound4.sdiv.Q[9] ),
    .C1(_2189_),
    .X(_0010_));
 sky130_fd_sc_hd__and2_1 _5718_ (.A(\sound4.count[3] ),
    .B(_2186_),
    .X(_2190_));
 sky130_fd_sc_hd__a221o_1 _5719_ (.A1(\sound4.sdiv.Q[11] ),
    .A2(_2182_),
    .B1(_2185_),
    .B2(\sound4.sdiv.Q[10] ),
    .C1(_2190_),
    .X(_0011_));
 sky130_fd_sc_hd__and2_1 _5720_ (.A(\sound4.count[4] ),
    .B(_2186_),
    .X(_2191_));
 sky130_fd_sc_hd__a221o_1 _5721_ (.A1(\sound4.sdiv.Q[12] ),
    .A2(_2182_),
    .B1(_2185_),
    .B2(\sound4.sdiv.Q[11] ),
    .C1(_2191_),
    .X(_0012_));
 sky130_fd_sc_hd__and2_1 _5722_ (.A(\sound4.count[5] ),
    .B(_2186_),
    .X(_2192_));
 sky130_fd_sc_hd__a221o_1 _5723_ (.A1(\sound4.sdiv.Q[13] ),
    .A2(_2182_),
    .B1(_2185_),
    .B2(\sound4.sdiv.Q[12] ),
    .C1(_2192_),
    .X(_0013_));
 sky130_fd_sc_hd__and2_1 _5724_ (.A(\sound4.count[6] ),
    .B(_2186_),
    .X(_2193_));
 sky130_fd_sc_hd__a221o_1 _5725_ (.A1(\sound4.sdiv.Q[14] ),
    .A2(_2182_),
    .B1(_2185_),
    .B2(\sound4.sdiv.Q[13] ),
    .C1(_2193_),
    .X(_0014_));
 sky130_fd_sc_hd__and2_1 _5726_ (.A(\sound4.count[7] ),
    .B(_2186_),
    .X(_2194_));
 sky130_fd_sc_hd__a221o_1 _5727_ (.A1(\sound4.sdiv.Q[15] ),
    .A2(_2182_),
    .B1(_2185_),
    .B2(\sound4.sdiv.Q[14] ),
    .C1(_2194_),
    .X(_0015_));
 sky130_fd_sc_hd__and2_1 _5728_ (.A(\sound4.count[8] ),
    .B(_2186_),
    .X(_2195_));
 sky130_fd_sc_hd__a221o_1 _5729_ (.A1(\sound4.sdiv.Q[16] ),
    .A2(_2182_),
    .B1(_2185_),
    .B2(\sound4.sdiv.Q[15] ),
    .C1(_2195_),
    .X(_0016_));
 sky130_fd_sc_hd__and2_1 _5730_ (.A(\sound4.count[9] ),
    .B(_2186_),
    .X(_2196_));
 sky130_fd_sc_hd__a221o_1 _5731_ (.A1(\sound4.sdiv.Q[17] ),
    .A2(_2182_),
    .B1(_2185_),
    .B2(\sound4.sdiv.Q[16] ),
    .C1(_2196_),
    .X(_0017_));
 sky130_fd_sc_hd__and2_1 _5732_ (.A(\sound4.count[10] ),
    .B(_2186_),
    .X(_2197_));
 sky130_fd_sc_hd__a221o_1 _5733_ (.A1(\sound4.sdiv.Q[18] ),
    .A2(_2182_),
    .B1(_2185_),
    .B2(\sound4.sdiv.Q[17] ),
    .C1(_2197_),
    .X(_0018_));
 sky130_fd_sc_hd__and2_1 _5734_ (.A(\sound4.count[11] ),
    .B(_2186_),
    .X(_2198_));
 sky130_fd_sc_hd__a221o_1 _5735_ (.A1(\sound4.sdiv.Q[19] ),
    .A2(_2182_),
    .B1(_2185_),
    .B2(\sound4.sdiv.Q[18] ),
    .C1(_2198_),
    .X(_0019_));
 sky130_fd_sc_hd__and2_1 _5736_ (.A(\sound4.count[12] ),
    .B(_2186_),
    .X(_2199_));
 sky130_fd_sc_hd__a221o_1 _5737_ (.A1(\sound4.sdiv.Q[20] ),
    .A2(_2182_),
    .B1(_2185_),
    .B2(\sound4.sdiv.Q[19] ),
    .C1(_2199_),
    .X(_0020_));
 sky130_fd_sc_hd__and2_1 _5738_ (.A(\sound4.count[13] ),
    .B(_2186_),
    .X(_2200_));
 sky130_fd_sc_hd__a221o_1 _5739_ (.A1(\sound4.sdiv.Q[21] ),
    .A2(_2182_),
    .B1(_2185_),
    .B2(\sound4.sdiv.Q[20] ),
    .C1(_2200_),
    .X(_0021_));
 sky130_fd_sc_hd__clkbuf_8 _5740_ (.A(_0575_),
    .X(_2201_));
 sky130_fd_sc_hd__and2_1 _5741_ (.A(\sound4.count[14] ),
    .B(_2201_),
    .X(_2202_));
 sky130_fd_sc_hd__a221o_1 _5742_ (.A1(\sound4.sdiv.Q[22] ),
    .A2(_2182_),
    .B1(_2185_),
    .B2(\sound4.sdiv.Q[21] ),
    .C1(_2202_),
    .X(_0022_));
 sky130_fd_sc_hd__and2_1 _5743_ (.A(\sound4.count[15] ),
    .B(_2201_),
    .X(_2203_));
 sky130_fd_sc_hd__a221o_1 _5744_ (.A1(\sound4.sdiv.Q[23] ),
    .A2(_2182_),
    .B1(_2185_),
    .B2(\sound4.sdiv.Q[22] ),
    .C1(_2203_),
    .X(_0023_));
 sky130_fd_sc_hd__and2_1 _5745_ (.A(\sound4.count[16] ),
    .B(_2201_),
    .X(_2204_));
 sky130_fd_sc_hd__a221o_1 _5746_ (.A1(\sound4.sdiv.Q[24] ),
    .A2(_2182_),
    .B1(_2185_),
    .B2(\sound4.sdiv.Q[23] ),
    .C1(_2204_),
    .X(_0024_));
 sky130_fd_sc_hd__and2_1 _5747_ (.A(\sound4.count[17] ),
    .B(_2201_),
    .X(_2205_));
 sky130_fd_sc_hd__a221o_1 _5748_ (.A1(\sound4.sdiv.Q[25] ),
    .A2(_2182_),
    .B1(_2185_),
    .B2(\sound4.sdiv.Q[24] ),
    .C1(_2205_),
    .X(_0025_));
 sky130_fd_sc_hd__and2_1 _5749_ (.A(\sound4.count[18] ),
    .B(_2201_),
    .X(_2206_));
 sky130_fd_sc_hd__a221o_1 _5750_ (.A1(\sound4.sdiv.Q[26] ),
    .A2(_2182_),
    .B1(_2185_),
    .B2(\sound4.sdiv.Q[25] ),
    .C1(_2206_),
    .X(_0026_));
 sky130_fd_sc_hd__a22o_1 _5751_ (.A1(\sound4.sdiv.Q[27] ),
    .A2(_2183_),
    .B1(\sound4.sdiv.next_dived ),
    .B2(\sound4.sdiv.Q[26] ),
    .X(_0027_));
 sky130_fd_sc_hd__nand2_1 _5752_ (.A(\wave_comb.u1.M[0] ),
    .B(\wave_comb.u1.Q[11] ),
    .Y(_2207_));
 sky130_fd_sc_hd__or2_1 _5753_ (.A(\wave_comb.u1.M[0] ),
    .B(\wave_comb.u1.Q[11] ),
    .X(_2208_));
 sky130_fd_sc_hd__a32o_1 _5754_ (.A1(\wave_comb.u1.next_dived ),
    .A2(_2207_),
    .A3(_2208_),
    .B1(_0573_),
    .B2(\wave_comb.u1.A[0] ),
    .X(_0028_));
 sky130_fd_sc_hd__inv_2 _5755_ (.A(\wave_comb.u1.A[10] ),
    .Y(_2209_));
 sky130_fd_sc_hd__nand2_1 _5756_ (.A(\wave_comb.u1.M[0] ),
    .B(_2209_),
    .Y(_2210_));
 sky130_fd_sc_hd__xnor2_1 _5757_ (.A(\wave_comb.u1.M[1] ),
    .B(_2210_),
    .Y(_2211_));
 sky130_fd_sc_hd__xnor2_1 _5758_ (.A(\wave_comb.u1.A[0] ),
    .B(_2211_),
    .Y(_2212_));
 sky130_fd_sc_hd__or2_1 _5759_ (.A(_2207_),
    .B(_2212_),
    .X(_2213_));
 sky130_fd_sc_hd__nand2_1 _5760_ (.A(_2207_),
    .B(_2212_),
    .Y(_2214_));
 sky130_fd_sc_hd__a32o_1 _5761_ (.A1(\wave_comb.u1.next_dived ),
    .A2(_2213_),
    .A3(_2214_),
    .B1(_0573_),
    .B2(\wave_comb.u1.A[1] ),
    .X(_0029_));
 sky130_fd_sc_hd__a21bo_1 _5762_ (.A1(\wave_comb.u1.A[0] ),
    .A2(_2211_),
    .B1_N(_2213_),
    .X(_2215_));
 sky130_fd_sc_hd__inv_2 _5763_ (.A(\wave_comb.u1.A[1] ),
    .Y(_2216_));
 sky130_fd_sc_hd__o21a_1 _5764_ (.A1(\wave_comb.u1.M[0] ),
    .A2(\wave_comb.u1.M[1] ),
    .B1(_2209_),
    .X(_2217_));
 sky130_fd_sc_hd__xnor2_1 _5765_ (.A(\wave_comb.u1.M[2] ),
    .B(_2217_),
    .Y(_2218_));
 sky130_fd_sc_hd__xnor2_1 _5766_ (.A(_2216_),
    .B(_2218_),
    .Y(_2219_));
 sky130_fd_sc_hd__xnor2_1 _5767_ (.A(_2215_),
    .B(_2219_),
    .Y(_2220_));
 sky130_fd_sc_hd__a22o_1 _5768_ (.A1(\wave_comb.u1.A[2] ),
    .A2(_0573_),
    .B1(\wave_comb.u1.next_dived ),
    .B2(_2220_),
    .X(_0030_));
 sky130_fd_sc_hd__and2b_1 _5769_ (.A_N(_2219_),
    .B(_2215_),
    .X(_2221_));
 sky130_fd_sc_hd__o21bai_1 _5770_ (.A1(_2216_),
    .A2(_2218_),
    .B1_N(_2221_),
    .Y(_2222_));
 sky130_fd_sc_hd__o31a_1 _5771_ (.A1(\wave_comb.u1.M[0] ),
    .A2(\wave_comb.u1.M[1] ),
    .A3(\wave_comb.u1.M[2] ),
    .B1(_2209_),
    .X(_2223_));
 sky130_fd_sc_hd__buf_4 _5772_ (.A(_2223_),
    .X(_2224_));
 sky130_fd_sc_hd__xnor2_1 _5773_ (.A(\wave_comb.u1.A[2] ),
    .B(_2224_),
    .Y(_2225_));
 sky130_fd_sc_hd__xnor2_1 _5774_ (.A(_2222_),
    .B(_2225_),
    .Y(_2226_));
 sky130_fd_sc_hd__a22o_1 _5775_ (.A1(\wave_comb.u1.A[3] ),
    .A2(_0573_),
    .B1(\wave_comb.u1.next_dived ),
    .B2(_2226_),
    .X(_0031_));
 sky130_fd_sc_hd__or2_1 _5776_ (.A(\wave_comb.u1.A[3] ),
    .B(_2224_),
    .X(_2227_));
 sky130_fd_sc_hd__nand2_1 _5777_ (.A(\wave_comb.u1.A[3] ),
    .B(_2224_),
    .Y(_2228_));
 sky130_fd_sc_hd__nand2_1 _5778_ (.A(_2227_),
    .B(_2228_),
    .Y(_2229_));
 sky130_fd_sc_hd__or2b_1 _5779_ (.A(_2225_),
    .B_N(_2222_),
    .X(_2230_));
 sky130_fd_sc_hd__a21bo_1 _5780_ (.A1(\wave_comb.u1.A[2] ),
    .A2(_2224_),
    .B1_N(_2230_),
    .X(_2231_));
 sky130_fd_sc_hd__xnor2_1 _5781_ (.A(_2229_),
    .B(_2231_),
    .Y(_2232_));
 sky130_fd_sc_hd__a22o_1 _5782_ (.A1(\wave_comb.u1.A[4] ),
    .A2(_0573_),
    .B1(\wave_comb.u1.next_dived ),
    .B2(_2232_),
    .X(_0032_));
 sky130_fd_sc_hd__or2b_1 _5783_ (.A(_2229_),
    .B_N(_2231_),
    .X(_2233_));
 sky130_fd_sc_hd__xnor2_1 _5784_ (.A(\wave_comb.u1.A[4] ),
    .B(_2224_),
    .Y(_2234_));
 sky130_fd_sc_hd__a21o_1 _5785_ (.A1(_2228_),
    .A2(_2233_),
    .B1(_2234_),
    .X(_2235_));
 sky130_fd_sc_hd__nand3_1 _5786_ (.A(_2228_),
    .B(_2233_),
    .C(_2234_),
    .Y(_2236_));
 sky130_fd_sc_hd__a32o_1 _5787_ (.A1(\wave_comb.u1.next_dived ),
    .A2(_2235_),
    .A3(_2236_),
    .B1(_0573_),
    .B2(\wave_comb.u1.A[5] ),
    .X(_0033_));
 sky130_fd_sc_hd__or2_1 _5788_ (.A(\wave_comb.u1.A[5] ),
    .B(_2224_),
    .X(_2237_));
 sky130_fd_sc_hd__nand2_1 _5789_ (.A(\wave_comb.u1.A[5] ),
    .B(_2224_),
    .Y(_2238_));
 sky130_fd_sc_hd__nand2_1 _5790_ (.A(_2237_),
    .B(_2238_),
    .Y(_2239_));
 sky130_fd_sc_hd__o21ai_1 _5791_ (.A1(\wave_comb.u1.A[4] ),
    .A2(\wave_comb.u1.A[3] ),
    .B1(_2224_),
    .Y(_2240_));
 sky130_fd_sc_hd__or2_1 _5792_ (.A(_2233_),
    .B(_2234_),
    .X(_2241_));
 sky130_fd_sc_hd__nand3_1 _5793_ (.A(_2239_),
    .B(_2240_),
    .C(_2241_),
    .Y(_2242_));
 sky130_fd_sc_hd__a21o_1 _5794_ (.A1(_2240_),
    .A2(_2241_),
    .B1(_2239_),
    .X(_2243_));
 sky130_fd_sc_hd__a32o_1 _5795_ (.A1(\wave_comb.u1.next_dived ),
    .A2(_2242_),
    .A3(_2243_),
    .B1(_0573_),
    .B2(\wave_comb.u1.A[6] ),
    .X(_0034_));
 sky130_fd_sc_hd__xnor2_1 _5796_ (.A(\wave_comb.u1.A[6] ),
    .B(_2224_),
    .Y(_2244_));
 sky130_fd_sc_hd__nand3_1 _5797_ (.A(_2238_),
    .B(_2243_),
    .C(_2244_),
    .Y(_2245_));
 sky130_fd_sc_hd__a21o_1 _5798_ (.A1(_2238_),
    .A2(_2243_),
    .B1(_2244_),
    .X(_2246_));
 sky130_fd_sc_hd__a32o_1 _5799_ (.A1(\wave_comb.u1.next_dived ),
    .A2(_2245_),
    .A3(_2246_),
    .B1(_0573_),
    .B2(\wave_comb.u1.A[7] ),
    .X(_0035_));
 sky130_fd_sc_hd__nand2_1 _5800_ (.A(\wave_comb.u1.A[7] ),
    .B(_2224_),
    .Y(_2247_));
 sky130_fd_sc_hd__or2_1 _5801_ (.A(\wave_comb.u1.A[7] ),
    .B(_2224_),
    .X(_2248_));
 sky130_fd_sc_hd__nand2_1 _5802_ (.A(_2247_),
    .B(_2248_),
    .Y(_2249_));
 sky130_fd_sc_hd__nor3_1 _5803_ (.A(_2239_),
    .B(_2241_),
    .C(_2244_),
    .Y(_2250_));
 sky130_fd_sc_hd__o21a_1 _5804_ (.A1(\wave_comb.u1.A[6] ),
    .A2(\wave_comb.u1.A[5] ),
    .B1(_2224_),
    .X(_2251_));
 sky130_fd_sc_hd__or3b_1 _5805_ (.A(_2250_),
    .B(_2251_),
    .C_N(_2240_),
    .X(_2252_));
 sky130_fd_sc_hd__xnor2_1 _5806_ (.A(_2249_),
    .B(_2252_),
    .Y(_2253_));
 sky130_fd_sc_hd__a22o_1 _5807_ (.A1(\wave_comb.u1.A[8] ),
    .A2(_0573_),
    .B1(\wave_comb.u1.next_dived ),
    .B2(_2253_),
    .X(_0036_));
 sky130_fd_sc_hd__nand2_1 _5808_ (.A(\wave_comb.u1.A[8] ),
    .B(_2224_),
    .Y(_2254_));
 sky130_fd_sc_hd__or2_1 _5809_ (.A(\wave_comb.u1.A[8] ),
    .B(_2224_),
    .X(_2255_));
 sky130_fd_sc_hd__nand2_1 _5810_ (.A(_2254_),
    .B(_2255_),
    .Y(_2256_));
 sky130_fd_sc_hd__a21boi_1 _5811_ (.A1(_2248_),
    .A2(_2252_),
    .B1_N(_2247_),
    .Y(_2257_));
 sky130_fd_sc_hd__xor2_1 _5812_ (.A(_2256_),
    .B(_2257_),
    .X(_2258_));
 sky130_fd_sc_hd__a22o_1 _5813_ (.A1(\wave_comb.u1.A[9] ),
    .A2(_0573_),
    .B1(\wave_comb.u1.next_dived ),
    .B2(_2258_),
    .X(_0037_));
 sky130_fd_sc_hd__o21bai_1 _5814_ (.A1(\wave_comb.u1.A[8] ),
    .A2(_2224_),
    .B1_N(_2257_),
    .Y(_2259_));
 sky130_fd_sc_hd__xnor2_1 _5815_ (.A(\wave_comb.u1.A[9] ),
    .B(_2224_),
    .Y(_2260_));
 sky130_fd_sc_hd__a21oi_1 _5816_ (.A1(_2254_),
    .A2(_2259_),
    .B1(_2260_),
    .Y(_2261_));
 sky130_fd_sc_hd__a311o_1 _5817_ (.A1(_2254_),
    .A2(_2260_),
    .A3(_2259_),
    .B1(_0573_),
    .C1(_0645_),
    .X(_2262_));
 sky130_fd_sc_hd__a2bb2o_1 _5818_ (.A1_N(_2261_),
    .A2_N(_2262_),
    .B1(\wave_comb.u1.A[10] ),
    .B2(_0573_),
    .X(_0038_));
 sky130_fd_sc_hd__mux2_1 _5819_ (.A0(_0646_),
    .A1(_0573_),
    .S(\wave_comb.u1.C[0] ),
    .X(_2263_));
 sky130_fd_sc_hd__clkbuf_1 _5820_ (.A(_2263_),
    .X(_0039_));
 sky130_fd_sc_hd__nand2_1 _5821_ (.A(\wave_comb.u1.C[0] ),
    .B(\wave_comb.u1.C[1] ),
    .Y(_2264_));
 sky130_fd_sc_hd__or2_1 _5822_ (.A(\wave_comb.u1.C[0] ),
    .B(\wave_comb.u1.C[1] ),
    .X(_2265_));
 sky130_fd_sc_hd__a32o_1 _5823_ (.A1(_0646_),
    .A2(_2264_),
    .A3(_2265_),
    .B1(_0573_),
    .B2(\wave_comb.u1.C[1] ),
    .X(_0040_));
 sky130_fd_sc_hd__a21o_1 _5824_ (.A1(\wave_comb.u1.C[0] ),
    .A2(\wave_comb.u1.C[1] ),
    .B1(\wave_comb.u1.C[2] ),
    .X(_2266_));
 sky130_fd_sc_hd__nand3_1 _5825_ (.A(\wave_comb.u1.C[2] ),
    .B(\wave_comb.u1.C[0] ),
    .C(\wave_comb.u1.C[1] ),
    .Y(_2267_));
 sky130_fd_sc_hd__a32o_1 _5826_ (.A1(_0646_),
    .A2(_2266_),
    .A3(_2267_),
    .B1(_0573_),
    .B2(\wave_comb.u1.C[2] ),
    .X(_0041_));
 sky130_fd_sc_hd__o21bai_1 _5827_ (.A1(_0571_),
    .A2(_2267_),
    .B1_N(\wave_comb.u1.C[3] ),
    .Y(_2268_));
 sky130_fd_sc_hd__and2_1 _5828_ (.A(_0569_),
    .B(_2268_),
    .X(_2269_));
 sky130_fd_sc_hd__clkbuf_1 _5829_ (.A(_2269_),
    .X(_0042_));
 sky130_fd_sc_hd__and2_1 _5830_ (.A(\wave_comb.u1.C[4] ),
    .B(_0569_),
    .X(_2270_));
 sky130_fd_sc_hd__clkbuf_1 _5831_ (.A(_2270_),
    .X(_0043_));
 sky130_fd_sc_hd__and2_1 _5832_ (.A(\wave_comb.u1.C[5] ),
    .B(_0569_),
    .X(_2271_));
 sky130_fd_sc_hd__clkbuf_1 _5833_ (.A(_2271_),
    .X(_0044_));
 sky130_fd_sc_hd__nor4_1 _5834_ (.A(\wave_comb.u1.M[0] ),
    .B(\wave_comb.u1.M[1] ),
    .C(\wave_comb.u1.M[2] ),
    .D(\wave_comb.u1.A[10] ),
    .Y(_2272_));
 sky130_fd_sc_hd__a211o_1 _5835_ (.A1(\wave_comb.u1.A[9] ),
    .A2(_2224_),
    .B1(_2261_),
    .C1(_2272_),
    .X(_2273_));
 sky130_fd_sc_hd__and3_1 _5836_ (.A(\wave_comb.u1.Q[0] ),
    .B(_0569_),
    .C(_0571_),
    .X(_2274_));
 sky130_fd_sc_hd__nand2_2 _5837_ (.A(\sound3.sdiv.Q[0] ),
    .B(_0577_),
    .Y(_2275_));
 sky130_fd_sc_hd__nand2_1 _5838_ (.A(\sound2.sdiv.Q[0] ),
    .B(_0578_),
    .Y(_2276_));
 sky130_fd_sc_hd__nand2_2 _5839_ (.A(\sound1.sdiv.Q[0] ),
    .B(_0579_),
    .Y(_2277_));
 sky130_fd_sc_hd__or3b_1 _5840_ (.A(\wave.mode[0] ),
    .B(net1),
    .C_N(\wave.mode[1] ),
    .X(_2278_));
 sky130_fd_sc_hd__buf_4 _5841_ (.A(_2278_),
    .X(_2279_));
 sky130_fd_sc_hd__nor2_1 _5842_ (.A(_2279_),
    .B(_2277_),
    .Y(_2280_));
 sky130_fd_sc_hd__and3_1 _5843_ (.A(\sound2.sdiv.Q[0] ),
    .B(_0578_),
    .C(_2280_),
    .X(_2281_));
 sky130_fd_sc_hd__a21o_1 _5844_ (.A1(_2276_),
    .A2(_2277_),
    .B1(_2281_),
    .X(_2282_));
 sky130_fd_sc_hd__nor3_1 _5845_ (.A(_2275_),
    .B(_2279_),
    .C(_2282_),
    .Y(_2283_));
 sky130_fd_sc_hd__a21oi_1 _5846_ (.A1(_2275_),
    .A2(_2282_),
    .B1(_2283_),
    .Y(_2284_));
 sky130_fd_sc_hd__nand2_1 _5847_ (.A(_2181_),
    .B(_2284_),
    .Y(_2285_));
 sky130_fd_sc_hd__and2b_1 _5848_ (.A_N(net30),
    .B(net31),
    .X(_2286_));
 sky130_fd_sc_hd__o2111a_1 _5849_ (.A1(_2181_),
    .A2(_2284_),
    .B1(_2285_),
    .C1(_2286_),
    .D1(_0645_),
    .X(_2287_));
 sky130_fd_sc_hd__a211o_1 _5850_ (.A1(\wave_comb.u1.next_dived ),
    .A2(_2273_),
    .B1(_2274_),
    .C1(_2287_),
    .X(_0045_));
 sky130_fd_sc_hd__and2_1 _5851_ (.A(net30),
    .B(net31),
    .X(_2288_));
 sky130_fd_sc_hd__buf_4 _5852_ (.A(_2288_),
    .X(_2289_));
 sky130_fd_sc_hd__nor2_2 _5853_ (.A(\sound4.sdiv.next_start ),
    .B(_2279_),
    .Y(_2290_));
 sky130_fd_sc_hd__a22o_1 _5854_ (.A1(_2181_),
    .A2(_2289_),
    .B1(_2290_),
    .B2(\sound4.sdiv.Q[1] ),
    .X(_2291_));
 sky130_fd_sc_hd__nand2_8 _5855_ (.A(net30),
    .B(net31),
    .Y(_2292_));
 sky130_fd_sc_hd__nor2_2 _5856_ (.A(\sound1.sdiv.next_start ),
    .B(_2279_),
    .Y(_2293_));
 sky130_fd_sc_hd__a2bb2o_1 _5857_ (.A1_N(_2277_),
    .A2_N(_2292_),
    .B1(_2293_),
    .B2(\sound1.sdiv.Q[1] ),
    .X(_2294_));
 sky130_fd_sc_hd__nor2_1 _5858_ (.A(\sound2.sdiv.next_start ),
    .B(_2279_),
    .Y(_2295_));
 sky130_fd_sc_hd__a2bb2o_1 _5859_ (.A1_N(_2276_),
    .A2_N(_2292_),
    .B1(_2295_),
    .B2(\sound2.sdiv.Q[1] ),
    .X(_2296_));
 sky130_fd_sc_hd__and2_1 _5860_ (.A(_2294_),
    .B(_2296_),
    .X(_2297_));
 sky130_fd_sc_hd__nor2_1 _5861_ (.A(_2294_),
    .B(_2296_),
    .Y(_2298_));
 sky130_fd_sc_hd__nor2_1 _5862_ (.A(_2297_),
    .B(_2298_),
    .Y(_2299_));
 sky130_fd_sc_hd__xnor2_1 _5863_ (.A(_2281_),
    .B(_2299_),
    .Y(_2300_));
 sky130_fd_sc_hd__nor2_2 _5864_ (.A(\sound3.sdiv.next_start ),
    .B(_2279_),
    .Y(_2301_));
 sky130_fd_sc_hd__a2bb2o_1 _5865_ (.A1_N(_2275_),
    .A2_N(_2292_),
    .B1(_2301_),
    .B2(\sound3.sdiv.Q[1] ),
    .X(_2302_));
 sky130_fd_sc_hd__and2b_1 _5866_ (.A_N(_2300_),
    .B(_2302_),
    .X(_2303_));
 sky130_fd_sc_hd__and2b_1 _5867_ (.A_N(_2302_),
    .B(_2300_),
    .X(_2304_));
 sky130_fd_sc_hd__nor2_1 _5868_ (.A(_2303_),
    .B(_2304_),
    .Y(_2305_));
 sky130_fd_sc_hd__xnor2_1 _5869_ (.A(_2291_),
    .B(_2305_),
    .Y(_2306_));
 sky130_fd_sc_hd__a31o_1 _5870_ (.A1(_2181_),
    .A2(_2286_),
    .A3(_2284_),
    .B1(_2283_),
    .X(_2307_));
 sky130_fd_sc_hd__xnor2_1 _5871_ (.A(_2306_),
    .B(_2307_),
    .Y(_2308_));
 sky130_fd_sc_hd__mux2_1 _5872_ (.A0(\wave_comb.u1.Q[0] ),
    .A1(_2308_),
    .S(_0645_),
    .X(_2309_));
 sky130_fd_sc_hd__and3_1 _5873_ (.A(\wave_comb.u1.Q[1] ),
    .B(_0569_),
    .C(_0571_),
    .X(_2310_));
 sky130_fd_sc_hd__a21o_1 _5874_ (.A1(\wave_comb.u1.next_start ),
    .A2(_2309_),
    .B1(_2310_),
    .X(_0046_));
 sky130_fd_sc_hd__or2b_1 _5875_ (.A(_2306_),
    .B_N(_2307_),
    .X(_2311_));
 sky130_fd_sc_hd__inv_2 _5876_ (.A(\sound4.count_m[4] ),
    .Y(_2312_));
 sky130_fd_sc_hd__inv_2 _5877_ (.A(\sound4.count_m[3] ),
    .Y(_2313_));
 sky130_fd_sc_hd__o22a_1 _5878_ (.A1(\sound4.divisor_m[5] ),
    .A2(_2312_),
    .B1(_2313_),
    .B2(\sound4.divisor_m[4] ),
    .X(_2314_));
 sky130_fd_sc_hd__inv_2 _5879_ (.A(\sound4.count_m[7] ),
    .Y(_2315_));
 sky130_fd_sc_hd__inv_2 _5880_ (.A(\sound4.count_m[6] ),
    .Y(_2316_));
 sky130_fd_sc_hd__a22o_1 _5881_ (.A1(_2315_),
    .A2(\sound4.divisor_m[8] ),
    .B1(_2316_),
    .B2(\sound4.divisor_m[7] ),
    .X(_2317_));
 sky130_fd_sc_hd__inv_2 _5882_ (.A(\sound4.count_m[5] ),
    .Y(_2318_));
 sky130_fd_sc_hd__a22o_1 _5883_ (.A1(_2318_),
    .A2(\sound4.divisor_m[6] ),
    .B1(\sound4.divisor_m[5] ),
    .B2(_2312_),
    .X(_2319_));
 sky130_fd_sc_hd__and2b_1 _5884_ (.A_N(\sound4.count_m[2] ),
    .B(\sound4.divisor_m[3] ),
    .X(_2320_));
 sky130_fd_sc_hd__a2111oi_1 _5885_ (.A1(_2313_),
    .A2(\sound4.divisor_m[4] ),
    .B1(_2317_),
    .C1(_2319_),
    .D1(_2320_),
    .Y(_2321_));
 sky130_fd_sc_hd__inv_2 _5886_ (.A(\sound4.count_m[16] ),
    .Y(_2322_));
 sky130_fd_sc_hd__or2_1 _5887_ (.A(_2322_),
    .B(\sound4.divisor_m[17] ),
    .X(_2323_));
 sky130_fd_sc_hd__inv_2 _5888_ (.A(\sound4.count_m[12] ),
    .Y(_2324_));
 sky130_fd_sc_hd__a2bb2o_1 _5889_ (.A1_N(\sound4.count_m[13] ),
    .A2_N(_2142_),
    .B1(\sound4.divisor_m[13] ),
    .B2(_2324_),
    .X(_2325_));
 sky130_fd_sc_hd__inv_2 _5890_ (.A(\sound4.count_m[11] ),
    .Y(_2326_));
 sky130_fd_sc_hd__inv_2 _5891_ (.A(\sound4.count_m[10] ),
    .Y(_2327_));
 sky130_fd_sc_hd__a22o_1 _5892_ (.A1(_2326_),
    .A2(\sound4.divisor_m[12] ),
    .B1(_2327_),
    .B2(\sound4.divisor_m[11] ),
    .X(_2328_));
 sky130_fd_sc_hd__nor2_1 _5893_ (.A(_2326_),
    .B(\sound4.divisor_m[12] ),
    .Y(_2329_));
 sky130_fd_sc_hd__nor2_1 _5894_ (.A(\sound4.divisor_m[13] ),
    .B(_2324_),
    .Y(_2330_));
 sky130_fd_sc_hd__inv_2 _5895_ (.A(\sound4.divisor_m[15] ),
    .Y(_2331_));
 sky130_fd_sc_hd__a22o_1 _5896_ (.A1(\sound4.count_m[14] ),
    .A2(_2331_),
    .B1(\sound4.count_m[13] ),
    .B2(_2142_),
    .X(_2332_));
 sky130_fd_sc_hd__inv_2 _5897_ (.A(\sound4.count_m[9] ),
    .Y(_2333_));
 sky130_fd_sc_hd__inv_2 _5898_ (.A(\sound4.count_m[8] ),
    .Y(_2334_));
 sky130_fd_sc_hd__a22o_1 _5899_ (.A1(_2333_),
    .A2(\sound4.divisor_m[10] ),
    .B1(\sound4.divisor_m[9] ),
    .B2(_2334_),
    .X(_2335_));
 sky130_fd_sc_hd__and2b_1 _5900_ (.A_N(\sound4.divisor_m[10] ),
    .B(\sound4.count_m[9] ),
    .X(_2336_));
 sky130_fd_sc_hd__and2b_1 _5901_ (.A_N(\sound4.divisor_m[11] ),
    .B(\sound4.count_m[10] ),
    .X(_2337_));
 sky130_fd_sc_hd__or3_1 _5902_ (.A(_2335_),
    .B(_2336_),
    .C(_2337_),
    .X(_2338_));
 sky130_fd_sc_hd__or4_1 _5903_ (.A(_2329_),
    .B(_2330_),
    .C(_2332_),
    .D(_2338_),
    .X(_2339_));
 sky130_fd_sc_hd__inv_2 _5904_ (.A(\sound4.count_m[15] ),
    .Y(_2340_));
 sky130_fd_sc_hd__inv_2 _5905_ (.A(\sound4.divisor_m[16] ),
    .Y(_2341_));
 sky130_fd_sc_hd__o22a_1 _5906_ (.A1(\sound4.count_m[15] ),
    .A2(_2341_),
    .B1(\sound4.count_m[14] ),
    .B2(_2331_),
    .X(_2342_));
 sky130_fd_sc_hd__o221a_1 _5907_ (.A1(_2340_),
    .A2(\sound4.divisor_m[16] ),
    .B1(\sound4.divisor_m[9] ),
    .B2(_2334_),
    .C1(_2342_),
    .X(_2343_));
 sky130_fd_sc_hd__nor4b_1 _5908_ (.A(_2325_),
    .B(_2328_),
    .C(_2339_),
    .D_N(_2343_),
    .Y(_2344_));
 sky130_fd_sc_hd__or2_1 _5909_ (.A(_2315_),
    .B(\sound4.divisor_m[8] ),
    .X(_2345_));
 sky130_fd_sc_hd__inv_2 _5910_ (.A(\sound4.divisor_m[1] ),
    .Y(_2346_));
 sky130_fd_sc_hd__o22a_1 _5911_ (.A1(_2316_),
    .A2(\sound4.divisor_m[7] ),
    .B1(_2318_),
    .B2(\sound4.divisor_m[6] ),
    .X(_2347_));
 sky130_fd_sc_hd__or2b_1 _5912_ (.A(\sound4.divisor_m[3] ),
    .B_N(\sound4.count_m[2] ),
    .X(_2348_));
 sky130_fd_sc_hd__inv_2 _5913_ (.A(\sound4.divisor_m[18] ),
    .Y(_2349_));
 sky130_fd_sc_hd__a2bb2o_1 _5914_ (.A1_N(\sound4.count_m[17] ),
    .A2_N(_2349_),
    .B1(_2322_),
    .B2(\sound4.divisor_m[17] ),
    .X(_2350_));
 sky130_fd_sc_hd__and2b_1 _5915_ (.A_N(\sound4.count_m[1] ),
    .B(\sound4.divisor_m[2] ),
    .X(_2351_));
 sky130_fd_sc_hd__and2b_1 _5916_ (.A_N(\sound4.divisor_m[2] ),
    .B(\sound4.count_m[1] ),
    .X(_2352_));
 sky130_fd_sc_hd__a211o_1 _5917_ (.A1(_2346_),
    .A2(\sound4.count_m[0] ),
    .B1(_2351_),
    .C1(_2352_),
    .X(_2353_));
 sky130_fd_sc_hd__nor2_1 _5918_ (.A(_2350_),
    .B(_2353_),
    .Y(_2354_));
 sky130_fd_sc_hd__o2111a_1 _5919_ (.A1(_2346_),
    .A2(\sound4.count_m[0] ),
    .B1(_2347_),
    .C1(_2348_),
    .D1(_2354_),
    .X(_2355_));
 sky130_fd_sc_hd__and4_1 _5920_ (.A(_2323_),
    .B(net61),
    .C(_2345_),
    .D(_2355_),
    .X(_2356_));
 sky130_fd_sc_hd__or2b_1 _5921_ (.A(_2351_),
    .B_N(_2353_),
    .X(_2357_));
 sky130_fd_sc_hd__a221o_1 _5922_ (.A1(_2313_),
    .A2(\sound4.divisor_m[4] ),
    .B1(_2348_),
    .B2(_2357_),
    .C1(_2320_),
    .X(_2358_));
 sky130_fd_sc_hd__a21o_1 _5923_ (.A1(_2314_),
    .A2(_2358_),
    .B1(_2319_),
    .X(_2359_));
 sky130_fd_sc_hd__a21o_1 _5924_ (.A1(_2347_),
    .A2(_2359_),
    .B1(_2317_),
    .X(_2360_));
 sky130_fd_sc_hd__nor2_1 _5925_ (.A(_2336_),
    .B(_2337_),
    .Y(_2361_));
 sky130_fd_sc_hd__a21oi_1 _5926_ (.A1(_2335_),
    .A2(_2361_),
    .B1(_2328_),
    .Y(_2362_));
 sky130_fd_sc_hd__inv_2 _5927_ (.A(_2325_),
    .Y(_2363_));
 sky130_fd_sc_hd__o31a_1 _5928_ (.A1(_2362_),
    .A2(_2329_),
    .A3(_2330_),
    .B1(_2363_),
    .X(_2364_));
 sky130_fd_sc_hd__o21a_1 _5929_ (.A1(_2364_),
    .A2(_2332_),
    .B1(_2342_),
    .X(_2365_));
 sky130_fd_sc_hd__a21oi_1 _5930_ (.A1(\sound4.count_m[15] ),
    .A2(_2341_),
    .B1(_2365_),
    .Y(_2366_));
 sky130_fd_sc_hd__a31o_1 _5931_ (.A1(_2360_),
    .A2(net61),
    .A3(_2345_),
    .B1(_2366_),
    .X(_2367_));
 sky130_fd_sc_hd__a21oi_1 _5932_ (.A1(_2323_),
    .A2(_2367_),
    .B1(_2350_),
    .Y(_2368_));
 sky130_fd_sc_hd__a211o_1 _5933_ (.A1(\sound4.count_m[17] ),
    .A2(_2349_),
    .B1(\sound4.count_m[18] ),
    .C1(_2368_),
    .X(_2369_));
 sky130_fd_sc_hd__a31o_1 _5934_ (.A1(_2314_),
    .A2(_2321_),
    .A3(_2356_),
    .B1(_2369_),
    .X(_2370_));
 sky130_fd_sc_hd__nand2_1 _5935_ (.A(\sound4.sdiv.Q[1] ),
    .B(_0576_),
    .Y(_2371_));
 sky130_fd_sc_hd__a21bo_1 _5936_ (.A1(_2181_),
    .A2(_2370_),
    .B1_N(_2371_),
    .X(_2372_));
 sky130_fd_sc_hd__nand3_1 _5937_ (.A(\sound4.sdiv.Q[1] ),
    .B(_2181_),
    .C(_2370_),
    .Y(_2373_));
 sky130_fd_sc_hd__a32o_1 _5938_ (.A1(_2289_),
    .A2(_2372_),
    .A3(_2373_),
    .B1(_2290_),
    .B2(\sound4.sdiv.Q[2] ),
    .X(_2374_));
 sky130_fd_sc_hd__inv_2 _5939_ (.A(\sound1.divisor_m[15] ),
    .Y(_2375_));
 sky130_fd_sc_hd__inv_2 _5940_ (.A(\sound1.divisor_m[14] ),
    .Y(_2376_));
 sky130_fd_sc_hd__a22o_1 _5941_ (.A1(\sound1.count_m[14] ),
    .A2(_2375_),
    .B1(\sound1.count_m[13] ),
    .B2(_2376_),
    .X(_2377_));
 sky130_fd_sc_hd__inv_2 _5942_ (.A(\sound1.divisor_m[11] ),
    .Y(_2378_));
 sky130_fd_sc_hd__and2b_1 _5943_ (.A_N(\sound1.divisor_m[10] ),
    .B(\sound1.count_m[9] ),
    .X(_2379_));
 sky130_fd_sc_hd__a21o_1 _5944_ (.A1(\sound1.count_m[10] ),
    .A2(_2378_),
    .B1(_2379_),
    .X(_2380_));
 sky130_fd_sc_hd__inv_2 _5945_ (.A(\sound1.divisor_m[16] ),
    .Y(_2381_));
 sky130_fd_sc_hd__o22a_1 _5946_ (.A1(\sound1.count_m[15] ),
    .A2(_2381_),
    .B1(\sound1.count_m[14] ),
    .B2(_2375_),
    .X(_2382_));
 sky130_fd_sc_hd__inv_2 _5947_ (.A(\sound1.divisor_m[13] ),
    .Y(_2383_));
 sky130_fd_sc_hd__o22a_1 _5948_ (.A1(\sound1.count_m[13] ),
    .A2(_2376_),
    .B1(_2383_),
    .B2(\sound1.count_m[12] ),
    .X(_2384_));
 sky130_fd_sc_hd__inv_2 _5949_ (.A(\sound1.count_m[11] ),
    .Y(_2385_));
 sky130_fd_sc_hd__o2bb2a_1 _5950_ (.A1_N(_2383_),
    .A2_N(\sound1.count_m[12] ),
    .B1(_2385_),
    .B2(\sound1.divisor_m[12] ),
    .X(_2386_));
 sky130_fd_sc_hd__o2bb2a_1 _5951_ (.A1_N(_2385_),
    .A2_N(\sound1.divisor_m[12] ),
    .B1(\sound1.count_m[10] ),
    .B2(_2378_),
    .X(_2387_));
 sky130_fd_sc_hd__and4_1 _5952_ (.A(_2382_),
    .B(_2384_),
    .C(_2386_),
    .D(_2387_),
    .X(_2388_));
 sky130_fd_sc_hd__and2_1 _5953_ (.A(\sound1.count_m[15] ),
    .B(_2381_),
    .X(_2389_));
 sky130_fd_sc_hd__or2b_1 _5954_ (.A(\sound1.count_m[8] ),
    .B_N(\sound1.divisor_m[9] ),
    .X(_2390_));
 sky130_fd_sc_hd__or2b_1 _5955_ (.A(\sound1.count_m[9] ),
    .B_N(\sound1.divisor_m[10] ),
    .X(_2391_));
 sky130_fd_sc_hd__or2b_1 _5956_ (.A(\sound1.divisor_m[9] ),
    .B_N(\sound1.count_m[8] ),
    .X(_2392_));
 sky130_fd_sc_hd__and4b_1 _5957_ (.A_N(_2389_),
    .B(_2390_),
    .C(_2391_),
    .D(_2392_),
    .X(_2393_));
 sky130_fd_sc_hd__and4bb_1 _5958_ (.A_N(_2377_),
    .B_N(_2380_),
    .C(_2388_),
    .D(_2393_),
    .X(_2394_));
 sky130_fd_sc_hd__inv_2 _5959_ (.A(\sound1.divisor_m[8] ),
    .Y(_2395_));
 sky130_fd_sc_hd__inv_2 _5960_ (.A(\sound1.count_m[6] ),
    .Y(_2396_));
 sky130_fd_sc_hd__a2bb2o_1 _5961_ (.A1_N(\sound1.count_m[7] ),
    .A2_N(_2395_),
    .B1(_2396_),
    .B2(\sound1.divisor_m[7] ),
    .X(_2397_));
 sky130_fd_sc_hd__inv_2 _5962_ (.A(\sound1.count_m[5] ),
    .Y(_2398_));
 sky130_fd_sc_hd__inv_2 _5963_ (.A(\sound1.count_m[4] ),
    .Y(_2399_));
 sky130_fd_sc_hd__a22o_1 _5964_ (.A1(_2398_),
    .A2(\sound1.divisor_m[6] ),
    .B1(\sound1.divisor_m[5] ),
    .B2(_2399_),
    .X(_2400_));
 sky130_fd_sc_hd__o22a_1 _5965_ (.A1(_2396_),
    .A2(\sound1.divisor_m[7] ),
    .B1(_2398_),
    .B2(\sound1.divisor_m[6] ),
    .X(_2401_));
 sky130_fd_sc_hd__or2b_1 _5966_ (.A(\sound1.divisor_m[8] ),
    .B_N(\sound1.count_m[7] ),
    .X(_2402_));
 sky130_fd_sc_hd__o21a_1 _5967_ (.A1(\sound1.divisor_m[5] ),
    .A2(_2399_),
    .B1(_2402_),
    .X(_2403_));
 sky130_fd_sc_hd__and4bb_1 _5968_ (.A_N(_2397_),
    .B_N(_2400_),
    .C(_2401_),
    .D(_2403_),
    .X(_2404_));
 sky130_fd_sc_hd__inv_2 _5969_ (.A(\sound1.divisor_m[18] ),
    .Y(_2405_));
 sky130_fd_sc_hd__inv_2 _5970_ (.A(\sound1.divisor_m[17] ),
    .Y(_2406_));
 sky130_fd_sc_hd__o22a_1 _5971_ (.A1(\sound1.count_m[17] ),
    .A2(_2405_),
    .B1(\sound1.count_m[16] ),
    .B2(_2406_),
    .X(_2407_));
 sky130_fd_sc_hd__inv_2 _5972_ (.A(_2407_),
    .Y(_2408_));
 sky130_fd_sc_hd__inv_2 _5973_ (.A(\sound1.count_m[3] ),
    .Y(_2409_));
 sky130_fd_sc_hd__inv_2 _5974_ (.A(\sound1.count_m[2] ),
    .Y(_2410_));
 sky130_fd_sc_hd__a22o_1 _5975_ (.A1(_2409_),
    .A2(\sound1.divisor_m[4] ),
    .B1(_2410_),
    .B2(\sound1.divisor_m[3] ),
    .X(_2411_));
 sky130_fd_sc_hd__a21o_1 _5976_ (.A1(\sound1.count_m[17] ),
    .A2(_2405_),
    .B1(\sound1.count_m[18] ),
    .X(_2412_));
 sky130_fd_sc_hd__inv_2 _5977_ (.A(\sound1.divisor_m[3] ),
    .Y(_2413_));
 sky130_fd_sc_hd__and2_1 _5978_ (.A(\sound1.count_m[16] ),
    .B(_2406_),
    .X(_2414_));
 sky130_fd_sc_hd__inv_2 _5979_ (.A(\sound1.count_m[0] ),
    .Y(_2415_));
 sky130_fd_sc_hd__or2b_1 _5980_ (.A(\sound1.count_m[1] ),
    .B_N(\sound1.divisor_m[2] ),
    .X(_2416_));
 sky130_fd_sc_hd__or2b_1 _5981_ (.A(\sound1.divisor_m[2] ),
    .B_N(\sound1.count_m[1] ),
    .X(_2417_));
 sky130_fd_sc_hd__o211ai_1 _5982_ (.A1(\sound1.divisor_m[1] ),
    .A2(_2415_),
    .B1(_2416_),
    .C1(_2417_),
    .Y(_2418_));
 sky130_fd_sc_hd__inv_2 _5983_ (.A(\sound1.divisor_m[4] ),
    .Y(_2419_));
 sky130_fd_sc_hd__a22o_1 _5984_ (.A1(\sound1.count_m[3] ),
    .A2(_2419_),
    .B1(\sound1.divisor_m[1] ),
    .B2(_2415_),
    .X(_2420_));
 sky130_fd_sc_hd__a2111o_1 _5985_ (.A1(\sound1.count_m[2] ),
    .A2(_2413_),
    .B1(_2414_),
    .C1(_2418_),
    .D1(_2420_),
    .X(_2421_));
 sky130_fd_sc_hd__nor4_1 _5986_ (.A(_2408_),
    .B(_2411_),
    .C(_2412_),
    .D(_2421_),
    .Y(_2422_));
 sky130_fd_sc_hd__a221o_1 _5987_ (.A1(\sound1.count_m[10] ),
    .A2(_2378_),
    .B1(_2390_),
    .B2(_2391_),
    .C1(_2379_),
    .X(_2423_));
 sky130_fd_sc_hd__a21bo_1 _5988_ (.A1(_2387_),
    .A2(_2423_),
    .B1_N(_2386_),
    .X(_2424_));
 sky130_fd_sc_hd__a21o_1 _5989_ (.A1(_2384_),
    .A2(_2424_),
    .B1(_2377_),
    .X(_2425_));
 sky130_fd_sc_hd__a21o_1 _5990_ (.A1(_2382_),
    .A2(_2425_),
    .B1(_2389_),
    .X(_2426_));
 sky130_fd_sc_hd__a21o_1 _5991_ (.A1(_2400_),
    .A2(_2401_),
    .B1(_2397_),
    .X(_2427_));
 sky130_fd_sc_hd__and2_1 _5992_ (.A(_2402_),
    .B(_2427_),
    .X(_2428_));
 sky130_fd_sc_hd__o2bb2a_1 _5993_ (.A1_N(_2416_),
    .A2_N(_2418_),
    .B1(_2410_),
    .B2(\sound1.divisor_m[3] ),
    .X(_2429_));
 sky130_fd_sc_hd__o221a_1 _5994_ (.A1(_2409_),
    .A2(\sound1.divisor_m[4] ),
    .B1(_2411_),
    .B2(_2429_),
    .C1(_2404_),
    .X(_2430_));
 sky130_fd_sc_hd__o21ai_1 _5995_ (.A1(_2428_),
    .A2(_2430_),
    .B1(_2394_),
    .Y(_2431_));
 sky130_fd_sc_hd__a21o_1 _5996_ (.A1(_2426_),
    .A2(_2431_),
    .B1(_2414_),
    .X(_2432_));
 sky130_fd_sc_hd__a21o_1 _5997_ (.A1(_2407_),
    .A2(_2432_),
    .B1(_2412_),
    .X(_2433_));
 sky130_fd_sc_hd__a31o_2 _5998_ (.A1(_2394_),
    .A2(_2404_),
    .A3(_2422_),
    .B1(_2433_),
    .X(_2434_));
 sky130_fd_sc_hd__inv_2 _5999_ (.A(\sound1.sdiv.Q[1] ),
    .Y(_2435_));
 sky130_fd_sc_hd__nor2_1 _6000_ (.A(_2435_),
    .B(\sound1.sdiv.next_start ),
    .Y(_2436_));
 sky130_fd_sc_hd__a31o_1 _6001_ (.A1(\sound1.sdiv.Q[0] ),
    .A2(_0579_),
    .A3(_2434_),
    .B1(_2436_),
    .X(_2437_));
 sky130_fd_sc_hd__or3b_1 _6002_ (.A(_2435_),
    .B(_2277_),
    .C_N(_2434_),
    .X(_2438_));
 sky130_fd_sc_hd__a32o_1 _6003_ (.A1(_2289_),
    .A2(_2437_),
    .A3(_2438_),
    .B1(_2293_),
    .B2(\sound1.sdiv.Q[2] ),
    .X(_2439_));
 sky130_fd_sc_hd__inv_2 _6004_ (.A(\sound2.divisor_m[15] ),
    .Y(_2440_));
 sky130_fd_sc_hd__inv_2 _6005_ (.A(\sound2.divisor_m[14] ),
    .Y(_2441_));
 sky130_fd_sc_hd__a22o_1 _6006_ (.A1(\sound2.count_m[14] ),
    .A2(_2440_),
    .B1(\sound2.count_m[13] ),
    .B2(_2441_),
    .X(_2442_));
 sky130_fd_sc_hd__inv_2 _6007_ (.A(\sound2.divisor_m[11] ),
    .Y(_2443_));
 sky130_fd_sc_hd__and2b_1 _6008_ (.A_N(\sound2.divisor_m[10] ),
    .B(\sound2.count_m[9] ),
    .X(_2444_));
 sky130_fd_sc_hd__a21o_1 _6009_ (.A1(\sound2.count_m[10] ),
    .A2(_2443_),
    .B1(_2444_),
    .X(_2445_));
 sky130_fd_sc_hd__inv_2 _6010_ (.A(\sound2.divisor_m[16] ),
    .Y(_2446_));
 sky130_fd_sc_hd__o22a_1 _6011_ (.A1(\sound2.count_m[15] ),
    .A2(_2446_),
    .B1(\sound2.count_m[14] ),
    .B2(_2440_),
    .X(_2447_));
 sky130_fd_sc_hd__inv_2 _6012_ (.A(\sound2.divisor_m[13] ),
    .Y(_2448_));
 sky130_fd_sc_hd__o22a_1 _6013_ (.A1(\sound2.count_m[13] ),
    .A2(_2441_),
    .B1(_2448_),
    .B2(\sound2.count_m[12] ),
    .X(_2449_));
 sky130_fd_sc_hd__inv_2 _6014_ (.A(\sound2.count_m[11] ),
    .Y(_2450_));
 sky130_fd_sc_hd__o2bb2a_1 _6015_ (.A1_N(_2448_),
    .A2_N(\sound2.count_m[12] ),
    .B1(_2450_),
    .B2(\sound2.divisor_m[12] ),
    .X(_2451_));
 sky130_fd_sc_hd__o2bb2a_1 _6016_ (.A1_N(_2450_),
    .A2_N(\sound2.divisor_m[12] ),
    .B1(\sound2.count_m[10] ),
    .B2(_2443_),
    .X(_2452_));
 sky130_fd_sc_hd__and4_1 _6017_ (.A(_2447_),
    .B(_2449_),
    .C(_2451_),
    .D(_2452_),
    .X(_2453_));
 sky130_fd_sc_hd__and2_1 _6018_ (.A(\sound2.count_m[15] ),
    .B(_2446_),
    .X(_2454_));
 sky130_fd_sc_hd__or2b_1 _6019_ (.A(\sound2.count_m[8] ),
    .B_N(\sound2.divisor_m[9] ),
    .X(_2455_));
 sky130_fd_sc_hd__or2b_1 _6020_ (.A(\sound2.count_m[9] ),
    .B_N(\sound2.divisor_m[10] ),
    .X(_2456_));
 sky130_fd_sc_hd__or2b_1 _6021_ (.A(\sound2.divisor_m[9] ),
    .B_N(\sound2.count_m[8] ),
    .X(_2457_));
 sky130_fd_sc_hd__and4b_1 _6022_ (.A_N(_2454_),
    .B(_2455_),
    .C(_2456_),
    .D(_2457_),
    .X(_2458_));
 sky130_fd_sc_hd__and4bb_1 _6023_ (.A_N(_2442_),
    .B_N(_2445_),
    .C(_2453_),
    .D(_2458_),
    .X(_2459_));
 sky130_fd_sc_hd__inv_2 _6024_ (.A(\sound2.divisor_m[8] ),
    .Y(_2460_));
 sky130_fd_sc_hd__inv_2 _6025_ (.A(\sound2.count_m[6] ),
    .Y(_2461_));
 sky130_fd_sc_hd__a2bb2o_1 _6026_ (.A1_N(\sound2.count_m[7] ),
    .A2_N(_2460_),
    .B1(_2461_),
    .B2(\sound2.divisor_m[7] ),
    .X(_2462_));
 sky130_fd_sc_hd__inv_2 _6027_ (.A(\sound2.count_m[5] ),
    .Y(_2463_));
 sky130_fd_sc_hd__inv_2 _6028_ (.A(\sound2.count_m[4] ),
    .Y(_2464_));
 sky130_fd_sc_hd__a22o_1 _6029_ (.A1(_2463_),
    .A2(\sound2.divisor_m[6] ),
    .B1(\sound2.divisor_m[5] ),
    .B2(_2464_),
    .X(_2465_));
 sky130_fd_sc_hd__o22a_1 _6030_ (.A1(_2461_),
    .A2(\sound2.divisor_m[7] ),
    .B1(_2463_),
    .B2(\sound2.divisor_m[6] ),
    .X(_2466_));
 sky130_fd_sc_hd__or2b_1 _6031_ (.A(\sound2.divisor_m[8] ),
    .B_N(\sound2.count_m[7] ),
    .X(_2467_));
 sky130_fd_sc_hd__o21a_1 _6032_ (.A1(\sound2.divisor_m[5] ),
    .A2(_2464_),
    .B1(_2467_),
    .X(_2468_));
 sky130_fd_sc_hd__and4bb_1 _6033_ (.A_N(_2462_),
    .B_N(_2465_),
    .C(_2466_),
    .D(_2468_),
    .X(_2469_));
 sky130_fd_sc_hd__inv_2 _6034_ (.A(\sound2.divisor_m[18] ),
    .Y(_2470_));
 sky130_fd_sc_hd__inv_2 _6035_ (.A(\sound2.divisor_m[17] ),
    .Y(_2471_));
 sky130_fd_sc_hd__o22a_1 _6036_ (.A1(\sound2.count_m[17] ),
    .A2(_2470_),
    .B1(\sound2.count_m[16] ),
    .B2(_2471_),
    .X(_2472_));
 sky130_fd_sc_hd__inv_2 _6037_ (.A(_2472_),
    .Y(_2473_));
 sky130_fd_sc_hd__inv_2 _6038_ (.A(\sound2.count_m[3] ),
    .Y(_2474_));
 sky130_fd_sc_hd__inv_2 _6039_ (.A(\sound2.count_m[2] ),
    .Y(_2475_));
 sky130_fd_sc_hd__a22o_1 _6040_ (.A1(_2474_),
    .A2(\sound2.divisor_m[4] ),
    .B1(_2475_),
    .B2(\sound2.divisor_m[3] ),
    .X(_2476_));
 sky130_fd_sc_hd__a21o_1 _6041_ (.A1(\sound2.count_m[17] ),
    .A2(_2470_),
    .B1(\sound2.count_m[18] ),
    .X(_2477_));
 sky130_fd_sc_hd__inv_2 _6042_ (.A(\sound2.divisor_m[3] ),
    .Y(_2478_));
 sky130_fd_sc_hd__and2_1 _6043_ (.A(\sound2.count_m[16] ),
    .B(_2471_),
    .X(_2479_));
 sky130_fd_sc_hd__inv_2 _6044_ (.A(\sound2.count_m[0] ),
    .Y(_2480_));
 sky130_fd_sc_hd__or2b_1 _6045_ (.A(\sound2.count_m[1] ),
    .B_N(\sound2.divisor_m[2] ),
    .X(_2481_));
 sky130_fd_sc_hd__or2b_1 _6046_ (.A(\sound2.divisor_m[2] ),
    .B_N(\sound2.count_m[1] ),
    .X(_2482_));
 sky130_fd_sc_hd__o211ai_1 _6047_ (.A1(\sound2.divisor_m[1] ),
    .A2(_2480_),
    .B1(_2481_),
    .C1(_2482_),
    .Y(_2483_));
 sky130_fd_sc_hd__inv_2 _6048_ (.A(\sound2.divisor_m[4] ),
    .Y(_2484_));
 sky130_fd_sc_hd__a22o_1 _6049_ (.A1(\sound2.count_m[3] ),
    .A2(_2484_),
    .B1(\sound2.divisor_m[1] ),
    .B2(_2480_),
    .X(_2485_));
 sky130_fd_sc_hd__a2111o_1 _6050_ (.A1(\sound2.count_m[2] ),
    .A2(_2478_),
    .B1(_2479_),
    .C1(_2483_),
    .D1(_2485_),
    .X(_2486_));
 sky130_fd_sc_hd__nor4_1 _6051_ (.A(_2473_),
    .B(_2476_),
    .C(_2477_),
    .D(_2486_),
    .Y(_2487_));
 sky130_fd_sc_hd__a221o_1 _6052_ (.A1(\sound2.count_m[10] ),
    .A2(_2443_),
    .B1(_2455_),
    .B2(_2456_),
    .C1(_2444_),
    .X(_2488_));
 sky130_fd_sc_hd__a21bo_1 _6053_ (.A1(_2452_),
    .A2(_2488_),
    .B1_N(_2451_),
    .X(_2489_));
 sky130_fd_sc_hd__a21o_1 _6054_ (.A1(_2449_),
    .A2(_2489_),
    .B1(_2442_),
    .X(_2490_));
 sky130_fd_sc_hd__a21o_1 _6055_ (.A1(_2447_),
    .A2(_2490_),
    .B1(_2454_),
    .X(_2491_));
 sky130_fd_sc_hd__a21o_1 _6056_ (.A1(_2465_),
    .A2(_2466_),
    .B1(_2462_),
    .X(_2492_));
 sky130_fd_sc_hd__and2_1 _6057_ (.A(_2467_),
    .B(_2492_),
    .X(_2493_));
 sky130_fd_sc_hd__o2bb2a_1 _6058_ (.A1_N(_2481_),
    .A2_N(_2483_),
    .B1(_2475_),
    .B2(\sound2.divisor_m[3] ),
    .X(_2494_));
 sky130_fd_sc_hd__o221a_1 _6059_ (.A1(_2474_),
    .A2(\sound2.divisor_m[4] ),
    .B1(_2476_),
    .B2(_2494_),
    .C1(_2469_),
    .X(_2495_));
 sky130_fd_sc_hd__o21ai_1 _6060_ (.A1(_2493_),
    .A2(_2495_),
    .B1(_2459_),
    .Y(_2496_));
 sky130_fd_sc_hd__a21o_1 _6061_ (.A1(_2491_),
    .A2(_2496_),
    .B1(_2479_),
    .X(_2497_));
 sky130_fd_sc_hd__a21o_1 _6062_ (.A1(_2472_),
    .A2(_2497_),
    .B1(_2477_),
    .X(_2498_));
 sky130_fd_sc_hd__a31o_2 _6063_ (.A1(_2459_),
    .A2(_2469_),
    .A3(_2487_),
    .B1(_2498_),
    .X(_2499_));
 sky130_fd_sc_hd__inv_2 _6064_ (.A(\sound2.sdiv.Q[1] ),
    .Y(_2500_));
 sky130_fd_sc_hd__nor2_1 _6065_ (.A(_2500_),
    .B(\sound2.sdiv.next_start ),
    .Y(_2501_));
 sky130_fd_sc_hd__a31o_1 _6066_ (.A1(\sound2.sdiv.Q[0] ),
    .A2(_0578_),
    .A3(_2499_),
    .B1(_2501_),
    .X(_2502_));
 sky130_fd_sc_hd__or3b_1 _6067_ (.A(_2500_),
    .B(_2276_),
    .C_N(_2499_),
    .X(_2503_));
 sky130_fd_sc_hd__a32o_1 _6068_ (.A1(_2289_),
    .A2(_2502_),
    .A3(_2503_),
    .B1(_2295_),
    .B2(\sound2.sdiv.Q[2] ),
    .X(_2504_));
 sky130_fd_sc_hd__xnor2_1 _6069_ (.A(_2439_),
    .B(_2504_),
    .Y(_2505_));
 sky130_fd_sc_hd__a21o_1 _6070_ (.A1(_2281_),
    .A2(_2299_),
    .B1(_2297_),
    .X(_2506_));
 sky130_fd_sc_hd__xnor2_1 _6071_ (.A(_2505_),
    .B(_2506_),
    .Y(_2507_));
 sky130_fd_sc_hd__inv_2 _6072_ (.A(\sound3.count_m[3] ),
    .Y(_2508_));
 sky130_fd_sc_hd__inv_2 _6073_ (.A(\sound3.count_m[2] ),
    .Y(_2509_));
 sky130_fd_sc_hd__a22o_1 _6074_ (.A1(_2508_),
    .A2(\sound3.divisor_m[4] ),
    .B1(_2509_),
    .B2(\sound3.divisor_m[3] ),
    .X(_2510_));
 sky130_fd_sc_hd__inv_2 _6075_ (.A(\sound3.count_m[4] ),
    .Y(_2511_));
 sky130_fd_sc_hd__o22a_1 _6076_ (.A1(\sound3.divisor_m[5] ),
    .A2(_2511_),
    .B1(_2508_),
    .B2(\sound3.divisor_m[4] ),
    .X(_2512_));
 sky130_fd_sc_hd__inv_2 _6077_ (.A(\sound3.count_m[6] ),
    .Y(_2513_));
 sky130_fd_sc_hd__inv_2 _6078_ (.A(\sound3.count_m[5] ),
    .Y(_2514_));
 sky130_fd_sc_hd__o22a_1 _6079_ (.A1(_2513_),
    .A2(\sound3.divisor_m[7] ),
    .B1(_2514_),
    .B2(\sound3.divisor_m[6] ),
    .X(_2515_));
 sky130_fd_sc_hd__nand3b_1 _6080_ (.A_N(_2510_),
    .B(_2512_),
    .C(_2515_),
    .Y(_2516_));
 sky130_fd_sc_hd__inv_2 _6081_ (.A(\sound3.count_m[0] ),
    .Y(_2517_));
 sky130_fd_sc_hd__or2b_1 _6082_ (.A(\sound3.count_m[1] ),
    .B_N(\sound3.divisor_m[2] ),
    .X(_2518_));
 sky130_fd_sc_hd__or2b_1 _6083_ (.A(\sound3.divisor_m[2] ),
    .B_N(\sound3.count_m[1] ),
    .X(_2519_));
 sky130_fd_sc_hd__o211ai_1 _6084_ (.A1(\sound3.divisor_m[1] ),
    .A2(_2517_),
    .B1(_2518_),
    .C1(_2519_),
    .Y(_2520_));
 sky130_fd_sc_hd__inv_2 _6085_ (.A(\sound3.count_m[13] ),
    .Y(_2521_));
 sky130_fd_sc_hd__inv_2 _6086_ (.A(\sound3.count_m[12] ),
    .Y(_2522_));
 sky130_fd_sc_hd__a22o_1 _6087_ (.A1(_2521_),
    .A2(\sound3.divisor_m[14] ),
    .B1(\sound3.divisor_m[13] ),
    .B2(_2522_),
    .X(_2523_));
 sky130_fd_sc_hd__inv_2 _6088_ (.A(\sound3.count_m[11] ),
    .Y(_2524_));
 sky130_fd_sc_hd__inv_2 _6089_ (.A(\sound3.count_m[10] ),
    .Y(_2525_));
 sky130_fd_sc_hd__a22o_1 _6090_ (.A1(_2524_),
    .A2(\sound3.divisor_m[12] ),
    .B1(_2525_),
    .B2(\sound3.divisor_m[11] ),
    .X(_2526_));
 sky130_fd_sc_hd__nor2_1 _6091_ (.A(_2524_),
    .B(\sound3.divisor_m[12] ),
    .Y(_2527_));
 sky130_fd_sc_hd__nor2_1 _6092_ (.A(\sound3.divisor_m[13] ),
    .B(_2522_),
    .Y(_2528_));
 sky130_fd_sc_hd__inv_2 _6093_ (.A(\sound3.divisor_m[15] ),
    .Y(_2529_));
 sky130_fd_sc_hd__a2bb2o_1 _6094_ (.A1_N(\sound3.divisor_m[14] ),
    .A2_N(_2521_),
    .B1(_2529_),
    .B2(\sound3.count_m[14] ),
    .X(_2530_));
 sky130_fd_sc_hd__inv_2 _6095_ (.A(\sound3.count_m[9] ),
    .Y(_2531_));
 sky130_fd_sc_hd__inv_2 _6096_ (.A(\sound3.count_m[8] ),
    .Y(_2532_));
 sky130_fd_sc_hd__a22o_1 _6097_ (.A1(_2531_),
    .A2(\sound3.divisor_m[10] ),
    .B1(\sound3.divisor_m[9] ),
    .B2(_2532_),
    .X(_2533_));
 sky130_fd_sc_hd__and2b_1 _6098_ (.A_N(\sound3.divisor_m[10] ),
    .B(\sound3.count_m[9] ),
    .X(_2534_));
 sky130_fd_sc_hd__and2b_1 _6099_ (.A_N(\sound3.divisor_m[11] ),
    .B(\sound3.count_m[10] ),
    .X(_2535_));
 sky130_fd_sc_hd__or3_1 _6100_ (.A(_2533_),
    .B(_2534_),
    .C(_2535_),
    .X(_2536_));
 sky130_fd_sc_hd__or4_1 _6101_ (.A(_2527_),
    .B(_2528_),
    .C(_2530_),
    .D(_2536_),
    .X(_2537_));
 sky130_fd_sc_hd__inv_2 _6102_ (.A(\sound3.count_m[15] ),
    .Y(_2538_));
 sky130_fd_sc_hd__o2bb2a_1 _6103_ (.A1_N(_2538_),
    .A2_N(\sound3.divisor_m[16] ),
    .B1(\sound3.count_m[14] ),
    .B2(_2529_),
    .X(_2539_));
 sky130_fd_sc_hd__o221a_1 _6104_ (.A1(_2538_),
    .A2(\sound3.divisor_m[16] ),
    .B1(\sound3.divisor_m[9] ),
    .B2(_2532_),
    .C1(_2539_),
    .X(_2540_));
 sky130_fd_sc_hd__nor4b_1 _6105_ (.A(_2523_),
    .B(_2526_),
    .C(_2537_),
    .D_N(_2540_),
    .Y(_2541_));
 sky130_fd_sc_hd__inv_2 _6106_ (.A(net59),
    .Y(_2542_));
 sky130_fd_sc_hd__inv_2 _6107_ (.A(\sound3.divisor_m[18] ),
    .Y(_2543_));
 sky130_fd_sc_hd__a21o_1 _6108_ (.A1(\sound3.count_m[17] ),
    .A2(_2543_),
    .B1(\sound3.count_m[18] ),
    .X(_2544_));
 sky130_fd_sc_hd__inv_2 _6109_ (.A(\sound3.count_m[16] ),
    .Y(_2545_));
 sky130_fd_sc_hd__a2bb2o_1 _6110_ (.A1_N(\sound3.count_m[17] ),
    .A2_N(_2543_),
    .B1(_2545_),
    .B2(\sound3.divisor_m[17] ),
    .X(_2546_));
 sky130_fd_sc_hd__inv_2 _6111_ (.A(\sound3.count_m[7] ),
    .Y(_2547_));
 sky130_fd_sc_hd__a22o_1 _6112_ (.A1(_2547_),
    .A2(\sound3.divisor_m[8] ),
    .B1(_2513_),
    .B2(\sound3.divisor_m[7] ),
    .X(_2548_));
 sky130_fd_sc_hd__a22o_1 _6113_ (.A1(_2514_),
    .A2(\sound3.divisor_m[6] ),
    .B1(\sound3.divisor_m[5] ),
    .B2(_2511_),
    .X(_2549_));
 sky130_fd_sc_hd__or4_1 _6114_ (.A(_2544_),
    .B(_2546_),
    .C(_2548_),
    .D(_2549_),
    .X(_2550_));
 sky130_fd_sc_hd__inv_2 _6115_ (.A(\sound3.divisor_m[1] ),
    .Y(_2551_));
 sky130_fd_sc_hd__or2_1 _6116_ (.A(_2545_),
    .B(\sound3.divisor_m[17] ),
    .X(_2552_));
 sky130_fd_sc_hd__or2_1 _6117_ (.A(_2509_),
    .B(\sound3.divisor_m[3] ),
    .X(_2553_));
 sky130_fd_sc_hd__or2_1 _6118_ (.A(_2547_),
    .B(\sound3.divisor_m[8] ),
    .X(_2554_));
 sky130_fd_sc_hd__o2111a_1 _6119_ (.A1(_2551_),
    .A2(\sound3.count_m[0] ),
    .B1(_2552_),
    .C1(_2553_),
    .D1(_2554_),
    .X(_2555_));
 sky130_fd_sc_hd__or4b_1 _6120_ (.A(_2520_),
    .B(_2542_),
    .C(_2550_),
    .D_N(_2555_),
    .X(_2556_));
 sky130_fd_sc_hd__nand2_1 _6121_ (.A(_2518_),
    .B(_2520_),
    .Y(_2557_));
 sky130_fd_sc_hd__a21o_1 _6122_ (.A1(_2553_),
    .A2(_2557_),
    .B1(_2510_),
    .X(_2558_));
 sky130_fd_sc_hd__a21o_1 _6123_ (.A1(_2558_),
    .A2(_2512_),
    .B1(_2549_),
    .X(_2559_));
 sky130_fd_sc_hd__a21o_1 _6124_ (.A1(_2559_),
    .A2(_2515_),
    .B1(_2548_),
    .X(_2560_));
 sky130_fd_sc_hd__nor2_1 _6125_ (.A(_2534_),
    .B(_2535_),
    .Y(_2561_));
 sky130_fd_sc_hd__a21oi_1 _6126_ (.A1(_2533_),
    .A2(_2561_),
    .B1(_2526_),
    .Y(_2562_));
 sky130_fd_sc_hd__inv_2 _6127_ (.A(_2523_),
    .Y(_2563_));
 sky130_fd_sc_hd__o31a_1 _6128_ (.A1(_2562_),
    .A2(_2527_),
    .A3(_2528_),
    .B1(_2563_),
    .X(_2564_));
 sky130_fd_sc_hd__or2_1 _6129_ (.A(_2564_),
    .B(_2530_),
    .X(_2565_));
 sky130_fd_sc_hd__o2bb2a_1 _6130_ (.A1_N(_2565_),
    .A2_N(_2539_),
    .B1(\sound3.divisor_m[16] ),
    .B2(_2538_),
    .X(_2566_));
 sky130_fd_sc_hd__a31o_1 _6131_ (.A1(_2560_),
    .A2(net60),
    .A3(_2554_),
    .B1(_2566_),
    .X(_2567_));
 sky130_fd_sc_hd__a21oi_1 _6132_ (.A1(_2552_),
    .A2(_2567_),
    .B1(_2546_),
    .Y(_2568_));
 sky130_fd_sc_hd__nor2_1 _6133_ (.A(_2544_),
    .B(_2568_),
    .Y(_2569_));
 sky130_fd_sc_hd__o21a_1 _6134_ (.A1(_2516_),
    .A2(_2556_),
    .B1(_2569_),
    .X(_2570_));
 sky130_fd_sc_hd__a2bb2o_1 _6135_ (.A1_N(_2275_),
    .A2_N(_2570_),
    .B1(\sound3.sdiv.Q[1] ),
    .B2(_0577_),
    .X(_2571_));
 sky130_fd_sc_hd__or3b_1 _6136_ (.A(_2570_),
    .B(_2275_),
    .C_N(\sound3.sdiv.Q[1] ),
    .X(_2572_));
 sky130_fd_sc_hd__a32o_1 _6137_ (.A1(_2289_),
    .A2(_2571_),
    .A3(_2572_),
    .B1(_2301_),
    .B2(\sound3.sdiv.Q[2] ),
    .X(_2573_));
 sky130_fd_sc_hd__xor2_1 _6138_ (.A(_2507_),
    .B(_2573_),
    .X(_2574_));
 sky130_fd_sc_hd__xnor2_1 _6139_ (.A(_2374_),
    .B(_2574_),
    .Y(_2575_));
 sky130_fd_sc_hd__a21oi_1 _6140_ (.A1(_2291_),
    .A2(_2305_),
    .B1(_2303_),
    .Y(_2576_));
 sky130_fd_sc_hd__xnor2_1 _6141_ (.A(_2575_),
    .B(_2576_),
    .Y(_2577_));
 sky130_fd_sc_hd__or2_1 _6142_ (.A(_2311_),
    .B(_2577_),
    .X(_2578_));
 sky130_fd_sc_hd__a21oi_1 _6143_ (.A1(_2311_),
    .A2(_2577_),
    .B1(_0569_),
    .Y(_2579_));
 sky130_fd_sc_hd__a22o_1 _6144_ (.A1(\wave_comb.u1.Q[1] ),
    .A2(_0569_),
    .B1(_2578_),
    .B2(_2579_),
    .X(_2580_));
 sky130_fd_sc_hd__and3_1 _6145_ (.A(\wave_comb.u1.Q[2] ),
    .B(_0569_),
    .C(_0571_),
    .X(_2581_));
 sky130_fd_sc_hd__a21o_1 _6146_ (.A1(\wave_comb.u1.next_start ),
    .A2(_2580_),
    .B1(_2581_),
    .X(_0047_));
 sky130_fd_sc_hd__o211a_1 _6147_ (.A1(\sound4.sdiv.Q[0] ),
    .A2(\sound4.sdiv.Q[1] ),
    .B1(_0576_),
    .C1(_2370_),
    .X(_2582_));
 sky130_fd_sc_hd__nand2_1 _6148_ (.A(\sound4.sdiv.Q[2] ),
    .B(_2582_),
    .Y(_2583_));
 sky130_fd_sc_hd__a21o_1 _6149_ (.A1(\sound4.sdiv.Q[2] ),
    .A2(_0576_),
    .B1(_2582_),
    .X(_2584_));
 sky130_fd_sc_hd__a32o_1 _6150_ (.A1(_2289_),
    .A2(_2583_),
    .A3(_2584_),
    .B1(_2290_),
    .B2(\sound4.sdiv.Q[3] ),
    .X(_2585_));
 sky130_fd_sc_hd__nand2_1 _6151_ (.A(\sound1.sdiv.Q[3] ),
    .B(_0579_),
    .Y(_2586_));
 sky130_fd_sc_hd__o211a_1 _6152_ (.A1(\sound1.sdiv.Q[0] ),
    .A2(\sound1.sdiv.Q[1] ),
    .B1(_0579_),
    .C1(_2434_),
    .X(_2587_));
 sky130_fd_sc_hd__nand2_1 _6153_ (.A(\sound1.sdiv.Q[2] ),
    .B(_0579_),
    .Y(_2588_));
 sky130_fd_sc_hd__xnor2_1 _6154_ (.A(_2587_),
    .B(_2588_),
    .Y(_2589_));
 sky130_fd_sc_hd__a2bb2o_2 _6155_ (.A1_N(_2279_),
    .A2_N(_2586_),
    .B1(_2589_),
    .B2(_2289_),
    .X(_2590_));
 sky130_fd_sc_hd__o211a_1 _6156_ (.A1(\sound2.sdiv.Q[0] ),
    .A2(\sound2.sdiv.Q[1] ),
    .B1(_0578_),
    .C1(_2499_),
    .X(_2591_));
 sky130_fd_sc_hd__and3_1 _6157_ (.A(\sound2.sdiv.Q[2] ),
    .B(_0578_),
    .C(_2591_),
    .X(_2592_));
 sky130_fd_sc_hd__a21oi_2 _6158_ (.A1(\sound2.sdiv.Q[2] ),
    .A2(_0578_),
    .B1(_2591_),
    .Y(_2593_));
 sky130_fd_sc_hd__nand2_1 _6159_ (.A(\sound2.sdiv.Q[3] ),
    .B(_0578_),
    .Y(_2594_));
 sky130_fd_sc_hd__o32ai_4 _6160_ (.A1(_2292_),
    .A2(_2592_),
    .A3(_2593_),
    .B1(_2594_),
    .B2(_2279_),
    .Y(_2595_));
 sky130_fd_sc_hd__xor2_1 _6161_ (.A(_2590_),
    .B(_2595_),
    .X(_2596_));
 sky130_fd_sc_hd__or2_1 _6162_ (.A(_2439_),
    .B(_2504_),
    .X(_2597_));
 sky130_fd_sc_hd__and2_1 _6163_ (.A(_2439_),
    .B(_2504_),
    .X(_2598_));
 sky130_fd_sc_hd__a21oi_1 _6164_ (.A1(_2597_),
    .A2(_2506_),
    .B1(_2598_),
    .Y(_2599_));
 sky130_fd_sc_hd__xnor2_1 _6165_ (.A(_2596_),
    .B(_2599_),
    .Y(_2600_));
 sky130_fd_sc_hd__o21ai_1 _6166_ (.A1(\sound3.sdiv.Q[0] ),
    .A2(\sound3.sdiv.Q[1] ),
    .B1(_0577_),
    .Y(_2601_));
 sky130_fd_sc_hd__nor2_1 _6167_ (.A(_2570_),
    .B(_2601_),
    .Y(_2602_));
 sky130_fd_sc_hd__a21oi_1 _6168_ (.A1(\sound3.sdiv.Q[2] ),
    .A2(_0577_),
    .B1(_2602_),
    .Y(_2603_));
 sky130_fd_sc_hd__a21o_1 _6169_ (.A1(\sound3.sdiv.Q[2] ),
    .A2(_2602_),
    .B1(_2292_),
    .X(_2604_));
 sky130_fd_sc_hd__o2bb2a_1 _6170_ (.A1_N(\sound3.sdiv.Q[3] ),
    .A2_N(_2301_),
    .B1(_2603_),
    .B2(_2604_),
    .X(_2605_));
 sky130_fd_sc_hd__xnor2_1 _6171_ (.A(_2600_),
    .B(_2605_),
    .Y(_2606_));
 sky130_fd_sc_hd__xnor2_1 _6172_ (.A(_2585_),
    .B(_2606_),
    .Y(_2607_));
 sky130_fd_sc_hd__and2_1 _6173_ (.A(_2507_),
    .B(_2573_),
    .X(_2608_));
 sky130_fd_sc_hd__a21o_1 _6174_ (.A1(_2374_),
    .A2(_2574_),
    .B1(_2608_),
    .X(_2609_));
 sky130_fd_sc_hd__xnor2_1 _6175_ (.A(_2607_),
    .B(_2609_),
    .Y(_2610_));
 sky130_fd_sc_hd__or2_1 _6176_ (.A(_2575_),
    .B(_2576_),
    .X(_2611_));
 sky130_fd_sc_hd__o21ai_2 _6177_ (.A1(_2311_),
    .A2(_2577_),
    .B1(_2611_),
    .Y(_2612_));
 sky130_fd_sc_hd__nor2_1 _6178_ (.A(_2610_),
    .B(_2612_),
    .Y(_2613_));
 sky130_fd_sc_hd__a21o_1 _6179_ (.A1(_2610_),
    .A2(_2612_),
    .B1(_0569_),
    .X(_2614_));
 sky130_fd_sc_hd__a2bb2o_1 _6180_ (.A1_N(_2613_),
    .A2_N(_2614_),
    .B1(\wave_comb.u1.Q[2] ),
    .B2(_0569_),
    .X(_2615_));
 sky130_fd_sc_hd__and3_1 _6181_ (.A(\wave_comb.u1.Q[3] ),
    .B(_0569_),
    .C(_0571_),
    .X(_2616_));
 sky130_fd_sc_hd__a21o_1 _6182_ (.A1(\wave_comb.u1.next_start ),
    .A2(_2615_),
    .B1(_2616_),
    .X(_0048_));
 sky130_fd_sc_hd__nor2_1 _6183_ (.A(_2590_),
    .B(_2595_),
    .Y(_2617_));
 sky130_fd_sc_hd__nand2_1 _6184_ (.A(_2590_),
    .B(_2595_),
    .Y(_2618_));
 sky130_fd_sc_hd__o21ai_1 _6185_ (.A1(_2617_),
    .A2(_2599_),
    .B1(_2618_),
    .Y(_2619_));
 sky130_fd_sc_hd__nand2_1 _6186_ (.A(\sound1.sdiv.Q[4] ),
    .B(_0579_),
    .Y(_2620_));
 sky130_fd_sc_hd__o311a_1 _6187_ (.A1(\sound1.sdiv.Q[0] ),
    .A2(\sound1.sdiv.Q[1] ),
    .A3(\sound1.sdiv.Q[2] ),
    .B1(_0579_),
    .C1(_2434_),
    .X(_2621_));
 sky130_fd_sc_hd__xor2_1 _6188_ (.A(_2586_),
    .B(_2621_),
    .X(_2622_));
 sky130_fd_sc_hd__o22a_1 _6189_ (.A1(_2279_),
    .A2(_2620_),
    .B1(_2622_),
    .B2(_2292_),
    .X(_2623_));
 sky130_fd_sc_hd__nand2_1 _6190_ (.A(\sound2.sdiv.Q[4] ),
    .B(_0578_),
    .Y(_2624_));
 sky130_fd_sc_hd__o311a_1 _6191_ (.A1(\sound2.sdiv.Q[0] ),
    .A2(\sound2.sdiv.Q[1] ),
    .A3(\sound2.sdiv.Q[2] ),
    .B1(_0578_),
    .C1(_2499_),
    .X(_2625_));
 sky130_fd_sc_hd__xor2_1 _6192_ (.A(_2594_),
    .B(_2625_),
    .X(_2626_));
 sky130_fd_sc_hd__o22a_1 _6193_ (.A1(_2279_),
    .A2(_2624_),
    .B1(_2626_),
    .B2(_2292_),
    .X(_2627_));
 sky130_fd_sc_hd__nor2_1 _6194_ (.A(_2623_),
    .B(_2627_),
    .Y(_2628_));
 sky130_fd_sc_hd__nand2_1 _6195_ (.A(_2623_),
    .B(_2627_),
    .Y(_2629_));
 sky130_fd_sc_hd__and2b_1 _6196_ (.A_N(_2628_),
    .B(_2629_),
    .X(_2630_));
 sky130_fd_sc_hd__xnor2_1 _6197_ (.A(_2619_),
    .B(_2630_),
    .Y(_2631_));
 sky130_fd_sc_hd__nor2_1 _6198_ (.A(\sound3.sdiv.next_start ),
    .B(_2570_),
    .Y(_2632_));
 sky130_fd_sc_hd__a21o_1 _6199_ (.A1(\sound3.sdiv.Q[2] ),
    .A2(_2632_),
    .B1(_2602_),
    .X(_2633_));
 sky130_fd_sc_hd__and3_1 _6200_ (.A(\sound3.sdiv.Q[3] ),
    .B(_0577_),
    .C(_2633_),
    .X(_2634_));
 sky130_fd_sc_hd__a21oi_1 _6201_ (.A1(\sound3.sdiv.Q[3] ),
    .A2(_0577_),
    .B1(_2633_),
    .Y(_2635_));
 sky130_fd_sc_hd__nand2_1 _6202_ (.A(\sound3.sdiv.Q[4] ),
    .B(_0577_),
    .Y(_2636_));
 sky130_fd_sc_hd__o32a_1 _6203_ (.A1(_2292_),
    .A2(_2634_),
    .A3(_2635_),
    .B1(_2636_),
    .B2(_2279_),
    .X(_2637_));
 sky130_fd_sc_hd__xnor2_1 _6204_ (.A(_2631_),
    .B(_2637_),
    .Y(_2638_));
 sky130_fd_sc_hd__nand2_1 _6205_ (.A(\sound4.sdiv.Q[4] ),
    .B(_0576_),
    .Y(_2639_));
 sky130_fd_sc_hd__nand2_1 _6206_ (.A(\sound4.sdiv.Q[3] ),
    .B(_0576_),
    .Y(_2640_));
 sky130_fd_sc_hd__and2_1 _6207_ (.A(_0576_),
    .B(_2370_),
    .X(_2641_));
 sky130_fd_sc_hd__a21o_1 _6208_ (.A1(\sound4.sdiv.Q[2] ),
    .A2(_2641_),
    .B1(_2582_),
    .X(_2642_));
 sky130_fd_sc_hd__xor2_1 _6209_ (.A(_2640_),
    .B(_2642_),
    .X(_2643_));
 sky130_fd_sc_hd__o22a_1 _6210_ (.A1(_2639_),
    .A2(_2279_),
    .B1(_2292_),
    .B2(_2643_),
    .X(_2644_));
 sky130_fd_sc_hd__xnor2_1 _6211_ (.A(_2638_),
    .B(_2644_),
    .Y(_2645_));
 sky130_fd_sc_hd__and2b_1 _6212_ (.A_N(_2605_),
    .B(_2600_),
    .X(_2646_));
 sky130_fd_sc_hd__a21oi_1 _6213_ (.A1(_2585_),
    .A2(_2606_),
    .B1(_2646_),
    .Y(_2647_));
 sky130_fd_sc_hd__nor2_1 _6214_ (.A(_2645_),
    .B(_2647_),
    .Y(_2648_));
 sky130_fd_sc_hd__nand2_1 _6215_ (.A(_2645_),
    .B(_2647_),
    .Y(_2649_));
 sky130_fd_sc_hd__or2b_1 _6216_ (.A(_2648_),
    .B_N(_2649_),
    .X(_2650_));
 sky130_fd_sc_hd__or2b_1 _6217_ (.A(_2607_),
    .B_N(_2609_),
    .X(_2651_));
 sky130_fd_sc_hd__a21bo_1 _6218_ (.A1(_2610_),
    .A2(_2612_),
    .B1_N(_2651_),
    .X(_2652_));
 sky130_fd_sc_hd__xnor2_1 _6219_ (.A(_2650_),
    .B(_2652_),
    .Y(_2653_));
 sky130_fd_sc_hd__mux2_1 _6220_ (.A0(\wave_comb.u1.Q[3] ),
    .A1(_2653_),
    .S(_0645_),
    .X(_2654_));
 sky130_fd_sc_hd__nand2_1 _6221_ (.A(\wave_comb.u1.Q[4] ),
    .B(_0573_),
    .Y(_2655_));
 sky130_fd_sc_hd__a21bo_1 _6222_ (.A1(\wave_comb.u1.next_start ),
    .A2(_2654_),
    .B1_N(_2655_),
    .X(_0049_));
 sky130_fd_sc_hd__and2_1 _6223_ (.A(_0579_),
    .B(_2434_),
    .X(_2656_));
 sky130_fd_sc_hd__a21oi_1 _6224_ (.A1(\sound1.sdiv.Q[3] ),
    .A2(_2656_),
    .B1(_2621_),
    .Y(_2657_));
 sky130_fd_sc_hd__xnor2_1 _6225_ (.A(_2620_),
    .B(_2657_),
    .Y(_2658_));
 sky130_fd_sc_hd__o2bb2a_1 _6226_ (.A1_N(\sound1.sdiv.Q[5] ),
    .A2_N(_2293_),
    .B1(_2658_),
    .B2(_2292_),
    .X(_2659_));
 sky130_fd_sc_hd__and2_1 _6227_ (.A(_0578_),
    .B(_2499_),
    .X(_2660_));
 sky130_fd_sc_hd__a21oi_1 _6228_ (.A1(\sound2.sdiv.Q[3] ),
    .A2(_2660_),
    .B1(_2625_),
    .Y(_2661_));
 sky130_fd_sc_hd__xnor2_1 _6229_ (.A(_2624_),
    .B(_2661_),
    .Y(_2662_));
 sky130_fd_sc_hd__o2bb2a_1 _6230_ (.A1_N(\sound2.sdiv.Q[5] ),
    .A2_N(_2295_),
    .B1(_2662_),
    .B2(_2292_),
    .X(_2663_));
 sky130_fd_sc_hd__nor2_1 _6231_ (.A(_2659_),
    .B(_2663_),
    .Y(_2664_));
 sky130_fd_sc_hd__nand2_1 _6232_ (.A(_2659_),
    .B(_2663_),
    .Y(_2665_));
 sky130_fd_sc_hd__and2b_1 _6233_ (.A_N(_2664_),
    .B(_2665_),
    .X(_2666_));
 sky130_fd_sc_hd__a21o_1 _6234_ (.A1(_2619_),
    .A2(_2629_),
    .B1(_2628_),
    .X(_2667_));
 sky130_fd_sc_hd__xnor2_1 _6235_ (.A(_2666_),
    .B(_2667_),
    .Y(_2668_));
 sky130_fd_sc_hd__a21o_1 _6236_ (.A1(\sound3.sdiv.Q[3] ),
    .A2(_2632_),
    .B1(_2633_),
    .X(_2669_));
 sky130_fd_sc_hd__xor2_1 _6237_ (.A(_2636_),
    .B(_2669_),
    .X(_2670_));
 sky130_fd_sc_hd__o2bb2a_1 _6238_ (.A1_N(\sound3.sdiv.Q[5] ),
    .A2_N(_2301_),
    .B1(_2670_),
    .B2(_2292_),
    .X(_2671_));
 sky130_fd_sc_hd__xnor2_1 _6239_ (.A(_2668_),
    .B(_2671_),
    .Y(_2672_));
 sky130_fd_sc_hd__a21o_1 _6240_ (.A1(\sound4.sdiv.Q[3] ),
    .A2(_2641_),
    .B1(_2642_),
    .X(_2673_));
 sky130_fd_sc_hd__xor2_1 _6241_ (.A(_2639_),
    .B(_2673_),
    .X(_2674_));
 sky130_fd_sc_hd__o2bb2a_1 _6242_ (.A1_N(\sound4.sdiv.Q[5] ),
    .A2_N(_2290_),
    .B1(_2674_),
    .B2(_2292_),
    .X(_2675_));
 sky130_fd_sc_hd__xnor2_1 _6243_ (.A(_2672_),
    .B(_2675_),
    .Y(_2676_));
 sky130_fd_sc_hd__o22ai_2 _6244_ (.A1(_2631_),
    .A2(_2637_),
    .B1(_2638_),
    .B2(_2644_),
    .Y(_2677_));
 sky130_fd_sc_hd__xor2_1 _6245_ (.A(_2676_),
    .B(_2677_),
    .X(_2678_));
 sky130_fd_sc_hd__a21oi_1 _6246_ (.A1(_2649_),
    .A2(_2652_),
    .B1(_2648_),
    .Y(_2679_));
 sky130_fd_sc_hd__xor2_1 _6247_ (.A(_2678_),
    .B(_2679_),
    .X(_2680_));
 sky130_fd_sc_hd__mux2_1 _6248_ (.A0(\wave_comb.u1.Q[4] ),
    .A1(_2680_),
    .S(_0645_),
    .X(_2681_));
 sky130_fd_sc_hd__nand2_1 _6249_ (.A(\wave_comb.u1.Q[5] ),
    .B(_0572_),
    .Y(_2682_));
 sky130_fd_sc_hd__a21bo_1 _6250_ (.A1(\wave_comb.u1.next_start ),
    .A2(_2681_),
    .B1_N(_2682_),
    .X(_0050_));
 sky130_fd_sc_hd__or2b_1 _6251_ (.A(_2676_),
    .B_N(_2677_),
    .X(_2683_));
 sky130_fd_sc_hd__o21ai_1 _6252_ (.A1(_2678_),
    .A2(_2679_),
    .B1(_2683_),
    .Y(_2684_));
 sky130_fd_sc_hd__nand2_1 _6253_ (.A(\sound2.sdiv.Q[6] ),
    .B(_2295_),
    .Y(_2685_));
 sky130_fd_sc_hd__a21bo_1 _6254_ (.A1(\sound2.sdiv.Q[4] ),
    .A2(_2660_),
    .B1_N(_2661_),
    .X(_2686_));
 sky130_fd_sc_hd__a21o_1 _6255_ (.A1(\sound2.sdiv.Q[5] ),
    .A2(_0578_),
    .B1(_2686_),
    .X(_2687_));
 sky130_fd_sc_hd__a21oi_1 _6256_ (.A1(\sound2.sdiv.Q[5] ),
    .A2(_2686_),
    .B1(_2292_),
    .Y(_2688_));
 sky130_fd_sc_hd__nand2_1 _6257_ (.A(_2687_),
    .B(_2688_),
    .Y(_2689_));
 sky130_fd_sc_hd__a21bo_1 _6258_ (.A1(\sound1.sdiv.Q[4] ),
    .A2(_2656_),
    .B1_N(_2657_),
    .X(_2690_));
 sky130_fd_sc_hd__nand2_1 _6259_ (.A(\sound1.sdiv.Q[5] ),
    .B(_2690_),
    .Y(_2691_));
 sky130_fd_sc_hd__a21o_1 _6260_ (.A1(\sound1.sdiv.Q[5] ),
    .A2(_0579_),
    .B1(_2690_),
    .X(_2692_));
 sky130_fd_sc_hd__a32o_1 _6261_ (.A1(_2289_),
    .A2(_2691_),
    .A3(_2692_),
    .B1(_2293_),
    .B2(\sound1.sdiv.Q[6] ),
    .X(_2693_));
 sky130_fd_sc_hd__a21boi_1 _6262_ (.A1(_2685_),
    .A2(_2689_),
    .B1_N(_2693_),
    .Y(_2694_));
 sky130_fd_sc_hd__nand3b_1 _6263_ (.A_N(_2693_),
    .B(_2685_),
    .C(_2689_),
    .Y(_2695_));
 sky130_fd_sc_hd__and2b_1 _6264_ (.A_N(_2694_),
    .B(_2695_),
    .X(_2696_));
 sky130_fd_sc_hd__a21o_1 _6265_ (.A1(_2665_),
    .A2(_2667_),
    .B1(_2664_),
    .X(_2697_));
 sky130_fd_sc_hd__xor2_1 _6266_ (.A(_2696_),
    .B(_2697_),
    .X(_2698_));
 sky130_fd_sc_hd__a21o_1 _6267_ (.A1(\sound3.sdiv.Q[4] ),
    .A2(_2632_),
    .B1(_2669_),
    .X(_2699_));
 sky130_fd_sc_hd__nand2_1 _6268_ (.A(\sound3.sdiv.Q[5] ),
    .B(_2699_),
    .Y(_2700_));
 sky130_fd_sc_hd__a21o_1 _6269_ (.A1(\sound3.sdiv.Q[5] ),
    .A2(_0577_),
    .B1(_2699_),
    .X(_2701_));
 sky130_fd_sc_hd__a32o_1 _6270_ (.A1(_2289_),
    .A2(_2700_),
    .A3(_2701_),
    .B1(_2301_),
    .B2(\sound3.sdiv.Q[6] ),
    .X(_2702_));
 sky130_fd_sc_hd__xor2_1 _6271_ (.A(_2698_),
    .B(_2702_),
    .X(_2703_));
 sky130_fd_sc_hd__a21o_1 _6272_ (.A1(\sound4.sdiv.Q[4] ),
    .A2(_2641_),
    .B1(_2673_),
    .X(_2704_));
 sky130_fd_sc_hd__a21o_1 _6273_ (.A1(\sound4.sdiv.Q[5] ),
    .A2(_0576_),
    .B1(_2704_),
    .X(_2705_));
 sky130_fd_sc_hd__nand2_1 _6274_ (.A(\sound4.sdiv.Q[5] ),
    .B(_2704_),
    .Y(_2706_));
 sky130_fd_sc_hd__a32o_1 _6275_ (.A1(_2289_),
    .A2(_2705_),
    .A3(_2706_),
    .B1(_2290_),
    .B2(\sound4.sdiv.Q[6] ),
    .X(_2707_));
 sky130_fd_sc_hd__xor2_1 _6276_ (.A(_2703_),
    .B(_2707_),
    .X(_2708_));
 sky130_fd_sc_hd__or2_1 _6277_ (.A(_2668_),
    .B(_2671_),
    .X(_2709_));
 sky130_fd_sc_hd__o21a_1 _6278_ (.A1(_2672_),
    .A2(_2675_),
    .B1(_2709_),
    .X(_2710_));
 sky130_fd_sc_hd__xnor2_1 _6279_ (.A(_2708_),
    .B(_2710_),
    .Y(_2711_));
 sky130_fd_sc_hd__nand2_1 _6280_ (.A(_2684_),
    .B(_2711_),
    .Y(_2712_));
 sky130_fd_sc_hd__or2_1 _6281_ (.A(_2684_),
    .B(_2711_),
    .X(_2713_));
 sky130_fd_sc_hd__a21o_1 _6282_ (.A1(_2712_),
    .A2(_2713_),
    .B1(_0569_),
    .X(_2714_));
 sky130_fd_sc_hd__or2_1 _6283_ (.A(\wave_comb.u1.Q[5] ),
    .B(_0645_),
    .X(_2715_));
 sky130_fd_sc_hd__and3_1 _6284_ (.A(\wave_comb.u1.Q[6] ),
    .B(_0569_),
    .C(_0571_),
    .X(_2716_));
 sky130_fd_sc_hd__a31o_1 _6285_ (.A1(\wave_comb.u1.next_start ),
    .A2(_2714_),
    .A3(_2715_),
    .B1(_2716_),
    .X(_0051_));
 sky130_fd_sc_hd__and3_1 _6286_ (.A(\sound2.sdiv.Q[7] ),
    .B(_0578_),
    .C(_2286_),
    .X(_2717_));
 sky130_fd_sc_hd__a21o_1 _6287_ (.A1(\sound2.sdiv.Q[5] ),
    .A2(_2660_),
    .B1(_2686_),
    .X(_2718_));
 sky130_fd_sc_hd__nand2_1 _6288_ (.A(\sound2.sdiv.Q[6] ),
    .B(_2718_),
    .Y(_2719_));
 sky130_fd_sc_hd__a21o_1 _6289_ (.A1(\sound2.sdiv.Q[6] ),
    .A2(_0578_),
    .B1(_2718_),
    .X(_2720_));
 sky130_fd_sc_hd__and3_1 _6290_ (.A(_2289_),
    .B(_2719_),
    .C(_2720_),
    .X(_2721_));
 sky130_fd_sc_hd__a21o_1 _6291_ (.A1(\sound1.sdiv.Q[5] ),
    .A2(_2656_),
    .B1(_2690_),
    .X(_2722_));
 sky130_fd_sc_hd__nand2_1 _6292_ (.A(\sound1.sdiv.Q[6] ),
    .B(_2722_),
    .Y(_2723_));
 sky130_fd_sc_hd__a21o_1 _6293_ (.A1(\sound1.sdiv.Q[6] ),
    .A2(_0579_),
    .B1(_2722_),
    .X(_2724_));
 sky130_fd_sc_hd__a32o_1 _6294_ (.A1(_2289_),
    .A2(_2723_),
    .A3(_2724_),
    .B1(_2293_),
    .B2(\sound1.sdiv.Q[7] ),
    .X(_2725_));
 sky130_fd_sc_hd__o21ai_1 _6295_ (.A1(_2717_),
    .A2(_2721_),
    .B1(_2725_),
    .Y(_2726_));
 sky130_fd_sc_hd__or3_1 _6296_ (.A(_2725_),
    .B(_2717_),
    .C(_2721_),
    .X(_2727_));
 sky130_fd_sc_hd__nand2_1 _6297_ (.A(_2726_),
    .B(_2727_),
    .Y(_2728_));
 sky130_fd_sc_hd__a21oi_2 _6298_ (.A1(_2695_),
    .A2(_2697_),
    .B1(_2694_),
    .Y(_2729_));
 sky130_fd_sc_hd__xnor2_2 _6299_ (.A(_2728_),
    .B(_2729_),
    .Y(_2730_));
 sky130_fd_sc_hd__a21o_1 _6300_ (.A1(\sound3.sdiv.Q[5] ),
    .A2(_2632_),
    .B1(_2699_),
    .X(_2731_));
 sky130_fd_sc_hd__a21oi_1 _6301_ (.A1(\sound3.sdiv.Q[6] ),
    .A2(_0577_),
    .B1(_2731_),
    .Y(_2732_));
 sky130_fd_sc_hd__a21o_1 _6302_ (.A1(\sound3.sdiv.Q[6] ),
    .A2(_2731_),
    .B1(_2292_),
    .X(_2733_));
 sky130_fd_sc_hd__o2bb2a_1 _6303_ (.A1_N(\sound3.sdiv.Q[7] ),
    .A2_N(_2301_),
    .B1(_2732_),
    .B2(_2733_),
    .X(_2734_));
 sky130_fd_sc_hd__xor2_1 _6304_ (.A(_2730_),
    .B(_2734_),
    .X(_2735_));
 sky130_fd_sc_hd__a21o_1 _6305_ (.A1(\sound4.sdiv.Q[5] ),
    .A2(_2641_),
    .B1(_2704_),
    .X(_2736_));
 sky130_fd_sc_hd__a21o_1 _6306_ (.A1(\sound4.sdiv.Q[6] ),
    .A2(_0576_),
    .B1(_2736_),
    .X(_2737_));
 sky130_fd_sc_hd__nand2_1 _6307_ (.A(\sound4.sdiv.Q[6] ),
    .B(_2736_),
    .Y(_2738_));
 sky130_fd_sc_hd__a32o_1 _6308_ (.A1(_2289_),
    .A2(_2737_),
    .A3(_2738_),
    .B1(_2290_),
    .B2(\sound4.sdiv.Q[7] ),
    .X(_2739_));
 sky130_fd_sc_hd__xnor2_1 _6309_ (.A(_2735_),
    .B(_2739_),
    .Y(_2740_));
 sky130_fd_sc_hd__and2_1 _6310_ (.A(_2698_),
    .B(_2702_),
    .X(_2741_));
 sky130_fd_sc_hd__a21o_1 _6311_ (.A1(_2703_),
    .A2(_2707_),
    .B1(_2741_),
    .X(_2742_));
 sky130_fd_sc_hd__xor2_1 _6312_ (.A(_2740_),
    .B(_2742_),
    .X(_2743_));
 sky130_fd_sc_hd__and2b_1 _6313_ (.A_N(_2710_),
    .B(_2708_),
    .X(_2744_));
 sky130_fd_sc_hd__a21o_1 _6314_ (.A1(_2684_),
    .A2(_2711_),
    .B1(_2744_),
    .X(_2745_));
 sky130_fd_sc_hd__xnor2_1 _6315_ (.A(_2743_),
    .B(_2745_),
    .Y(_2746_));
 sky130_fd_sc_hd__mux2_1 _6316_ (.A0(\wave_comb.u1.Q[6] ),
    .A1(_2746_),
    .S(_0645_),
    .X(_2747_));
 sky130_fd_sc_hd__and3_1 _6317_ (.A(\wave_comb.u1.Q[7] ),
    .B(_0569_),
    .C(_0571_),
    .X(_2748_));
 sky130_fd_sc_hd__a21o_1 _6318_ (.A1(\wave_comb.u1.next_start ),
    .A2(_2747_),
    .B1(_2748_),
    .X(_0052_));
 sky130_fd_sc_hd__a21o_1 _6319_ (.A1(\sound1.sdiv.Q[6] ),
    .A2(_2656_),
    .B1(_2722_),
    .X(_2749_));
 sky130_fd_sc_hd__nand2_1 _6320_ (.A(\sound1.sdiv.Q[7] ),
    .B(_0579_),
    .Y(_2750_));
 sky130_fd_sc_hd__xor2_1 _6321_ (.A(_2749_),
    .B(_2750_),
    .X(_2751_));
 sky130_fd_sc_hd__a21oi_2 _6322_ (.A1(_2407_),
    .A2(_2432_),
    .B1(_2412_),
    .Y(_2752_));
 sky130_fd_sc_hd__or3b_2 _6323_ (.A(net1),
    .B(\wave.mode[1] ),
    .C_N(\wave.mode[0] ),
    .X(_2753_));
 sky130_fd_sc_hd__o2bb2a_1 _6324_ (.A1_N(\sound1.sdiv.Q[8] ),
    .A2_N(_2293_),
    .B1(_2752_),
    .B2(_2753_),
    .X(_2754_));
 sky130_fd_sc_hd__o21a_1 _6325_ (.A1(_2292_),
    .A2(_2751_),
    .B1(_2754_),
    .X(_2755_));
 sky130_fd_sc_hd__a21oi_1 _6326_ (.A1(\sound2.sdiv.Q[6] ),
    .A2(_2660_),
    .B1(_2718_),
    .Y(_2756_));
 sky130_fd_sc_hd__nand2_1 _6327_ (.A(\sound2.sdiv.Q[7] ),
    .B(_0578_),
    .Y(_2757_));
 sky130_fd_sc_hd__xor2_1 _6328_ (.A(_2756_),
    .B(_2757_),
    .X(_2758_));
 sky130_fd_sc_hd__a21oi_2 _6329_ (.A1(_2472_),
    .A2(_2497_),
    .B1(_2477_),
    .Y(_2759_));
 sky130_fd_sc_hd__a2bb2o_1 _6330_ (.A1_N(_2759_),
    .A2_N(_2753_),
    .B1(\sound2.sdiv.Q[8] ),
    .B2(_2295_),
    .X(_2760_));
 sky130_fd_sc_hd__a21oi_1 _6331_ (.A1(_2289_),
    .A2(_2758_),
    .B1(_2760_),
    .Y(_2761_));
 sky130_fd_sc_hd__nor2_1 _6332_ (.A(_2755_),
    .B(_2761_),
    .Y(_2762_));
 sky130_fd_sc_hd__and2_1 _6333_ (.A(_2755_),
    .B(_2761_),
    .X(_2763_));
 sky130_fd_sc_hd__or2_1 _6334_ (.A(_2762_),
    .B(_2763_),
    .X(_2764_));
 sky130_fd_sc_hd__o21a_1 _6335_ (.A1(_2728_),
    .A2(_2729_),
    .B1(_2726_),
    .X(_2765_));
 sky130_fd_sc_hd__xnor2_1 _6336_ (.A(_2764_),
    .B(_2765_),
    .Y(_2766_));
 sky130_fd_sc_hd__a21o_1 _6337_ (.A1(\sound3.sdiv.Q[6] ),
    .A2(_2632_),
    .B1(_2731_),
    .X(_2767_));
 sky130_fd_sc_hd__nand2_1 _6338_ (.A(\sound3.sdiv.Q[7] ),
    .B(_0577_),
    .Y(_2768_));
 sky130_fd_sc_hd__xnor2_1 _6339_ (.A(_2767_),
    .B(_2768_),
    .Y(_2769_));
 sky130_fd_sc_hd__a2bb2o_1 _6340_ (.A1_N(_2569_),
    .A2_N(_2753_),
    .B1(\sound3.sdiv.Q[8] ),
    .B2(_2301_),
    .X(_2770_));
 sky130_fd_sc_hd__a21oi_2 _6341_ (.A1(_2289_),
    .A2(_2769_),
    .B1(_2770_),
    .Y(_2771_));
 sky130_fd_sc_hd__xnor2_1 _6342_ (.A(_2766_),
    .B(_2771_),
    .Y(_2772_));
 sky130_fd_sc_hd__and2b_1 _6343_ (.A_N(net31),
    .B(net30),
    .X(_2773_));
 sky130_fd_sc_hd__nand2_1 _6344_ (.A(\sound4.sdiv.Q[7] ),
    .B(_0576_),
    .Y(_2774_));
 sky130_fd_sc_hd__a21oi_1 _6345_ (.A1(\sound4.sdiv.Q[6] ),
    .A2(_2641_),
    .B1(_2736_),
    .Y(_2775_));
 sky130_fd_sc_hd__xnor2_1 _6346_ (.A(_2774_),
    .B(_2775_),
    .Y(_2776_));
 sky130_fd_sc_hd__nor2_1 _6347_ (.A(_2292_),
    .B(_2776_),
    .Y(_2777_));
 sky130_fd_sc_hd__a221oi_2 _6348_ (.A1(\sound4.sdiv.Q[8] ),
    .A2(_2290_),
    .B1(_2369_),
    .B2(_2773_),
    .C1(_2777_),
    .Y(_2778_));
 sky130_fd_sc_hd__xnor2_1 _6349_ (.A(_2772_),
    .B(_2778_),
    .Y(_2779_));
 sky130_fd_sc_hd__nand2_1 _6350_ (.A(_2730_),
    .B(_2734_),
    .Y(_2780_));
 sky130_fd_sc_hd__nor2_1 _6351_ (.A(_2730_),
    .B(_2734_),
    .Y(_2781_));
 sky130_fd_sc_hd__a21oi_1 _6352_ (.A1(_2780_),
    .A2(_2739_),
    .B1(_2781_),
    .Y(_2782_));
 sky130_fd_sc_hd__xor2_1 _6353_ (.A(_2779_),
    .B(_2782_),
    .X(_2783_));
 sky130_fd_sc_hd__or2b_1 _6354_ (.A(_2742_),
    .B_N(_2740_),
    .X(_2784_));
 sky130_fd_sc_hd__and2b_1 _6355_ (.A_N(_2740_),
    .B(_2742_),
    .X(_2785_));
 sky130_fd_sc_hd__a21o_1 _6356_ (.A1(_2784_),
    .A2(_2745_),
    .B1(_2785_),
    .X(_2786_));
 sky130_fd_sc_hd__or2_1 _6357_ (.A(_2783_),
    .B(_2786_),
    .X(_2787_));
 sky130_fd_sc_hd__a21oi_1 _6358_ (.A1(_2783_),
    .A2(_2786_),
    .B1(_0569_),
    .Y(_2788_));
 sky130_fd_sc_hd__a22o_1 _6359_ (.A1(\wave_comb.u1.Q[7] ),
    .A2(_0569_),
    .B1(_2787_),
    .B2(_2788_),
    .X(_2789_));
 sky130_fd_sc_hd__nand2_1 _6360_ (.A(\wave_comb.u1.Q[8] ),
    .B(_0572_),
    .Y(_2790_));
 sky130_fd_sc_hd__a21bo_1 _6361_ (.A1(\wave_comb.u1.next_start ),
    .A2(_2789_),
    .B1_N(_2790_),
    .X(_0053_));
 sky130_fd_sc_hd__nor2_1 _6362_ (.A(_2764_),
    .B(_2765_),
    .Y(_2791_));
 sky130_fd_sc_hd__nor2_1 _6363_ (.A(_2766_),
    .B(_2771_),
    .Y(_2792_));
 sky130_fd_sc_hd__nor2_1 _6364_ (.A(_2772_),
    .B(_2778_),
    .Y(_2793_));
 sky130_fd_sc_hd__o22a_1 _6365_ (.A1(_2762_),
    .A2(_2791_),
    .B1(_2792_),
    .B2(_2793_),
    .X(_2794_));
 sky130_fd_sc_hd__nor2_1 _6366_ (.A(_2779_),
    .B(_2782_),
    .Y(_2795_));
 sky130_fd_sc_hd__a21oi_1 _6367_ (.A1(_2783_),
    .A2(_2786_),
    .B1(_2795_),
    .Y(_2796_));
 sky130_fd_sc_hd__nor4_1 _6368_ (.A(_2762_),
    .B(_2791_),
    .C(_2792_),
    .D(_2793_),
    .Y(_2797_));
 sky130_fd_sc_hd__or3_1 _6369_ (.A(_2794_),
    .B(_2796_),
    .C(net53),
    .X(_2798_));
 sky130_fd_sc_hd__o21ai_1 _6370_ (.A1(_2794_),
    .A2(net54),
    .B1(_2796_),
    .Y(_2799_));
 sky130_fd_sc_hd__a22o_1 _6371_ (.A1(\wave_comb.u1.Q[9] ),
    .A2(_0573_),
    .B1(_0646_),
    .B2(\wave_comb.u1.Q[8] ),
    .X(_2800_));
 sky130_fd_sc_hd__a31o_1 _6372_ (.A1(_0645_),
    .A2(_2798_),
    .A3(_2799_),
    .B1(_2800_),
    .X(_0054_));
 sky130_fd_sc_hd__mux2_1 _6373_ (.A0(\wave_comb.u1.Q[9] ),
    .A1(\wave_comb.u1.Q[10] ),
    .S(_0571_),
    .X(_2801_));
 sky130_fd_sc_hd__or2_1 _6374_ (.A(_0569_),
    .B(_2794_),
    .X(_2802_));
 sky130_fd_sc_hd__nor2_1 _6375_ (.A(_2796_),
    .B(net53),
    .Y(_2803_));
 sky130_fd_sc_hd__o22a_1 _6376_ (.A1(_0645_),
    .A2(_2801_),
    .B1(_2802_),
    .B2(_2803_),
    .X(_0055_));
 sky130_fd_sc_hd__a22o_1 _6377_ (.A1(\wave_comb.u1.Q[11] ),
    .A2(_0573_),
    .B1(\wave_comb.u1.next_dived ),
    .B2(\wave_comb.u1.Q[10] ),
    .X(_0056_));
 sky130_fd_sc_hd__nand2_1 _6378_ (.A(_0632_),
    .B(_0643_),
    .Y(_2804_));
 sky130_fd_sc_hd__o21a_4 _6379_ (.A1(net34),
    .A2(_2804_),
    .B1(_0700_),
    .X(_2805_));
 sky130_fd_sc_hd__mux2_1 _6380_ (.A0(_2280_),
    .A1(_2274_),
    .S(_2805_),
    .X(_2806_));
 sky130_fd_sc_hd__and3_1 _6381_ (.A(\wave_comb.u1.dived ),
    .B(_0569_),
    .C(_0571_),
    .X(_2807_));
 sky130_fd_sc_hd__clkbuf_4 _6382_ (.A(_2807_),
    .X(_2808_));
 sky130_fd_sc_hd__mux2_1 _6383_ (.A0(\pm.current_waveform[0] ),
    .A1(_2806_),
    .S(_2808_),
    .X(_2809_));
 sky130_fd_sc_hd__clkbuf_1 _6384_ (.A(_2809_),
    .X(_0057_));
 sky130_fd_sc_hd__mux2_1 _6385_ (.A0(_2294_),
    .A1(_2310_),
    .S(_2805_),
    .X(_2810_));
 sky130_fd_sc_hd__mux2_1 _6386_ (.A0(\pm.current_waveform[1] ),
    .A1(_2810_),
    .S(_2808_),
    .X(_2811_));
 sky130_fd_sc_hd__clkbuf_1 _6387_ (.A(_2811_),
    .X(_0058_));
 sky130_fd_sc_hd__mux2_1 _6388_ (.A0(_2439_),
    .A1(_2581_),
    .S(_2805_),
    .X(_2812_));
 sky130_fd_sc_hd__mux2_1 _6389_ (.A0(\pm.current_waveform[2] ),
    .A1(_2812_),
    .S(_2808_),
    .X(_2813_));
 sky130_fd_sc_hd__clkbuf_1 _6390_ (.A(_2813_),
    .X(_0059_));
 sky130_fd_sc_hd__mux2_1 _6391_ (.A0(_2590_),
    .A1(_2616_),
    .S(_2805_),
    .X(_2814_));
 sky130_fd_sc_hd__mux2_1 _6392_ (.A0(\pm.current_waveform[3] ),
    .A1(_2814_),
    .S(_2808_),
    .X(_2815_));
 sky130_fd_sc_hd__clkbuf_1 _6393_ (.A(_2815_),
    .X(_0060_));
 sky130_fd_sc_hd__mux2_1 _6394_ (.A0(_2623_),
    .A1(_2655_),
    .S(_2805_),
    .X(_2816_));
 sky130_fd_sc_hd__inv_2 _6395_ (.A(_2816_),
    .Y(_2817_));
 sky130_fd_sc_hd__mux2_1 _6396_ (.A0(\pm.current_waveform[4] ),
    .A1(_2817_),
    .S(_2808_),
    .X(_2818_));
 sky130_fd_sc_hd__clkbuf_1 _6397_ (.A(_2818_),
    .X(_0061_));
 sky130_fd_sc_hd__mux2_1 _6398_ (.A0(_2659_),
    .A1(_2682_),
    .S(_2805_),
    .X(_2819_));
 sky130_fd_sc_hd__inv_2 _6399_ (.A(_2819_),
    .Y(_2820_));
 sky130_fd_sc_hd__mux2_1 _6400_ (.A0(\pm.current_waveform[5] ),
    .A1(_2820_),
    .S(_2808_),
    .X(_2821_));
 sky130_fd_sc_hd__clkbuf_1 _6401_ (.A(_2821_),
    .X(_0062_));
 sky130_fd_sc_hd__mux2_1 _6402_ (.A0(_2693_),
    .A1(_2716_),
    .S(_2805_),
    .X(_2822_));
 sky130_fd_sc_hd__mux2_1 _6403_ (.A0(\pm.current_waveform[6] ),
    .A1(_2822_),
    .S(_2808_),
    .X(_2823_));
 sky130_fd_sc_hd__clkbuf_1 _6404_ (.A(_2823_),
    .X(_0063_));
 sky130_fd_sc_hd__mux2_1 _6405_ (.A0(_2725_),
    .A1(_2748_),
    .S(_2805_),
    .X(_2824_));
 sky130_fd_sc_hd__mux2_1 _6406_ (.A0(\pm.current_waveform[7] ),
    .A1(_2824_),
    .S(_2808_),
    .X(_2825_));
 sky130_fd_sc_hd__clkbuf_1 _6407_ (.A(_2825_),
    .X(_0064_));
 sky130_fd_sc_hd__mux2_1 _6408_ (.A0(_2755_),
    .A1(_2790_),
    .S(_2805_),
    .X(_2826_));
 sky130_fd_sc_hd__inv_2 _6409_ (.A(_2826_),
    .Y(_2827_));
 sky130_fd_sc_hd__mux2_1 _6410_ (.A0(\pm.current_waveform[8] ),
    .A1(_2827_),
    .S(_2808_),
    .X(_2828_));
 sky130_fd_sc_hd__clkbuf_1 _6411_ (.A(_2828_),
    .X(_0065_));
 sky130_fd_sc_hd__nand2_1 _6412_ (.A(_0719_),
    .B(\seq.encode.play ),
    .Y(_2829_));
 sky130_fd_sc_hd__nor2_1 _6413_ (.A(_0811_),
    .B(_2829_),
    .Y(_2830_));
 sky130_fd_sc_hd__xor2_1 _6414_ (.A(\seq.beat[0] ),
    .B(_2830_),
    .X(_0066_));
 sky130_fd_sc_hd__a21oi_1 _6415_ (.A1(\seq.beat[0] ),
    .A2(_2830_),
    .B1(\seq.beat[1] ),
    .Y(_2831_));
 sky130_fd_sc_hd__and3_1 _6416_ (.A(\seq.beat[1] ),
    .B(\seq.beat[0] ),
    .C(_2830_),
    .X(_2832_));
 sky130_fd_sc_hd__nor2_1 _6417_ (.A(_2831_),
    .B(_2832_),
    .Y(_0067_));
 sky130_fd_sc_hd__or2_1 _6418_ (.A(\seq.beat[2] ),
    .B(_2832_),
    .X(_2833_));
 sky130_fd_sc_hd__nand2_1 _6419_ (.A(\seq.beat[2] ),
    .B(_2832_),
    .Y(_2834_));
 sky130_fd_sc_hd__and2_1 _6420_ (.A(_2833_),
    .B(_2834_),
    .X(_2835_));
 sky130_fd_sc_hd__clkbuf_1 _6421_ (.A(_2835_),
    .X(_0068_));
 sky130_fd_sc_hd__xnor2_1 _6422_ (.A(\seq.beat[3] ),
    .B(_2834_),
    .Y(_0069_));
 sky130_fd_sc_hd__buf_4 _6423_ (.A(_0554_),
    .X(_2836_));
 sky130_fd_sc_hd__and2_1 _6424_ (.A(\sound1.count[0] ),
    .B(_2201_),
    .X(_2837_));
 sky130_fd_sc_hd__a21o_1 _6425_ (.A1(\sound1.count_m[0] ),
    .A2(_2836_),
    .B1(_2837_),
    .X(_0070_));
 sky130_fd_sc_hd__and2_1 _6426_ (.A(\sound1.count[1] ),
    .B(_2201_),
    .X(_2838_));
 sky130_fd_sc_hd__a21o_1 _6427_ (.A1(\sound1.count_m[1] ),
    .A2(_2836_),
    .B1(_2838_),
    .X(_0071_));
 sky130_fd_sc_hd__and2_1 _6428_ (.A(\sound1.count[2] ),
    .B(_2201_),
    .X(_2839_));
 sky130_fd_sc_hd__a21o_1 _6429_ (.A1(\sound1.count_m[2] ),
    .A2(_2836_),
    .B1(_2839_),
    .X(_0072_));
 sky130_fd_sc_hd__and2_1 _6430_ (.A(\sound1.count[3] ),
    .B(_2201_),
    .X(_2840_));
 sky130_fd_sc_hd__a21o_1 _6431_ (.A1(\sound1.count_m[3] ),
    .A2(_2836_),
    .B1(_2840_),
    .X(_0073_));
 sky130_fd_sc_hd__and2_1 _6432_ (.A(\sound1.count[4] ),
    .B(_2201_),
    .X(_2841_));
 sky130_fd_sc_hd__a21o_1 _6433_ (.A1(\sound1.count_m[4] ),
    .A2(_2836_),
    .B1(_2841_),
    .X(_0074_));
 sky130_fd_sc_hd__and2_1 _6434_ (.A(\sound1.count[5] ),
    .B(_2201_),
    .X(_2842_));
 sky130_fd_sc_hd__a21o_1 _6435_ (.A1(\sound1.count_m[5] ),
    .A2(_2836_),
    .B1(_2842_),
    .X(_0075_));
 sky130_fd_sc_hd__clkbuf_16 _6436_ (.A(_0554_),
    .X(_2843_));
 sky130_fd_sc_hd__nor2_1 _6437_ (.A(_1237_),
    .B(_2843_),
    .Y(_2844_));
 sky130_fd_sc_hd__a21o_1 _6438_ (.A1(\sound1.count_m[6] ),
    .A2(_2836_),
    .B1(_2844_),
    .X(_0076_));
 sky130_fd_sc_hd__nor2_1 _6439_ (.A(_1073_),
    .B(_2843_),
    .Y(_2845_));
 sky130_fd_sc_hd__a21o_1 _6440_ (.A1(\sound1.count_m[7] ),
    .A2(_2836_),
    .B1(_2845_),
    .X(_0077_));
 sky130_fd_sc_hd__and2_1 _6441_ (.A(\sound1.count[8] ),
    .B(_2201_),
    .X(_2846_));
 sky130_fd_sc_hd__a21o_1 _6442_ (.A1(\sound1.count_m[8] ),
    .A2(_2836_),
    .B1(_2846_),
    .X(_0078_));
 sky130_fd_sc_hd__and2_1 _6443_ (.A(\sound1.count[9] ),
    .B(_2201_),
    .X(_2847_));
 sky130_fd_sc_hd__a21o_1 _6444_ (.A1(\sound1.count_m[9] ),
    .A2(_2836_),
    .B1(_2847_),
    .X(_0079_));
 sky130_fd_sc_hd__and2_1 _6445_ (.A(\sound1.count[10] ),
    .B(_2201_),
    .X(_2848_));
 sky130_fd_sc_hd__a21o_1 _6446_ (.A1(\sound1.count_m[10] ),
    .A2(_2836_),
    .B1(_2848_),
    .X(_0080_));
 sky130_fd_sc_hd__and2_1 _6447_ (.A(\sound1.count[11] ),
    .B(_2201_),
    .X(_2849_));
 sky130_fd_sc_hd__a21o_1 _6448_ (.A1(\sound1.count_m[11] ),
    .A2(_2836_),
    .B1(_2849_),
    .X(_0081_));
 sky130_fd_sc_hd__and2_1 _6449_ (.A(\sound1.count[12] ),
    .B(_2201_),
    .X(_2850_));
 sky130_fd_sc_hd__a21o_1 _6450_ (.A1(\sound1.count_m[12] ),
    .A2(_2836_),
    .B1(_2850_),
    .X(_0082_));
 sky130_fd_sc_hd__and2_1 _6451_ (.A(\sound1.count[13] ),
    .B(_2201_),
    .X(_2851_));
 sky130_fd_sc_hd__a21o_1 _6452_ (.A1(\sound1.count_m[13] ),
    .A2(_2836_),
    .B1(_2851_),
    .X(_0083_));
 sky130_fd_sc_hd__and2_1 _6453_ (.A(\sound1.count[14] ),
    .B(_2201_),
    .X(_2852_));
 sky130_fd_sc_hd__a21o_1 _6454_ (.A1(\sound1.count_m[14] ),
    .A2(_2836_),
    .B1(_2852_),
    .X(_0084_));
 sky130_fd_sc_hd__and2_1 _6455_ (.A(\sound1.count[15] ),
    .B(_2201_),
    .X(_2853_));
 sky130_fd_sc_hd__a21o_1 _6456_ (.A1(\sound1.count_m[15] ),
    .A2(_2836_),
    .B1(_2853_),
    .X(_0085_));
 sky130_fd_sc_hd__and2_1 _6457_ (.A(\sound1.count[16] ),
    .B(_2201_),
    .X(_2854_));
 sky130_fd_sc_hd__a21o_1 _6458_ (.A1(\sound1.count_m[16] ),
    .A2(_2836_),
    .B1(_2854_),
    .X(_0086_));
 sky130_fd_sc_hd__buf_6 _6459_ (.A(_0575_),
    .X(_2855_));
 sky130_fd_sc_hd__and2_1 _6460_ (.A(\sound1.count[17] ),
    .B(_2855_),
    .X(_2856_));
 sky130_fd_sc_hd__a21o_1 _6461_ (.A1(\sound1.count_m[17] ),
    .A2(_2836_),
    .B1(_2856_),
    .X(_0087_));
 sky130_fd_sc_hd__buf_6 _6462_ (.A(_0554_),
    .X(_2857_));
 sky130_fd_sc_hd__and2_1 _6463_ (.A(\sound1.count[18] ),
    .B(_2855_),
    .X(_2858_));
 sky130_fd_sc_hd__a21o_1 _6464_ (.A1(\sound1.count_m[18] ),
    .A2(_2857_),
    .B1(_2858_),
    .X(_0088_));
 sky130_fd_sc_hd__inv_2 _6465_ (.A(_1104_),
    .Y(_2859_));
 sky130_fd_sc_hd__mux2_1 _6466_ (.A0(\sound1.divisor_m[0] ),
    .A1(_2859_),
    .S(_2005_),
    .X(_2860_));
 sky130_fd_sc_hd__clkbuf_1 _6467_ (.A(_2860_),
    .X(_0089_));
 sky130_fd_sc_hd__mux2_1 _6468_ (.A0(\sound1.divisor_m[1] ),
    .A1(_1008_),
    .S(_2005_),
    .X(_2861_));
 sky130_fd_sc_hd__clkbuf_1 _6469_ (.A(_2861_),
    .X(_0090_));
 sky130_fd_sc_hd__inv_2 _6470_ (.A(_1032_),
    .Y(_2862_));
 sky130_fd_sc_hd__clkbuf_8 _6471_ (.A(_0575_),
    .X(_2863_));
 sky130_fd_sc_hd__clkbuf_16 _6472_ (.A(_2863_),
    .X(_2864_));
 sky130_fd_sc_hd__mux2_1 _6473_ (.A0(\sound1.divisor_m[2] ),
    .A1(_2862_),
    .S(_2864_),
    .X(_2865_));
 sky130_fd_sc_hd__clkbuf_1 _6474_ (.A(_2865_),
    .X(_0091_));
 sky130_fd_sc_hd__nor2_1 _6475_ (.A(\sound1.divisor_m[3] ),
    .B(_2005_),
    .Y(_2866_));
 sky130_fd_sc_hd__a21oi_1 _6476_ (.A1(_2005_),
    .A2(_1208_),
    .B1(_2866_),
    .Y(_0092_));
 sky130_fd_sc_hd__inv_2 _6477_ (.A(_1145_),
    .Y(_2867_));
 sky130_fd_sc_hd__mux2_1 _6478_ (.A0(\sound1.divisor_m[4] ),
    .A1(_2867_),
    .S(_2864_),
    .X(_2868_));
 sky130_fd_sc_hd__clkbuf_1 _6479_ (.A(_2868_),
    .X(_0093_));
 sky130_fd_sc_hd__mux2_1 _6480_ (.A0(\sound1.divisor_m[5] ),
    .A1(_1186_),
    .S(_2864_),
    .X(_2869_));
 sky130_fd_sc_hd__clkbuf_1 _6481_ (.A(_2869_),
    .X(_0094_));
 sky130_fd_sc_hd__mux2_1 _6482_ (.A0(\sound1.divisor_m[6] ),
    .A1(_1071_),
    .S(_2864_),
    .X(_2870_));
 sky130_fd_sc_hd__clkbuf_1 _6483_ (.A(_2870_),
    .X(_0095_));
 sky130_fd_sc_hd__mux2_1 _6484_ (.A0(\sound1.divisor_m[7] ),
    .A1(_1089_),
    .S(_2864_),
    .X(_2871_));
 sky130_fd_sc_hd__clkbuf_1 _6485_ (.A(_2871_),
    .X(_0096_));
 sky130_fd_sc_hd__inv_2 _6486_ (.A(_1170_),
    .Y(_2872_));
 sky130_fd_sc_hd__mux2_1 _6487_ (.A0(\sound1.divisor_m[8] ),
    .A1(_2872_),
    .S(_2864_),
    .X(_2873_));
 sky130_fd_sc_hd__clkbuf_1 _6488_ (.A(_2873_),
    .X(_0097_));
 sky130_fd_sc_hd__nor2_1 _6489_ (.A(\sound1.divisor_m[9] ),
    .B(_2005_),
    .Y(_2874_));
 sky130_fd_sc_hd__a21oi_1 _6490_ (.A1(_2005_),
    .A2(_1196_),
    .B1(_2874_),
    .Y(_0098_));
 sky130_fd_sc_hd__inv_2 _6491_ (.A(_1157_),
    .Y(_2875_));
 sky130_fd_sc_hd__mux2_1 _6492_ (.A0(\sound1.divisor_m[10] ),
    .A1(_2875_),
    .S(_2864_),
    .X(_2876_));
 sky130_fd_sc_hd__clkbuf_1 _6493_ (.A(_2876_),
    .X(_0099_));
 sky130_fd_sc_hd__inv_2 _6494_ (.A(_1050_),
    .Y(_2877_));
 sky130_fd_sc_hd__mux2_1 _6495_ (.A0(\sound1.divisor_m[11] ),
    .A1(_2877_),
    .S(_2864_),
    .X(_2878_));
 sky130_fd_sc_hd__clkbuf_1 _6496_ (.A(_2878_),
    .X(_0100_));
 sky130_fd_sc_hd__inv_2 _6497_ (.A(_1249_),
    .Y(_2879_));
 sky130_fd_sc_hd__mux2_1 _6498_ (.A0(\sound1.divisor_m[12] ),
    .A1(_2879_),
    .S(_2864_),
    .X(_2880_));
 sky130_fd_sc_hd__clkbuf_1 _6499_ (.A(_2880_),
    .X(_0101_));
 sky130_fd_sc_hd__mux2_1 _6500_ (.A0(\sound1.divisor_m[13] ),
    .A1(_1120_),
    .S(_2864_),
    .X(_2881_));
 sky130_fd_sc_hd__clkbuf_1 _6501_ (.A(_2881_),
    .X(_0102_));
 sky130_fd_sc_hd__inv_2 _6502_ (.A(_1235_),
    .Y(_2882_));
 sky130_fd_sc_hd__mux2_1 _6503_ (.A0(\sound1.divisor_m[14] ),
    .A1(_2882_),
    .S(_2864_),
    .X(_2883_));
 sky130_fd_sc_hd__clkbuf_1 _6504_ (.A(_2883_),
    .X(_0103_));
 sky130_fd_sc_hd__inv_2 _6505_ (.A(_1215_),
    .Y(_2884_));
 sky130_fd_sc_hd__mux2_1 _6506_ (.A0(\sound1.divisor_m[15] ),
    .A1(_2884_),
    .S(_2864_),
    .X(_2885_));
 sky130_fd_sc_hd__clkbuf_1 _6507_ (.A(_2885_),
    .X(_0104_));
 sky130_fd_sc_hd__inv_2 _6508_ (.A(_1219_),
    .Y(_2886_));
 sky130_fd_sc_hd__mux2_1 _6509_ (.A0(\sound1.divisor_m[16] ),
    .A1(_2886_),
    .S(_2864_),
    .X(_2887_));
 sky130_fd_sc_hd__clkbuf_1 _6510_ (.A(_2887_),
    .X(_0105_));
 sky130_fd_sc_hd__mux2_1 _6511_ (.A0(\sound1.divisor_m[17] ),
    .A1(_1225_),
    .S(_2864_),
    .X(_2888_));
 sky130_fd_sc_hd__clkbuf_1 _6512_ (.A(_2888_),
    .X(_0106_));
 sky130_fd_sc_hd__mux2_1 _6513_ (.A0(\sound1.divisor_m[18] ),
    .A1(_1223_),
    .S(_2864_),
    .X(_2889_));
 sky130_fd_sc_hd__clkbuf_1 _6514_ (.A(_2889_),
    .X(_0107_));
 sky130_fd_sc_hd__buf_8 _6515_ (.A(_0867_),
    .X(_2890_));
 sky130_fd_sc_hd__nand2_1 _6516_ (.A(\sound1.divisor_m[0] ),
    .B(\sound1.sdiv.Q[27] ),
    .Y(_2891_));
 sky130_fd_sc_hd__or2_1 _6517_ (.A(\sound1.divisor_m[0] ),
    .B(\sound1.sdiv.Q[27] ),
    .X(_2892_));
 sky130_fd_sc_hd__buf_6 _6518_ (.A(_0579_),
    .X(_2893_));
 sky130_fd_sc_hd__buf_6 _6519_ (.A(_2893_),
    .X(_2894_));
 sky130_fd_sc_hd__a32o_1 _6520_ (.A1(_2890_),
    .A2(_2891_),
    .A3(_2892_),
    .B1(_2894_),
    .B2(\sound1.sdiv.A[0] ),
    .X(_0108_));
 sky130_fd_sc_hd__clkbuf_8 _6521_ (.A(_2893_),
    .X(_2895_));
 sky130_fd_sc_hd__and2b_1 _6522_ (.A_N(\sound1.sdiv.A[26] ),
    .B(\sound1.divisor_m[0] ),
    .X(_2896_));
 sky130_fd_sc_hd__xnor2_1 _6523_ (.A(\sound1.divisor_m[1] ),
    .B(_2896_),
    .Y(_2897_));
 sky130_fd_sc_hd__xnor2_1 _6524_ (.A(\sound1.sdiv.A[0] ),
    .B(_2897_),
    .Y(_2898_));
 sky130_fd_sc_hd__xnor2_1 _6525_ (.A(_2891_),
    .B(_2898_),
    .Y(_2899_));
 sky130_fd_sc_hd__a22o_1 _6526_ (.A1(\sound1.sdiv.A[1] ),
    .A2(_2895_),
    .B1(\sound1.sdiv.next_dived ),
    .B2(_2899_),
    .X(_0109_));
 sky130_fd_sc_hd__and2b_1 _6527_ (.A_N(_2897_),
    .B(\sound1.sdiv.A[0] ),
    .X(_2900_));
 sky130_fd_sc_hd__a31oi_2 _6528_ (.A1(\sound1.divisor_m[0] ),
    .A2(\sound1.sdiv.Q[27] ),
    .A3(_2898_),
    .B1(_2900_),
    .Y(_2901_));
 sky130_fd_sc_hd__inv_2 _6529_ (.A(\sound1.sdiv.A[1] ),
    .Y(_2902_));
 sky130_fd_sc_hd__clkinv_4 _6530_ (.A(\sound1.sdiv.A[26] ),
    .Y(_2903_));
 sky130_fd_sc_hd__o21a_1 _6531_ (.A1(\sound1.divisor_m[1] ),
    .A2(\sound1.divisor_m[0] ),
    .B1(_2903_),
    .X(_2904_));
 sky130_fd_sc_hd__xnor2_1 _6532_ (.A(\sound1.divisor_m[2] ),
    .B(_2904_),
    .Y(_2905_));
 sky130_fd_sc_hd__xnor2_1 _6533_ (.A(_2902_),
    .B(_2905_),
    .Y(_2906_));
 sky130_fd_sc_hd__xor2_1 _6534_ (.A(_2901_),
    .B(_2906_),
    .X(_2907_));
 sky130_fd_sc_hd__a22o_1 _6535_ (.A1(\sound1.sdiv.A[2] ),
    .A2(_2895_),
    .B1(\sound1.sdiv.next_dived ),
    .B2(_2907_),
    .X(_0110_));
 sky130_fd_sc_hd__or2_1 _6536_ (.A(_2902_),
    .B(_2905_),
    .X(_2908_));
 sky130_fd_sc_hd__o21a_1 _6537_ (.A1(_2901_),
    .A2(_2906_),
    .B1(_2908_),
    .X(_2909_));
 sky130_fd_sc_hd__inv_2 _6538_ (.A(\sound1.sdiv.A[2] ),
    .Y(_2910_));
 sky130_fd_sc_hd__o31a_1 _6539_ (.A1(\sound1.divisor_m[2] ),
    .A2(\sound1.divisor_m[1] ),
    .A3(\sound1.divisor_m[0] ),
    .B1(_2903_),
    .X(_2911_));
 sky130_fd_sc_hd__xnor2_1 _6540_ (.A(\sound1.divisor_m[3] ),
    .B(_2911_),
    .Y(_2912_));
 sky130_fd_sc_hd__or2_1 _6541_ (.A(_2910_),
    .B(_2912_),
    .X(_2913_));
 sky130_fd_sc_hd__nand2_1 _6542_ (.A(_2910_),
    .B(_2912_),
    .Y(_2914_));
 sky130_fd_sc_hd__nand2_1 _6543_ (.A(_2913_),
    .B(_2914_),
    .Y(_2915_));
 sky130_fd_sc_hd__or2_1 _6544_ (.A(_2909_),
    .B(_2915_),
    .X(_2916_));
 sky130_fd_sc_hd__a21oi_1 _6545_ (.A1(_2909_),
    .A2(_2915_),
    .B1(_0866_),
    .Y(_2917_));
 sky130_fd_sc_hd__a22o_1 _6546_ (.A1(\sound1.sdiv.A[3] ),
    .A2(_2895_),
    .B1(_2916_),
    .B2(_2917_),
    .X(_0111_));
 sky130_fd_sc_hd__inv_2 _6547_ (.A(\sound1.sdiv.A[3] ),
    .Y(_2918_));
 sky130_fd_sc_hd__or4_1 _6548_ (.A(\sound1.divisor_m[3] ),
    .B(\sound1.divisor_m[2] ),
    .C(\sound1.divisor_m[1] ),
    .D(\sound1.divisor_m[0] ),
    .X(_2919_));
 sky130_fd_sc_hd__nand2_1 _6549_ (.A(_2903_),
    .B(_2919_),
    .Y(_2920_));
 sky130_fd_sc_hd__xnor2_1 _6550_ (.A(_2419_),
    .B(_2920_),
    .Y(_2921_));
 sky130_fd_sc_hd__nor2_1 _6551_ (.A(_2918_),
    .B(_2921_),
    .Y(_2922_));
 sky130_fd_sc_hd__nand2_1 _6552_ (.A(_2918_),
    .B(_2921_),
    .Y(_2923_));
 sky130_fd_sc_hd__or2b_1 _6553_ (.A(_2922_),
    .B_N(_2923_),
    .X(_2924_));
 sky130_fd_sc_hd__o21ai_1 _6554_ (.A1(_2909_),
    .A2(_2915_),
    .B1(_2913_),
    .Y(_2925_));
 sky130_fd_sc_hd__xnor2_1 _6555_ (.A(_2924_),
    .B(_2925_),
    .Y(_2926_));
 sky130_fd_sc_hd__a22o_1 _6556_ (.A1(\sound1.sdiv.A[4] ),
    .A2(_2895_),
    .B1(\sound1.sdiv.next_dived ),
    .B2(_2926_),
    .X(_0112_));
 sky130_fd_sc_hd__inv_2 _6557_ (.A(\sound1.sdiv.A[4] ),
    .Y(_2927_));
 sky130_fd_sc_hd__o21a_1 _6558_ (.A1(\sound1.divisor_m[4] ),
    .A2(_2919_),
    .B1(_2903_),
    .X(_2928_));
 sky130_fd_sc_hd__xnor2_1 _6559_ (.A(\sound1.divisor_m[5] ),
    .B(_2928_),
    .Y(_2929_));
 sky130_fd_sc_hd__or2_1 _6560_ (.A(_2927_),
    .B(_2929_),
    .X(_2930_));
 sky130_fd_sc_hd__nand2_1 _6561_ (.A(_2927_),
    .B(_2929_),
    .Y(_2931_));
 sky130_fd_sc_hd__nand2_1 _6562_ (.A(_2930_),
    .B(_2931_),
    .Y(_2932_));
 sky130_fd_sc_hd__a21oi_1 _6563_ (.A1(_2923_),
    .A2(_2925_),
    .B1(_2922_),
    .Y(_2933_));
 sky130_fd_sc_hd__or2_1 _6564_ (.A(_2932_),
    .B(_2933_),
    .X(_2934_));
 sky130_fd_sc_hd__nand2_1 _6565_ (.A(_2932_),
    .B(_2933_),
    .Y(_2935_));
 sky130_fd_sc_hd__a32o_1 _6566_ (.A1(_2890_),
    .A2(_2934_),
    .A3(_2935_),
    .B1(_2894_),
    .B2(\sound1.sdiv.A[5] ),
    .X(_0113_));
 sky130_fd_sc_hd__inv_2 _6567_ (.A(\sound1.sdiv.A[5] ),
    .Y(_2936_));
 sky130_fd_sc_hd__or3_1 _6568_ (.A(\sound1.divisor_m[5] ),
    .B(\sound1.divisor_m[4] ),
    .C(_2919_),
    .X(_2937_));
 sky130_fd_sc_hd__and2_1 _6569_ (.A(_2903_),
    .B(_2937_),
    .X(_2938_));
 sky130_fd_sc_hd__xnor2_1 _6570_ (.A(\sound1.divisor_m[6] ),
    .B(_2938_),
    .Y(_2939_));
 sky130_fd_sc_hd__or2_1 _6571_ (.A(_2936_),
    .B(_2939_),
    .X(_2940_));
 sky130_fd_sc_hd__nand2_1 _6572_ (.A(_2936_),
    .B(_2939_),
    .Y(_2941_));
 sky130_fd_sc_hd__nand2_1 _6573_ (.A(_2940_),
    .B(_2941_),
    .Y(_2942_));
 sky130_fd_sc_hd__o21a_1 _6574_ (.A1(_2932_),
    .A2(_2933_),
    .B1(_2930_),
    .X(_2943_));
 sky130_fd_sc_hd__nor2_1 _6575_ (.A(_2942_),
    .B(_2943_),
    .Y(_2944_));
 sky130_fd_sc_hd__a21o_1 _6576_ (.A1(_2942_),
    .A2(_2943_),
    .B1(_0866_),
    .X(_2945_));
 sky130_fd_sc_hd__a2bb2o_1 _6577_ (.A1_N(_2944_),
    .A2_N(_2945_),
    .B1(\sound1.sdiv.A[6] ),
    .B2(_2895_),
    .X(_0114_));
 sky130_fd_sc_hd__o21a_1 _6578_ (.A1(_2942_),
    .A2(_2943_),
    .B1(_2940_),
    .X(_2946_));
 sky130_fd_sc_hd__inv_2 _6579_ (.A(\sound1.sdiv.A[6] ),
    .Y(_2947_));
 sky130_fd_sc_hd__or2_1 _6580_ (.A(\sound1.divisor_m[6] ),
    .B(_2937_),
    .X(_2948_));
 sky130_fd_sc_hd__and2_1 _6581_ (.A(_2903_),
    .B(_2948_),
    .X(_2949_));
 sky130_fd_sc_hd__xnor2_1 _6582_ (.A(\sound1.divisor_m[7] ),
    .B(_2949_),
    .Y(_2950_));
 sky130_fd_sc_hd__or2_1 _6583_ (.A(_2947_),
    .B(_2950_),
    .X(_2951_));
 sky130_fd_sc_hd__nand2_1 _6584_ (.A(_2947_),
    .B(_2950_),
    .Y(_2952_));
 sky130_fd_sc_hd__nand2_1 _6585_ (.A(_2951_),
    .B(_2952_),
    .Y(_2953_));
 sky130_fd_sc_hd__nor2_1 _6586_ (.A(_2946_),
    .B(_2953_),
    .Y(_2954_));
 sky130_fd_sc_hd__a21o_1 _6587_ (.A1(_2946_),
    .A2(_2953_),
    .B1(_0866_),
    .X(_2955_));
 sky130_fd_sc_hd__a2bb2o_1 _6588_ (.A1_N(_2954_),
    .A2_N(_2955_),
    .B1(\sound1.sdiv.A[7] ),
    .B2(_2895_),
    .X(_0115_));
 sky130_fd_sc_hd__inv_2 _6589_ (.A(\sound1.sdiv.A[7] ),
    .Y(_2956_));
 sky130_fd_sc_hd__nor2_1 _6590_ (.A(\sound1.divisor_m[7] ),
    .B(_2948_),
    .Y(_2957_));
 sky130_fd_sc_hd__nor2_1 _6591_ (.A(\sound1.sdiv.A[26] ),
    .B(_2957_),
    .Y(_2958_));
 sky130_fd_sc_hd__xnor2_1 _6592_ (.A(\sound1.divisor_m[8] ),
    .B(_2958_),
    .Y(_2959_));
 sky130_fd_sc_hd__nor2_1 _6593_ (.A(_2956_),
    .B(_2959_),
    .Y(_2960_));
 sky130_fd_sc_hd__and2_1 _6594_ (.A(_2956_),
    .B(_2959_),
    .X(_2961_));
 sky130_fd_sc_hd__or2_1 _6595_ (.A(_2960_),
    .B(_2961_),
    .X(_2962_));
 sky130_fd_sc_hd__o21a_1 _6596_ (.A1(_2946_),
    .A2(_2953_),
    .B1(_2951_),
    .X(_2963_));
 sky130_fd_sc_hd__or2_1 _6597_ (.A(_2962_),
    .B(_2963_),
    .X(_2964_));
 sky130_fd_sc_hd__a21oi_1 _6598_ (.A1(_2962_),
    .A2(_2963_),
    .B1(_0866_),
    .Y(_2965_));
 sky130_fd_sc_hd__a22o_1 _6599_ (.A1(\sound1.sdiv.A[8] ),
    .A2(_2895_),
    .B1(_2964_),
    .B2(_2965_),
    .X(_0116_));
 sky130_fd_sc_hd__inv_2 _6600_ (.A(_2960_),
    .Y(_2966_));
 sky130_fd_sc_hd__a21o_1 _6601_ (.A1(_2395_),
    .A2(_2957_),
    .B1(\sound1.sdiv.A[26] ),
    .X(_2967_));
 sky130_fd_sc_hd__xnor2_1 _6602_ (.A(\sound1.divisor_m[9] ),
    .B(_2967_),
    .Y(_2968_));
 sky130_fd_sc_hd__and2_1 _6603_ (.A(\sound1.sdiv.A[8] ),
    .B(_2968_),
    .X(_2969_));
 sky130_fd_sc_hd__nor2_1 _6604_ (.A(\sound1.sdiv.A[8] ),
    .B(_2968_),
    .Y(_2970_));
 sky130_fd_sc_hd__or2_1 _6605_ (.A(_2969_),
    .B(_2970_),
    .X(_2971_));
 sky130_fd_sc_hd__and3_1 _6606_ (.A(_2966_),
    .B(_2964_),
    .C(_2971_),
    .X(_2972_));
 sky130_fd_sc_hd__a21oi_1 _6607_ (.A1(_2966_),
    .A2(_2964_),
    .B1(_2971_),
    .Y(_2973_));
 sky130_fd_sc_hd__inv_2 _6608_ (.A(\sound1.sdiv.A[9] ),
    .Y(_2974_));
 sky130_fd_sc_hd__o32ai_1 _6609_ (.A1(_0866_),
    .A2(_2972_),
    .A3(_2973_),
    .B1(\sound1.sdiv.next_start ),
    .B2(_2974_),
    .Y(_0117_));
 sky130_fd_sc_hd__inv_2 _6610_ (.A(_2969_),
    .Y(_2975_));
 sky130_fd_sc_hd__o211a_1 _6611_ (.A1(_2962_),
    .A2(_2963_),
    .B1(_2975_),
    .C1(_2966_),
    .X(_2976_));
 sky130_fd_sc_hd__or4_1 _6612_ (.A(\sound1.divisor_m[9] ),
    .B(\sound1.divisor_m[8] ),
    .C(\sound1.divisor_m[7] ),
    .D(_2948_),
    .X(_2977_));
 sky130_fd_sc_hd__and2_1 _6613_ (.A(_2903_),
    .B(_2977_),
    .X(_2978_));
 sky130_fd_sc_hd__xnor2_1 _6614_ (.A(\sound1.divisor_m[10] ),
    .B(_2978_),
    .Y(_2979_));
 sky130_fd_sc_hd__xnor2_1 _6615_ (.A(_2974_),
    .B(_2979_),
    .Y(_2980_));
 sky130_fd_sc_hd__o21ai_1 _6616_ (.A1(_2970_),
    .A2(_2976_),
    .B1(_2980_),
    .Y(_2981_));
 sky130_fd_sc_hd__or3_1 _6617_ (.A(_2970_),
    .B(_2980_),
    .C(_2976_),
    .X(_2982_));
 sky130_fd_sc_hd__a32o_1 _6618_ (.A1(_2890_),
    .A2(_2981_),
    .A3(_2982_),
    .B1(_2894_),
    .B2(\sound1.sdiv.A[10] ),
    .X(_0118_));
 sky130_fd_sc_hd__inv_2 _6619_ (.A(\sound1.sdiv.A[10] ),
    .Y(_2983_));
 sky130_fd_sc_hd__or2_1 _6620_ (.A(\sound1.divisor_m[10] ),
    .B(_2977_),
    .X(_2984_));
 sky130_fd_sc_hd__and2_1 _6621_ (.A(_2903_),
    .B(_2984_),
    .X(_2985_));
 sky130_fd_sc_hd__xnor2_1 _6622_ (.A(\sound1.divisor_m[11] ),
    .B(_2985_),
    .Y(_2986_));
 sky130_fd_sc_hd__nor2_1 _6623_ (.A(_2983_),
    .B(_2986_),
    .Y(_2987_));
 sky130_fd_sc_hd__and2_1 _6624_ (.A(_2983_),
    .B(_2986_),
    .X(_2988_));
 sky130_fd_sc_hd__or2_1 _6625_ (.A(_2987_),
    .B(_2988_),
    .X(_2989_));
 sky130_fd_sc_hd__o32a_1 _6626_ (.A1(_2970_),
    .A2(_2980_),
    .A3(_2976_),
    .B1(_2979_),
    .B2(_2974_),
    .X(_2990_));
 sky130_fd_sc_hd__nor2_1 _6627_ (.A(_2989_),
    .B(_2990_),
    .Y(_2991_));
 sky130_fd_sc_hd__a21o_1 _6628_ (.A1(_2989_),
    .A2(_2990_),
    .B1(_0866_),
    .X(_2992_));
 sky130_fd_sc_hd__a2bb2o_1 _6629_ (.A1_N(_2991_),
    .A2_N(_2992_),
    .B1(\sound1.sdiv.A[11] ),
    .B2(_2895_),
    .X(_0119_));
 sky130_fd_sc_hd__inv_2 _6630_ (.A(\sound1.sdiv.A[11] ),
    .Y(_2993_));
 sky130_fd_sc_hd__o21a_1 _6631_ (.A1(\sound1.divisor_m[11] ),
    .A2(_2984_),
    .B1(_2903_),
    .X(_2994_));
 sky130_fd_sc_hd__xnor2_1 _6632_ (.A(\sound1.divisor_m[12] ),
    .B(_2994_),
    .Y(_2995_));
 sky130_fd_sc_hd__or2_1 _6633_ (.A(_2993_),
    .B(_2995_),
    .X(_2996_));
 sky130_fd_sc_hd__nand2_1 _6634_ (.A(_2993_),
    .B(_2995_),
    .Y(_2997_));
 sky130_fd_sc_hd__nand2_1 _6635_ (.A(_2996_),
    .B(_2997_),
    .Y(_2998_));
 sky130_fd_sc_hd__or3b_1 _6636_ (.A(_2987_),
    .B(_2991_),
    .C_N(_2998_),
    .X(_2999_));
 sky130_fd_sc_hd__o21bai_2 _6637_ (.A1(_2987_),
    .A2(_2991_),
    .B1_N(_2998_),
    .Y(_3000_));
 sky130_fd_sc_hd__a32o_1 _6638_ (.A1(_2890_),
    .A2(_2999_),
    .A3(_3000_),
    .B1(_2894_),
    .B2(\sound1.sdiv.A[12] ),
    .X(_0120_));
 sky130_fd_sc_hd__inv_2 _6639_ (.A(\sound1.sdiv.A[12] ),
    .Y(_3001_));
 sky130_fd_sc_hd__or3_1 _6640_ (.A(\sound1.divisor_m[12] ),
    .B(\sound1.divisor_m[11] ),
    .C(_2984_),
    .X(_3002_));
 sky130_fd_sc_hd__and2_1 _6641_ (.A(_2903_),
    .B(_3002_),
    .X(_3003_));
 sky130_fd_sc_hd__xnor2_1 _6642_ (.A(\sound1.divisor_m[13] ),
    .B(_3003_),
    .Y(_3004_));
 sky130_fd_sc_hd__or2_1 _6643_ (.A(_3001_),
    .B(_3004_),
    .X(_3005_));
 sky130_fd_sc_hd__nand2_1 _6644_ (.A(_3001_),
    .B(_3004_),
    .Y(_3006_));
 sky130_fd_sc_hd__nand2_1 _6645_ (.A(_3005_),
    .B(_3006_),
    .Y(_3007_));
 sky130_fd_sc_hd__a21o_1 _6646_ (.A1(_2996_),
    .A2(_3000_),
    .B1(_3007_),
    .X(_3008_));
 sky130_fd_sc_hd__nand3_1 _6647_ (.A(_2996_),
    .B(_3000_),
    .C(_3007_),
    .Y(_3009_));
 sky130_fd_sc_hd__a32o_1 _6648_ (.A1(_2890_),
    .A2(_3008_),
    .A3(_3009_),
    .B1(_2894_),
    .B2(\sound1.sdiv.A[13] ),
    .X(_0121_));
 sky130_fd_sc_hd__inv_2 _6649_ (.A(\sound1.sdiv.A[13] ),
    .Y(_3010_));
 sky130_fd_sc_hd__or2_1 _6650_ (.A(\sound1.divisor_m[13] ),
    .B(_3002_),
    .X(_3011_));
 sky130_fd_sc_hd__nand2_1 _6651_ (.A(_2903_),
    .B(_3011_),
    .Y(_3012_));
 sky130_fd_sc_hd__xnor2_1 _6652_ (.A(_2376_),
    .B(_3012_),
    .Y(_3013_));
 sky130_fd_sc_hd__or2_1 _6653_ (.A(_3010_),
    .B(_3013_),
    .X(_3014_));
 sky130_fd_sc_hd__nand2_1 _6654_ (.A(_3010_),
    .B(_3013_),
    .Y(_3015_));
 sky130_fd_sc_hd__nand2_1 _6655_ (.A(_3014_),
    .B(_3015_),
    .Y(_3016_));
 sky130_fd_sc_hd__nand3_1 _6656_ (.A(_3005_),
    .B(_3008_),
    .C(_3016_),
    .Y(_3017_));
 sky130_fd_sc_hd__a21o_1 _6657_ (.A1(_3005_),
    .A2(_3008_),
    .B1(_3016_),
    .X(_3018_));
 sky130_fd_sc_hd__a32o_1 _6658_ (.A1(_2890_),
    .A2(_3017_),
    .A3(_3018_),
    .B1(_2894_),
    .B2(\sound1.sdiv.A[14] ),
    .X(_0122_));
 sky130_fd_sc_hd__inv_2 _6659_ (.A(\sound1.sdiv.A[14] ),
    .Y(_3019_));
 sky130_fd_sc_hd__o21a_1 _6660_ (.A1(\sound1.divisor_m[14] ),
    .A2(_3011_),
    .B1(_2903_),
    .X(_3020_));
 sky130_fd_sc_hd__xnor2_1 _6661_ (.A(\sound1.divisor_m[15] ),
    .B(_3020_),
    .Y(_3021_));
 sky130_fd_sc_hd__or2_1 _6662_ (.A(_3019_),
    .B(_3021_),
    .X(_3022_));
 sky130_fd_sc_hd__nand2_1 _6663_ (.A(_3019_),
    .B(_3021_),
    .Y(_3023_));
 sky130_fd_sc_hd__nand2_1 _6664_ (.A(_3022_),
    .B(_3023_),
    .Y(_3024_));
 sky130_fd_sc_hd__nand3_1 _6665_ (.A(_3014_),
    .B(_3018_),
    .C(_3024_),
    .Y(_3025_));
 sky130_fd_sc_hd__a21o_1 _6666_ (.A1(_3014_),
    .A2(_3018_),
    .B1(_3024_),
    .X(_3026_));
 sky130_fd_sc_hd__a32o_1 _6667_ (.A1(_2890_),
    .A2(_3025_),
    .A3(_3026_),
    .B1(_2894_),
    .B2(\sound1.sdiv.A[15] ),
    .X(_0123_));
 sky130_fd_sc_hd__inv_2 _6668_ (.A(\sound1.sdiv.A[15] ),
    .Y(_3027_));
 sky130_fd_sc_hd__or3_1 _6669_ (.A(\sound1.divisor_m[15] ),
    .B(\sound1.divisor_m[14] ),
    .C(_3011_),
    .X(_3028_));
 sky130_fd_sc_hd__and2_1 _6670_ (.A(_2903_),
    .B(_3028_),
    .X(_3029_));
 sky130_fd_sc_hd__xnor2_1 _6671_ (.A(\sound1.divisor_m[16] ),
    .B(_3029_),
    .Y(_3030_));
 sky130_fd_sc_hd__or2_1 _6672_ (.A(_3027_),
    .B(_3030_),
    .X(_3031_));
 sky130_fd_sc_hd__nand2_1 _6673_ (.A(_3027_),
    .B(_3030_),
    .Y(_3032_));
 sky130_fd_sc_hd__nand2_1 _6674_ (.A(_3031_),
    .B(_3032_),
    .Y(_3033_));
 sky130_fd_sc_hd__nand3_1 _6675_ (.A(_3022_),
    .B(_3026_),
    .C(_3033_),
    .Y(_3034_));
 sky130_fd_sc_hd__a21o_1 _6676_ (.A1(_3022_),
    .A2(_3026_),
    .B1(_3033_),
    .X(_3035_));
 sky130_fd_sc_hd__a32o_1 _6677_ (.A1(_2890_),
    .A2(_3034_),
    .A3(_3035_),
    .B1(_2894_),
    .B2(\sound1.sdiv.A[16] ),
    .X(_0124_));
 sky130_fd_sc_hd__or2_1 _6678_ (.A(\sound1.divisor_m[16] ),
    .B(_3028_),
    .X(_3036_));
 sky130_fd_sc_hd__and2_1 _6679_ (.A(_2903_),
    .B(_3036_),
    .X(_3037_));
 sky130_fd_sc_hd__xnor2_1 _6680_ (.A(\sound1.divisor_m[17] ),
    .B(_3037_),
    .Y(_3038_));
 sky130_fd_sc_hd__inv_2 _6681_ (.A(_3038_),
    .Y(_3039_));
 sky130_fd_sc_hd__nand2_1 _6682_ (.A(\sound1.sdiv.A[16] ),
    .B(_3039_),
    .Y(_3040_));
 sky130_fd_sc_hd__or2_1 _6683_ (.A(\sound1.sdiv.A[16] ),
    .B(_3039_),
    .X(_3041_));
 sky130_fd_sc_hd__nand2_1 _6684_ (.A(_3040_),
    .B(_3041_),
    .Y(_3042_));
 sky130_fd_sc_hd__nand2_1 _6685_ (.A(_3031_),
    .B(_3035_),
    .Y(_3043_));
 sky130_fd_sc_hd__xnor2_1 _6686_ (.A(_3042_),
    .B(_3043_),
    .Y(_3044_));
 sky130_fd_sc_hd__a22o_1 _6687_ (.A1(\sound1.sdiv.A[17] ),
    .A2(_2895_),
    .B1(\sound1.sdiv.next_dived ),
    .B2(_3044_),
    .X(_0125_));
 sky130_fd_sc_hd__inv_2 _6688_ (.A(\sound1.sdiv.A[17] ),
    .Y(_3045_));
 sky130_fd_sc_hd__o21a_1 _6689_ (.A1(\sound1.divisor_m[17] ),
    .A2(_3036_),
    .B1(_2903_),
    .X(_3046_));
 sky130_fd_sc_hd__xnor2_1 _6690_ (.A(\sound1.divisor_m[18] ),
    .B(_3046_),
    .Y(_3047_));
 sky130_fd_sc_hd__or2_1 _6691_ (.A(_3045_),
    .B(_3047_),
    .X(_3048_));
 sky130_fd_sc_hd__nand2_1 _6692_ (.A(_3045_),
    .B(_3047_),
    .Y(_3049_));
 sky130_fd_sc_hd__nand2_1 _6693_ (.A(_3048_),
    .B(_3049_),
    .Y(_3050_));
 sky130_fd_sc_hd__a21boi_1 _6694_ (.A1(_3041_),
    .A2(_3043_),
    .B1_N(_3040_),
    .Y(_3051_));
 sky130_fd_sc_hd__nand2_1 _6695_ (.A(_3050_),
    .B(_3051_),
    .Y(_3052_));
 sky130_fd_sc_hd__or2_1 _6696_ (.A(_3050_),
    .B(_3051_),
    .X(_3053_));
 sky130_fd_sc_hd__a32o_1 _6697_ (.A1(_2890_),
    .A2(_3052_),
    .A3(_3053_),
    .B1(_2894_),
    .B2(\sound1.sdiv.A[18] ),
    .X(_0126_));
 sky130_fd_sc_hd__o31a_1 _6698_ (.A1(\sound1.divisor_m[18] ),
    .A2(\sound1.divisor_m[17] ),
    .A3(_3036_),
    .B1(_2903_),
    .X(_3054_));
 sky130_fd_sc_hd__buf_4 _6699_ (.A(_3054_),
    .X(_3055_));
 sky130_fd_sc_hd__nor2_1 _6700_ (.A(\sound1.sdiv.A[18] ),
    .B(_3055_),
    .Y(_3056_));
 sky130_fd_sc_hd__nand2_1 _6701_ (.A(\sound1.sdiv.A[18] ),
    .B(_3055_),
    .Y(_3057_));
 sky130_fd_sc_hd__or2b_1 _6702_ (.A(_3056_),
    .B_N(_3057_),
    .X(_3058_));
 sky130_fd_sc_hd__o21ai_1 _6703_ (.A1(_3050_),
    .A2(_3051_),
    .B1(_3048_),
    .Y(_3059_));
 sky130_fd_sc_hd__xnor2_1 _6704_ (.A(_3058_),
    .B(_3059_),
    .Y(_3060_));
 sky130_fd_sc_hd__a22o_1 _6705_ (.A1(\sound1.sdiv.A[19] ),
    .A2(_2895_),
    .B1(\sound1.sdiv.next_dived ),
    .B2(_3060_),
    .X(_0127_));
 sky130_fd_sc_hd__a21bo_1 _6706_ (.A1(_3031_),
    .A2(_3040_),
    .B1_N(_3041_),
    .X(_3061_));
 sky130_fd_sc_hd__o21a_1 _6707_ (.A1(_3048_),
    .A2(_3056_),
    .B1(_3057_),
    .X(_3062_));
 sky130_fd_sc_hd__o31a_1 _6708_ (.A1(_3050_),
    .A2(_3061_),
    .A3(_3058_),
    .B1(_3062_),
    .X(_3063_));
 sky130_fd_sc_hd__or2_1 _6709_ (.A(_3050_),
    .B(_3058_),
    .X(_3064_));
 sky130_fd_sc_hd__a2111o_1 _6710_ (.A1(_3022_),
    .A2(_3026_),
    .B1(_3033_),
    .C1(_3042_),
    .D1(_3064_),
    .X(_3065_));
 sky130_fd_sc_hd__or2_1 _6711_ (.A(\sound1.sdiv.A[19] ),
    .B(_3055_),
    .X(_3066_));
 sky130_fd_sc_hd__nand2_1 _6712_ (.A(\sound1.sdiv.A[19] ),
    .B(_3055_),
    .Y(_3067_));
 sky130_fd_sc_hd__nand2_1 _6713_ (.A(_3066_),
    .B(_3067_),
    .Y(_3068_));
 sky130_fd_sc_hd__a21o_1 _6714_ (.A1(_3063_),
    .A2(_3065_),
    .B1(_3068_),
    .X(_3069_));
 sky130_fd_sc_hd__and3_1 _6715_ (.A(_3068_),
    .B(_3063_),
    .C(_3065_),
    .X(_3070_));
 sky130_fd_sc_hd__nor2_1 _6716_ (.A(_0866_),
    .B(_3070_),
    .Y(_3071_));
 sky130_fd_sc_hd__a22o_1 _6717_ (.A1(\sound1.sdiv.A[20] ),
    .A2(_2895_),
    .B1(_3069_),
    .B2(_3071_),
    .X(_0128_));
 sky130_fd_sc_hd__xor2_1 _6718_ (.A(\sound1.sdiv.A[20] ),
    .B(_3055_),
    .X(_3072_));
 sky130_fd_sc_hd__inv_2 _6719_ (.A(_3072_),
    .Y(_3073_));
 sky130_fd_sc_hd__a21oi_1 _6720_ (.A1(_3067_),
    .A2(_3069_),
    .B1(_3073_),
    .Y(_3074_));
 sky130_fd_sc_hd__a31o_1 _6721_ (.A1(_3067_),
    .A2(_3069_),
    .A3(_3073_),
    .B1(_0866_),
    .X(_3075_));
 sky130_fd_sc_hd__a2bb2o_1 _6722_ (.A1_N(_3074_),
    .A2_N(_3075_),
    .B1(\sound1.sdiv.A[21] ),
    .B2(_2895_),
    .X(_0129_));
 sky130_fd_sc_hd__o21bai_1 _6723_ (.A1(\sound1.sdiv.A[20] ),
    .A2(_3055_),
    .B1_N(_3069_),
    .Y(_3076_));
 sky130_fd_sc_hd__o21ai_1 _6724_ (.A1(\sound1.sdiv.A[20] ),
    .A2(\sound1.sdiv.A[19] ),
    .B1(_3055_),
    .Y(_3077_));
 sky130_fd_sc_hd__xnor2_1 _6725_ (.A(\sound1.sdiv.A[21] ),
    .B(_3055_),
    .Y(_3078_));
 sky130_fd_sc_hd__a21oi_1 _6726_ (.A1(_3076_),
    .A2(_3077_),
    .B1(_3078_),
    .Y(_3079_));
 sky130_fd_sc_hd__a31o_1 _6727_ (.A1(_3078_),
    .A2(_3076_),
    .A3(_3077_),
    .B1(_0866_),
    .X(_3080_));
 sky130_fd_sc_hd__a2bb2o_1 _6728_ (.A1_N(_3079_),
    .A2_N(_3080_),
    .B1(\sound1.sdiv.A[22] ),
    .B2(_2895_),
    .X(_0130_));
 sky130_fd_sc_hd__xor2_1 _6729_ (.A(\sound1.sdiv.A[22] ),
    .B(_3055_),
    .X(_3081_));
 sky130_fd_sc_hd__a21oi_1 _6730_ (.A1(\sound1.sdiv.A[21] ),
    .A2(_3055_),
    .B1(_3079_),
    .Y(_3082_));
 sky130_fd_sc_hd__xnor2_1 _6731_ (.A(_3081_),
    .B(_3082_),
    .Y(_3083_));
 sky130_fd_sc_hd__a22o_1 _6732_ (.A1(\sound1.sdiv.A[23] ),
    .A2(_2895_),
    .B1(\sound1.sdiv.next_dived ),
    .B2(_3083_),
    .X(_0131_));
 sky130_fd_sc_hd__or2_1 _6733_ (.A(\sound1.sdiv.A[23] ),
    .B(_3055_),
    .X(_3084_));
 sky130_fd_sc_hd__nand2_1 _6734_ (.A(\sound1.sdiv.A[23] ),
    .B(_3055_),
    .Y(_3085_));
 sky130_fd_sc_hd__nor4b_1 _6735_ (.A(_3069_),
    .B(_3073_),
    .C(_3078_),
    .D_N(_3081_),
    .Y(_3086_));
 sky130_fd_sc_hd__o41a_1 _6736_ (.A1(\sound1.sdiv.A[22] ),
    .A2(\sound1.sdiv.A[21] ),
    .A3(\sound1.sdiv.A[20] ),
    .A4(\sound1.sdiv.A[19] ),
    .B1(_3055_),
    .X(_3087_));
 sky130_fd_sc_hd__a211o_1 _6737_ (.A1(_3084_),
    .A2(_3085_),
    .B1(net55),
    .C1(_3087_),
    .X(_3088_));
 sky130_fd_sc_hd__o211a_1 _6738_ (.A1(net55),
    .A2(_3087_),
    .B1(_3084_),
    .C1(_3085_),
    .X(_3089_));
 sky130_fd_sc_hd__nor2_1 _6739_ (.A(_0866_),
    .B(_3089_),
    .Y(_3090_));
 sky130_fd_sc_hd__a22o_1 _6740_ (.A1(\sound1.sdiv.A[24] ),
    .A2(_2895_),
    .B1(_3088_),
    .B2(_3090_),
    .X(_0132_));
 sky130_fd_sc_hd__a21oi_1 _6741_ (.A1(\sound1.sdiv.A[23] ),
    .A2(_3055_),
    .B1(_3089_),
    .Y(_3091_));
 sky130_fd_sc_hd__or2_1 _6742_ (.A(\sound1.sdiv.A[24] ),
    .B(_3055_),
    .X(_3092_));
 sky130_fd_sc_hd__nand2_1 _6743_ (.A(\sound1.sdiv.A[24] ),
    .B(_3055_),
    .Y(_3093_));
 sky130_fd_sc_hd__and2_1 _6744_ (.A(_3092_),
    .B(_3093_),
    .X(_3094_));
 sky130_fd_sc_hd__xnor2_1 _6745_ (.A(_3091_),
    .B(_3094_),
    .Y(_3095_));
 sky130_fd_sc_hd__a22o_1 _6746_ (.A1(\sound1.sdiv.A[25] ),
    .A2(_2895_),
    .B1(\sound1.sdiv.next_dived ),
    .B2(_3095_),
    .X(_0133_));
 sky130_fd_sc_hd__nand2_1 _6747_ (.A(\sound1.sdiv.A[25] ),
    .B(_3055_),
    .Y(_3096_));
 sky130_fd_sc_hd__or2_1 _6748_ (.A(\sound1.sdiv.A[25] ),
    .B(_3055_),
    .X(_3097_));
 sky130_fd_sc_hd__nand2_1 _6749_ (.A(_3096_),
    .B(_3097_),
    .Y(_3098_));
 sky130_fd_sc_hd__o21a_1 _6750_ (.A1(\sound1.sdiv.A[24] ),
    .A2(\sound1.sdiv.A[23] ),
    .B1(_3055_),
    .X(_3099_));
 sky130_fd_sc_hd__a21oi_1 _6751_ (.A1(_3089_),
    .A2(_3092_),
    .B1(_3099_),
    .Y(_3100_));
 sky130_fd_sc_hd__xor2_1 _6752_ (.A(_3098_),
    .B(_3100_),
    .X(_3101_));
 sky130_fd_sc_hd__a22o_1 _6753_ (.A1(\sound1.sdiv.A[26] ),
    .A2(_2895_),
    .B1(\sound1.sdiv.next_dived ),
    .B2(_3101_),
    .X(_0134_));
 sky130_fd_sc_hd__mux2_1 _6754_ (.A0(_0867_),
    .A1(_2893_),
    .S(\sound1.sdiv.C[0] ),
    .X(_3102_));
 sky130_fd_sc_hd__clkbuf_1 _6755_ (.A(_3102_),
    .X(_0135_));
 sky130_fd_sc_hd__nand2_1 _6756_ (.A(\sound1.sdiv.C[1] ),
    .B(\sound1.sdiv.C[0] ),
    .Y(_3103_));
 sky130_fd_sc_hd__or2_1 _6757_ (.A(\sound1.sdiv.C[1] ),
    .B(\sound1.sdiv.C[0] ),
    .X(_3104_));
 sky130_fd_sc_hd__a32o_1 _6758_ (.A1(_2890_),
    .A2(_3103_),
    .A3(_3104_),
    .B1(_2894_),
    .B2(\sound1.sdiv.C[1] ),
    .X(_0136_));
 sky130_fd_sc_hd__a21o_1 _6759_ (.A1(\sound1.sdiv.C[1] ),
    .A2(\sound1.sdiv.C[0] ),
    .B1(\sound1.sdiv.C[2] ),
    .X(_3105_));
 sky130_fd_sc_hd__and3_1 _6760_ (.A(\sound1.sdiv.C[2] ),
    .B(\sound1.sdiv.C[1] ),
    .C(\sound1.sdiv.C[0] ),
    .X(_3106_));
 sky130_fd_sc_hd__inv_2 _6761_ (.A(_3106_),
    .Y(_3107_));
 sky130_fd_sc_hd__a32o_1 _6762_ (.A1(_2890_),
    .A2(_3105_),
    .A3(_3107_),
    .B1(_2894_),
    .B2(\sound1.sdiv.C[2] ),
    .X(_0137_));
 sky130_fd_sc_hd__and3_1 _6763_ (.A(\sound1.sdiv.C[3] ),
    .B(_0565_),
    .C(_3106_),
    .X(_3108_));
 sky130_fd_sc_hd__a21oi_1 _6764_ (.A1(_0565_),
    .A2(_3106_),
    .B1(\sound1.sdiv.C[3] ),
    .Y(_3109_));
 sky130_fd_sc_hd__nor3_1 _6765_ (.A(_2005_),
    .B(_3108_),
    .C(_3109_),
    .Y(_0138_));
 sky130_fd_sc_hd__a31o_1 _6766_ (.A1(\sound1.sdiv.C[3] ),
    .A2(_0565_),
    .A3(_3106_),
    .B1(\sound1.sdiv.C[4] ),
    .X(_3110_));
 sky130_fd_sc_hd__and2_1 _6767_ (.A(_2843_),
    .B(_3110_),
    .X(_3111_));
 sky130_fd_sc_hd__clkbuf_1 _6768_ (.A(_3111_),
    .X(_0139_));
 sky130_fd_sc_hd__and2_1 _6769_ (.A(\sound1.sdiv.C[5] ),
    .B(_2843_),
    .X(_3112_));
 sky130_fd_sc_hd__clkbuf_1 _6770_ (.A(_3112_),
    .X(_0140_));
 sky130_fd_sc_hd__or4_1 _6771_ (.A(\sound1.divisor_m[18] ),
    .B(\sound1.divisor_m[17] ),
    .C(\sound1.sdiv.A[26] ),
    .D(_3036_),
    .X(_3113_));
 sky130_fd_sc_hd__o211a_1 _6772_ (.A1(_3098_),
    .A2(_3100_),
    .B1(_3113_),
    .C1(_3096_),
    .X(_3114_));
 sky130_fd_sc_hd__o21ai_1 _6773_ (.A1(_0866_),
    .A2(_3114_),
    .B1(_2277_),
    .Y(_0141_));
 sky130_fd_sc_hd__a21o_1 _6774_ (.A1(\sound1.sdiv.Q[0] ),
    .A2(\sound1.sdiv.next_dived ),
    .B1(_2436_),
    .X(_0142_));
 sky130_fd_sc_hd__o21ai_1 _6775_ (.A1(_2435_),
    .A2(_0866_),
    .B1(_2588_),
    .Y(_0143_));
 sky130_fd_sc_hd__a22o_1 _6776_ (.A1(\sound1.sdiv.Q[3] ),
    .A2(_2895_),
    .B1(\sound1.sdiv.next_dived ),
    .B2(\sound1.sdiv.Q[2] ),
    .X(_0144_));
 sky130_fd_sc_hd__a22o_1 _6777_ (.A1(\sound1.sdiv.Q[4] ),
    .A2(_2894_),
    .B1(\sound1.sdiv.next_dived ),
    .B2(\sound1.sdiv.Q[3] ),
    .X(_0145_));
 sky130_fd_sc_hd__a22o_1 _6778_ (.A1(\sound1.sdiv.Q[5] ),
    .A2(_2894_),
    .B1(\sound1.sdiv.next_dived ),
    .B2(\sound1.sdiv.Q[4] ),
    .X(_0146_));
 sky130_fd_sc_hd__a22o_1 _6779_ (.A1(\sound1.sdiv.Q[6] ),
    .A2(_2894_),
    .B1(_2890_),
    .B2(\sound1.sdiv.Q[5] ),
    .X(_0147_));
 sky130_fd_sc_hd__a22o_1 _6780_ (.A1(\sound1.sdiv.Q[7] ),
    .A2(_2894_),
    .B1(_2890_),
    .B2(\sound1.sdiv.Q[6] ),
    .X(_0148_));
 sky130_fd_sc_hd__a221o_1 _6781_ (.A1(\sound1.sdiv.Q[8] ),
    .A2(_2894_),
    .B1(_2890_),
    .B2(\sound1.sdiv.Q[7] ),
    .C1(_2837_),
    .X(_0149_));
 sky130_fd_sc_hd__a221o_1 _6782_ (.A1(\sound1.sdiv.Q[9] ),
    .A2(_2894_),
    .B1(_2890_),
    .B2(\sound1.sdiv.Q[8] ),
    .C1(_2838_),
    .X(_0150_));
 sky130_fd_sc_hd__a221o_1 _6783_ (.A1(\sound1.sdiv.Q[10] ),
    .A2(_2894_),
    .B1(_2890_),
    .B2(\sound1.sdiv.Q[9] ),
    .C1(_2839_),
    .X(_0151_));
 sky130_fd_sc_hd__a221o_1 _6784_ (.A1(\sound1.sdiv.Q[11] ),
    .A2(_2893_),
    .B1(_2890_),
    .B2(\sound1.sdiv.Q[10] ),
    .C1(_2840_),
    .X(_0152_));
 sky130_fd_sc_hd__a221o_1 _6785_ (.A1(\sound1.sdiv.Q[12] ),
    .A2(_2893_),
    .B1(_2890_),
    .B2(\sound1.sdiv.Q[11] ),
    .C1(_2841_),
    .X(_0153_));
 sky130_fd_sc_hd__a221o_1 _6786_ (.A1(\sound1.sdiv.Q[13] ),
    .A2(_2893_),
    .B1(_2890_),
    .B2(\sound1.sdiv.Q[12] ),
    .C1(_2842_),
    .X(_0154_));
 sky130_fd_sc_hd__a221o_1 _6787_ (.A1(\sound1.sdiv.Q[14] ),
    .A2(_2893_),
    .B1(_0867_),
    .B2(\sound1.sdiv.Q[13] ),
    .C1(_2844_),
    .X(_0155_));
 sky130_fd_sc_hd__a221o_1 _6788_ (.A1(\sound1.sdiv.Q[15] ),
    .A2(_2893_),
    .B1(_0867_),
    .B2(\sound1.sdiv.Q[14] ),
    .C1(_2845_),
    .X(_0156_));
 sky130_fd_sc_hd__a221o_1 _6789_ (.A1(\sound1.sdiv.Q[16] ),
    .A2(_2893_),
    .B1(_0867_),
    .B2(\sound1.sdiv.Q[15] ),
    .C1(_2846_),
    .X(_0157_));
 sky130_fd_sc_hd__a221o_1 _6790_ (.A1(\sound1.sdiv.Q[17] ),
    .A2(_2893_),
    .B1(_0867_),
    .B2(\sound1.sdiv.Q[16] ),
    .C1(_2847_),
    .X(_0158_));
 sky130_fd_sc_hd__a221o_1 _6791_ (.A1(\sound1.sdiv.Q[18] ),
    .A2(_2893_),
    .B1(_0867_),
    .B2(\sound1.sdiv.Q[17] ),
    .C1(_2848_),
    .X(_0159_));
 sky130_fd_sc_hd__a221o_1 _6792_ (.A1(\sound1.sdiv.Q[19] ),
    .A2(_2893_),
    .B1(_0867_),
    .B2(\sound1.sdiv.Q[18] ),
    .C1(_2849_),
    .X(_0160_));
 sky130_fd_sc_hd__a221o_1 _6793_ (.A1(\sound1.sdiv.Q[20] ),
    .A2(_2893_),
    .B1(_0867_),
    .B2(\sound1.sdiv.Q[19] ),
    .C1(_2850_),
    .X(_0161_));
 sky130_fd_sc_hd__a221o_1 _6794_ (.A1(\sound1.sdiv.Q[21] ),
    .A2(_2893_),
    .B1(_0867_),
    .B2(\sound1.sdiv.Q[20] ),
    .C1(_2851_),
    .X(_0162_));
 sky130_fd_sc_hd__a221o_1 _6795_ (.A1(\sound1.sdiv.Q[22] ),
    .A2(_2893_),
    .B1(_0867_),
    .B2(\sound1.sdiv.Q[21] ),
    .C1(_2852_),
    .X(_0163_));
 sky130_fd_sc_hd__a221o_1 _6796_ (.A1(\sound1.sdiv.Q[23] ),
    .A2(_2893_),
    .B1(_0867_),
    .B2(\sound1.sdiv.Q[22] ),
    .C1(_2853_),
    .X(_0164_));
 sky130_fd_sc_hd__a221o_1 _6797_ (.A1(\sound1.sdiv.Q[24] ),
    .A2(_2893_),
    .B1(_0867_),
    .B2(\sound1.sdiv.Q[23] ),
    .C1(_2854_),
    .X(_0165_));
 sky130_fd_sc_hd__a221o_1 _6798_ (.A1(\sound1.sdiv.Q[25] ),
    .A2(_2893_),
    .B1(_0867_),
    .B2(\sound1.sdiv.Q[24] ),
    .C1(_2856_),
    .X(_0166_));
 sky130_fd_sc_hd__a221o_1 _6799_ (.A1(\sound1.sdiv.Q[26] ),
    .A2(_2893_),
    .B1(_0867_),
    .B2(\sound1.sdiv.Q[25] ),
    .C1(_2858_),
    .X(_0167_));
 sky130_fd_sc_hd__a22o_1 _6800_ (.A1(\sound1.sdiv.Q[27] ),
    .A2(_2894_),
    .B1(_2890_),
    .B2(\sound1.sdiv.Q[26] ),
    .X(_0168_));
 sky130_fd_sc_hd__and2_1 _6801_ (.A(\sound2.count[0] ),
    .B(_2855_),
    .X(_3115_));
 sky130_fd_sc_hd__a21o_1 _6802_ (.A1(\sound2.count_m[0] ),
    .A2(_2857_),
    .B1(_3115_),
    .X(_0169_));
 sky130_fd_sc_hd__and2_1 _6803_ (.A(\sound2.count[1] ),
    .B(_2855_),
    .X(_3116_));
 sky130_fd_sc_hd__a21o_1 _6804_ (.A1(\sound2.count_m[1] ),
    .A2(_2857_),
    .B1(_3116_),
    .X(_0170_));
 sky130_fd_sc_hd__nor2_1 _6805_ (.A(_1470_),
    .B(_2843_),
    .Y(_3117_));
 sky130_fd_sc_hd__a21o_1 _6806_ (.A1(\sound2.count_m[2] ),
    .A2(_2857_),
    .B1(_3117_),
    .X(_0171_));
 sky130_fd_sc_hd__nor2_1 _6807_ (.A(_1318_),
    .B(_2843_),
    .Y(_3118_));
 sky130_fd_sc_hd__a21o_1 _6808_ (.A1(\sound2.count_m[3] ),
    .A2(_2857_),
    .B1(_3118_),
    .X(_0172_));
 sky130_fd_sc_hd__and2_1 _6809_ (.A(\sound2.count[4] ),
    .B(_2855_),
    .X(_3119_));
 sky130_fd_sc_hd__a21o_1 _6810_ (.A1(\sound2.count_m[4] ),
    .A2(_2857_),
    .B1(_3119_),
    .X(_0173_));
 sky130_fd_sc_hd__and2_1 _6811_ (.A(\sound2.count[5] ),
    .B(_2855_),
    .X(_3120_));
 sky130_fd_sc_hd__a21o_1 _6812_ (.A1(\sound2.count_m[5] ),
    .A2(_2857_),
    .B1(_3120_),
    .X(_0174_));
 sky130_fd_sc_hd__and2_1 _6813_ (.A(\sound2.count[6] ),
    .B(_2855_),
    .X(_3121_));
 sky130_fd_sc_hd__a21o_1 _6814_ (.A1(\sound2.count_m[6] ),
    .A2(_2857_),
    .B1(_3121_),
    .X(_0175_));
 sky130_fd_sc_hd__and2_1 _6815_ (.A(\sound2.count[7] ),
    .B(_2855_),
    .X(_3122_));
 sky130_fd_sc_hd__a21o_1 _6816_ (.A1(\sound2.count_m[7] ),
    .A2(_2857_),
    .B1(_3122_),
    .X(_0176_));
 sky130_fd_sc_hd__and2_1 _6817_ (.A(\sound2.count[8] ),
    .B(_2855_),
    .X(_3123_));
 sky130_fd_sc_hd__a21o_1 _6818_ (.A1(\sound2.count_m[8] ),
    .A2(_2857_),
    .B1(_3123_),
    .X(_0177_));
 sky130_fd_sc_hd__and2_1 _6819_ (.A(\sound2.count[9] ),
    .B(_2855_),
    .X(_3124_));
 sky130_fd_sc_hd__a21o_1 _6820_ (.A1(\sound2.count_m[9] ),
    .A2(_2857_),
    .B1(_3124_),
    .X(_0178_));
 sky130_fd_sc_hd__and2_1 _6821_ (.A(\sound2.count[10] ),
    .B(_2855_),
    .X(_3125_));
 sky130_fd_sc_hd__a21o_1 _6822_ (.A1(\sound2.count_m[10] ),
    .A2(_2857_),
    .B1(_3125_),
    .X(_0179_));
 sky130_fd_sc_hd__and2_1 _6823_ (.A(\sound2.count[11] ),
    .B(_2855_),
    .X(_3126_));
 sky130_fd_sc_hd__a21o_1 _6824_ (.A1(\sound2.count_m[11] ),
    .A2(_2857_),
    .B1(_3126_),
    .X(_0180_));
 sky130_fd_sc_hd__and2_1 _6825_ (.A(\sound2.count[12] ),
    .B(_2855_),
    .X(_3127_));
 sky130_fd_sc_hd__a21o_1 _6826_ (.A1(\sound2.count_m[12] ),
    .A2(_2857_),
    .B1(_3127_),
    .X(_0181_));
 sky130_fd_sc_hd__and2_1 _6827_ (.A(\sound2.count[13] ),
    .B(_2855_),
    .X(_3128_));
 sky130_fd_sc_hd__a21o_1 _6828_ (.A1(\sound2.count_m[13] ),
    .A2(_2857_),
    .B1(_3128_),
    .X(_0182_));
 sky130_fd_sc_hd__and2_1 _6829_ (.A(\sound2.count[14] ),
    .B(_2855_),
    .X(_3129_));
 sky130_fd_sc_hd__a21o_1 _6830_ (.A1(\sound2.count_m[14] ),
    .A2(_2857_),
    .B1(_3129_),
    .X(_0183_));
 sky130_fd_sc_hd__and2_1 _6831_ (.A(\sound2.count[15] ),
    .B(_2855_),
    .X(_3130_));
 sky130_fd_sc_hd__a21o_1 _6832_ (.A1(\sound2.count_m[15] ),
    .A2(_2857_),
    .B1(_3130_),
    .X(_0184_));
 sky130_fd_sc_hd__and2_1 _6833_ (.A(\sound2.count[16] ),
    .B(_2855_),
    .X(_3131_));
 sky130_fd_sc_hd__a21o_1 _6834_ (.A1(\sound2.count_m[16] ),
    .A2(_2857_),
    .B1(_3131_),
    .X(_0185_));
 sky130_fd_sc_hd__buf_6 _6835_ (.A(_0554_),
    .X(_3132_));
 sky130_fd_sc_hd__and2_1 _6836_ (.A(\sound2.count[17] ),
    .B(_2855_),
    .X(_3133_));
 sky130_fd_sc_hd__a21o_1 _6837_ (.A1(\sound2.count_m[17] ),
    .A2(_3132_),
    .B1(_3133_),
    .X(_0186_));
 sky130_fd_sc_hd__and2_1 _6838_ (.A(\sound2.count[18] ),
    .B(_2855_),
    .X(_3134_));
 sky130_fd_sc_hd__a21o_1 _6839_ (.A1(\sound2.count_m[18] ),
    .A2(_3132_),
    .B1(_3134_),
    .X(_0187_));
 sky130_fd_sc_hd__mux2_1 _6840_ (.A0(\sound2.divisor_m[0] ),
    .A1(_1477_),
    .S(_2864_),
    .X(_3135_));
 sky130_fd_sc_hd__clkbuf_1 _6841_ (.A(_3135_),
    .X(_0188_));
 sky130_fd_sc_hd__inv_2 _6842_ (.A(_1404_),
    .Y(_3136_));
 sky130_fd_sc_hd__mux2_1 _6843_ (.A0(\sound2.divisor_m[1] ),
    .A1(_3136_),
    .S(_2864_),
    .X(_3137_));
 sky130_fd_sc_hd__clkbuf_1 _6844_ (.A(_3137_),
    .X(_0189_));
 sky130_fd_sc_hd__mux2_1 _6845_ (.A0(\sound2.divisor_m[2] ),
    .A1(_1469_),
    .S(_2864_),
    .X(_3138_));
 sky130_fd_sc_hd__clkbuf_1 _6846_ (.A(_3138_),
    .X(_0190_));
 sky130_fd_sc_hd__mux2_1 _6847_ (.A0(\sound2.divisor_m[3] ),
    .A1(_1352_),
    .S(_2864_),
    .X(_3139_));
 sky130_fd_sc_hd__clkbuf_1 _6848_ (.A(_3139_),
    .X(_0191_));
 sky130_fd_sc_hd__mux2_1 _6849_ (.A0(\sound2.divisor_m[4] ),
    .A1(_1441_),
    .S(_2864_),
    .X(_3140_));
 sky130_fd_sc_hd__clkbuf_1 _6850_ (.A(_3140_),
    .X(_0192_));
 sky130_fd_sc_hd__inv_2 _6851_ (.A(_1396_),
    .Y(_3141_));
 sky130_fd_sc_hd__buf_8 _6852_ (.A(_2863_),
    .X(_3142_));
 sky130_fd_sc_hd__mux2_1 _6853_ (.A0(\sound2.divisor_m[5] ),
    .A1(_3141_),
    .S(_3142_),
    .X(_3143_));
 sky130_fd_sc_hd__clkbuf_1 _6854_ (.A(_3143_),
    .X(_0193_));
 sky130_fd_sc_hd__mux2_1 _6855_ (.A0(\sound2.divisor_m[6] ),
    .A1(_1378_),
    .S(_3142_),
    .X(_3144_));
 sky130_fd_sc_hd__clkbuf_1 _6856_ (.A(_3144_),
    .X(_0194_));
 sky130_fd_sc_hd__inv_2 _6857_ (.A(_1368_),
    .Y(_3145_));
 sky130_fd_sc_hd__mux2_1 _6858_ (.A0(\sound2.divisor_m[7] ),
    .A1(_3145_),
    .S(_3142_),
    .X(_3146_));
 sky130_fd_sc_hd__clkbuf_1 _6859_ (.A(_3146_),
    .X(_0195_));
 sky130_fd_sc_hd__inv_2 _6860_ (.A(_1412_),
    .Y(_3147_));
 sky130_fd_sc_hd__mux2_1 _6861_ (.A0(\sound2.divisor_m[8] ),
    .A1(_3147_),
    .S(_3142_),
    .X(_3148_));
 sky130_fd_sc_hd__clkbuf_1 _6862_ (.A(_3148_),
    .X(_0196_));
 sky130_fd_sc_hd__inv_2 _6863_ (.A(_1495_),
    .Y(_3149_));
 sky130_fd_sc_hd__mux2_1 _6864_ (.A0(\sound2.divisor_m[9] ),
    .A1(_3149_),
    .S(_3142_),
    .X(_3150_));
 sky130_fd_sc_hd__clkbuf_1 _6865_ (.A(_3150_),
    .X(_0197_));
 sky130_fd_sc_hd__inv_2 _6866_ (.A(_1387_),
    .Y(_3151_));
 sky130_fd_sc_hd__mux2_1 _6867_ (.A0(\sound2.divisor_m[10] ),
    .A1(_3151_),
    .S(_3142_),
    .X(_3152_));
 sky130_fd_sc_hd__clkbuf_1 _6868_ (.A(_3152_),
    .X(_0198_));
 sky130_fd_sc_hd__inv_2 _6869_ (.A(_1488_),
    .Y(_3153_));
 sky130_fd_sc_hd__mux2_1 _6870_ (.A0(\sound2.divisor_m[11] ),
    .A1(_3153_),
    .S(_3142_),
    .X(_3154_));
 sky130_fd_sc_hd__clkbuf_1 _6871_ (.A(_3154_),
    .X(_0199_));
 sky130_fd_sc_hd__inv_2 _6872_ (.A(_1360_),
    .Y(_3155_));
 sky130_fd_sc_hd__mux2_1 _6873_ (.A0(\sound2.divisor_m[12] ),
    .A1(_3155_),
    .S(_3142_),
    .X(_3156_));
 sky130_fd_sc_hd__clkbuf_1 _6874_ (.A(_3156_),
    .X(_0200_));
 sky130_fd_sc_hd__inv_2 _6875_ (.A(_1434_),
    .Y(_3157_));
 sky130_fd_sc_hd__mux2_1 _6876_ (.A0(\sound2.divisor_m[13] ),
    .A1(_3157_),
    .S(_3142_),
    .X(_3158_));
 sky130_fd_sc_hd__clkbuf_1 _6877_ (.A(_3158_),
    .X(_0201_));
 sky130_fd_sc_hd__mux2_1 _6878_ (.A0(\sound2.divisor_m[14] ),
    .A1(_1422_),
    .S(_3142_),
    .X(_3159_));
 sky130_fd_sc_hd__clkbuf_1 _6879_ (.A(_3159_),
    .X(_0202_));
 sky130_fd_sc_hd__mux2_1 _6880_ (.A0(\sound2.divisor_m[15] ),
    .A1(_1454_),
    .S(_3142_),
    .X(_3160_));
 sky130_fd_sc_hd__clkbuf_1 _6881_ (.A(_3160_),
    .X(_0203_));
 sky130_fd_sc_hd__mux2_1 _6882_ (.A0(\sound2.divisor_m[16] ),
    .A1(_1459_),
    .S(_3142_),
    .X(_3161_));
 sky130_fd_sc_hd__clkbuf_1 _6883_ (.A(_3161_),
    .X(_0204_));
 sky130_fd_sc_hd__mux2_1 _6884_ (.A0(\sound2.divisor_m[17] ),
    .A1(_1446_),
    .S(_3142_),
    .X(_3162_));
 sky130_fd_sc_hd__clkbuf_1 _6885_ (.A(_3162_),
    .X(_0205_));
 sky130_fd_sc_hd__or2_1 _6886_ (.A(_2470_),
    .B(_2005_),
    .X(_3163_));
 sky130_fd_sc_hd__o21ai_1 _6887_ (.A1(_2843_),
    .A2(_1445_),
    .B1(_3163_),
    .Y(_0206_));
 sky130_fd_sc_hd__buf_6 _6888_ (.A(_1311_),
    .X(_3164_));
 sky130_fd_sc_hd__nand2_1 _6889_ (.A(\sound2.divisor_m[0] ),
    .B(\sound2.sdiv.Q[27] ),
    .Y(_3165_));
 sky130_fd_sc_hd__or2_1 _6890_ (.A(\sound2.divisor_m[0] ),
    .B(\sound2.sdiv.Q[27] ),
    .X(_3166_));
 sky130_fd_sc_hd__buf_6 _6891_ (.A(_0578_),
    .X(_3167_));
 sky130_fd_sc_hd__clkbuf_8 _6892_ (.A(_3167_),
    .X(_3168_));
 sky130_fd_sc_hd__a32o_1 _6893_ (.A1(_3164_),
    .A2(_3165_),
    .A3(_3166_),
    .B1(_3168_),
    .B2(\sound2.sdiv.A[0] ),
    .X(_0207_));
 sky130_fd_sc_hd__and2b_1 _6894_ (.A_N(\sound2.sdiv.A[26] ),
    .B(\sound2.divisor_m[0] ),
    .X(_3169_));
 sky130_fd_sc_hd__xnor2_1 _6895_ (.A(\sound2.divisor_m[1] ),
    .B(_3169_),
    .Y(_3170_));
 sky130_fd_sc_hd__xnor2_1 _6896_ (.A(\sound2.sdiv.A[0] ),
    .B(_3170_),
    .Y(_3171_));
 sky130_fd_sc_hd__or2b_1 _6897_ (.A(_3165_),
    .B_N(_3171_),
    .X(_3172_));
 sky130_fd_sc_hd__a21o_1 _6898_ (.A1(\sound2.divisor_m[0] ),
    .A2(\sound2.sdiv.Q[27] ),
    .B1(_3171_),
    .X(_3173_));
 sky130_fd_sc_hd__buf_6 _6899_ (.A(_0578_),
    .X(_3174_));
 sky130_fd_sc_hd__a32o_1 _6900_ (.A1(_3164_),
    .A2(_3172_),
    .A3(_3173_),
    .B1(_3174_),
    .B2(\sound2.sdiv.A[1] ),
    .X(_0208_));
 sky130_fd_sc_hd__or2b_1 _6901_ (.A(_3170_),
    .B_N(\sound2.sdiv.A[0] ),
    .X(_3175_));
 sky130_fd_sc_hd__inv_2 _6902_ (.A(\sound2.sdiv.A[1] ),
    .Y(_3176_));
 sky130_fd_sc_hd__clkinv_4 _6903_ (.A(\sound2.sdiv.A[26] ),
    .Y(_3177_));
 sky130_fd_sc_hd__o21a_1 _6904_ (.A1(\sound2.divisor_m[1] ),
    .A2(\sound2.divisor_m[0] ),
    .B1(_3177_),
    .X(_3178_));
 sky130_fd_sc_hd__xnor2_1 _6905_ (.A(\sound2.divisor_m[2] ),
    .B(_3178_),
    .Y(_3179_));
 sky130_fd_sc_hd__xnor2_1 _6906_ (.A(_3176_),
    .B(_3179_),
    .Y(_3180_));
 sky130_fd_sc_hd__a21o_1 _6907_ (.A1(_3175_),
    .A2(_3172_),
    .B1(_3180_),
    .X(_3181_));
 sky130_fd_sc_hd__nand3_1 _6908_ (.A(_3175_),
    .B(_3172_),
    .C(_3180_),
    .Y(_3182_));
 sky130_fd_sc_hd__a32o_1 _6909_ (.A1(_3164_),
    .A2(_3181_),
    .A3(_3182_),
    .B1(_3174_),
    .B2(\sound2.sdiv.A[2] ),
    .X(_0209_));
 sky130_fd_sc_hd__or2_1 _6910_ (.A(_3176_),
    .B(_3179_),
    .X(_3183_));
 sky130_fd_sc_hd__inv_2 _6911_ (.A(\sound2.sdiv.A[2] ),
    .Y(_3184_));
 sky130_fd_sc_hd__o31a_1 _6912_ (.A1(\sound2.divisor_m[2] ),
    .A2(\sound2.divisor_m[1] ),
    .A3(\sound2.divisor_m[0] ),
    .B1(_3177_),
    .X(_3185_));
 sky130_fd_sc_hd__xnor2_1 _6913_ (.A(\sound2.divisor_m[3] ),
    .B(_3185_),
    .Y(_3186_));
 sky130_fd_sc_hd__nor2_1 _6914_ (.A(_3184_),
    .B(_3186_),
    .Y(_3187_));
 sky130_fd_sc_hd__and2_1 _6915_ (.A(_3184_),
    .B(_3186_),
    .X(_3188_));
 sky130_fd_sc_hd__or2_1 _6916_ (.A(_3187_),
    .B(_3188_),
    .X(_3189_));
 sky130_fd_sc_hd__and3_1 _6917_ (.A(_3183_),
    .B(_3181_),
    .C(_3189_),
    .X(_3190_));
 sky130_fd_sc_hd__a21oi_1 _6918_ (.A1(_3183_),
    .A2(_3181_),
    .B1(_3189_),
    .Y(_3191_));
 sky130_fd_sc_hd__nor2_1 _6919_ (.A(_3190_),
    .B(_3191_),
    .Y(_3192_));
 sky130_fd_sc_hd__a22o_1 _6920_ (.A1(\sound2.sdiv.A[3] ),
    .A2(_3168_),
    .B1(\sound2.sdiv.next_dived ),
    .B2(_3192_),
    .X(_0210_));
 sky130_fd_sc_hd__inv_2 _6921_ (.A(\sound2.sdiv.A[3] ),
    .Y(_3193_));
 sky130_fd_sc_hd__or4_1 _6922_ (.A(\sound2.divisor_m[3] ),
    .B(\sound2.divisor_m[2] ),
    .C(\sound2.divisor_m[1] ),
    .D(\sound2.divisor_m[0] ),
    .X(_3194_));
 sky130_fd_sc_hd__nand2_1 _6923_ (.A(_3177_),
    .B(_3194_),
    .Y(_3195_));
 sky130_fd_sc_hd__xnor2_1 _6924_ (.A(_2484_),
    .B(_3195_),
    .Y(_3196_));
 sky130_fd_sc_hd__nor2_1 _6925_ (.A(_3193_),
    .B(_3196_),
    .Y(_3197_));
 sky130_fd_sc_hd__and2_1 _6926_ (.A(_3193_),
    .B(_3196_),
    .X(_3198_));
 sky130_fd_sc_hd__or2_1 _6927_ (.A(_3197_),
    .B(_3198_),
    .X(_3199_));
 sky130_fd_sc_hd__o21ba_1 _6928_ (.A1(_3187_),
    .A2(_3191_),
    .B1_N(_3199_),
    .X(_3200_));
 sky130_fd_sc_hd__or3b_1 _6929_ (.A(_3187_),
    .B(_3191_),
    .C_N(_3199_),
    .X(_3201_));
 sky130_fd_sc_hd__nand2_1 _6930_ (.A(_1311_),
    .B(_3201_),
    .Y(_3202_));
 sky130_fd_sc_hd__a2bb2o_1 _6931_ (.A1_N(_3200_),
    .A2_N(_3202_),
    .B1(\sound2.sdiv.A[4] ),
    .B2(_3168_),
    .X(_0211_));
 sky130_fd_sc_hd__inv_2 _6932_ (.A(\sound2.sdiv.A[4] ),
    .Y(_3203_));
 sky130_fd_sc_hd__o21a_1 _6933_ (.A1(\sound2.divisor_m[4] ),
    .A2(_3194_),
    .B1(_3177_),
    .X(_3204_));
 sky130_fd_sc_hd__xnor2_1 _6934_ (.A(\sound2.divisor_m[5] ),
    .B(_3204_),
    .Y(_3205_));
 sky130_fd_sc_hd__or2_1 _6935_ (.A(_3203_),
    .B(_3205_),
    .X(_3206_));
 sky130_fd_sc_hd__nand2_1 _6936_ (.A(_3203_),
    .B(_3205_),
    .Y(_3207_));
 sky130_fd_sc_hd__nand2_1 _6937_ (.A(_3206_),
    .B(_3207_),
    .Y(_3208_));
 sky130_fd_sc_hd__o21bai_1 _6938_ (.A1(_3197_),
    .A2(_3200_),
    .B1_N(_3208_),
    .Y(_3209_));
 sky130_fd_sc_hd__or3b_1 _6939_ (.A(_3197_),
    .B(_3200_),
    .C_N(_3208_),
    .X(_3210_));
 sky130_fd_sc_hd__a32o_1 _6940_ (.A1(_3164_),
    .A2(_3209_),
    .A3(_3210_),
    .B1(_3174_),
    .B2(\sound2.sdiv.A[5] ),
    .X(_0212_));
 sky130_fd_sc_hd__inv_2 _6941_ (.A(\sound2.sdiv.A[5] ),
    .Y(_3211_));
 sky130_fd_sc_hd__or3_1 _6942_ (.A(\sound2.divisor_m[5] ),
    .B(\sound2.divisor_m[4] ),
    .C(_3194_),
    .X(_3212_));
 sky130_fd_sc_hd__and2_1 _6943_ (.A(_3177_),
    .B(_3212_),
    .X(_3213_));
 sky130_fd_sc_hd__xnor2_1 _6944_ (.A(\sound2.divisor_m[6] ),
    .B(_3213_),
    .Y(_3214_));
 sky130_fd_sc_hd__or2_1 _6945_ (.A(_3211_),
    .B(_3214_),
    .X(_3215_));
 sky130_fd_sc_hd__nand2_1 _6946_ (.A(_3211_),
    .B(_3214_),
    .Y(_3216_));
 sky130_fd_sc_hd__nand2_1 _6947_ (.A(_3215_),
    .B(_3216_),
    .Y(_3217_));
 sky130_fd_sc_hd__nand3_1 _6948_ (.A(_3206_),
    .B(_3209_),
    .C(_3217_),
    .Y(_3218_));
 sky130_fd_sc_hd__a21o_1 _6949_ (.A1(_3206_),
    .A2(_3209_),
    .B1(_3217_),
    .X(_3219_));
 sky130_fd_sc_hd__a32o_1 _6950_ (.A1(_3164_),
    .A2(_3218_),
    .A3(_3219_),
    .B1(_3174_),
    .B2(\sound2.sdiv.A[6] ),
    .X(_0213_));
 sky130_fd_sc_hd__inv_2 _6951_ (.A(\sound2.sdiv.A[6] ),
    .Y(_3220_));
 sky130_fd_sc_hd__or2_1 _6952_ (.A(\sound2.divisor_m[6] ),
    .B(_3212_),
    .X(_3221_));
 sky130_fd_sc_hd__and2_1 _6953_ (.A(_3177_),
    .B(_3221_),
    .X(_3222_));
 sky130_fd_sc_hd__xnor2_1 _6954_ (.A(\sound2.divisor_m[7] ),
    .B(_3222_),
    .Y(_3223_));
 sky130_fd_sc_hd__or2_1 _6955_ (.A(_3220_),
    .B(_3223_),
    .X(_3224_));
 sky130_fd_sc_hd__nand2_1 _6956_ (.A(_3220_),
    .B(_3223_),
    .Y(_3225_));
 sky130_fd_sc_hd__nand2_1 _6957_ (.A(_3224_),
    .B(_3225_),
    .Y(_3226_));
 sky130_fd_sc_hd__nand3_1 _6958_ (.A(_3215_),
    .B(_3219_),
    .C(_3226_),
    .Y(_3227_));
 sky130_fd_sc_hd__a21o_1 _6959_ (.A1(_3215_),
    .A2(_3219_),
    .B1(_3226_),
    .X(_3228_));
 sky130_fd_sc_hd__a32o_1 _6960_ (.A1(_3164_),
    .A2(_3227_),
    .A3(_3228_),
    .B1(_3174_),
    .B2(\sound2.sdiv.A[7] ),
    .X(_0214_));
 sky130_fd_sc_hd__inv_2 _6961_ (.A(\sound2.sdiv.A[7] ),
    .Y(_3229_));
 sky130_fd_sc_hd__nor2_1 _6962_ (.A(\sound2.divisor_m[7] ),
    .B(_3221_),
    .Y(_3230_));
 sky130_fd_sc_hd__nor2_1 _6963_ (.A(\sound2.sdiv.A[26] ),
    .B(_3230_),
    .Y(_3231_));
 sky130_fd_sc_hd__xnor2_1 _6964_ (.A(\sound2.divisor_m[8] ),
    .B(_3231_),
    .Y(_3232_));
 sky130_fd_sc_hd__or2_2 _6965_ (.A(_3229_),
    .B(_3232_),
    .X(_3233_));
 sky130_fd_sc_hd__nand2_1 _6966_ (.A(_3229_),
    .B(_3232_),
    .Y(_3234_));
 sky130_fd_sc_hd__nand2_1 _6967_ (.A(_3233_),
    .B(_3234_),
    .Y(_3235_));
 sky130_fd_sc_hd__nand3_1 _6968_ (.A(_3224_),
    .B(_3228_),
    .C(_3235_),
    .Y(_3236_));
 sky130_fd_sc_hd__a21o_1 _6969_ (.A1(_3224_),
    .A2(_3228_),
    .B1(_3235_),
    .X(_3237_));
 sky130_fd_sc_hd__a32o_1 _6970_ (.A1(_3164_),
    .A2(_3236_),
    .A3(_3237_),
    .B1(_3174_),
    .B2(\sound2.sdiv.A[8] ),
    .X(_0215_));
 sky130_fd_sc_hd__a21o_1 _6971_ (.A1(_2460_),
    .A2(_3230_),
    .B1(\sound2.sdiv.A[26] ),
    .X(_3238_));
 sky130_fd_sc_hd__xnor2_1 _6972_ (.A(\sound2.divisor_m[9] ),
    .B(_3238_),
    .Y(_3239_));
 sky130_fd_sc_hd__and2_1 _6973_ (.A(\sound2.sdiv.A[8] ),
    .B(_3239_),
    .X(_3240_));
 sky130_fd_sc_hd__nor2_1 _6974_ (.A(\sound2.sdiv.A[8] ),
    .B(_3239_),
    .Y(_3241_));
 sky130_fd_sc_hd__o211ai_1 _6975_ (.A1(_3240_),
    .A2(_3241_),
    .B1(_3233_),
    .C1(_3237_),
    .Y(_3242_));
 sky130_fd_sc_hd__a211o_1 _6976_ (.A1(_3233_),
    .A2(_3237_),
    .B1(_3240_),
    .C1(_3241_),
    .X(_3243_));
 sky130_fd_sc_hd__a32o_1 _6977_ (.A1(_3164_),
    .A2(_3242_),
    .A3(_3243_),
    .B1(_3174_),
    .B2(\sound2.sdiv.A[9] ),
    .X(_0216_));
 sky130_fd_sc_hd__inv_2 _6978_ (.A(\sound2.sdiv.A[9] ),
    .Y(_3244_));
 sky130_fd_sc_hd__or4_1 _6979_ (.A(\sound2.divisor_m[9] ),
    .B(\sound2.divisor_m[8] ),
    .C(\sound2.divisor_m[7] ),
    .D(_3221_),
    .X(_3245_));
 sky130_fd_sc_hd__and2_1 _6980_ (.A(_3177_),
    .B(_3245_),
    .X(_3246_));
 sky130_fd_sc_hd__xnor2_1 _6981_ (.A(\sound2.divisor_m[10] ),
    .B(_3246_),
    .Y(_3247_));
 sky130_fd_sc_hd__or2_1 _6982_ (.A(_3244_),
    .B(_3247_),
    .X(_3248_));
 sky130_fd_sc_hd__nand2_1 _6983_ (.A(_3244_),
    .B(_3247_),
    .Y(_3249_));
 sky130_fd_sc_hd__nand2_1 _6984_ (.A(_3248_),
    .B(_3249_),
    .Y(_3250_));
 sky130_fd_sc_hd__inv_2 _6985_ (.A(_3240_),
    .Y(_3251_));
 sky130_fd_sc_hd__a31o_1 _6986_ (.A1(_3233_),
    .A2(_3237_),
    .A3(_3251_),
    .B1(_3241_),
    .X(_3252_));
 sky130_fd_sc_hd__nand2_1 _6987_ (.A(_3250_),
    .B(_3252_),
    .Y(_3253_));
 sky130_fd_sc_hd__a311o_1 _6988_ (.A1(_3233_),
    .A2(_3237_),
    .A3(_3251_),
    .B1(_3241_),
    .C1(_3250_),
    .X(_3254_));
 sky130_fd_sc_hd__a32o_1 _6989_ (.A1(_3164_),
    .A2(_3253_),
    .A3(_3254_),
    .B1(_3174_),
    .B2(\sound2.sdiv.A[10] ),
    .X(_0217_));
 sky130_fd_sc_hd__inv_2 _6990_ (.A(\sound2.sdiv.A[10] ),
    .Y(_3255_));
 sky130_fd_sc_hd__or2_1 _6991_ (.A(\sound2.divisor_m[10] ),
    .B(_3245_),
    .X(_3256_));
 sky130_fd_sc_hd__and2_1 _6992_ (.A(_3177_),
    .B(_3256_),
    .X(_3257_));
 sky130_fd_sc_hd__xnor2_1 _6993_ (.A(\sound2.divisor_m[11] ),
    .B(_3257_),
    .Y(_3258_));
 sky130_fd_sc_hd__nor2_1 _6994_ (.A(_3255_),
    .B(_3258_),
    .Y(_3259_));
 sky130_fd_sc_hd__and2_1 _6995_ (.A(_3255_),
    .B(_3258_),
    .X(_3260_));
 sky130_fd_sc_hd__or2_1 _6996_ (.A(_3259_),
    .B(_3260_),
    .X(_3261_));
 sky130_fd_sc_hd__a21oi_1 _6997_ (.A1(_3248_),
    .A2(_3254_),
    .B1(_3261_),
    .Y(_3262_));
 sky130_fd_sc_hd__and3_1 _6998_ (.A(_3248_),
    .B(_3254_),
    .C(_3261_),
    .X(_3263_));
 sky130_fd_sc_hd__nor2_1 _6999_ (.A(_3262_),
    .B(_3263_),
    .Y(_3264_));
 sky130_fd_sc_hd__a22o_1 _7000_ (.A1(\sound2.sdiv.A[11] ),
    .A2(_3168_),
    .B1(\sound2.sdiv.next_dived ),
    .B2(_3264_),
    .X(_0218_));
 sky130_fd_sc_hd__inv_2 _7001_ (.A(\sound2.sdiv.A[11] ),
    .Y(_3265_));
 sky130_fd_sc_hd__o21a_1 _7002_ (.A1(\sound2.divisor_m[11] ),
    .A2(_3256_),
    .B1(_3177_),
    .X(_3266_));
 sky130_fd_sc_hd__xnor2_1 _7003_ (.A(\sound2.divisor_m[12] ),
    .B(_3266_),
    .Y(_3267_));
 sky130_fd_sc_hd__or2_1 _7004_ (.A(_3265_),
    .B(_3267_),
    .X(_3268_));
 sky130_fd_sc_hd__nand2_1 _7005_ (.A(_3265_),
    .B(_3267_),
    .Y(_3269_));
 sky130_fd_sc_hd__nand2_1 _7006_ (.A(_3268_),
    .B(_3269_),
    .Y(_3270_));
 sky130_fd_sc_hd__or3b_1 _7007_ (.A(_3259_),
    .B(_3262_),
    .C_N(_3270_),
    .X(_3271_));
 sky130_fd_sc_hd__o21bai_1 _7008_ (.A1(_3259_),
    .A2(_3262_),
    .B1_N(_3270_),
    .Y(_3272_));
 sky130_fd_sc_hd__a32o_1 _7009_ (.A1(_3164_),
    .A2(_3271_),
    .A3(_3272_),
    .B1(_3174_),
    .B2(\sound2.sdiv.A[12] ),
    .X(_0219_));
 sky130_fd_sc_hd__inv_2 _7010_ (.A(\sound2.sdiv.A[12] ),
    .Y(_3273_));
 sky130_fd_sc_hd__or3_1 _7011_ (.A(\sound2.divisor_m[12] ),
    .B(\sound2.divisor_m[11] ),
    .C(_3256_),
    .X(_3274_));
 sky130_fd_sc_hd__and2_1 _7012_ (.A(_3177_),
    .B(_3274_),
    .X(_3275_));
 sky130_fd_sc_hd__xnor2_1 _7013_ (.A(\sound2.divisor_m[13] ),
    .B(_3275_),
    .Y(_3276_));
 sky130_fd_sc_hd__or2_1 _7014_ (.A(_3273_),
    .B(_3276_),
    .X(_3277_));
 sky130_fd_sc_hd__nand2_1 _7015_ (.A(_3273_),
    .B(_3276_),
    .Y(_3278_));
 sky130_fd_sc_hd__nand2_1 _7016_ (.A(_3277_),
    .B(_3278_),
    .Y(_3279_));
 sky130_fd_sc_hd__a21o_1 _7017_ (.A1(_3268_),
    .A2(_3272_),
    .B1(_3279_),
    .X(_3280_));
 sky130_fd_sc_hd__nand3_1 _7018_ (.A(_3268_),
    .B(_3272_),
    .C(_3279_),
    .Y(_3281_));
 sky130_fd_sc_hd__a32o_1 _7019_ (.A1(_3164_),
    .A2(_3280_),
    .A3(_3281_),
    .B1(_3174_),
    .B2(\sound2.sdiv.A[13] ),
    .X(_0220_));
 sky130_fd_sc_hd__inv_2 _7020_ (.A(\sound2.sdiv.A[13] ),
    .Y(_3282_));
 sky130_fd_sc_hd__or2_1 _7021_ (.A(\sound2.divisor_m[13] ),
    .B(_3274_),
    .X(_3283_));
 sky130_fd_sc_hd__nand2_1 _7022_ (.A(_3177_),
    .B(_3283_),
    .Y(_3284_));
 sky130_fd_sc_hd__xnor2_1 _7023_ (.A(_2441_),
    .B(_3284_),
    .Y(_3285_));
 sky130_fd_sc_hd__or2_1 _7024_ (.A(_3282_),
    .B(_3285_),
    .X(_3286_));
 sky130_fd_sc_hd__nand2_1 _7025_ (.A(_3282_),
    .B(_3285_),
    .Y(_3287_));
 sky130_fd_sc_hd__nand2_1 _7026_ (.A(_3286_),
    .B(_3287_),
    .Y(_3288_));
 sky130_fd_sc_hd__nand3_1 _7027_ (.A(_3277_),
    .B(_3280_),
    .C(_3288_),
    .Y(_3289_));
 sky130_fd_sc_hd__a21o_1 _7028_ (.A1(_3277_),
    .A2(_3280_),
    .B1(_3288_),
    .X(_3290_));
 sky130_fd_sc_hd__a32o_1 _7029_ (.A1(_3164_),
    .A2(_3289_),
    .A3(_3290_),
    .B1(_3174_),
    .B2(\sound2.sdiv.A[14] ),
    .X(_0221_));
 sky130_fd_sc_hd__inv_2 _7030_ (.A(\sound2.sdiv.A[14] ),
    .Y(_3291_));
 sky130_fd_sc_hd__o21a_1 _7031_ (.A1(\sound2.divisor_m[14] ),
    .A2(_3283_),
    .B1(_3177_),
    .X(_3292_));
 sky130_fd_sc_hd__xnor2_1 _7032_ (.A(\sound2.divisor_m[15] ),
    .B(_3292_),
    .Y(_3293_));
 sky130_fd_sc_hd__or2_1 _7033_ (.A(_3291_),
    .B(_3293_),
    .X(_3294_));
 sky130_fd_sc_hd__nand2_1 _7034_ (.A(_3291_),
    .B(_3293_),
    .Y(_3295_));
 sky130_fd_sc_hd__nand2_1 _7035_ (.A(_3294_),
    .B(_3295_),
    .Y(_3296_));
 sky130_fd_sc_hd__nand3_1 _7036_ (.A(_3286_),
    .B(_3290_),
    .C(_3296_),
    .Y(_3297_));
 sky130_fd_sc_hd__a21o_1 _7037_ (.A1(_3286_),
    .A2(_3290_),
    .B1(_3296_),
    .X(_3298_));
 sky130_fd_sc_hd__a32o_1 _7038_ (.A1(_3164_),
    .A2(_3297_),
    .A3(_3298_),
    .B1(_3174_),
    .B2(\sound2.sdiv.A[15] ),
    .X(_0222_));
 sky130_fd_sc_hd__inv_2 _7039_ (.A(\sound2.sdiv.A[15] ),
    .Y(_3299_));
 sky130_fd_sc_hd__o31a_1 _7040_ (.A1(\sound2.divisor_m[15] ),
    .A2(\sound2.divisor_m[14] ),
    .A3(_3283_),
    .B1(_3177_),
    .X(_3300_));
 sky130_fd_sc_hd__xnor2_1 _7041_ (.A(\sound2.divisor_m[16] ),
    .B(_3300_),
    .Y(_3301_));
 sky130_fd_sc_hd__nor2_1 _7042_ (.A(_3299_),
    .B(_3301_),
    .Y(_3302_));
 sky130_fd_sc_hd__and2_1 _7043_ (.A(_3299_),
    .B(_3301_),
    .X(_3303_));
 sky130_fd_sc_hd__or2_1 _7044_ (.A(_3302_),
    .B(_3303_),
    .X(_3304_));
 sky130_fd_sc_hd__and3_1 _7045_ (.A(_3294_),
    .B(_3298_),
    .C(_3304_),
    .X(_3305_));
 sky130_fd_sc_hd__a21oi_2 _7046_ (.A1(_3294_),
    .A2(_3298_),
    .B1(_3304_),
    .Y(_3306_));
 sky130_fd_sc_hd__nor2_1 _7047_ (.A(_3305_),
    .B(_3306_),
    .Y(_3307_));
 sky130_fd_sc_hd__a22o_1 _7048_ (.A1(\sound2.sdiv.A[16] ),
    .A2(_3168_),
    .B1(\sound2.sdiv.next_dived ),
    .B2(_3307_),
    .X(_0223_));
 sky130_fd_sc_hd__or4_1 _7049_ (.A(\sound2.divisor_m[16] ),
    .B(\sound2.divisor_m[15] ),
    .C(\sound2.divisor_m[14] ),
    .D(_3283_),
    .X(_3308_));
 sky130_fd_sc_hd__and2_1 _7050_ (.A(_3177_),
    .B(_3308_),
    .X(_3309_));
 sky130_fd_sc_hd__xnor2_1 _7051_ (.A(\sound2.divisor_m[17] ),
    .B(_3309_),
    .Y(_3310_));
 sky130_fd_sc_hd__inv_2 _7052_ (.A(_3310_),
    .Y(_3311_));
 sky130_fd_sc_hd__nand2_1 _7053_ (.A(\sound2.sdiv.A[16] ),
    .B(_3311_),
    .Y(_3312_));
 sky130_fd_sc_hd__inv_2 _7054_ (.A(_3312_),
    .Y(_3313_));
 sky130_fd_sc_hd__nor2_1 _7055_ (.A(\sound2.sdiv.A[16] ),
    .B(_3311_),
    .Y(_3314_));
 sky130_fd_sc_hd__nor2_1 _7056_ (.A(_3313_),
    .B(_3314_),
    .Y(_3315_));
 sky130_fd_sc_hd__o21ai_1 _7057_ (.A1(_3302_),
    .A2(_3306_),
    .B1(_3315_),
    .Y(_3316_));
 sky130_fd_sc_hd__or3_1 _7058_ (.A(_3302_),
    .B(_3306_),
    .C(_3315_),
    .X(_3317_));
 sky130_fd_sc_hd__a32o_1 _7059_ (.A1(_3164_),
    .A2(_3316_),
    .A3(_3317_),
    .B1(_3174_),
    .B2(\sound2.sdiv.A[17] ),
    .X(_0224_));
 sky130_fd_sc_hd__o21a_1 _7060_ (.A1(\sound2.divisor_m[17] ),
    .A2(_3308_),
    .B1(_3177_),
    .X(_3318_));
 sky130_fd_sc_hd__xnor2_1 _7061_ (.A(\sound2.divisor_m[18] ),
    .B(_3318_),
    .Y(_3319_));
 sky130_fd_sc_hd__inv_2 _7062_ (.A(_3319_),
    .Y(_3320_));
 sky130_fd_sc_hd__nand2_1 _7063_ (.A(\sound2.sdiv.A[17] ),
    .B(_3320_),
    .Y(_3321_));
 sky130_fd_sc_hd__or2_1 _7064_ (.A(\sound2.sdiv.A[17] ),
    .B(_3320_),
    .X(_3322_));
 sky130_fd_sc_hd__nand2_1 _7065_ (.A(_3321_),
    .B(_3322_),
    .Y(_3323_));
 sky130_fd_sc_hd__o21ba_1 _7066_ (.A1(_3302_),
    .A2(_3313_),
    .B1_N(_3314_),
    .X(_3324_));
 sky130_fd_sc_hd__a21o_1 _7067_ (.A1(_3306_),
    .A2(_3315_),
    .B1(_3324_),
    .X(_3325_));
 sky130_fd_sc_hd__xnor2_1 _7068_ (.A(_3323_),
    .B(_3325_),
    .Y(_3326_));
 sky130_fd_sc_hd__a22o_1 _7069_ (.A1(\sound2.sdiv.A[18] ),
    .A2(_3168_),
    .B1(\sound2.sdiv.next_dived ),
    .B2(_3326_),
    .X(_0225_));
 sky130_fd_sc_hd__and3b_1 _7070_ (.A_N(_3308_),
    .B(_2471_),
    .C(_2470_),
    .X(_3327_));
 sky130_fd_sc_hd__nor2_1 _7071_ (.A(\sound2.sdiv.A[26] ),
    .B(_3327_),
    .Y(_3328_));
 sky130_fd_sc_hd__buf_4 _7072_ (.A(_3328_),
    .X(_3329_));
 sky130_fd_sc_hd__nor2_1 _7073_ (.A(\sound2.sdiv.A[18] ),
    .B(_3329_),
    .Y(_3330_));
 sky130_fd_sc_hd__nand2_1 _7074_ (.A(\sound2.sdiv.A[18] ),
    .B(_3329_),
    .Y(_3331_));
 sky130_fd_sc_hd__or2b_1 _7075_ (.A(_3330_),
    .B_N(_3331_),
    .X(_3332_));
 sky130_fd_sc_hd__a21bo_1 _7076_ (.A1(_3322_),
    .A2(_3325_),
    .B1_N(_3321_),
    .X(_3333_));
 sky130_fd_sc_hd__xnor2_1 _7077_ (.A(_3332_),
    .B(_3333_),
    .Y(_3334_));
 sky130_fd_sc_hd__a22o_1 _7078_ (.A1(\sound2.sdiv.A[19] ),
    .A2(_3168_),
    .B1(\sound2.sdiv.next_dived ),
    .B2(_3334_),
    .X(_0226_));
 sky130_fd_sc_hd__or2_1 _7079_ (.A(\sound2.sdiv.A[19] ),
    .B(_3329_),
    .X(_3335_));
 sky130_fd_sc_hd__nand2_1 _7080_ (.A(\sound2.sdiv.A[19] ),
    .B(_3329_),
    .Y(_3336_));
 sky130_fd_sc_hd__nand2_1 _7081_ (.A(_3335_),
    .B(_3336_),
    .Y(_3337_));
 sky130_fd_sc_hd__or3_1 _7082_ (.A(_3304_),
    .B(_3313_),
    .C(_3314_),
    .X(_3338_));
 sky130_fd_sc_hd__a2111o_1 _7083_ (.A1(_3294_),
    .A2(_3298_),
    .B1(_3323_),
    .C1(_3338_),
    .D1(_3332_),
    .X(_3339_));
 sky130_fd_sc_hd__or4bb_1 _7084_ (.A(_3323_),
    .B(_3330_),
    .C_N(_3331_),
    .D_N(_3324_),
    .X(_3340_));
 sky130_fd_sc_hd__o211a_1 _7085_ (.A1(_3321_),
    .A2(_3330_),
    .B1(_3331_),
    .C1(_3340_),
    .X(_3341_));
 sky130_fd_sc_hd__and3_1 _7086_ (.A(_3337_),
    .B(_3339_),
    .C(_3341_),
    .X(_3342_));
 sky130_fd_sc_hd__a21o_1 _7087_ (.A1(_3339_),
    .A2(_3341_),
    .B1(_3337_),
    .X(_3343_));
 sky130_fd_sc_hd__nand2_1 _7088_ (.A(_1311_),
    .B(_3343_),
    .Y(_3344_));
 sky130_fd_sc_hd__a2bb2o_1 _7089_ (.A1_N(_3342_),
    .A2_N(_3344_),
    .B1(\sound2.sdiv.A[20] ),
    .B2(_3168_),
    .X(_0227_));
 sky130_fd_sc_hd__xor2_1 _7090_ (.A(\sound2.sdiv.A[20] ),
    .B(_3329_),
    .X(_3345_));
 sky130_fd_sc_hd__inv_2 _7091_ (.A(_3345_),
    .Y(_3346_));
 sky130_fd_sc_hd__a21o_1 _7092_ (.A1(_3336_),
    .A2(_3343_),
    .B1(_3346_),
    .X(_3347_));
 sky130_fd_sc_hd__nand3_1 _7093_ (.A(_3336_),
    .B(_3343_),
    .C(_3346_),
    .Y(_3348_));
 sky130_fd_sc_hd__a32o_1 _7094_ (.A1(_3164_),
    .A2(_3347_),
    .A3(_3348_),
    .B1(_3174_),
    .B2(\sound2.sdiv.A[21] ),
    .X(_0228_));
 sky130_fd_sc_hd__buf_6 _7095_ (.A(_1311_),
    .X(_3349_));
 sky130_fd_sc_hd__xnor2_1 _7096_ (.A(\sound2.sdiv.A[21] ),
    .B(_3329_),
    .Y(_3350_));
 sky130_fd_sc_hd__o21bai_1 _7097_ (.A1(\sound2.sdiv.A[20] ),
    .A2(_3329_),
    .B1_N(_3343_),
    .Y(_3351_));
 sky130_fd_sc_hd__o21ai_1 _7098_ (.A1(\sound2.sdiv.A[20] ),
    .A2(\sound2.sdiv.A[19] ),
    .B1(_3329_),
    .Y(_3352_));
 sky130_fd_sc_hd__nand3_1 _7099_ (.A(_3350_),
    .B(_3351_),
    .C(_3352_),
    .Y(_3353_));
 sky130_fd_sc_hd__a21o_1 _7100_ (.A1(_3351_),
    .A2(_3352_),
    .B1(_3350_),
    .X(_3354_));
 sky130_fd_sc_hd__a32o_1 _7101_ (.A1(_3349_),
    .A2(_3353_),
    .A3(_3354_),
    .B1(_3174_),
    .B2(\sound2.sdiv.A[22] ),
    .X(_0229_));
 sky130_fd_sc_hd__xor2_1 _7102_ (.A(\sound2.sdiv.A[22] ),
    .B(_3329_),
    .X(_3355_));
 sky130_fd_sc_hd__a21boi_1 _7103_ (.A1(\sound2.sdiv.A[21] ),
    .A2(_3329_),
    .B1_N(_3354_),
    .Y(_3356_));
 sky130_fd_sc_hd__xnor2_1 _7104_ (.A(_3355_),
    .B(_3356_),
    .Y(_3357_));
 sky130_fd_sc_hd__a22o_1 _7105_ (.A1(\sound2.sdiv.A[23] ),
    .A2(_3168_),
    .B1(\sound2.sdiv.next_dived ),
    .B2(_3357_),
    .X(_0230_));
 sky130_fd_sc_hd__or2_1 _7106_ (.A(\sound2.sdiv.A[23] ),
    .B(_3329_),
    .X(_3358_));
 sky130_fd_sc_hd__nand2_1 _7107_ (.A(\sound2.sdiv.A[23] ),
    .B(_3329_),
    .Y(_3359_));
 sky130_fd_sc_hd__nand2_1 _7108_ (.A(_3358_),
    .B(_3359_),
    .Y(_3360_));
 sky130_fd_sc_hd__or3b_1 _7109_ (.A(_3346_),
    .B(_3350_),
    .C_N(_3355_),
    .X(_3361_));
 sky130_fd_sc_hd__o21ai_1 _7110_ (.A1(\sound2.sdiv.A[22] ),
    .A2(\sound2.sdiv.A[21] ),
    .B1(_3329_),
    .Y(_3362_));
 sky130_fd_sc_hd__o211a_1 _7111_ (.A1(_3343_),
    .A2(_3361_),
    .B1(_3362_),
    .C1(_3352_),
    .X(_3363_));
 sky130_fd_sc_hd__xor2_1 _7112_ (.A(_3360_),
    .B(_3363_),
    .X(_3364_));
 sky130_fd_sc_hd__a22o_1 _7113_ (.A1(\sound2.sdiv.A[24] ),
    .A2(_3168_),
    .B1(\sound2.sdiv.next_dived ),
    .B2(_3364_),
    .X(_0231_));
 sky130_fd_sc_hd__o21a_1 _7114_ (.A1(_3360_),
    .A2(_3363_),
    .B1(_3359_),
    .X(_3365_));
 sky130_fd_sc_hd__nor2_1 _7115_ (.A(\sound2.sdiv.A[24] ),
    .B(_3329_),
    .Y(_3366_));
 sky130_fd_sc_hd__nand2_1 _7116_ (.A(\sound2.sdiv.A[24] ),
    .B(_3329_),
    .Y(_3367_));
 sky130_fd_sc_hd__and2b_1 _7117_ (.A_N(_3366_),
    .B(_3367_),
    .X(_3368_));
 sky130_fd_sc_hd__xnor2_1 _7118_ (.A(_3365_),
    .B(_3368_),
    .Y(_3369_));
 sky130_fd_sc_hd__a22o_1 _7119_ (.A1(\sound2.sdiv.A[25] ),
    .A2(_3168_),
    .B1(\sound2.sdiv.next_dived ),
    .B2(_3369_),
    .X(_0232_));
 sky130_fd_sc_hd__xnor2_1 _7120_ (.A(\sound2.sdiv.A[25] ),
    .B(_3329_),
    .Y(_3370_));
 sky130_fd_sc_hd__o211ai_1 _7121_ (.A1(_3365_),
    .A2(_3366_),
    .B1(_3367_),
    .C1(_3370_),
    .Y(_3371_));
 sky130_fd_sc_hd__or3_1 _7122_ (.A(_3360_),
    .B(_3363_),
    .C(_3366_),
    .X(_3372_));
 sky130_fd_sc_hd__a31o_1 _7123_ (.A1(_3359_),
    .A2(_3367_),
    .A3(_3372_),
    .B1(_3370_),
    .X(_3373_));
 sky130_fd_sc_hd__a32o_1 _7124_ (.A1(_3349_),
    .A2(_3371_),
    .A3(_3373_),
    .B1(_3174_),
    .B2(\sound2.sdiv.A[26] ),
    .X(_0233_));
 sky130_fd_sc_hd__mux2_1 _7125_ (.A0(_1311_),
    .A1(_3167_),
    .S(\sound2.sdiv.C[0] ),
    .X(_3374_));
 sky130_fd_sc_hd__clkbuf_1 _7126_ (.A(_3374_),
    .X(_0234_));
 sky130_fd_sc_hd__nand2_1 _7127_ (.A(\sound2.sdiv.C[1] ),
    .B(\sound2.sdiv.C[0] ),
    .Y(_3375_));
 sky130_fd_sc_hd__or2_1 _7128_ (.A(\sound2.sdiv.C[1] ),
    .B(\sound2.sdiv.C[0] ),
    .X(_3376_));
 sky130_fd_sc_hd__a32o_1 _7129_ (.A1(_3349_),
    .A2(_3375_),
    .A3(_3376_),
    .B1(_3174_),
    .B2(\sound2.sdiv.C[1] ),
    .X(_0235_));
 sky130_fd_sc_hd__a21o_1 _7130_ (.A1(\sound2.sdiv.C[1] ),
    .A2(\sound2.sdiv.C[0] ),
    .B1(\sound2.sdiv.C[2] ),
    .X(_3377_));
 sky130_fd_sc_hd__and3_1 _7131_ (.A(\sound2.sdiv.C[2] ),
    .B(\sound2.sdiv.C[1] ),
    .C(\sound2.sdiv.C[0] ),
    .X(_3378_));
 sky130_fd_sc_hd__inv_2 _7132_ (.A(_3378_),
    .Y(_3379_));
 sky130_fd_sc_hd__a32o_1 _7133_ (.A1(_3349_),
    .A2(_3377_),
    .A3(_3379_),
    .B1(_3174_),
    .B2(\sound2.sdiv.C[2] ),
    .X(_0236_));
 sky130_fd_sc_hd__and3_1 _7134_ (.A(\sound2.sdiv.C[3] ),
    .B(net66),
    .C(_3378_),
    .X(_3380_));
 sky130_fd_sc_hd__a21oi_1 _7135_ (.A1(_0559_),
    .A2(_3378_),
    .B1(\sound2.sdiv.C[3] ),
    .Y(_3381_));
 sky130_fd_sc_hd__nor3_1 _7136_ (.A(_2005_),
    .B(_3380_),
    .C(_3381_),
    .Y(_0237_));
 sky130_fd_sc_hd__a31o_1 _7137_ (.A1(\sound2.sdiv.C[3] ),
    .A2(_0559_),
    .A3(_3378_),
    .B1(\sound2.sdiv.C[4] ),
    .X(_3382_));
 sky130_fd_sc_hd__and2_1 _7138_ (.A(_2843_),
    .B(_3382_),
    .X(_3383_));
 sky130_fd_sc_hd__clkbuf_1 _7139_ (.A(_3383_),
    .X(_0238_));
 sky130_fd_sc_hd__and2_1 _7140_ (.A(\sound2.sdiv.C[5] ),
    .B(_0554_),
    .X(_3384_));
 sky130_fd_sc_hd__clkbuf_1 _7141_ (.A(_3384_),
    .X(_0239_));
 sky130_fd_sc_hd__o21ai_1 _7142_ (.A1(\sound2.sdiv.A[25] ),
    .A2(_3327_),
    .B1(_3177_),
    .Y(_3385_));
 sky130_fd_sc_hd__nand2_1 _7143_ (.A(_3373_),
    .B(_3385_),
    .Y(_3386_));
 sky130_fd_sc_hd__a21bo_1 _7144_ (.A1(\sound2.sdiv.next_dived ),
    .A2(_3386_),
    .B1_N(_2276_),
    .X(_0240_));
 sky130_fd_sc_hd__a21o_1 _7145_ (.A1(\sound2.sdiv.Q[0] ),
    .A2(\sound2.sdiv.next_dived ),
    .B1(_2501_),
    .X(_0241_));
 sky130_fd_sc_hd__a22o_1 _7146_ (.A1(\sound2.sdiv.Q[2] ),
    .A2(_3168_),
    .B1(\sound2.sdiv.next_dived ),
    .B2(\sound2.sdiv.Q[1] ),
    .X(_0242_));
 sky130_fd_sc_hd__a22o_1 _7147_ (.A1(\sound2.sdiv.Q[3] ),
    .A2(_3168_),
    .B1(\sound2.sdiv.next_dived ),
    .B2(\sound2.sdiv.Q[2] ),
    .X(_0243_));
 sky130_fd_sc_hd__a22o_1 _7148_ (.A1(\sound2.sdiv.Q[4] ),
    .A2(_3168_),
    .B1(_3164_),
    .B2(\sound2.sdiv.Q[3] ),
    .X(_0244_));
 sky130_fd_sc_hd__a22o_1 _7149_ (.A1(\sound2.sdiv.Q[5] ),
    .A2(_3168_),
    .B1(_3164_),
    .B2(\sound2.sdiv.Q[4] ),
    .X(_0245_));
 sky130_fd_sc_hd__a22o_1 _7150_ (.A1(\sound2.sdiv.Q[6] ),
    .A2(_3168_),
    .B1(_3164_),
    .B2(\sound2.sdiv.Q[5] ),
    .X(_0246_));
 sky130_fd_sc_hd__a22o_1 _7151_ (.A1(\sound2.sdiv.Q[7] ),
    .A2(_3168_),
    .B1(_3164_),
    .B2(\sound2.sdiv.Q[6] ),
    .X(_0247_));
 sky130_fd_sc_hd__a221o_1 _7152_ (.A1(\sound2.sdiv.Q[8] ),
    .A2(_3174_),
    .B1(_3349_),
    .B2(\sound2.sdiv.Q[7] ),
    .C1(_3115_),
    .X(_0248_));
 sky130_fd_sc_hd__a221o_1 _7153_ (.A1(\sound2.sdiv.Q[9] ),
    .A2(_3174_),
    .B1(_3349_),
    .B2(\sound2.sdiv.Q[8] ),
    .C1(_3116_),
    .X(_0249_));
 sky130_fd_sc_hd__a221o_1 _7154_ (.A1(\sound2.sdiv.Q[10] ),
    .A2(_3167_),
    .B1(_3349_),
    .B2(\sound2.sdiv.Q[9] ),
    .C1(_3117_),
    .X(_0250_));
 sky130_fd_sc_hd__a221o_1 _7155_ (.A1(\sound2.sdiv.Q[11] ),
    .A2(_3167_),
    .B1(_3349_),
    .B2(\sound2.sdiv.Q[10] ),
    .C1(_3118_),
    .X(_0251_));
 sky130_fd_sc_hd__a221o_1 _7156_ (.A1(\sound2.sdiv.Q[12] ),
    .A2(_3167_),
    .B1(_3349_),
    .B2(\sound2.sdiv.Q[11] ),
    .C1(_3119_),
    .X(_0252_));
 sky130_fd_sc_hd__a221o_1 _7157_ (.A1(\sound2.sdiv.Q[13] ),
    .A2(_3167_),
    .B1(_3349_),
    .B2(\sound2.sdiv.Q[12] ),
    .C1(_3120_),
    .X(_0253_));
 sky130_fd_sc_hd__a221o_1 _7158_ (.A1(\sound2.sdiv.Q[14] ),
    .A2(_3167_),
    .B1(_3349_),
    .B2(\sound2.sdiv.Q[13] ),
    .C1(_3121_),
    .X(_0254_));
 sky130_fd_sc_hd__a221o_1 _7159_ (.A1(\sound2.sdiv.Q[15] ),
    .A2(_3167_),
    .B1(_3349_),
    .B2(\sound2.sdiv.Q[14] ),
    .C1(_3122_),
    .X(_0255_));
 sky130_fd_sc_hd__a221o_1 _7160_ (.A1(\sound2.sdiv.Q[16] ),
    .A2(_3167_),
    .B1(_3349_),
    .B2(\sound2.sdiv.Q[15] ),
    .C1(_3123_),
    .X(_0256_));
 sky130_fd_sc_hd__a221o_1 _7161_ (.A1(\sound2.sdiv.Q[17] ),
    .A2(_3167_),
    .B1(_3349_),
    .B2(\sound2.sdiv.Q[16] ),
    .C1(_3124_),
    .X(_0257_));
 sky130_fd_sc_hd__a221o_1 _7162_ (.A1(\sound2.sdiv.Q[18] ),
    .A2(_3167_),
    .B1(_3349_),
    .B2(\sound2.sdiv.Q[17] ),
    .C1(_3125_),
    .X(_0258_));
 sky130_fd_sc_hd__a221o_1 _7163_ (.A1(\sound2.sdiv.Q[19] ),
    .A2(_3167_),
    .B1(_3349_),
    .B2(\sound2.sdiv.Q[18] ),
    .C1(_3126_),
    .X(_0259_));
 sky130_fd_sc_hd__a221o_1 _7164_ (.A1(\sound2.sdiv.Q[20] ),
    .A2(_3167_),
    .B1(_3349_),
    .B2(\sound2.sdiv.Q[19] ),
    .C1(_3127_),
    .X(_0260_));
 sky130_fd_sc_hd__a221o_1 _7165_ (.A1(\sound2.sdiv.Q[21] ),
    .A2(_3167_),
    .B1(_3349_),
    .B2(\sound2.sdiv.Q[20] ),
    .C1(_3128_),
    .X(_0261_));
 sky130_fd_sc_hd__a221o_1 _7166_ (.A1(\sound2.sdiv.Q[22] ),
    .A2(_3167_),
    .B1(_3349_),
    .B2(\sound2.sdiv.Q[21] ),
    .C1(_3129_),
    .X(_0262_));
 sky130_fd_sc_hd__a221o_1 _7167_ (.A1(\sound2.sdiv.Q[23] ),
    .A2(_3167_),
    .B1(_3349_),
    .B2(\sound2.sdiv.Q[22] ),
    .C1(_3130_),
    .X(_0263_));
 sky130_fd_sc_hd__a221o_1 _7168_ (.A1(\sound2.sdiv.Q[24] ),
    .A2(_3167_),
    .B1(_1311_),
    .B2(\sound2.sdiv.Q[23] ),
    .C1(_3131_),
    .X(_0264_));
 sky130_fd_sc_hd__a221o_1 _7169_ (.A1(\sound2.sdiv.Q[25] ),
    .A2(_3167_),
    .B1(_1311_),
    .B2(\sound2.sdiv.Q[24] ),
    .C1(_3133_),
    .X(_0265_));
 sky130_fd_sc_hd__a221o_1 _7170_ (.A1(\sound2.sdiv.Q[26] ),
    .A2(_3167_),
    .B1(_1311_),
    .B2(\sound2.sdiv.Q[25] ),
    .C1(_3134_),
    .X(_0266_));
 sky130_fd_sc_hd__a22o_1 _7171_ (.A1(\sound2.sdiv.Q[27] ),
    .A2(_3168_),
    .B1(_3164_),
    .B2(\sound2.sdiv.Q[26] ),
    .X(_0267_));
 sky130_fd_sc_hd__and2_1 _7172_ (.A(\sound3.count[0] ),
    .B(_2855_),
    .X(_3387_));
 sky130_fd_sc_hd__a21o_1 _7173_ (.A1(\sound3.count_m[0] ),
    .A2(_3132_),
    .B1(_3387_),
    .X(_0268_));
 sky130_fd_sc_hd__and2_1 _7174_ (.A(\sound3.count[1] ),
    .B(_2863_),
    .X(_3388_));
 sky130_fd_sc_hd__a21o_1 _7175_ (.A1(\sound3.count_m[1] ),
    .A2(_3132_),
    .B1(_3388_),
    .X(_0269_));
 sky130_fd_sc_hd__and2_1 _7176_ (.A(\sound3.count[2] ),
    .B(_2863_),
    .X(_3389_));
 sky130_fd_sc_hd__a21o_1 _7177_ (.A1(\sound3.count_m[2] ),
    .A2(_3132_),
    .B1(_3389_),
    .X(_0270_));
 sky130_fd_sc_hd__and2_1 _7178_ (.A(\sound3.count[3] ),
    .B(_2863_),
    .X(_3390_));
 sky130_fd_sc_hd__a21o_1 _7179_ (.A1(\sound3.count_m[3] ),
    .A2(_3132_),
    .B1(_3390_),
    .X(_0271_));
 sky130_fd_sc_hd__and2_1 _7180_ (.A(\sound3.count[4] ),
    .B(_2863_),
    .X(_3391_));
 sky130_fd_sc_hd__a21o_1 _7181_ (.A1(\sound3.count_m[4] ),
    .A2(_3132_),
    .B1(_3391_),
    .X(_0272_));
 sky130_fd_sc_hd__and2_1 _7182_ (.A(\sound3.count[5] ),
    .B(_2863_),
    .X(_3392_));
 sky130_fd_sc_hd__a21o_1 _7183_ (.A1(\sound3.count_m[5] ),
    .A2(_3132_),
    .B1(_3392_),
    .X(_0273_));
 sky130_fd_sc_hd__and2_1 _7184_ (.A(\sound3.count[6] ),
    .B(_2863_),
    .X(_3393_));
 sky130_fd_sc_hd__a21o_1 _7185_ (.A1(\sound3.count_m[6] ),
    .A2(_3132_),
    .B1(_3393_),
    .X(_0274_));
 sky130_fd_sc_hd__nor2_1 _7186_ (.A(_1642_),
    .B(_2843_),
    .Y(_3394_));
 sky130_fd_sc_hd__a21o_1 _7187_ (.A1(\sound3.count_m[7] ),
    .A2(_3132_),
    .B1(_3394_),
    .X(_0275_));
 sky130_fd_sc_hd__and2_1 _7188_ (.A(\sound3.count[8] ),
    .B(_2863_),
    .X(_3395_));
 sky130_fd_sc_hd__a21o_1 _7189_ (.A1(\sound3.count_m[8] ),
    .A2(_3132_),
    .B1(_3395_),
    .X(_0276_));
 sky130_fd_sc_hd__and2_1 _7190_ (.A(\sound3.count[9] ),
    .B(_2863_),
    .X(_3396_));
 sky130_fd_sc_hd__a21o_1 _7191_ (.A1(\sound3.count_m[9] ),
    .A2(_3132_),
    .B1(_3396_),
    .X(_0277_));
 sky130_fd_sc_hd__and2_1 _7192_ (.A(\sound3.count[10] ),
    .B(_2863_),
    .X(_3397_));
 sky130_fd_sc_hd__a21o_1 _7193_ (.A1(\sound3.count_m[10] ),
    .A2(_3132_),
    .B1(_3397_),
    .X(_0278_));
 sky130_fd_sc_hd__and2_1 _7194_ (.A(\sound3.count[11] ),
    .B(_2863_),
    .X(_3398_));
 sky130_fd_sc_hd__a21o_1 _7195_ (.A1(\sound3.count_m[11] ),
    .A2(_3132_),
    .B1(_3398_),
    .X(_0279_));
 sky130_fd_sc_hd__and2_1 _7196_ (.A(\sound3.count[12] ),
    .B(_2863_),
    .X(_3399_));
 sky130_fd_sc_hd__a21o_1 _7197_ (.A1(\sound3.count_m[12] ),
    .A2(_3132_),
    .B1(_3399_),
    .X(_0280_));
 sky130_fd_sc_hd__nor2_1 _7198_ (.A(_1658_),
    .B(_2843_),
    .Y(_3400_));
 sky130_fd_sc_hd__a21o_1 _7199_ (.A1(\sound3.count_m[13] ),
    .A2(_3132_),
    .B1(_3400_),
    .X(_0281_));
 sky130_fd_sc_hd__and2_1 _7200_ (.A(\sound3.count[14] ),
    .B(_2863_),
    .X(_3401_));
 sky130_fd_sc_hd__a21o_1 _7201_ (.A1(\sound3.count_m[14] ),
    .A2(_3132_),
    .B1(_3401_),
    .X(_0282_));
 sky130_fd_sc_hd__and2_1 _7202_ (.A(\sound3.count[15] ),
    .B(_2863_),
    .X(_3402_));
 sky130_fd_sc_hd__a21o_1 _7203_ (.A1(\sound3.count_m[15] ),
    .A2(_3132_),
    .B1(_3402_),
    .X(_0283_));
 sky130_fd_sc_hd__clkbuf_8 _7204_ (.A(_0554_),
    .X(_3403_));
 sky130_fd_sc_hd__and2_1 _7205_ (.A(\sound3.count[16] ),
    .B(_2863_),
    .X(_3404_));
 sky130_fd_sc_hd__a21o_1 _7206_ (.A1(\sound3.count_m[16] ),
    .A2(_3403_),
    .B1(_3404_),
    .X(_0284_));
 sky130_fd_sc_hd__and2_1 _7207_ (.A(\sound3.count[17] ),
    .B(_2863_),
    .X(_3405_));
 sky130_fd_sc_hd__a21o_1 _7208_ (.A1(\sound3.count_m[17] ),
    .A2(_3403_),
    .B1(_3405_),
    .X(_0285_));
 sky130_fd_sc_hd__and2_1 _7209_ (.A(\sound3.count[18] ),
    .B(_2863_),
    .X(_3406_));
 sky130_fd_sc_hd__a21o_1 _7210_ (.A1(\sound3.count_m[18] ),
    .A2(_3403_),
    .B1(_3406_),
    .X(_0286_));
 sky130_fd_sc_hd__mux2_1 _7211_ (.A0(\sound3.divisor_m[0] ),
    .A1(_1583_),
    .S(_3142_),
    .X(_3407_));
 sky130_fd_sc_hd__clkbuf_1 _7212_ (.A(_3407_),
    .X(_0287_));
 sky130_fd_sc_hd__inv_2 _7213_ (.A(_1673_),
    .Y(_3408_));
 sky130_fd_sc_hd__mux2_1 _7214_ (.A0(\sound3.divisor_m[1] ),
    .A1(_3408_),
    .S(_3142_),
    .X(_3409_));
 sky130_fd_sc_hd__clkbuf_1 _7215_ (.A(_3409_),
    .X(_0288_));
 sky130_fd_sc_hd__inv_2 _7216_ (.A(_1655_),
    .Y(_3410_));
 sky130_fd_sc_hd__mux2_1 _7217_ (.A0(\sound3.divisor_m[2] ),
    .A1(_3410_),
    .S(_3142_),
    .X(_3411_));
 sky130_fd_sc_hd__clkbuf_1 _7218_ (.A(_3411_),
    .X(_0289_));
 sky130_fd_sc_hd__inv_2 _7219_ (.A(_1641_),
    .Y(_3412_));
 sky130_fd_sc_hd__mux2_1 _7220_ (.A0(\sound3.divisor_m[3] ),
    .A1(_3412_),
    .S(_3142_),
    .X(_3413_));
 sky130_fd_sc_hd__clkbuf_1 _7221_ (.A(_3413_),
    .X(_0290_));
 sky130_fd_sc_hd__inv_2 _7222_ (.A(_1601_),
    .Y(_3414_));
 sky130_fd_sc_hd__mux2_1 _7223_ (.A0(\sound3.divisor_m[4] ),
    .A1(_3414_),
    .S(_3142_),
    .X(_3415_));
 sky130_fd_sc_hd__clkbuf_1 _7224_ (.A(_3415_),
    .X(_0291_));
 sky130_fd_sc_hd__inv_2 _7225_ (.A(_1635_),
    .Y(_3416_));
 sky130_fd_sc_hd__mux2_1 _7226_ (.A0(\sound3.divisor_m[5] ),
    .A1(_3416_),
    .S(_3142_),
    .X(_3417_));
 sky130_fd_sc_hd__clkbuf_1 _7227_ (.A(_3417_),
    .X(_0292_));
 sky130_fd_sc_hd__mux2_1 _7228_ (.A0(\sound3.divisor_m[6] ),
    .A1(_1594_),
    .S(_3142_),
    .X(_3418_));
 sky130_fd_sc_hd__clkbuf_1 _7229_ (.A(_3418_),
    .X(_0293_));
 sky130_fd_sc_hd__buf_8 _7230_ (.A(_2863_),
    .X(_3419_));
 sky130_fd_sc_hd__mux2_1 _7231_ (.A0(\sound3.divisor_m[7] ),
    .A1(_1649_),
    .S(_3419_),
    .X(_3420_));
 sky130_fd_sc_hd__clkbuf_1 _7232_ (.A(_3420_),
    .X(_0294_));
 sky130_fd_sc_hd__nand2_1 _7233_ (.A(\sound3.divisor_m[8] ),
    .B(_2843_),
    .Y(_3421_));
 sky130_fd_sc_hd__o21ai_1 _7234_ (.A1(_2843_),
    .A2(_1706_),
    .B1(_3421_),
    .Y(_0295_));
 sky130_fd_sc_hd__inv_2 _7235_ (.A(_1714_),
    .Y(_3422_));
 sky130_fd_sc_hd__mux2_1 _7236_ (.A0(\sound3.divisor_m[9] ),
    .A1(_3422_),
    .S(_3419_),
    .X(_3423_));
 sky130_fd_sc_hd__clkbuf_1 _7237_ (.A(_3423_),
    .X(_0296_));
 sky130_fd_sc_hd__mux2_1 _7238_ (.A0(\sound3.divisor_m[10] ),
    .A1(_1690_),
    .S(_3419_),
    .X(_3424_));
 sky130_fd_sc_hd__clkbuf_1 _7239_ (.A(_3424_),
    .X(_0297_));
 sky130_fd_sc_hd__inv_2 _7240_ (.A(_1699_),
    .Y(_3425_));
 sky130_fd_sc_hd__mux2_1 _7241_ (.A0(\sound3.divisor_m[11] ),
    .A1(_3425_),
    .S(_3419_),
    .X(_3426_));
 sky130_fd_sc_hd__clkbuf_1 _7242_ (.A(_3426_),
    .X(_0298_));
 sky130_fd_sc_hd__inv_2 _7243_ (.A(_1681_),
    .Y(_3427_));
 sky130_fd_sc_hd__mux2_1 _7244_ (.A0(\sound3.divisor_m[12] ),
    .A1(_3427_),
    .S(_3419_),
    .X(_3428_));
 sky130_fd_sc_hd__clkbuf_1 _7245_ (.A(_3428_),
    .X(_0299_));
 sky130_fd_sc_hd__mux2_1 _7246_ (.A0(\sound3.divisor_m[13] ),
    .A1(_1667_),
    .S(_3419_),
    .X(_3429_));
 sky130_fd_sc_hd__clkbuf_1 _7247_ (.A(_3429_),
    .X(_0300_));
 sky130_fd_sc_hd__mux2_1 _7248_ (.A0(\sound3.divisor_m[14] ),
    .A1(_1628_),
    .S(_3419_),
    .X(_3430_));
 sky130_fd_sc_hd__clkbuf_1 _7249_ (.A(_3430_),
    .X(_0301_));
 sky130_fd_sc_hd__inv_2 _7250_ (.A(_1615_),
    .Y(_3431_));
 sky130_fd_sc_hd__mux2_1 _7251_ (.A0(\sound3.divisor_m[15] ),
    .A1(_3431_),
    .S(_3419_),
    .X(_3432_));
 sky130_fd_sc_hd__clkbuf_1 _7252_ (.A(_3432_),
    .X(_0302_));
 sky130_fd_sc_hd__inv_2 _7253_ (.A(_1608_),
    .Y(_3433_));
 sky130_fd_sc_hd__mux2_1 _7254_ (.A0(\sound3.divisor_m[16] ),
    .A1(_3433_),
    .S(_3419_),
    .X(_3434_));
 sky130_fd_sc_hd__clkbuf_1 _7255_ (.A(_3434_),
    .X(_0303_));
 sky130_fd_sc_hd__mux2_1 _7256_ (.A0(\sound3.divisor_m[17] ),
    .A1(_1604_),
    .S(_3419_),
    .X(_3435_));
 sky130_fd_sc_hd__clkbuf_1 _7257_ (.A(_3435_),
    .X(_0304_));
 sky130_fd_sc_hd__or2_1 _7258_ (.A(_2543_),
    .B(_2005_),
    .X(_3436_));
 sky130_fd_sc_hd__o21ai_1 _7259_ (.A1(_2843_),
    .A2(_1618_),
    .B1(_3436_),
    .Y(_0305_));
 sky130_fd_sc_hd__buf_6 _7260_ (.A(_1545_),
    .X(_3437_));
 sky130_fd_sc_hd__nand2_1 _7261_ (.A(\sound3.divisor_m[0] ),
    .B(\sound3.sdiv.Q[27] ),
    .Y(_3438_));
 sky130_fd_sc_hd__or2_1 _7262_ (.A(\sound3.divisor_m[0] ),
    .B(\sound3.sdiv.Q[27] ),
    .X(_3439_));
 sky130_fd_sc_hd__clkbuf_8 _7263_ (.A(_0577_),
    .X(_3440_));
 sky130_fd_sc_hd__a32o_1 _7264_ (.A1(_3437_),
    .A2(_3438_),
    .A3(_3439_),
    .B1(_3440_),
    .B2(\sound3.sdiv.A[0] ),
    .X(_0306_));
 sky130_fd_sc_hd__and2b_1 _7265_ (.A_N(\sound3.sdiv.A[26] ),
    .B(\sound3.divisor_m[0] ),
    .X(_3441_));
 sky130_fd_sc_hd__xnor2_1 _7266_ (.A(\sound3.divisor_m[1] ),
    .B(_3441_),
    .Y(_3442_));
 sky130_fd_sc_hd__xnor2_1 _7267_ (.A(\sound3.sdiv.A[0] ),
    .B(_3442_),
    .Y(_3443_));
 sky130_fd_sc_hd__or2b_1 _7268_ (.A(_3438_),
    .B_N(_3443_),
    .X(_3444_));
 sky130_fd_sc_hd__a21o_1 _7269_ (.A1(\sound3.divisor_m[0] ),
    .A2(\sound3.sdiv.Q[27] ),
    .B1(_3443_),
    .X(_3445_));
 sky130_fd_sc_hd__a32o_1 _7270_ (.A1(_3437_),
    .A2(_3444_),
    .A3(_3445_),
    .B1(_3440_),
    .B2(\sound3.sdiv.A[1] ),
    .X(_0307_));
 sky130_fd_sc_hd__or2b_1 _7271_ (.A(_3442_),
    .B_N(\sound3.sdiv.A[0] ),
    .X(_3446_));
 sky130_fd_sc_hd__inv_2 _7272_ (.A(\sound3.sdiv.A[1] ),
    .Y(_3447_));
 sky130_fd_sc_hd__inv_4 _7273_ (.A(\sound3.sdiv.A[26] ),
    .Y(_3448_));
 sky130_fd_sc_hd__o21a_1 _7274_ (.A1(\sound3.divisor_m[1] ),
    .A2(\sound3.divisor_m[0] ),
    .B1(_3448_),
    .X(_3449_));
 sky130_fd_sc_hd__xnor2_1 _7275_ (.A(\sound3.divisor_m[2] ),
    .B(_3449_),
    .Y(_3450_));
 sky130_fd_sc_hd__xnor2_1 _7276_ (.A(_3447_),
    .B(_3450_),
    .Y(_3451_));
 sky130_fd_sc_hd__a21o_1 _7277_ (.A1(_3446_),
    .A2(_3444_),
    .B1(_3451_),
    .X(_3452_));
 sky130_fd_sc_hd__nand3_1 _7278_ (.A(_3446_),
    .B(_3444_),
    .C(_3451_),
    .Y(_3453_));
 sky130_fd_sc_hd__a32o_1 _7279_ (.A1(_3437_),
    .A2(_3452_),
    .A3(_3453_),
    .B1(_3440_),
    .B2(\sound3.sdiv.A[2] ),
    .X(_0308_));
 sky130_fd_sc_hd__or2_1 _7280_ (.A(_3447_),
    .B(_3450_),
    .X(_3454_));
 sky130_fd_sc_hd__inv_2 _7281_ (.A(\sound3.sdiv.A[2] ),
    .Y(_3455_));
 sky130_fd_sc_hd__o31a_1 _7282_ (.A1(\sound3.divisor_m[2] ),
    .A2(\sound3.divisor_m[1] ),
    .A3(\sound3.divisor_m[0] ),
    .B1(_3448_),
    .X(_3456_));
 sky130_fd_sc_hd__xnor2_1 _7283_ (.A(\sound3.divisor_m[3] ),
    .B(_3456_),
    .Y(_3457_));
 sky130_fd_sc_hd__nor2_1 _7284_ (.A(_3455_),
    .B(_3457_),
    .Y(_3458_));
 sky130_fd_sc_hd__and2_1 _7285_ (.A(_3455_),
    .B(_3457_),
    .X(_3459_));
 sky130_fd_sc_hd__or2_1 _7286_ (.A(_3458_),
    .B(_3459_),
    .X(_3460_));
 sky130_fd_sc_hd__a21oi_1 _7287_ (.A1(_3454_),
    .A2(_3452_),
    .B1(_3460_),
    .Y(_3461_));
 sky130_fd_sc_hd__a311o_1 _7288_ (.A1(_3454_),
    .A2(_3452_),
    .A3(_3460_),
    .B1(_0563_),
    .C1(_2005_),
    .X(_3462_));
 sky130_fd_sc_hd__clkbuf_8 _7289_ (.A(_0577_),
    .X(_3463_));
 sky130_fd_sc_hd__a2bb2o_1 _7290_ (.A1_N(_3461_),
    .A2_N(_3462_),
    .B1(\sound3.sdiv.A[3] ),
    .B2(_3463_),
    .X(_0309_));
 sky130_fd_sc_hd__inv_2 _7291_ (.A(\sound3.sdiv.A[3] ),
    .Y(_3464_));
 sky130_fd_sc_hd__or4_1 _7292_ (.A(\sound3.divisor_m[3] ),
    .B(\sound3.divisor_m[2] ),
    .C(\sound3.divisor_m[1] ),
    .D(\sound3.divisor_m[0] ),
    .X(_3465_));
 sky130_fd_sc_hd__nand2_1 _7293_ (.A(_3448_),
    .B(_3465_),
    .Y(_3466_));
 sky130_fd_sc_hd__xor2_1 _7294_ (.A(\sound3.divisor_m[4] ),
    .B(_3466_),
    .X(_3467_));
 sky130_fd_sc_hd__nor2_1 _7295_ (.A(_3464_),
    .B(_3467_),
    .Y(_3468_));
 sky130_fd_sc_hd__and2_1 _7296_ (.A(_3464_),
    .B(_3467_),
    .X(_3469_));
 sky130_fd_sc_hd__or2_1 _7297_ (.A(_3468_),
    .B(_3469_),
    .X(_3470_));
 sky130_fd_sc_hd__o21ba_1 _7298_ (.A1(_3458_),
    .A2(_3461_),
    .B1_N(_3470_),
    .X(_3471_));
 sky130_fd_sc_hd__or3b_1 _7299_ (.A(_3458_),
    .B(_3461_),
    .C_N(_3470_),
    .X(_3472_));
 sky130_fd_sc_hd__nand2_1 _7300_ (.A(_1545_),
    .B(_3472_),
    .Y(_3473_));
 sky130_fd_sc_hd__a2bb2o_1 _7301_ (.A1_N(_3471_),
    .A2_N(_3473_),
    .B1(\sound3.sdiv.A[4] ),
    .B2(_3463_),
    .X(_0310_));
 sky130_fd_sc_hd__inv_2 _7302_ (.A(\sound3.sdiv.A[4] ),
    .Y(_3474_));
 sky130_fd_sc_hd__o21a_1 _7303_ (.A1(\sound3.divisor_m[4] ),
    .A2(_3465_),
    .B1(_3448_),
    .X(_3475_));
 sky130_fd_sc_hd__xnor2_1 _7304_ (.A(\sound3.divisor_m[5] ),
    .B(_3475_),
    .Y(_3476_));
 sky130_fd_sc_hd__or2_1 _7305_ (.A(_3474_),
    .B(_3476_),
    .X(_3477_));
 sky130_fd_sc_hd__nand2_1 _7306_ (.A(_3474_),
    .B(_3476_),
    .Y(_3478_));
 sky130_fd_sc_hd__nand2_1 _7307_ (.A(_3477_),
    .B(_3478_),
    .Y(_3479_));
 sky130_fd_sc_hd__o21bai_2 _7308_ (.A1(_3468_),
    .A2(_3471_),
    .B1_N(_3479_),
    .Y(_3480_));
 sky130_fd_sc_hd__or3b_1 _7309_ (.A(_3468_),
    .B(_3471_),
    .C_N(_3479_),
    .X(_3481_));
 sky130_fd_sc_hd__a32o_1 _7310_ (.A1(_3437_),
    .A2(_3480_),
    .A3(_3481_),
    .B1(_3440_),
    .B2(\sound3.sdiv.A[5] ),
    .X(_0311_));
 sky130_fd_sc_hd__inv_2 _7311_ (.A(\sound3.sdiv.A[5] ),
    .Y(_3482_));
 sky130_fd_sc_hd__or3_1 _7312_ (.A(\sound3.divisor_m[5] ),
    .B(\sound3.divisor_m[4] ),
    .C(_3465_),
    .X(_3483_));
 sky130_fd_sc_hd__and2_1 _7313_ (.A(_3448_),
    .B(_3483_),
    .X(_3484_));
 sky130_fd_sc_hd__xnor2_1 _7314_ (.A(\sound3.divisor_m[6] ),
    .B(_3484_),
    .Y(_3485_));
 sky130_fd_sc_hd__or2_1 _7315_ (.A(_3482_),
    .B(_3485_),
    .X(_3486_));
 sky130_fd_sc_hd__nand2_1 _7316_ (.A(_3482_),
    .B(_3485_),
    .Y(_3487_));
 sky130_fd_sc_hd__nand2_1 _7317_ (.A(_3486_),
    .B(_3487_),
    .Y(_3488_));
 sky130_fd_sc_hd__nand3_1 _7318_ (.A(_3477_),
    .B(_3480_),
    .C(_3488_),
    .Y(_3489_));
 sky130_fd_sc_hd__a21o_1 _7319_ (.A1(_3477_),
    .A2(_3480_),
    .B1(_3488_),
    .X(_3490_));
 sky130_fd_sc_hd__a32o_1 _7320_ (.A1(_3437_),
    .A2(_3489_),
    .A3(_3490_),
    .B1(_3440_),
    .B2(\sound3.sdiv.A[6] ),
    .X(_0312_));
 sky130_fd_sc_hd__inv_2 _7321_ (.A(\sound3.sdiv.A[6] ),
    .Y(_3491_));
 sky130_fd_sc_hd__or2_1 _7322_ (.A(\sound3.divisor_m[6] ),
    .B(_3483_),
    .X(_3492_));
 sky130_fd_sc_hd__and2_1 _7323_ (.A(_3448_),
    .B(_3492_),
    .X(_3493_));
 sky130_fd_sc_hd__xnor2_1 _7324_ (.A(\sound3.divisor_m[7] ),
    .B(_3493_),
    .Y(_3494_));
 sky130_fd_sc_hd__or2_1 _7325_ (.A(_3491_),
    .B(_3494_),
    .X(_3495_));
 sky130_fd_sc_hd__nand2_1 _7326_ (.A(_3491_),
    .B(_3494_),
    .Y(_3496_));
 sky130_fd_sc_hd__nand2_1 _7327_ (.A(_3495_),
    .B(_3496_),
    .Y(_3497_));
 sky130_fd_sc_hd__nand3_1 _7328_ (.A(_3486_),
    .B(_3490_),
    .C(_3497_),
    .Y(_3498_));
 sky130_fd_sc_hd__a21o_1 _7329_ (.A1(_3486_),
    .A2(_3490_),
    .B1(_3497_),
    .X(_3499_));
 sky130_fd_sc_hd__a32o_1 _7330_ (.A1(_3437_),
    .A2(_3498_),
    .A3(_3499_),
    .B1(_3440_),
    .B2(\sound3.sdiv.A[7] ),
    .X(_0313_));
 sky130_fd_sc_hd__inv_2 _7331_ (.A(\sound3.sdiv.A[7] ),
    .Y(_3500_));
 sky130_fd_sc_hd__o21a_1 _7332_ (.A1(\sound3.divisor_m[7] ),
    .A2(_3492_),
    .B1(_3448_),
    .X(_3501_));
 sky130_fd_sc_hd__xnor2_1 _7333_ (.A(\sound3.divisor_m[8] ),
    .B(_3501_),
    .Y(_3502_));
 sky130_fd_sc_hd__or2_2 _7334_ (.A(_3500_),
    .B(_3502_),
    .X(_3503_));
 sky130_fd_sc_hd__nand2_1 _7335_ (.A(_3500_),
    .B(_3502_),
    .Y(_3504_));
 sky130_fd_sc_hd__nand2_1 _7336_ (.A(_3503_),
    .B(_3504_),
    .Y(_3505_));
 sky130_fd_sc_hd__nand3_1 _7337_ (.A(_3495_),
    .B(_3499_),
    .C(_3505_),
    .Y(_3506_));
 sky130_fd_sc_hd__a21o_1 _7338_ (.A1(_3495_),
    .A2(_3499_),
    .B1(_3505_),
    .X(_3507_));
 sky130_fd_sc_hd__a32o_1 _7339_ (.A1(_3437_),
    .A2(_3506_),
    .A3(_3507_),
    .B1(_3440_),
    .B2(\sound3.sdiv.A[8] ),
    .X(_0314_));
 sky130_fd_sc_hd__a21o_1 _7340_ (.A1(\sound3.divisor_m[8] ),
    .A2(_3448_),
    .B1(_3501_),
    .X(_3508_));
 sky130_fd_sc_hd__xor2_1 _7341_ (.A(\sound3.divisor_m[9] ),
    .B(_3508_),
    .X(_3509_));
 sky130_fd_sc_hd__and2_1 _7342_ (.A(\sound3.sdiv.A[8] ),
    .B(_3509_),
    .X(_3510_));
 sky130_fd_sc_hd__nor2_1 _7343_ (.A(\sound3.sdiv.A[8] ),
    .B(_3509_),
    .Y(_3511_));
 sky130_fd_sc_hd__o211ai_1 _7344_ (.A1(_3510_),
    .A2(_3511_),
    .B1(_3503_),
    .C1(_3507_),
    .Y(_3512_));
 sky130_fd_sc_hd__a211o_1 _7345_ (.A1(_3503_),
    .A2(_3507_),
    .B1(_3510_),
    .C1(_3511_),
    .X(_3513_));
 sky130_fd_sc_hd__a32o_1 _7346_ (.A1(_3437_),
    .A2(_3512_),
    .A3(_3513_),
    .B1(_3440_),
    .B2(\sound3.sdiv.A[9] ),
    .X(_0315_));
 sky130_fd_sc_hd__inv_2 _7347_ (.A(\sound3.sdiv.A[9] ),
    .Y(_3514_));
 sky130_fd_sc_hd__or4_1 _7348_ (.A(\sound3.divisor_m[9] ),
    .B(\sound3.divisor_m[8] ),
    .C(\sound3.divisor_m[7] ),
    .D(_3492_),
    .X(_3515_));
 sky130_fd_sc_hd__and2_1 _7349_ (.A(_3448_),
    .B(_3515_),
    .X(_3516_));
 sky130_fd_sc_hd__xnor2_1 _7350_ (.A(\sound3.divisor_m[10] ),
    .B(_3516_),
    .Y(_3517_));
 sky130_fd_sc_hd__or2_1 _7351_ (.A(_3514_),
    .B(_3517_),
    .X(_3518_));
 sky130_fd_sc_hd__nand2_1 _7352_ (.A(_3514_),
    .B(_3517_),
    .Y(_3519_));
 sky130_fd_sc_hd__nand2_1 _7353_ (.A(_3518_),
    .B(_3519_),
    .Y(_3520_));
 sky130_fd_sc_hd__inv_2 _7354_ (.A(_3510_),
    .Y(_3521_));
 sky130_fd_sc_hd__a31o_1 _7355_ (.A1(_3503_),
    .A2(_3507_),
    .A3(_3521_),
    .B1(_3511_),
    .X(_3522_));
 sky130_fd_sc_hd__nand2_1 _7356_ (.A(_3520_),
    .B(_3522_),
    .Y(_3523_));
 sky130_fd_sc_hd__a311o_1 _7357_ (.A1(_3503_),
    .A2(_3507_),
    .A3(_3521_),
    .B1(_3511_),
    .C1(_3520_),
    .X(_3524_));
 sky130_fd_sc_hd__a32o_1 _7358_ (.A1(_3437_),
    .A2(_3523_),
    .A3(_3524_),
    .B1(_3440_),
    .B2(\sound3.sdiv.A[10] ),
    .X(_0316_));
 sky130_fd_sc_hd__inv_2 _7359_ (.A(\sound3.sdiv.A[10] ),
    .Y(_3525_));
 sky130_fd_sc_hd__or2_1 _7360_ (.A(\sound3.divisor_m[10] ),
    .B(_3515_),
    .X(_3526_));
 sky130_fd_sc_hd__and2_1 _7361_ (.A(_3448_),
    .B(_3526_),
    .X(_3527_));
 sky130_fd_sc_hd__xnor2_1 _7362_ (.A(\sound3.divisor_m[11] ),
    .B(_3527_),
    .Y(_3528_));
 sky130_fd_sc_hd__nor2_1 _7363_ (.A(_3525_),
    .B(_3528_),
    .Y(_3529_));
 sky130_fd_sc_hd__and2_1 _7364_ (.A(_3525_),
    .B(_3528_),
    .X(_3530_));
 sky130_fd_sc_hd__or2_1 _7365_ (.A(_3529_),
    .B(_3530_),
    .X(_3531_));
 sky130_fd_sc_hd__a21oi_1 _7366_ (.A1(_3518_),
    .A2(_3524_),
    .B1(_3531_),
    .Y(_3532_));
 sky130_fd_sc_hd__a311o_1 _7367_ (.A1(_3518_),
    .A2(_3524_),
    .A3(_3531_),
    .B1(_0563_),
    .C1(_2005_),
    .X(_3533_));
 sky130_fd_sc_hd__a2bb2o_1 _7368_ (.A1_N(_3532_),
    .A2_N(_3533_),
    .B1(\sound3.sdiv.A[11] ),
    .B2(_3463_),
    .X(_0317_));
 sky130_fd_sc_hd__inv_2 _7369_ (.A(\sound3.sdiv.A[11] ),
    .Y(_3534_));
 sky130_fd_sc_hd__o21a_1 _7370_ (.A1(\sound3.divisor_m[11] ),
    .A2(_3526_),
    .B1(_3448_),
    .X(_3535_));
 sky130_fd_sc_hd__xnor2_1 _7371_ (.A(\sound3.divisor_m[12] ),
    .B(_3535_),
    .Y(_3536_));
 sky130_fd_sc_hd__or2_1 _7372_ (.A(_3534_),
    .B(_3536_),
    .X(_3537_));
 sky130_fd_sc_hd__nand2_1 _7373_ (.A(_3534_),
    .B(_3536_),
    .Y(_3538_));
 sky130_fd_sc_hd__nand2_1 _7374_ (.A(_3537_),
    .B(_3538_),
    .Y(_3539_));
 sky130_fd_sc_hd__or3b_1 _7375_ (.A(_3529_),
    .B(_3532_),
    .C_N(_3539_),
    .X(_3540_));
 sky130_fd_sc_hd__o21bai_1 _7376_ (.A1(_3529_),
    .A2(_3532_),
    .B1_N(_3539_),
    .Y(_3541_));
 sky130_fd_sc_hd__a32o_1 _7377_ (.A1(_3437_),
    .A2(_3540_),
    .A3(_3541_),
    .B1(_3440_),
    .B2(\sound3.sdiv.A[12] ),
    .X(_0318_));
 sky130_fd_sc_hd__inv_2 _7378_ (.A(\sound3.sdiv.A[12] ),
    .Y(_3542_));
 sky130_fd_sc_hd__or3_1 _7379_ (.A(\sound3.divisor_m[12] ),
    .B(\sound3.divisor_m[11] ),
    .C(_3526_),
    .X(_3543_));
 sky130_fd_sc_hd__and2_1 _7380_ (.A(_3448_),
    .B(_3543_),
    .X(_3544_));
 sky130_fd_sc_hd__xnor2_1 _7381_ (.A(\sound3.divisor_m[13] ),
    .B(_3544_),
    .Y(_3545_));
 sky130_fd_sc_hd__or2_1 _7382_ (.A(_3542_),
    .B(_3545_),
    .X(_3546_));
 sky130_fd_sc_hd__nand2_1 _7383_ (.A(_3542_),
    .B(_3545_),
    .Y(_3547_));
 sky130_fd_sc_hd__nand2_1 _7384_ (.A(_3546_),
    .B(_3547_),
    .Y(_3548_));
 sky130_fd_sc_hd__a21o_1 _7385_ (.A1(_3537_),
    .A2(_3541_),
    .B1(_3548_),
    .X(_3549_));
 sky130_fd_sc_hd__nand3_1 _7386_ (.A(_3537_),
    .B(_3541_),
    .C(_3548_),
    .Y(_3550_));
 sky130_fd_sc_hd__a32o_1 _7387_ (.A1(_3437_),
    .A2(_3549_),
    .A3(_3550_),
    .B1(_3440_),
    .B2(\sound3.sdiv.A[13] ),
    .X(_0319_));
 sky130_fd_sc_hd__inv_2 _7388_ (.A(\sound3.sdiv.A[13] ),
    .Y(_3551_));
 sky130_fd_sc_hd__or2_1 _7389_ (.A(\sound3.divisor_m[13] ),
    .B(_3543_),
    .X(_3552_));
 sky130_fd_sc_hd__and2_1 _7390_ (.A(_3448_),
    .B(_3552_),
    .X(_3553_));
 sky130_fd_sc_hd__xnor2_1 _7391_ (.A(\sound3.divisor_m[14] ),
    .B(_3553_),
    .Y(_3554_));
 sky130_fd_sc_hd__or2_1 _7392_ (.A(_3551_),
    .B(_3554_),
    .X(_3555_));
 sky130_fd_sc_hd__nand2_1 _7393_ (.A(_3551_),
    .B(_3554_),
    .Y(_3556_));
 sky130_fd_sc_hd__nand2_1 _7394_ (.A(_3555_),
    .B(_3556_),
    .Y(_3557_));
 sky130_fd_sc_hd__nand3_1 _7395_ (.A(_3546_),
    .B(_3549_),
    .C(_3557_),
    .Y(_3558_));
 sky130_fd_sc_hd__a21o_1 _7396_ (.A1(_3546_),
    .A2(_3549_),
    .B1(_3557_),
    .X(_3559_));
 sky130_fd_sc_hd__a32o_1 _7397_ (.A1(_3437_),
    .A2(_3558_),
    .A3(_3559_),
    .B1(_3440_),
    .B2(\sound3.sdiv.A[14] ),
    .X(_0320_));
 sky130_fd_sc_hd__inv_2 _7398_ (.A(\sound3.sdiv.A[14] ),
    .Y(_3560_));
 sky130_fd_sc_hd__or2_1 _7399_ (.A(\sound3.divisor_m[14] ),
    .B(_3552_),
    .X(_3561_));
 sky130_fd_sc_hd__and2_1 _7400_ (.A(_3448_),
    .B(_3561_),
    .X(_3562_));
 sky130_fd_sc_hd__xnor2_1 _7401_ (.A(\sound3.divisor_m[15] ),
    .B(_3562_),
    .Y(_3563_));
 sky130_fd_sc_hd__or2_1 _7402_ (.A(_3560_),
    .B(_3563_),
    .X(_3564_));
 sky130_fd_sc_hd__nand2_1 _7403_ (.A(_3560_),
    .B(_3563_),
    .Y(_3565_));
 sky130_fd_sc_hd__nand2_1 _7404_ (.A(_3564_),
    .B(_3565_),
    .Y(_3566_));
 sky130_fd_sc_hd__nand3_1 _7405_ (.A(_3555_),
    .B(_3559_),
    .C(_3566_),
    .Y(_3567_));
 sky130_fd_sc_hd__a21o_1 _7406_ (.A1(_3555_),
    .A2(_3559_),
    .B1(_3566_),
    .X(_3568_));
 sky130_fd_sc_hd__a32o_1 _7407_ (.A1(_3437_),
    .A2(_3567_),
    .A3(_3568_),
    .B1(_3440_),
    .B2(\sound3.sdiv.A[15] ),
    .X(_0321_));
 sky130_fd_sc_hd__and2_1 _7408_ (.A(_3564_),
    .B(_3568_),
    .X(_3569_));
 sky130_fd_sc_hd__inv_2 _7409_ (.A(\sound3.sdiv.A[15] ),
    .Y(_3570_));
 sky130_fd_sc_hd__o21a_1 _7410_ (.A1(\sound3.divisor_m[15] ),
    .A2(_3561_),
    .B1(_3448_),
    .X(_3571_));
 sky130_fd_sc_hd__xnor2_1 _7411_ (.A(\sound3.divisor_m[16] ),
    .B(_3571_),
    .Y(_3572_));
 sky130_fd_sc_hd__nor2_1 _7412_ (.A(_3570_),
    .B(_3572_),
    .Y(_3573_));
 sky130_fd_sc_hd__and2_1 _7413_ (.A(_3570_),
    .B(_3572_),
    .X(_3574_));
 sky130_fd_sc_hd__or2_1 _7414_ (.A(_3573_),
    .B(_3574_),
    .X(_3575_));
 sky130_fd_sc_hd__xor2_1 _7415_ (.A(_3569_),
    .B(_3575_),
    .X(_3576_));
 sky130_fd_sc_hd__a22o_1 _7416_ (.A1(\sound3.sdiv.A[16] ),
    .A2(_3463_),
    .B1(\sound3.sdiv.next_dived ),
    .B2(_3576_),
    .X(_0322_));
 sky130_fd_sc_hd__inv_2 _7417_ (.A(\sound3.sdiv.A[16] ),
    .Y(_3577_));
 sky130_fd_sc_hd__or3_1 _7418_ (.A(\sound3.divisor_m[16] ),
    .B(\sound3.divisor_m[15] ),
    .C(_3561_),
    .X(_3578_));
 sky130_fd_sc_hd__and2_1 _7419_ (.A(_3448_),
    .B(_3578_),
    .X(_3579_));
 sky130_fd_sc_hd__xnor2_1 _7420_ (.A(\sound3.divisor_m[17] ),
    .B(_3579_),
    .Y(_3580_));
 sky130_fd_sc_hd__nor2_1 _7421_ (.A(_3577_),
    .B(_3580_),
    .Y(_3581_));
 sky130_fd_sc_hd__nand2_1 _7422_ (.A(_3577_),
    .B(_3580_),
    .Y(_3582_));
 sky130_fd_sc_hd__or2b_1 _7423_ (.A(_3581_),
    .B_N(_3582_),
    .X(_3583_));
 sky130_fd_sc_hd__o21bai_1 _7424_ (.A1(_3569_),
    .A2(_3575_),
    .B1_N(_3573_),
    .Y(_3584_));
 sky130_fd_sc_hd__xnor2_1 _7425_ (.A(_3583_),
    .B(_3584_),
    .Y(_3585_));
 sky130_fd_sc_hd__a22o_1 _7426_ (.A1(\sound3.sdiv.A[17] ),
    .A2(_3463_),
    .B1(\sound3.sdiv.next_dived ),
    .B2(_3585_),
    .X(_0323_));
 sky130_fd_sc_hd__inv_2 _7427_ (.A(\sound3.sdiv.A[17] ),
    .Y(_3586_));
 sky130_fd_sc_hd__o21a_1 _7428_ (.A1(\sound3.divisor_m[17] ),
    .A2(_3578_),
    .B1(_3448_),
    .X(_3587_));
 sky130_fd_sc_hd__xnor2_1 _7429_ (.A(\sound3.divisor_m[18] ),
    .B(_3587_),
    .Y(_3588_));
 sky130_fd_sc_hd__nor2_1 _7430_ (.A(_3586_),
    .B(_3588_),
    .Y(_3589_));
 sky130_fd_sc_hd__nand2_1 _7431_ (.A(_3586_),
    .B(_3588_),
    .Y(_3590_));
 sky130_fd_sc_hd__or2b_1 _7432_ (.A(_3589_),
    .B_N(_3590_),
    .X(_3591_));
 sky130_fd_sc_hd__a21o_1 _7433_ (.A1(_3582_),
    .A2(_3584_),
    .B1(_3581_),
    .X(_3592_));
 sky130_fd_sc_hd__xnor2_1 _7434_ (.A(_3591_),
    .B(_3592_),
    .Y(_3593_));
 sky130_fd_sc_hd__a22o_1 _7435_ (.A1(\sound3.sdiv.A[18] ),
    .A2(_3463_),
    .B1(\sound3.sdiv.next_dived ),
    .B2(_3593_),
    .X(_0324_));
 sky130_fd_sc_hd__o31a_1 _7436_ (.A1(\sound3.divisor_m[18] ),
    .A2(\sound3.divisor_m[17] ),
    .A3(_3578_),
    .B1(_3448_),
    .X(_3594_));
 sky130_fd_sc_hd__clkbuf_8 _7437_ (.A(_3594_),
    .X(_3595_));
 sky130_fd_sc_hd__xnor2_1 _7438_ (.A(\sound3.sdiv.A[18] ),
    .B(_3595_),
    .Y(_3596_));
 sky130_fd_sc_hd__a21o_1 _7439_ (.A1(_3590_),
    .A2(_3592_),
    .B1(_3589_),
    .X(_3597_));
 sky130_fd_sc_hd__xnor2_1 _7440_ (.A(_3596_),
    .B(_3597_),
    .Y(_3598_));
 sky130_fd_sc_hd__a22o_1 _7441_ (.A1(\sound3.sdiv.A[19] ),
    .A2(_3463_),
    .B1(\sound3.sdiv.next_dived ),
    .B2(_3598_),
    .X(_0325_));
 sky130_fd_sc_hd__xnor2_1 _7442_ (.A(\sound3.sdiv.A[19] ),
    .B(_3595_),
    .Y(_3599_));
 sky130_fd_sc_hd__nor2_1 _7443_ (.A(_3591_),
    .B(_3596_),
    .Y(_3600_));
 sky130_fd_sc_hd__inv_2 _7444_ (.A(_3600_),
    .Y(_3601_));
 sky130_fd_sc_hd__a2111o_1 _7445_ (.A1(_3564_),
    .A2(_3568_),
    .B1(_3575_),
    .C1(_3583_),
    .D1(_3601_),
    .X(_3602_));
 sky130_fd_sc_hd__o21a_1 _7446_ (.A1(_3573_),
    .A2(_3581_),
    .B1(_3582_),
    .X(_3603_));
 sky130_fd_sc_hd__o21a_1 _7447_ (.A1(\sound3.sdiv.A[18] ),
    .A2(_3595_),
    .B1(_3589_),
    .X(_3604_));
 sky130_fd_sc_hd__a221oi_2 _7448_ (.A1(\sound3.sdiv.A[18] ),
    .A2(_3595_),
    .B1(_3600_),
    .B2(_3603_),
    .C1(_3604_),
    .Y(_3605_));
 sky130_fd_sc_hd__and3_1 _7449_ (.A(_3599_),
    .B(_3602_),
    .C(_3605_),
    .X(_3606_));
 sky130_fd_sc_hd__a21oi_2 _7450_ (.A1(_3602_),
    .A2(_3605_),
    .B1(_3599_),
    .Y(_3607_));
 sky130_fd_sc_hd__nor2_1 _7451_ (.A(_3606_),
    .B(_3607_),
    .Y(_3608_));
 sky130_fd_sc_hd__a22o_1 _7452_ (.A1(\sound3.sdiv.A[20] ),
    .A2(_3463_),
    .B1(\sound3.sdiv.next_dived ),
    .B2(_3608_),
    .X(_0326_));
 sky130_fd_sc_hd__xor2_1 _7453_ (.A(\sound3.sdiv.A[20] ),
    .B(_3595_),
    .X(_3609_));
 sky130_fd_sc_hd__a21oi_1 _7454_ (.A1(\sound3.sdiv.A[19] ),
    .A2(_3595_),
    .B1(_3607_),
    .Y(_3610_));
 sky130_fd_sc_hd__xnor2_1 _7455_ (.A(_3609_),
    .B(_3610_),
    .Y(_3611_));
 sky130_fd_sc_hd__a22o_1 _7456_ (.A1(\sound3.sdiv.A[21] ),
    .A2(_3463_),
    .B1(\sound3.sdiv.next_dived ),
    .B2(_3611_),
    .X(_0327_));
 sky130_fd_sc_hd__xnor2_1 _7457_ (.A(\sound3.sdiv.A[21] ),
    .B(_3595_),
    .Y(_3612_));
 sky130_fd_sc_hd__o21ai_1 _7458_ (.A1(\sound3.sdiv.A[20] ),
    .A2(_3595_),
    .B1(_3607_),
    .Y(_3613_));
 sky130_fd_sc_hd__o21ai_1 _7459_ (.A1(\sound3.sdiv.A[20] ),
    .A2(\sound3.sdiv.A[19] ),
    .B1(_3595_),
    .Y(_3614_));
 sky130_fd_sc_hd__and3_1 _7460_ (.A(_3612_),
    .B(_3613_),
    .C(_3614_),
    .X(_3615_));
 sky130_fd_sc_hd__a21oi_1 _7461_ (.A1(_3613_),
    .A2(_3614_),
    .B1(_3612_),
    .Y(_3616_));
 sky130_fd_sc_hd__or3_1 _7462_ (.A(_2863_),
    .B(_0563_),
    .C(_3616_),
    .X(_3617_));
 sky130_fd_sc_hd__a2bb2o_1 _7463_ (.A1_N(_3615_),
    .A2_N(_3617_),
    .B1(\sound3.sdiv.A[22] ),
    .B2(_3463_),
    .X(_0328_));
 sky130_fd_sc_hd__xor2_1 _7464_ (.A(\sound3.sdiv.A[22] ),
    .B(_3595_),
    .X(_3618_));
 sky130_fd_sc_hd__a21oi_1 _7465_ (.A1(\sound3.sdiv.A[21] ),
    .A2(_3595_),
    .B1(_3616_),
    .Y(_3619_));
 sky130_fd_sc_hd__xnor2_1 _7466_ (.A(_3618_),
    .B(_3619_),
    .Y(_3620_));
 sky130_fd_sc_hd__a22o_1 _7467_ (.A1(\sound3.sdiv.A[23] ),
    .A2(_3463_),
    .B1(\sound3.sdiv.next_dived ),
    .B2(_3620_),
    .X(_0329_));
 sky130_fd_sc_hd__or2_1 _7468_ (.A(\sound3.sdiv.A[23] ),
    .B(_3595_),
    .X(_3621_));
 sky130_fd_sc_hd__nand2_1 _7469_ (.A(\sound3.sdiv.A[23] ),
    .B(_3595_),
    .Y(_3622_));
 sky130_fd_sc_hd__nand2_1 _7470_ (.A(_3621_),
    .B(_3622_),
    .Y(_3623_));
 sky130_fd_sc_hd__inv_2 _7471_ (.A(_3609_),
    .Y(_3624_));
 sky130_fd_sc_hd__nor2_1 _7472_ (.A(_3624_),
    .B(_3612_),
    .Y(_3625_));
 sky130_fd_sc_hd__o41a_1 _7473_ (.A1(\sound3.sdiv.A[22] ),
    .A2(\sound3.sdiv.A[21] ),
    .A3(\sound3.sdiv.A[20] ),
    .A4(\sound3.sdiv.A[19] ),
    .B1(_3595_),
    .X(_3626_));
 sky130_fd_sc_hd__a31o_1 _7474_ (.A1(_3607_),
    .A2(_3618_),
    .A3(_3625_),
    .B1(_3626_),
    .X(_3627_));
 sky130_fd_sc_hd__xnor2_1 _7475_ (.A(_3623_),
    .B(_3627_),
    .Y(_3628_));
 sky130_fd_sc_hd__a22o_1 _7476_ (.A1(\sound3.sdiv.A[24] ),
    .A2(_3463_),
    .B1(\sound3.sdiv.next_dived ),
    .B2(_3628_),
    .X(_0330_));
 sky130_fd_sc_hd__a21boi_1 _7477_ (.A1(_3621_),
    .A2(_3627_),
    .B1_N(_3622_),
    .Y(_3629_));
 sky130_fd_sc_hd__nor2_1 _7478_ (.A(\sound3.sdiv.A[24] ),
    .B(_3595_),
    .Y(_3630_));
 sky130_fd_sc_hd__nand2_1 _7479_ (.A(\sound3.sdiv.A[24] ),
    .B(_3595_),
    .Y(_3631_));
 sky130_fd_sc_hd__and2b_1 _7480_ (.A_N(_3630_),
    .B(_3631_),
    .X(_3632_));
 sky130_fd_sc_hd__xnor2_1 _7481_ (.A(_3629_),
    .B(_3632_),
    .Y(_3633_));
 sky130_fd_sc_hd__a22o_1 _7482_ (.A1(\sound3.sdiv.A[25] ),
    .A2(_3463_),
    .B1(\sound3.sdiv.next_dived ),
    .B2(_3633_),
    .X(_0331_));
 sky130_fd_sc_hd__nand2_1 _7483_ (.A(\sound3.sdiv.A[25] ),
    .B(_3595_),
    .Y(_3634_));
 sky130_fd_sc_hd__or2_1 _7484_ (.A(\sound3.sdiv.A[25] ),
    .B(_3595_),
    .X(_3635_));
 sky130_fd_sc_hd__nand2_1 _7485_ (.A(_3634_),
    .B(_3635_),
    .Y(_3636_));
 sky130_fd_sc_hd__o211ai_1 _7486_ (.A1(_3629_),
    .A2(_3630_),
    .B1(_3631_),
    .C1(_3636_),
    .Y(_3637_));
 sky130_fd_sc_hd__or3b_1 _7487_ (.A(_3630_),
    .B(_3623_),
    .C_N(_3627_),
    .X(_3638_));
 sky130_fd_sc_hd__a31o_1 _7488_ (.A1(_3622_),
    .A2(_3631_),
    .A3(_3638_),
    .B1(_3636_),
    .X(_3639_));
 sky130_fd_sc_hd__a32o_1 _7489_ (.A1(_3437_),
    .A2(_3637_),
    .A3(_3639_),
    .B1(_3440_),
    .B2(\sound3.sdiv.A[26] ),
    .X(_0332_));
 sky130_fd_sc_hd__mux2_1 _7490_ (.A0(_1545_),
    .A1(_0577_),
    .S(\sound3.sdiv.C[0] ),
    .X(_3640_));
 sky130_fd_sc_hd__clkbuf_1 _7491_ (.A(_3640_),
    .X(_0333_));
 sky130_fd_sc_hd__nand2_1 _7492_ (.A(\sound3.sdiv.C[1] ),
    .B(\sound3.sdiv.C[0] ),
    .Y(_3641_));
 sky130_fd_sc_hd__or2_1 _7493_ (.A(\sound3.sdiv.C[1] ),
    .B(\sound3.sdiv.C[0] ),
    .X(_3642_));
 sky130_fd_sc_hd__a32o_1 _7494_ (.A1(_3437_),
    .A2(_3641_),
    .A3(_3642_),
    .B1(_3440_),
    .B2(\sound3.sdiv.C[1] ),
    .X(_0334_));
 sky130_fd_sc_hd__clkbuf_8 _7495_ (.A(_1545_),
    .X(_3643_));
 sky130_fd_sc_hd__a21o_1 _7496_ (.A1(\sound3.sdiv.C[1] ),
    .A2(\sound3.sdiv.C[0] ),
    .B1(\sound3.sdiv.C[2] ),
    .X(_3644_));
 sky130_fd_sc_hd__and3_1 _7497_ (.A(\sound3.sdiv.C[2] ),
    .B(\sound3.sdiv.C[1] ),
    .C(\sound3.sdiv.C[0] ),
    .X(_3645_));
 sky130_fd_sc_hd__inv_2 _7498_ (.A(_3645_),
    .Y(_3646_));
 sky130_fd_sc_hd__a32o_1 _7499_ (.A1(_3643_),
    .A2(_3644_),
    .A3(_3646_),
    .B1(_3440_),
    .B2(\sound3.sdiv.C[2] ),
    .X(_0335_));
 sky130_fd_sc_hd__and3_1 _7500_ (.A(\sound3.sdiv.C[3] ),
    .B(_0562_),
    .C(_3645_),
    .X(_3647_));
 sky130_fd_sc_hd__a21oi_1 _7501_ (.A1(_0562_),
    .A2(_3645_),
    .B1(\sound3.sdiv.C[3] ),
    .Y(_3648_));
 sky130_fd_sc_hd__nor3_1 _7502_ (.A(_2005_),
    .B(_3647_),
    .C(_3648_),
    .Y(_0336_));
 sky130_fd_sc_hd__a31o_1 _7503_ (.A1(\sound3.sdiv.C[3] ),
    .A2(_0562_),
    .A3(_3645_),
    .B1(\sound3.sdiv.C[4] ),
    .X(_3649_));
 sky130_fd_sc_hd__and2_1 _7504_ (.A(_2843_),
    .B(_3649_),
    .X(_3650_));
 sky130_fd_sc_hd__clkbuf_1 _7505_ (.A(_3650_),
    .X(_0337_));
 sky130_fd_sc_hd__and2_1 _7506_ (.A(\sound3.sdiv.C[5] ),
    .B(_0554_),
    .X(_3651_));
 sky130_fd_sc_hd__clkbuf_1 _7507_ (.A(_3651_),
    .X(_0338_));
 sky130_fd_sc_hd__or4_1 _7508_ (.A(\sound3.divisor_m[18] ),
    .B(\sound3.divisor_m[17] ),
    .C(\sound3.sdiv.A[26] ),
    .D(_3578_),
    .X(_3652_));
 sky130_fd_sc_hd__a311o_1 _7509_ (.A1(_3634_),
    .A2(_3639_),
    .A3(_3652_),
    .B1(_0563_),
    .C1(_2005_),
    .X(_3653_));
 sky130_fd_sc_hd__nand2_1 _7510_ (.A(_2275_),
    .B(_3653_),
    .Y(_0339_));
 sky130_fd_sc_hd__a22o_1 _7511_ (.A1(\sound3.sdiv.Q[1] ),
    .A2(_3463_),
    .B1(\sound3.sdiv.next_dived ),
    .B2(\sound3.sdiv.Q[0] ),
    .X(_0340_));
 sky130_fd_sc_hd__a22o_1 _7512_ (.A1(\sound3.sdiv.Q[2] ),
    .A2(_3463_),
    .B1(\sound3.sdiv.next_dived ),
    .B2(\sound3.sdiv.Q[1] ),
    .X(_0341_));
 sky130_fd_sc_hd__a22o_1 _7513_ (.A1(\sound3.sdiv.Q[3] ),
    .A2(_3463_),
    .B1(\sound3.sdiv.next_dived ),
    .B2(\sound3.sdiv.Q[2] ),
    .X(_0342_));
 sky130_fd_sc_hd__a22o_1 _7514_ (.A1(\sound3.sdiv.Q[4] ),
    .A2(_3463_),
    .B1(_3437_),
    .B2(\sound3.sdiv.Q[3] ),
    .X(_0343_));
 sky130_fd_sc_hd__a22o_1 _7515_ (.A1(\sound3.sdiv.Q[5] ),
    .A2(_3463_),
    .B1(_3437_),
    .B2(\sound3.sdiv.Q[4] ),
    .X(_0344_));
 sky130_fd_sc_hd__a22o_1 _7516_ (.A1(\sound3.sdiv.Q[6] ),
    .A2(_3440_),
    .B1(_3437_),
    .B2(\sound3.sdiv.Q[5] ),
    .X(_0345_));
 sky130_fd_sc_hd__a22o_1 _7517_ (.A1(\sound3.sdiv.Q[7] ),
    .A2(_3440_),
    .B1(_3437_),
    .B2(\sound3.sdiv.Q[6] ),
    .X(_0346_));
 sky130_fd_sc_hd__clkbuf_8 _7518_ (.A(_0577_),
    .X(_3654_));
 sky130_fd_sc_hd__a221o_1 _7519_ (.A1(\sound3.sdiv.Q[8] ),
    .A2(_3654_),
    .B1(_3643_),
    .B2(\sound3.sdiv.Q[7] ),
    .C1(_3387_),
    .X(_0347_));
 sky130_fd_sc_hd__a221o_1 _7520_ (.A1(\sound3.sdiv.Q[9] ),
    .A2(_3654_),
    .B1(_3643_),
    .B2(\sound3.sdiv.Q[8] ),
    .C1(_3388_),
    .X(_0348_));
 sky130_fd_sc_hd__a221o_1 _7521_ (.A1(\sound3.sdiv.Q[10] ),
    .A2(_3654_),
    .B1(_3643_),
    .B2(\sound3.sdiv.Q[9] ),
    .C1(_3389_),
    .X(_0349_));
 sky130_fd_sc_hd__a221o_1 _7522_ (.A1(\sound3.sdiv.Q[11] ),
    .A2(_3654_),
    .B1(_3643_),
    .B2(\sound3.sdiv.Q[10] ),
    .C1(_3390_),
    .X(_0350_));
 sky130_fd_sc_hd__a221o_1 _7523_ (.A1(\sound3.sdiv.Q[12] ),
    .A2(_3654_),
    .B1(_3643_),
    .B2(\sound3.sdiv.Q[11] ),
    .C1(_3391_),
    .X(_0351_));
 sky130_fd_sc_hd__a221o_1 _7524_ (.A1(\sound3.sdiv.Q[13] ),
    .A2(_3654_),
    .B1(_3643_),
    .B2(\sound3.sdiv.Q[12] ),
    .C1(_3392_),
    .X(_0352_));
 sky130_fd_sc_hd__a221o_1 _7525_ (.A1(\sound3.sdiv.Q[14] ),
    .A2(_3654_),
    .B1(_3643_),
    .B2(\sound3.sdiv.Q[13] ),
    .C1(_3393_),
    .X(_0353_));
 sky130_fd_sc_hd__a221o_1 _7526_ (.A1(\sound3.sdiv.Q[15] ),
    .A2(_3654_),
    .B1(_3643_),
    .B2(\sound3.sdiv.Q[14] ),
    .C1(_3394_),
    .X(_0354_));
 sky130_fd_sc_hd__a221o_1 _7527_ (.A1(\sound3.sdiv.Q[16] ),
    .A2(_3654_),
    .B1(_3643_),
    .B2(\sound3.sdiv.Q[15] ),
    .C1(_3395_),
    .X(_0355_));
 sky130_fd_sc_hd__a221o_1 _7528_ (.A1(\sound3.sdiv.Q[17] ),
    .A2(_3654_),
    .B1(_3643_),
    .B2(\sound3.sdiv.Q[16] ),
    .C1(_3396_),
    .X(_0356_));
 sky130_fd_sc_hd__a221o_1 _7529_ (.A1(\sound3.sdiv.Q[18] ),
    .A2(_3654_),
    .B1(_3643_),
    .B2(\sound3.sdiv.Q[17] ),
    .C1(_3397_),
    .X(_0357_));
 sky130_fd_sc_hd__a221o_1 _7530_ (.A1(\sound3.sdiv.Q[19] ),
    .A2(_3654_),
    .B1(_3643_),
    .B2(\sound3.sdiv.Q[18] ),
    .C1(_3398_),
    .X(_0358_));
 sky130_fd_sc_hd__a221o_1 _7531_ (.A1(\sound3.sdiv.Q[20] ),
    .A2(_3654_),
    .B1(_3643_),
    .B2(\sound3.sdiv.Q[19] ),
    .C1(_3399_),
    .X(_0359_));
 sky130_fd_sc_hd__a221o_1 _7532_ (.A1(\sound3.sdiv.Q[21] ),
    .A2(_3654_),
    .B1(_3643_),
    .B2(\sound3.sdiv.Q[20] ),
    .C1(_3400_),
    .X(_0360_));
 sky130_fd_sc_hd__a221o_1 _7533_ (.A1(\sound3.sdiv.Q[22] ),
    .A2(_3654_),
    .B1(_3643_),
    .B2(\sound3.sdiv.Q[21] ),
    .C1(_3401_),
    .X(_0361_));
 sky130_fd_sc_hd__a221o_1 _7534_ (.A1(\sound3.sdiv.Q[23] ),
    .A2(_3654_),
    .B1(_3643_),
    .B2(\sound3.sdiv.Q[22] ),
    .C1(_3402_),
    .X(_0362_));
 sky130_fd_sc_hd__a221o_1 _7535_ (.A1(\sound3.sdiv.Q[24] ),
    .A2(_3654_),
    .B1(_3643_),
    .B2(\sound3.sdiv.Q[23] ),
    .C1(_3404_),
    .X(_0363_));
 sky130_fd_sc_hd__a221o_1 _7536_ (.A1(\sound3.sdiv.Q[25] ),
    .A2(_3654_),
    .B1(_3643_),
    .B2(\sound3.sdiv.Q[24] ),
    .C1(_3405_),
    .X(_0364_));
 sky130_fd_sc_hd__a221o_1 _7537_ (.A1(\sound3.sdiv.Q[26] ),
    .A2(_3654_),
    .B1(_3643_),
    .B2(\sound3.sdiv.Q[25] ),
    .C1(_3406_),
    .X(_0365_));
 sky130_fd_sc_hd__a22o_1 _7538_ (.A1(\sound3.sdiv.Q[27] ),
    .A2(_3440_),
    .B1(_3437_),
    .B2(\sound3.sdiv.Q[26] ),
    .X(_0366_));
 sky130_fd_sc_hd__a21o_1 _7539_ (.A1(\sound4.count_m[0] ),
    .A2(_3403_),
    .B1(_2187_),
    .X(_0367_));
 sky130_fd_sc_hd__a21o_1 _7540_ (.A1(\sound4.count_m[1] ),
    .A2(_3403_),
    .B1(_2188_),
    .X(_0368_));
 sky130_fd_sc_hd__a21o_1 _7541_ (.A1(\sound4.count_m[2] ),
    .A2(_3403_),
    .B1(_2189_),
    .X(_0369_));
 sky130_fd_sc_hd__a21o_1 _7542_ (.A1(\sound4.count_m[3] ),
    .A2(_3403_),
    .B1(_2190_),
    .X(_0370_));
 sky130_fd_sc_hd__a21o_1 _7543_ (.A1(\sound4.count_m[4] ),
    .A2(_3403_),
    .B1(_2191_),
    .X(_0371_));
 sky130_fd_sc_hd__a21o_1 _7544_ (.A1(\sound4.count_m[5] ),
    .A2(_3403_),
    .B1(_2192_),
    .X(_0372_));
 sky130_fd_sc_hd__a21o_1 _7545_ (.A1(\sound4.count_m[6] ),
    .A2(_3403_),
    .B1(_2193_),
    .X(_0373_));
 sky130_fd_sc_hd__a21o_1 _7546_ (.A1(\sound4.count_m[7] ),
    .A2(_3403_),
    .B1(_2194_),
    .X(_0374_));
 sky130_fd_sc_hd__a21o_1 _7547_ (.A1(\sound4.count_m[8] ),
    .A2(_3403_),
    .B1(_2195_),
    .X(_0375_));
 sky130_fd_sc_hd__a21o_1 _7548_ (.A1(\sound4.count_m[9] ),
    .A2(_3403_),
    .B1(_2196_),
    .X(_0376_));
 sky130_fd_sc_hd__a21o_1 _7549_ (.A1(\sound4.count_m[10] ),
    .A2(_3403_),
    .B1(_2197_),
    .X(_0377_));
 sky130_fd_sc_hd__a21o_1 _7550_ (.A1(\sound4.count_m[11] ),
    .A2(_3403_),
    .B1(_2198_),
    .X(_0378_));
 sky130_fd_sc_hd__a21o_1 _7551_ (.A1(\sound4.count_m[12] ),
    .A2(_3403_),
    .B1(_2199_),
    .X(_0379_));
 sky130_fd_sc_hd__a21o_1 _7552_ (.A1(\sound4.count_m[13] ),
    .A2(_3403_),
    .B1(_2200_),
    .X(_0380_));
 sky130_fd_sc_hd__a21o_1 _7553_ (.A1(\sound4.count_m[14] ),
    .A2(_3403_),
    .B1(_2202_),
    .X(_0381_));
 sky130_fd_sc_hd__a21o_1 _7554_ (.A1(\sound4.count_m[15] ),
    .A2(_2843_),
    .B1(_2203_),
    .X(_0382_));
 sky130_fd_sc_hd__a21o_1 _7555_ (.A1(\sound4.count_m[16] ),
    .A2(_2843_),
    .B1(_2204_),
    .X(_0383_));
 sky130_fd_sc_hd__a21o_1 _7556_ (.A1(\sound4.count_m[17] ),
    .A2(_2843_),
    .B1(_2205_),
    .X(_0384_));
 sky130_fd_sc_hd__a21o_1 _7557_ (.A1(\sound4.count_m[18] ),
    .A2(_2843_),
    .B1(_2206_),
    .X(_0385_));
 sky130_fd_sc_hd__mux2_1 _7558_ (.A0(\sound4.divisor_m[0] ),
    .A1(_1859_),
    .S(_3419_),
    .X(_3655_));
 sky130_fd_sc_hd__clkbuf_1 _7559_ (.A(_3655_),
    .X(_0386_));
 sky130_fd_sc_hd__inv_2 _7560_ (.A(_1931_),
    .Y(_3656_));
 sky130_fd_sc_hd__mux2_1 _7561_ (.A0(\sound4.divisor_m[1] ),
    .A1(_3656_),
    .S(_3419_),
    .X(_3657_));
 sky130_fd_sc_hd__clkbuf_1 _7562_ (.A(_3657_),
    .X(_0387_));
 sky130_fd_sc_hd__inv_2 _7563_ (.A(_1903_),
    .Y(_3658_));
 sky130_fd_sc_hd__mux2_1 _7564_ (.A0(\sound4.divisor_m[2] ),
    .A1(_3658_),
    .S(_3419_),
    .X(_3659_));
 sky130_fd_sc_hd__clkbuf_1 _7565_ (.A(_3659_),
    .X(_0388_));
 sky130_fd_sc_hd__mux2_1 _7566_ (.A0(\sound4.divisor_m[3] ),
    .A1(_1850_),
    .S(_3419_),
    .X(_3660_));
 sky130_fd_sc_hd__clkbuf_1 _7567_ (.A(_3660_),
    .X(_0389_));
 sky130_fd_sc_hd__mux2_1 _7568_ (.A0(\sound4.divisor_m[4] ),
    .A1(_1866_),
    .S(_3419_),
    .X(_3661_));
 sky130_fd_sc_hd__clkbuf_1 _7569_ (.A(_3661_),
    .X(_0390_));
 sky130_fd_sc_hd__mux2_1 _7570_ (.A0(\sound4.divisor_m[5] ),
    .A1(_1810_),
    .S(_3419_),
    .X(_3662_));
 sky130_fd_sc_hd__clkbuf_1 _7571_ (.A(_3662_),
    .X(_0391_));
 sky130_fd_sc_hd__mux2_1 _7572_ (.A0(\sound4.divisor_m[6] ),
    .A1(_1884_),
    .S(_3419_),
    .X(_3663_));
 sky130_fd_sc_hd__clkbuf_1 _7573_ (.A(_3663_),
    .X(_0392_));
 sky130_fd_sc_hd__inv_2 _7574_ (.A(_1897_),
    .Y(_3664_));
 sky130_fd_sc_hd__mux2_1 _7575_ (.A0(\sound4.divisor_m[7] ),
    .A1(_3664_),
    .S(_3419_),
    .X(_3665_));
 sky130_fd_sc_hd__clkbuf_1 _7576_ (.A(_3665_),
    .X(_0393_));
 sky130_fd_sc_hd__inv_2 _7577_ (.A(_1829_),
    .Y(_3666_));
 sky130_fd_sc_hd__mux2_1 _7578_ (.A0(\sound4.divisor_m[8] ),
    .A1(_3666_),
    .S(_3419_),
    .X(_3667_));
 sky130_fd_sc_hd__clkbuf_1 _7579_ (.A(_3667_),
    .X(_0394_));
 sky130_fd_sc_hd__nor2_1 _7580_ (.A(\sound4.divisor_m[9] ),
    .B(_2005_),
    .Y(_3668_));
 sky130_fd_sc_hd__a21oi_1 _7581_ (.A1(_2005_),
    .A2(_1840_),
    .B1(_3668_),
    .Y(_0395_));
 sky130_fd_sc_hd__mux2_1 _7582_ (.A0(\sound4.divisor_m[10] ),
    .A1(_1803_),
    .S(_3419_),
    .X(_3669_));
 sky130_fd_sc_hd__clkbuf_1 _7583_ (.A(_3669_),
    .X(_0396_));
 sky130_fd_sc_hd__inv_2 _7584_ (.A(_1909_),
    .Y(_3670_));
 sky130_fd_sc_hd__mux2_1 _7585_ (.A0(\sound4.divisor_m[11] ),
    .A1(_3670_),
    .S(_2186_),
    .X(_3671_));
 sky130_fd_sc_hd__clkbuf_1 _7586_ (.A(_3671_),
    .X(_0397_));
 sky130_fd_sc_hd__mux2_1 _7587_ (.A0(\sound4.divisor_m[12] ),
    .A1(_1924_),
    .S(_2186_),
    .X(_3672_));
 sky130_fd_sc_hd__clkbuf_1 _7588_ (.A(_3672_),
    .X(_0398_));
 sky130_fd_sc_hd__mux2_1 _7589_ (.A0(\sound4.divisor_m[13] ),
    .A1(_1875_),
    .S(_2186_),
    .X(_3673_));
 sky130_fd_sc_hd__clkbuf_1 _7590_ (.A(_3673_),
    .X(_0399_));
 sky130_fd_sc_hd__inv_2 _7591_ (.A(_1817_),
    .Y(_3674_));
 sky130_fd_sc_hd__mux2_1 _7592_ (.A0(\sound4.divisor_m[14] ),
    .A1(_3674_),
    .S(_2186_),
    .X(_3675_));
 sky130_fd_sc_hd__clkbuf_1 _7593_ (.A(_3675_),
    .X(_0400_));
 sky130_fd_sc_hd__inv_2 _7594_ (.A(_1891_),
    .Y(_3676_));
 sky130_fd_sc_hd__mux2_1 _7595_ (.A0(\sound4.divisor_m[15] ),
    .A1(_3676_),
    .S(_2186_),
    .X(_3677_));
 sky130_fd_sc_hd__clkbuf_1 _7596_ (.A(_3677_),
    .X(_0401_));
 sky130_fd_sc_hd__or2_1 _7597_ (.A(_2341_),
    .B(_2005_),
    .X(_3678_));
 sky130_fd_sc_hd__o21ai_1 _7598_ (.A1(_2843_),
    .A2(_1820_),
    .B1(_3678_),
    .Y(_0402_));
 sky130_fd_sc_hd__and2_1 _7599_ (.A(\sound4.divisor_m[17] ),
    .B(_0554_),
    .X(_3679_));
 sky130_fd_sc_hd__a31o_1 _7600_ (.A1(_2005_),
    .A2(_1018_),
    .A3(_1779_),
    .B1(_3679_),
    .X(_0403_));
 sky130_fd_sc_hd__mux2_1 _7601_ (.A0(\sound4.divisor_m[18] ),
    .A1(_1913_),
    .S(_2186_),
    .X(_3680_));
 sky130_fd_sc_hd__clkbuf_1 _7602_ (.A(_3680_),
    .X(_0404_));
 sky130_fd_sc_hd__buf_6 _7603_ (.A(_1764_),
    .X(_3681_));
 sky130_fd_sc_hd__nand2_1 _7604_ (.A(\sound4.divisor_m[0] ),
    .B(\sound4.sdiv.Q[27] ),
    .Y(_3682_));
 sky130_fd_sc_hd__or2_1 _7605_ (.A(\sound4.divisor_m[0] ),
    .B(\sound4.sdiv.Q[27] ),
    .X(_3683_));
 sky130_fd_sc_hd__a32o_1 _7606_ (.A1(_3681_),
    .A2(_3682_),
    .A3(_3683_),
    .B1(_2184_),
    .B2(\sound4.sdiv.A[0] ),
    .X(_0405_));
 sky130_fd_sc_hd__xnor2_1 _7607_ (.A(_2123_),
    .B(_3682_),
    .Y(_3684_));
 sky130_fd_sc_hd__a22o_1 _7608_ (.A1(\sound4.sdiv.A[1] ),
    .A2(_2183_),
    .B1(\sound4.sdiv.next_dived ),
    .B2(_3684_),
    .X(_0406_));
 sky130_fd_sc_hd__or2_1 _7609_ (.A(_2120_),
    .B(_2125_),
    .X(_3685_));
 sky130_fd_sc_hd__nand2_1 _7610_ (.A(_2120_),
    .B(_2125_),
    .Y(_3686_));
 sky130_fd_sc_hd__a32o_1 _7611_ (.A1(_3681_),
    .A2(_3685_),
    .A3(_3686_),
    .B1(_2184_),
    .B2(\sound4.sdiv.A[2] ),
    .X(_0407_));
 sky130_fd_sc_hd__or2_1 _7612_ (.A(_2116_),
    .B(_2127_),
    .X(_3687_));
 sky130_fd_sc_hd__nand2_1 _7613_ (.A(_2116_),
    .B(_2127_),
    .Y(_3688_));
 sky130_fd_sc_hd__a32o_1 _7614_ (.A1(_3681_),
    .A2(_3687_),
    .A3(_3688_),
    .B1(_2184_),
    .B2(\sound4.sdiv.A[3] ),
    .X(_0408_));
 sky130_fd_sc_hd__and2_1 _7615_ (.A(_2110_),
    .B(_2128_),
    .X(_3689_));
 sky130_fd_sc_hd__inv_2 _7616_ (.A(_3689_),
    .Y(_3690_));
 sky130_fd_sc_hd__or2_1 _7617_ (.A(_2110_),
    .B(_2128_),
    .X(_3691_));
 sky130_fd_sc_hd__a32o_1 _7618_ (.A1(_3681_),
    .A2(_3690_),
    .A3(_3691_),
    .B1(_2184_),
    .B2(\sound4.sdiv.A[4] ),
    .X(_0409_));
 sky130_fd_sc_hd__nand2_1 _7619_ (.A(_2130_),
    .B(_2103_),
    .Y(_3692_));
 sky130_fd_sc_hd__or2b_1 _7620_ (.A(_3692_),
    .B_N(_2129_),
    .X(_3693_));
 sky130_fd_sc_hd__or2b_1 _7621_ (.A(_2129_),
    .B_N(_3692_),
    .X(_3694_));
 sky130_fd_sc_hd__a32o_1 _7622_ (.A1(_3681_),
    .A2(_3693_),
    .A3(_3694_),
    .B1(_2184_),
    .B2(\sound4.sdiv.A[5] ),
    .X(_0410_));
 sky130_fd_sc_hd__and2_1 _7623_ (.A(_2099_),
    .B(_2131_),
    .X(_3695_));
 sky130_fd_sc_hd__o21ai_1 _7624_ (.A1(_2099_),
    .A2(_2131_),
    .B1(_2185_),
    .Y(_3696_));
 sky130_fd_sc_hd__a2bb2o_1 _7625_ (.A1_N(_3695_),
    .A2_N(_3696_),
    .B1(\sound4.sdiv.A[6] ),
    .B2(_2183_),
    .X(_0411_));
 sky130_fd_sc_hd__nand2_1 _7626_ (.A(_2133_),
    .B(_2093_),
    .Y(_3697_));
 sky130_fd_sc_hd__or2b_1 _7627_ (.A(_3697_),
    .B_N(_2132_),
    .X(_3698_));
 sky130_fd_sc_hd__or2b_1 _7628_ (.A(_2132_),
    .B_N(_3697_),
    .X(_3699_));
 sky130_fd_sc_hd__a32o_1 _7629_ (.A1(_3681_),
    .A2(_3698_),
    .A3(_3699_),
    .B1(_2184_),
    .B2(\sound4.sdiv.A[7] ),
    .X(_0412_));
 sky130_fd_sc_hd__and2_1 _7630_ (.A(_2089_),
    .B(_2134_),
    .X(_3700_));
 sky130_fd_sc_hd__o21ai_1 _7631_ (.A1(_2089_),
    .A2(_2134_),
    .B1(_1764_),
    .Y(_3701_));
 sky130_fd_sc_hd__a2bb2o_1 _7632_ (.A1_N(_3700_),
    .A2_N(_3701_),
    .B1(\sound4.sdiv.A[8] ),
    .B2(_2183_),
    .X(_0413_));
 sky130_fd_sc_hd__nand2_1 _7633_ (.A(_2136_),
    .B(_2083_),
    .Y(_3702_));
 sky130_fd_sc_hd__or2b_1 _7634_ (.A(_3702_),
    .B_N(_2135_),
    .X(_3703_));
 sky130_fd_sc_hd__or2b_1 _7635_ (.A(_2135_),
    .B_N(_3702_),
    .X(_3704_));
 sky130_fd_sc_hd__a32o_1 _7636_ (.A1(_3681_),
    .A2(_3703_),
    .A3(_3704_),
    .B1(_2184_),
    .B2(\sound4.sdiv.A[9] ),
    .X(_0414_));
 sky130_fd_sc_hd__nor2_1 _7637_ (.A(_2079_),
    .B(_2137_),
    .Y(_3705_));
 sky130_fd_sc_hd__and2_1 _7638_ (.A(_2079_),
    .B(_2137_),
    .X(_3706_));
 sky130_fd_sc_hd__o32ai_1 _7639_ (.A1(_1763_),
    .A2(_3705_),
    .A3(_3706_),
    .B1(\sound4.sdiv.next_start ),
    .B2(_2070_),
    .Y(_0415_));
 sky130_fd_sc_hd__or2b_1 _7640_ (.A(_2139_),
    .B_N(_2073_),
    .X(_3707_));
 sky130_fd_sc_hd__or2b_1 _7641_ (.A(_3707_),
    .B_N(_2138_),
    .X(_3708_));
 sky130_fd_sc_hd__or2b_1 _7642_ (.A(_2138_),
    .B_N(_3707_),
    .X(_3709_));
 sky130_fd_sc_hd__a32o_1 _7643_ (.A1(_3681_),
    .A2(_3708_),
    .A3(_3709_),
    .B1(_2184_),
    .B2(\sound4.sdiv.A[11] ),
    .X(_0416_));
 sky130_fd_sc_hd__nand2_1 _7644_ (.A(_2069_),
    .B(_2140_),
    .Y(_3710_));
 sky130_fd_sc_hd__or2_1 _7645_ (.A(_2069_),
    .B(_2140_),
    .X(_3711_));
 sky130_fd_sc_hd__a32o_1 _7646_ (.A1(_3681_),
    .A2(_3710_),
    .A3(_3711_),
    .B1(_2184_),
    .B2(\sound4.sdiv.A[12] ),
    .X(_0417_));
 sky130_fd_sc_hd__nand2_1 _7647_ (.A(_2066_),
    .B(_3710_),
    .Y(_3712_));
 sky130_fd_sc_hd__xnor2_1 _7648_ (.A(_2058_),
    .B(_2060_),
    .Y(_3713_));
 sky130_fd_sc_hd__xnor2_1 _7649_ (.A(_3712_),
    .B(_3713_),
    .Y(_3714_));
 sky130_fd_sc_hd__a22o_1 _7650_ (.A1(\sound4.sdiv.A[13] ),
    .A2(_2183_),
    .B1(\sound4.sdiv.next_dived ),
    .B2(_3714_),
    .X(_0418_));
 sky130_fd_sc_hd__nand3_1 _7651_ (.A(_2057_),
    .B(_2061_),
    .C(_2141_),
    .Y(_3715_));
 sky130_fd_sc_hd__a21o_1 _7652_ (.A1(_2061_),
    .A2(_2141_),
    .B1(_2057_),
    .X(_3716_));
 sky130_fd_sc_hd__a32o_1 _7653_ (.A1(_3681_),
    .A2(_3715_),
    .A3(_3716_),
    .B1(_2184_),
    .B2(\sound4.sdiv.A[14] ),
    .X(_0419_));
 sky130_fd_sc_hd__nand2_1 _7654_ (.A(_2150_),
    .B(_3715_),
    .Y(_3717_));
 sky130_fd_sc_hd__xor2_1 _7655_ (.A(_3717_),
    .B(_2148_),
    .X(_3718_));
 sky130_fd_sc_hd__a22o_1 _7656_ (.A1(\sound4.sdiv.A[15] ),
    .A2(_2183_),
    .B1(\sound4.sdiv.next_dived ),
    .B2(_3718_),
    .X(_0420_));
 sky130_fd_sc_hd__a31o_1 _7657_ (.A1(_2145_),
    .A2(_2150_),
    .A3(_3715_),
    .B1(_2147_),
    .X(_3719_));
 sky130_fd_sc_hd__or2_1 _7658_ (.A(_3719_),
    .B(_2154_),
    .X(_3720_));
 sky130_fd_sc_hd__nand2_1 _7659_ (.A(_3719_),
    .B(_2154_),
    .Y(_3721_));
 sky130_fd_sc_hd__a32o_1 _7660_ (.A1(_3681_),
    .A2(_3720_),
    .A3(_3721_),
    .B1(_2184_),
    .B2(\sound4.sdiv.A[16] ),
    .X(_0421_));
 sky130_fd_sc_hd__and2b_1 _7661_ (.A_N(_2053_),
    .B(_3720_),
    .X(_3722_));
 sky130_fd_sc_hd__xor2_1 _7662_ (.A(_3722_),
    .B(_2156_),
    .X(_3723_));
 sky130_fd_sc_hd__a22o_1 _7663_ (.A1(\sound4.sdiv.A[17] ),
    .A2(_2183_),
    .B1(\sound4.sdiv.next_dived ),
    .B2(_3723_),
    .X(_0422_));
 sky130_fd_sc_hd__xnor2_1 _7664_ (.A(_2158_),
    .B(_2164_),
    .Y(_3724_));
 sky130_fd_sc_hd__a22o_1 _7665_ (.A1(\sound4.sdiv.A[18] ),
    .A2(_2183_),
    .B1(_3681_),
    .B2(_3724_),
    .X(_0423_));
 sky130_fd_sc_hd__a21o_1 _7666_ (.A1(_2158_),
    .A2(_2163_),
    .B1(_2162_),
    .X(_3725_));
 sky130_fd_sc_hd__xnor2_1 _7667_ (.A(_3725_),
    .B(_2165_),
    .Y(_3726_));
 sky130_fd_sc_hd__a22o_1 _7668_ (.A1(\sound4.sdiv.A[19] ),
    .A2(_2183_),
    .B1(_3681_),
    .B2(_3726_),
    .X(_0424_));
 sky130_fd_sc_hd__and2b_1 _7669_ (.A_N(_2168_),
    .B(_2041_),
    .X(_3727_));
 sky130_fd_sc_hd__and2b_1 _7670_ (.A_N(_2041_),
    .B(_2168_),
    .X(_3728_));
 sky130_fd_sc_hd__nor2_1 _7671_ (.A(_3727_),
    .B(_3728_),
    .Y(_3729_));
 sky130_fd_sc_hd__a22o_1 _7672_ (.A1(\sound4.sdiv.A[20] ),
    .A2(_2183_),
    .B1(_3681_),
    .B2(_3729_),
    .X(_0425_));
 sky130_fd_sc_hd__a21oi_1 _7673_ (.A1(\sound4.sdiv.A[19] ),
    .A2(_2038_),
    .B1(_3728_),
    .Y(_3730_));
 sky130_fd_sc_hd__xor2_1 _7674_ (.A(_2040_),
    .B(_3730_),
    .X(_3731_));
 sky130_fd_sc_hd__a22o_1 _7675_ (.A1(\sound4.sdiv.A[21] ),
    .A2(_2184_),
    .B1(_3681_),
    .B2(_3731_),
    .X(_0426_));
 sky130_fd_sc_hd__or2b_1 _7676_ (.A(_2042_),
    .B_N(_2168_),
    .X(_3732_));
 sky130_fd_sc_hd__a21oi_1 _7677_ (.A1(_2171_),
    .A2(_3732_),
    .B1(_2045_),
    .Y(_3733_));
 sky130_fd_sc_hd__a31o_1 _7678_ (.A1(_2045_),
    .A2(_2171_),
    .A3(_3732_),
    .B1(_1763_),
    .X(_3734_));
 sky130_fd_sc_hd__a2bb2o_1 _7679_ (.A1_N(_3733_),
    .A2_N(_3734_),
    .B1(\sound4.sdiv.A[22] ),
    .B2(_2183_),
    .X(_0427_));
 sky130_fd_sc_hd__a21oi_1 _7680_ (.A1(\sound4.sdiv.A[21] ),
    .A2(_2038_),
    .B1(_3733_),
    .Y(_3735_));
 sky130_fd_sc_hd__xnor2_1 _7681_ (.A(_2043_),
    .B(_3735_),
    .Y(_3736_));
 sky130_fd_sc_hd__a22o_1 _7682_ (.A1(\sound4.sdiv.A[23] ),
    .A2(_2184_),
    .B1(_3681_),
    .B2(_3736_),
    .X(_0428_));
 sky130_fd_sc_hd__o2111a_1 _7683_ (.A1(_2173_),
    .A2(_2172_),
    .B1(_2169_),
    .C1(_2170_),
    .D1(_2171_),
    .X(_3737_));
 sky130_fd_sc_hd__nand2_1 _7684_ (.A(\sound4.sdiv.A[24] ),
    .B(_2182_),
    .Y(_3738_));
 sky130_fd_sc_hd__o31ai_1 _7685_ (.A1(_1763_),
    .A2(_2174_),
    .A3(_3737_),
    .B1(_3738_),
    .Y(_0429_));
 sky130_fd_sc_hd__xor2_1 _7686_ (.A(\sound4.sdiv.A[24] ),
    .B(_2038_),
    .X(_3739_));
 sky130_fd_sc_hd__or3_1 _7687_ (.A(_2173_),
    .B(_2174_),
    .C(_3739_),
    .X(_3740_));
 sky130_fd_sc_hd__o21ai_1 _7688_ (.A1(_2173_),
    .A2(_2174_),
    .B1(_3739_),
    .Y(_3741_));
 sky130_fd_sc_hd__a32o_1 _7689_ (.A1(_3681_),
    .A2(_3740_),
    .A3(_3741_),
    .B1(_2184_),
    .B2(\sound4.sdiv.A[25] ),
    .X(_0430_));
 sky130_fd_sc_hd__nand3_1 _7690_ (.A(_2178_),
    .B(_2175_),
    .C(_2176_),
    .Y(_3742_));
 sky130_fd_sc_hd__a32o_1 _7691_ (.A1(_3681_),
    .A2(_2179_),
    .A3(_3742_),
    .B1(_2184_),
    .B2(\sound4.sdiv.A[26] ),
    .X(_0431_));
 sky130_fd_sc_hd__mux2_1 _7692_ (.A0(_1764_),
    .A1(_2182_),
    .S(\sound4.sdiv.C[0] ),
    .X(_3743_));
 sky130_fd_sc_hd__clkbuf_1 _7693_ (.A(_3743_),
    .X(_0432_));
 sky130_fd_sc_hd__nand2_1 _7694_ (.A(\sound4.sdiv.C[1] ),
    .B(\sound4.sdiv.C[0] ),
    .Y(_3744_));
 sky130_fd_sc_hd__or2_1 _7695_ (.A(\sound4.sdiv.C[1] ),
    .B(\sound4.sdiv.C[0] ),
    .X(_3745_));
 sky130_fd_sc_hd__a32o_1 _7696_ (.A1(_3681_),
    .A2(_3744_),
    .A3(_3745_),
    .B1(_2184_),
    .B2(\sound4.sdiv.C[1] ),
    .X(_0433_));
 sky130_fd_sc_hd__a21o_1 _7697_ (.A1(\sound4.sdiv.C[1] ),
    .A2(\sound4.sdiv.C[0] ),
    .B1(\sound4.sdiv.C[2] ),
    .X(_3746_));
 sky130_fd_sc_hd__and3_1 _7698_ (.A(\sound4.sdiv.C[2] ),
    .B(\sound4.sdiv.C[1] ),
    .C(\sound4.sdiv.C[0] ),
    .X(_3747_));
 sky130_fd_sc_hd__inv_2 _7699_ (.A(_3747_),
    .Y(_3748_));
 sky130_fd_sc_hd__a32o_1 _7700_ (.A1(_3681_),
    .A2(_3746_),
    .A3(_3748_),
    .B1(_2184_),
    .B2(\sound4.sdiv.C[2] ),
    .X(_0434_));
 sky130_fd_sc_hd__and3_1 _7701_ (.A(\sound4.sdiv.C[3] ),
    .B(_0556_),
    .C(_3747_),
    .X(_3749_));
 sky130_fd_sc_hd__a21oi_1 _7702_ (.A1(_0556_),
    .A2(_3747_),
    .B1(\sound4.sdiv.C[3] ),
    .Y(_3750_));
 sky130_fd_sc_hd__nor3_1 _7703_ (.A(_2005_),
    .B(_3749_),
    .C(_3750_),
    .Y(_0435_));
 sky130_fd_sc_hd__a31o_1 _7704_ (.A1(\sound4.sdiv.C[3] ),
    .A2(_0556_),
    .A3(_3747_),
    .B1(\sound4.sdiv.C[4] ),
    .X(_3751_));
 sky130_fd_sc_hd__and2_1 _7705_ (.A(_2843_),
    .B(_3751_),
    .X(_3752_));
 sky130_fd_sc_hd__clkbuf_1 _7706_ (.A(_3752_),
    .X(_0436_));
 sky130_fd_sc_hd__and2_1 _7707_ (.A(\sound4.sdiv.C[5] ),
    .B(_0554_),
    .X(_3753_));
 sky130_fd_sc_hd__clkbuf_1 _7708_ (.A(_3753_),
    .X(_0437_));
 sky130_fd_sc_hd__mux2_1 _7709_ (.A0(\wave_comb.u1.M[0] ),
    .A1(net32),
    .S(_0645_),
    .X(_3754_));
 sky130_fd_sc_hd__clkbuf_1 _7710_ (.A(_3754_),
    .X(_0438_));
 sky130_fd_sc_hd__mux2_1 _7711_ (.A0(\wave_comb.u1.M[1] ),
    .A1(net33),
    .S(_0645_),
    .X(_3755_));
 sky130_fd_sc_hd__clkbuf_1 _7712_ (.A(_3755_),
    .X(_0439_));
 sky130_fd_sc_hd__mux2_1 _7713_ (.A0(\wave_comb.u1.M[2] ),
    .A1(net34),
    .S(_0645_),
    .X(_3756_));
 sky130_fd_sc_hd__clkbuf_1 _7714_ (.A(_3756_),
    .X(_0440_));
 sky130_fd_sc_hd__dfrtp_1 _7715_ (.CLK(net137),
    .D(_0000_),
    .RESET_B(net98),
    .Q(\sound4.sdiv.Q[0] ));
 sky130_fd_sc_hd__dfrtp_2 _7716_ (.CLK(net137),
    .D(_0001_),
    .RESET_B(net98),
    .Q(\sound4.sdiv.Q[1] ));
 sky130_fd_sc_hd__dfrtp_2 _7717_ (.CLK(net137),
    .D(_0002_),
    .RESET_B(net98),
    .Q(\sound4.sdiv.Q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7718_ (.CLK(net137),
    .D(_0003_),
    .RESET_B(net98),
    .Q(\sound4.sdiv.Q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7719_ (.CLK(net137),
    .D(_0004_),
    .RESET_B(net98),
    .Q(\sound4.sdiv.Q[4] ));
 sky130_fd_sc_hd__dfrtp_2 _7720_ (.CLK(net137),
    .D(_0005_),
    .RESET_B(net98),
    .Q(\sound4.sdiv.Q[5] ));
 sky130_fd_sc_hd__dfrtp_2 _7721_ (.CLK(net136),
    .D(_0006_),
    .RESET_B(net97),
    .Q(\sound4.sdiv.Q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _7722_ (.CLK(net137),
    .D(_0007_),
    .RESET_B(net98),
    .Q(\sound4.sdiv.Q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _7723_ (.CLK(net136),
    .D(_0008_),
    .RESET_B(net97),
    .Q(\sound4.sdiv.Q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _7724_ (.CLK(net120),
    .D(_0009_),
    .RESET_B(net81),
    .Q(\sound4.sdiv.Q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _7725_ (.CLK(net121),
    .D(_0010_),
    .RESET_B(net82),
    .Q(\sound4.sdiv.Q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _7726_ (.CLK(net121),
    .D(_0011_),
    .RESET_B(net82),
    .Q(\sound4.sdiv.Q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _7727_ (.CLK(net121),
    .D(_0012_),
    .RESET_B(net82),
    .Q(\sound4.sdiv.Q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _7728_ (.CLK(net120),
    .D(_0013_),
    .RESET_B(net81),
    .Q(\sound4.sdiv.Q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _7729_ (.CLK(net120),
    .D(_0014_),
    .RESET_B(net81),
    .Q(\sound4.sdiv.Q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _7730_ (.CLK(net120),
    .D(_0015_),
    .RESET_B(net81),
    .Q(\sound4.sdiv.Q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _7731_ (.CLK(net120),
    .D(_0016_),
    .RESET_B(net81),
    .Q(\sound4.sdiv.Q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _7732_ (.CLK(net120),
    .D(_0017_),
    .RESET_B(net81),
    .Q(\sound4.sdiv.Q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _7733_ (.CLK(net117),
    .D(_0018_),
    .RESET_B(net78),
    .Q(\sound4.sdiv.Q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _7734_ (.CLK(net118),
    .D(_0019_),
    .RESET_B(net79),
    .Q(\sound4.sdiv.Q[19] ));
 sky130_fd_sc_hd__dfrtp_1 _7735_ (.CLK(net122),
    .D(_0020_),
    .RESET_B(net83),
    .Q(\sound4.sdiv.Q[20] ));
 sky130_fd_sc_hd__dfrtp_1 _7736_ (.CLK(net122),
    .D(_0021_),
    .RESET_B(net83),
    .Q(\sound4.sdiv.Q[21] ));
 sky130_fd_sc_hd__dfrtp_1 _7737_ (.CLK(net122),
    .D(_0022_),
    .RESET_B(net83),
    .Q(\sound4.sdiv.Q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _7738_ (.CLK(net122),
    .D(_0023_),
    .RESET_B(net83),
    .Q(\sound4.sdiv.Q[23] ));
 sky130_fd_sc_hd__dfrtp_1 _7739_ (.CLK(net137),
    .D(_0024_),
    .RESET_B(net98),
    .Q(\sound4.sdiv.Q[24] ));
 sky130_fd_sc_hd__dfrtp_1 _7740_ (.CLK(net137),
    .D(_0025_),
    .RESET_B(net98),
    .Q(\sound4.sdiv.Q[25] ));
 sky130_fd_sc_hd__dfrtp_1 _7741_ (.CLK(net137),
    .D(_0026_),
    .RESET_B(net98),
    .Q(\sound4.sdiv.Q[26] ));
 sky130_fd_sc_hd__dfrtp_1 _7742_ (.CLK(net137),
    .D(_0027_),
    .RESET_B(net98),
    .Q(\sound4.sdiv.Q[27] ));
 sky130_fd_sc_hd__dfrtp_1 _7743_ (.CLK(net137),
    .D(_0028_),
    .RESET_B(net98),
    .Q(\wave_comb.u1.A[0] ));
 sky130_fd_sc_hd__dfrtp_1 _7744_ (.CLK(net137),
    .D(_0029_),
    .RESET_B(net98),
    .Q(\wave_comb.u1.A[1] ));
 sky130_fd_sc_hd__dfrtp_1 _7745_ (.CLK(net139),
    .D(_0030_),
    .RESET_B(net100),
    .Q(\wave_comb.u1.A[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7746_ (.CLK(net139),
    .D(_0031_),
    .RESET_B(net100),
    .Q(\wave_comb.u1.A[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7747_ (.CLK(net139),
    .D(_0032_),
    .RESET_B(net100),
    .Q(\wave_comb.u1.A[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7748_ (.CLK(net139),
    .D(_0033_),
    .RESET_B(net100),
    .Q(\wave_comb.u1.A[5] ));
 sky130_fd_sc_hd__dfrtp_1 _7749_ (.CLK(net143),
    .D(_0034_),
    .RESET_B(net104),
    .Q(\wave_comb.u1.A[6] ));
 sky130_fd_sc_hd__dfrtp_1 _7750_ (.CLK(net139),
    .D(_0035_),
    .RESET_B(net100),
    .Q(\wave_comb.u1.A[7] ));
 sky130_fd_sc_hd__dfrtp_1 _7751_ (.CLK(net139),
    .D(_0036_),
    .RESET_B(net100),
    .Q(\wave_comb.u1.A[8] ));
 sky130_fd_sc_hd__dfrtp_1 _7752_ (.CLK(net139),
    .D(_0037_),
    .RESET_B(net100),
    .Q(\wave_comb.u1.A[9] ));
 sky130_fd_sc_hd__dfrtp_1 _7753_ (.CLK(net139),
    .D(_0038_),
    .RESET_B(net100),
    .Q(\wave_comb.u1.A[10] ));
 sky130_fd_sc_hd__dfrtp_1 _7754_ (.CLK(net143),
    .D(_0039_),
    .RESET_B(net104),
    .Q(\wave_comb.u1.C[0] ));
 sky130_fd_sc_hd__dfrtp_1 _7755_ (.CLK(net143),
    .D(_0040_),
    .RESET_B(net104),
    .Q(\wave_comb.u1.C[1] ));
 sky130_fd_sc_hd__dfrtp_1 _7756_ (.CLK(net143),
    .D(_0041_),
    .RESET_B(net104),
    .Q(\wave_comb.u1.C[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7757_ (.CLK(net143),
    .D(_0042_),
    .RESET_B(net104),
    .Q(\wave_comb.u1.C[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7758_ (.CLK(net139),
    .D(_0043_),
    .RESET_B(net100),
    .Q(\wave_comb.u1.C[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7759_ (.CLK(net143),
    .D(_0044_),
    .RESET_B(net104),
    .Q(\wave_comb.u1.C[5] ));
 sky130_fd_sc_hd__dfrtp_1 _7760_ (.CLK(net143),
    .D(\wave_comb.u1.next_start ),
    .RESET_B(net104),
    .Q(\wave_comb.u1.start ));
 sky130_fd_sc_hd__dfrtp_1 _7761_ (.CLK(net144),
    .D(\pm.next_count[0] ),
    .RESET_B(net105),
    .Q(\pm.count[0] ));
 sky130_fd_sc_hd__dfrtp_2 _7762_ (.CLK(net144),
    .D(\pm.next_count[1] ),
    .RESET_B(net105),
    .Q(\pm.count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _7763_ (.CLK(net144),
    .D(\pm.next_count[2] ),
    .RESET_B(net105),
    .Q(\pm.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7764_ (.CLK(net144),
    .D(\pm.next_count[3] ),
    .RESET_B(net105),
    .Q(\pm.count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7765_ (.CLK(net144),
    .D(\pm.next_count[4] ),
    .RESET_B(net105),
    .Q(\pm.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7766_ (.CLK(net144),
    .D(\pm.next_count[5] ),
    .RESET_B(net105),
    .Q(\pm.count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _7767_ (.CLK(net144),
    .D(\pm.next_count[6] ),
    .RESET_B(net105),
    .Q(\pm.count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _7768_ (.CLK(net144),
    .D(\pm.next_count[7] ),
    .RESET_B(net105),
    .Q(\pm.count[7] ));
 sky130_fd_sc_hd__dfrtp_1 _7769_ (.CLK(net144),
    .D(\pm.next_count[8] ),
    .RESET_B(net105),
    .Q(\pm.count[8] ));
 sky130_fd_sc_hd__dfrtp_1 _7770_ (.CLK(net133),
    .D(\pm.next_pwm_o ),
    .RESET_B(net94),
    .Q(\pm.pwm_o ));
 sky130_fd_sc_hd__dfrtp_1 _7771_ (.CLK(net139),
    .D(_0045_),
    .RESET_B(net100),
    .Q(\wave_comb.u1.Q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _7772_ (.CLK(net139),
    .D(_0046_),
    .RESET_B(net100),
    .Q(\wave_comb.u1.Q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _7773_ (.CLK(net143),
    .D(_0047_),
    .RESET_B(net104),
    .Q(\wave_comb.u1.Q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7774_ (.CLK(net139),
    .D(_0048_),
    .RESET_B(net100),
    .Q(\wave_comb.u1.Q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7775_ (.CLK(net139),
    .D(_0049_),
    .RESET_B(net100),
    .Q(\wave_comb.u1.Q[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7776_ (.CLK(net139),
    .D(_0050_),
    .RESET_B(net100),
    .Q(\wave_comb.u1.Q[5] ));
 sky130_fd_sc_hd__dfrtp_1 _7777_ (.CLK(net139),
    .D(_0051_),
    .RESET_B(net100),
    .Q(\wave_comb.u1.Q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _7778_ (.CLK(net139),
    .D(_0052_),
    .RESET_B(net100),
    .Q(\wave_comb.u1.Q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _7779_ (.CLK(net139),
    .D(_0053_),
    .RESET_B(net100),
    .Q(\wave_comb.u1.Q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _7780_ (.CLK(net139),
    .D(_0054_),
    .RESET_B(net100),
    .Q(\wave_comb.u1.Q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _7781_ (.CLK(net137),
    .D(_0055_),
    .RESET_B(net98),
    .Q(\wave_comb.u1.Q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _7782_ (.CLK(net137),
    .D(_0056_),
    .RESET_B(net98),
    .Q(\wave_comb.u1.Q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _7783_ (.CLK(net142),
    .D(\inputcont.INTERNAL_MODE ),
    .RESET_B(net103),
    .Q(\inputcont.u3.next_in ));
 sky130_fd_sc_hd__dfrtp_1 _7784_ (.CLK(net118),
    .D(\inputcont.INTERNAL_OCTAVE_INPUT ),
    .RESET_B(net79),
    .Q(\inputcont.u2.next_in ));
 sky130_fd_sc_hd__dfrtp_1 _7785_ (.CLK(net142),
    .D(\inputcont.u1.ff_intermediate[14] ),
    .RESET_B(net103),
    .Q(\inputcont.INTERNAL_MODE ));
 sky130_fd_sc_hd__dfrtp_4 _7786_ (.CLK(net113),
    .D(\inputcont.u1.ff_intermediate[8] ),
    .RESET_B(net74),
    .Q(\inputcont.INTERNAL_SYNCED_I[8] ));
 sky130_fd_sc_hd__dfrtp_4 _7787_ (.CLK(net113),
    .D(\inputcont.u1.ff_intermediate[9] ),
    .RESET_B(net74),
    .Q(\inputcont.INTERNAL_SYNCED_I[9] ));
 sky130_fd_sc_hd__dfrtp_4 _7788_ (.CLK(net128),
    .D(\inputcont.u1.ff_intermediate[10] ),
    .RESET_B(net89),
    .Q(\inputcont.INTERNAL_SYNCED_I[10] ));
 sky130_fd_sc_hd__dfrtp_2 _7789_ (.CLK(net107),
    .D(\inputcont.u1.ff_intermediate[11] ),
    .RESET_B(net68),
    .Q(\inputcont.INTERNAL_SYNCED_I[11] ));
 sky130_fd_sc_hd__dfrtp_4 _7790_ (.CLK(net122),
    .D(\inputcont.u1.ff_intermediate[12] ),
    .RESET_B(net83),
    .Q(\inputcont.INTERNAL_SYNCED_I[12] ));
 sky130_fd_sc_hd__dfrtp_1 _7791_ (.CLK(net118),
    .D(\inputcont.u1.ff_intermediate[13] ),
    .RESET_B(net79),
    .Q(\inputcont.INTERNAL_OCTAVE_INPUT ));
 sky130_fd_sc_hd__dfrtp_4 _7792_ (.CLK(net144),
    .D(net17),
    .RESET_B(net105),
    .Q(\inputcont.u1.ff_intermediate[8] ));
 sky130_fd_sc_hd__dfrtp_2 _7793_ (.CLK(net130),
    .D(net18),
    .RESET_B(net91),
    .Q(\inputcont.u1.ff_intermediate[9] ));
 sky130_fd_sc_hd__dfrtp_2 _7794_ (.CLK(net139),
    .D(net5),
    .RESET_B(net100),
    .Q(\inputcont.u1.ff_intermediate[10] ));
 sky130_fd_sc_hd__dfrtp_1 _7795_ (.CLK(net110),
    .D(net6),
    .RESET_B(net71),
    .Q(\inputcont.u1.ff_intermediate[11] ));
 sky130_fd_sc_hd__dfrtp_1 _7796_ (.CLK(net138),
    .D(net7),
    .RESET_B(net99),
    .Q(\inputcont.u1.ff_intermediate[12] ));
 sky130_fd_sc_hd__dfrtp_1 _7797_ (.CLK(net118),
    .D(net8),
    .RESET_B(net79),
    .Q(\inputcont.u1.ff_intermediate[13] ));
 sky130_fd_sc_hd__dfrtp_1 _7798_ (.CLK(net142),
    .D(net9),
    .RESET_B(net103),
    .Q(\inputcont.u1.ff_intermediate[14] ));
 sky130_fd_sc_hd__dfstp_4 _7799_ (.CLK(net113),
    .D(\oct.next_state[0] ),
    .SET_B(net74),
    .Q(\oct.state[0] ));
 sky130_fd_sc_hd__dfstp_1 _7800_ (.CLK(net113),
    .D(\oct.next_state[1] ),
    .SET_B(net74),
    .Q(\oct.state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _7801_ (.CLK(net113),
    .D(\oct.next_state[2] ),
    .RESET_B(net74),
    .Q(\oct.state[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7802_ (.CLK(net107),
    .D(\seq.player_8.next_state[0] ),
    .RESET_B(net68),
    .Q(\seq.player_8.state[0] ));
 sky130_fd_sc_hd__dfrtp_1 _7803_ (.CLK(net107),
    .D(\seq.player_8.next_state[1] ),
    .RESET_B(net68),
    .Q(\seq.player_8.state[1] ));
 sky130_fd_sc_hd__dfrtp_4 _7804_ (.CLK(net107),
    .D(\seq.player_8.next_state[2] ),
    .RESET_B(net68),
    .Q(\seq.player_8.state[2] ));
 sky130_fd_sc_hd__dfrtp_2 _7805_ (.CLK(net107),
    .D(\seq.player_8.next_state[3] ),
    .RESET_B(net68),
    .Q(\seq.player_8.state[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7806_ (.CLK(net107),
    .D(\seq.player_7.next_state[0] ),
    .RESET_B(net68),
    .Q(\seq.player_7.state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _7807_ (.CLK(net107),
    .D(\seq.player_7.next_state[1] ),
    .RESET_B(net68),
    .Q(\seq.player_7.state[1] ));
 sky130_fd_sc_hd__dfrtp_4 _7808_ (.CLK(net108),
    .D(\seq.player_7.next_state[2] ),
    .RESET_B(net69),
    .Q(\seq.player_7.state[2] ));
 sky130_fd_sc_hd__dfrtp_2 _7809_ (.CLK(net107),
    .D(\seq.player_7.next_state[3] ),
    .RESET_B(net68),
    .Q(\seq.player_7.state[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7810_ (.CLK(net107),
    .D(\seq.player_6.next_state[0] ),
    .RESET_B(net68),
    .Q(\seq.player_6.state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _7811_ (.CLK(net107),
    .D(\seq.player_6.next_state[1] ),
    .RESET_B(net68),
    .Q(\seq.player_6.state[1] ));
 sky130_fd_sc_hd__dfrtp_4 _7812_ (.CLK(net107),
    .D(\seq.player_6.next_state[2] ),
    .RESET_B(net68),
    .Q(\seq.player_6.state[2] ));
 sky130_fd_sc_hd__dfrtp_2 _7813_ (.CLK(net107),
    .D(\seq.player_6.next_state[3] ),
    .RESET_B(net68),
    .Q(\seq.player_6.state[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7814_ (.CLK(net114),
    .D(\seq.player_5.next_state[0] ),
    .RESET_B(net75),
    .Q(\seq.player_5.state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _7815_ (.CLK(net114),
    .D(\seq.player_5.next_state[1] ),
    .RESET_B(net75),
    .Q(\seq.player_5.state[1] ));
 sky130_fd_sc_hd__dfrtp_4 _7816_ (.CLK(net114),
    .D(\seq.player_5.next_state[2] ),
    .RESET_B(net75),
    .Q(\seq.player_5.state[2] ));
 sky130_fd_sc_hd__dfrtp_2 _7817_ (.CLK(net114),
    .D(\seq.player_5.next_state[3] ),
    .RESET_B(net75),
    .Q(\seq.player_5.state[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7818_ (.CLK(net114),
    .D(\seq.player_4.next_state[0] ),
    .RESET_B(net75),
    .Q(\seq.player_4.state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _7819_ (.CLK(net114),
    .D(\seq.player_4.next_state[1] ),
    .RESET_B(net75),
    .Q(\seq.player_4.state[1] ));
 sky130_fd_sc_hd__dfrtp_4 _7820_ (.CLK(net114),
    .D(\seq.player_4.next_state[2] ),
    .RESET_B(net75),
    .Q(\seq.player_4.state[2] ));
 sky130_fd_sc_hd__dfrtp_2 _7821_ (.CLK(net114),
    .D(\seq.player_4.next_state[3] ),
    .RESET_B(net75),
    .Q(\seq.player_4.state[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7822_ (.CLK(net114),
    .D(\seq.player_3.next_state[0] ),
    .RESET_B(net75),
    .Q(\seq.player_3.state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _7823_ (.CLK(net114),
    .D(\seq.player_3.next_state[1] ),
    .RESET_B(net75),
    .Q(\seq.player_3.state[1] ));
 sky130_fd_sc_hd__dfrtp_4 _7824_ (.CLK(net113),
    .D(\seq.player_3.next_state[2] ),
    .RESET_B(net74),
    .Q(\seq.player_3.state[2] ));
 sky130_fd_sc_hd__dfrtp_2 _7825_ (.CLK(net113),
    .D(\seq.player_3.next_state[3] ),
    .RESET_B(net74),
    .Q(\seq.player_3.state[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7826_ (.CLK(net113),
    .D(\seq.player_2.next_state[0] ),
    .RESET_B(net74),
    .Q(\seq.player_2.state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _7827_ (.CLK(net113),
    .D(\seq.player_2.next_state[1] ),
    .RESET_B(net74),
    .Q(\seq.player_2.state[1] ));
 sky130_fd_sc_hd__dfrtp_4 _7828_ (.CLK(net113),
    .D(\seq.player_2.next_state[2] ),
    .RESET_B(net74),
    .Q(\seq.player_2.state[2] ));
 sky130_fd_sc_hd__dfrtp_2 _7829_ (.CLK(net113),
    .D(\seq.player_2.next_state[3] ),
    .RESET_B(net74),
    .Q(\seq.player_2.state[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7830_ (.CLK(net113),
    .D(\seq.player_1.next_state[0] ),
    .RESET_B(net74),
    .Q(\seq.player_1.state[0] ));
 sky130_fd_sc_hd__dfrtp_2 _7831_ (.CLK(net113),
    .D(\seq.player_1.next_state[1] ),
    .RESET_B(net74),
    .Q(\seq.player_1.state[1] ));
 sky130_fd_sc_hd__dfrtp_4 _7832_ (.CLK(net113),
    .D(\seq.player_1.next_state[2] ),
    .RESET_B(net74),
    .Q(\seq.player_1.state[2] ));
 sky130_fd_sc_hd__dfrtp_2 _7833_ (.CLK(net113),
    .D(\seq.player_1.next_state[3] ),
    .RESET_B(net74),
    .Q(\seq.player_1.state[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7834_ (.CLK(net144),
    .D(_0057_),
    .RESET_B(net105),
    .Q(\pm.current_waveform[0] ));
 sky130_fd_sc_hd__dfrtp_1 _7835_ (.CLK(net143),
    .D(_0058_),
    .RESET_B(net104),
    .Q(\pm.current_waveform[1] ));
 sky130_fd_sc_hd__dfrtp_1 _7836_ (.CLK(net143),
    .D(_0059_),
    .RESET_B(net104),
    .Q(\pm.current_waveform[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7837_ (.CLK(net143),
    .D(_0060_),
    .RESET_B(net104),
    .Q(\pm.current_waveform[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7838_ (.CLK(net143),
    .D(_0061_),
    .RESET_B(net104),
    .Q(\pm.current_waveform[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7839_ (.CLK(net143),
    .D(_0062_),
    .RESET_B(net104),
    .Q(\pm.current_waveform[5] ));
 sky130_fd_sc_hd__dfrtp_1 _7840_ (.CLK(net143),
    .D(_0063_),
    .RESET_B(net104),
    .Q(\pm.current_waveform[6] ));
 sky130_fd_sc_hd__dfrtp_1 _7841_ (.CLK(net143),
    .D(_0064_),
    .RESET_B(net104),
    .Q(\pm.current_waveform[7] ));
 sky130_fd_sc_hd__dfrtp_1 _7842_ (.CLK(net143),
    .D(_0065_),
    .RESET_B(net104),
    .Q(\pm.current_waveform[8] ));
 sky130_fd_sc_hd__dfrtp_1 _7843_ (.CLK(net107),
    .D(\seq.clk_div.next_count[0] ),
    .RESET_B(net68),
    .Q(\seq.clk_div.count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _7844_ (.CLK(net108),
    .D(\seq.clk_div.next_count[1] ),
    .RESET_B(net69),
    .Q(\seq.clk_div.count[1] ));
 sky130_fd_sc_hd__dfrtp_2 _7845_ (.CLK(net108),
    .D(\seq.clk_div.next_count[2] ),
    .RESET_B(net69),
    .Q(\seq.clk_div.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7846_ (.CLK(net108),
    .D(\seq.clk_div.next_count[3] ),
    .RESET_B(net69),
    .Q(\seq.clk_div.count[3] ));
 sky130_fd_sc_hd__dfrtp_2 _7847_ (.CLK(net108),
    .D(\seq.clk_div.next_count[4] ),
    .RESET_B(net69),
    .Q(\seq.clk_div.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7848_ (.CLK(net108),
    .D(\seq.clk_div.next_count[5] ),
    .RESET_B(net69),
    .Q(\seq.clk_div.count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _7849_ (.CLK(net108),
    .D(\seq.clk_div.next_count[6] ),
    .RESET_B(net69),
    .Q(\seq.clk_div.count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _7850_ (.CLK(net108),
    .D(\seq.clk_div.next_count[7] ),
    .RESET_B(net69),
    .Q(\seq.clk_div.count[7] ));
 sky130_fd_sc_hd__dfrtp_2 _7851_ (.CLK(net108),
    .D(\seq.clk_div.next_count[8] ),
    .RESET_B(net69),
    .Q(\seq.clk_div.count[8] ));
 sky130_fd_sc_hd__dfrtp_1 _7852_ (.CLK(net108),
    .D(\seq.clk_div.next_count[9] ),
    .RESET_B(net69),
    .Q(\seq.clk_div.count[9] ));
 sky130_fd_sc_hd__dfrtp_2 _7853_ (.CLK(net108),
    .D(\seq.clk_div.next_count[10] ),
    .RESET_B(net69),
    .Q(\seq.clk_div.count[10] ));
 sky130_fd_sc_hd__dfrtp_1 _7854_ (.CLK(net108),
    .D(\seq.clk_div.next_count[11] ),
    .RESET_B(net69),
    .Q(\seq.clk_div.count[11] ));
 sky130_fd_sc_hd__dfrtp_2 _7855_ (.CLK(net108),
    .D(\seq.clk_div.next_count[12] ),
    .RESET_B(net69),
    .Q(\seq.clk_div.count[12] ));
 sky130_fd_sc_hd__dfrtp_1 _7856_ (.CLK(net108),
    .D(\seq.clk_div.next_count[13] ),
    .RESET_B(net69),
    .Q(\seq.clk_div.count[13] ));
 sky130_fd_sc_hd__dfrtp_1 _7857_ (.CLK(net108),
    .D(\seq.clk_div.next_count[14] ),
    .RESET_B(net69),
    .Q(\seq.clk_div.count[14] ));
 sky130_fd_sc_hd__dfrtp_1 _7858_ (.CLK(net108),
    .D(\seq.clk_div.next_count[15] ),
    .RESET_B(net69),
    .Q(\seq.clk_div.count[15] ));
 sky130_fd_sc_hd__dfrtp_1 _7859_ (.CLK(net107),
    .D(\seq.clk_div.next_count[16] ),
    .RESET_B(net68),
    .Q(\seq.clk_div.count[16] ));
 sky130_fd_sc_hd__dfrtp_1 _7860_ (.CLK(net107),
    .D(\seq.clk_div.next_count[17] ),
    .RESET_B(net68),
    .Q(\seq.clk_div.count[17] ));
 sky130_fd_sc_hd__dfrtp_1 _7861_ (.CLK(net111),
    .D(\seq.clk_div.next_count[18] ),
    .RESET_B(net72),
    .Q(\seq.clk_div.count[18] ));
 sky130_fd_sc_hd__dfrtp_1 _7862_ (.CLK(net110),
    .D(\seq.clk_div.next_count[19] ),
    .RESET_B(net71),
    .Q(\seq.clk_div.count[19] ));
 sky130_fd_sc_hd__dfrtp_1 _7863_ (.CLK(net110),
    .D(\seq.clk_div.next_count[20] ),
    .RESET_B(net71),
    .Q(\seq.clk_div.count[20] ));
 sky130_fd_sc_hd__dfrtp_2 _7864_ (.CLK(net110),
    .D(\seq.clk_div.next_count[21] ),
    .RESET_B(net71),
    .Q(\seq.clk_div.count[21] ));
 sky130_fd_sc_hd__dfrtp_4 _7865_ (.CLK(net110),
    .D(\seq.tempo_select.next_state[0] ),
    .RESET_B(net71),
    .Q(\seq.tempo_select.state[0] ));
 sky130_fd_sc_hd__dfrtp_4 _7866_ (.CLK(net110),
    .D(\seq.tempo_select.next_state[1] ),
    .RESET_B(net71),
    .Q(\seq.tempo_select.state[1] ));
 sky130_fd_sc_hd__dfrtp_1 _7867_ (.CLK(net114),
    .D(\seq.encode.inter_keys[0] ),
    .RESET_B(net75),
    .Q(\seq.encode.keys_sync[0] ));
 sky130_fd_sc_hd__dfrtp_1 _7868_ (.CLK(net113),
    .D(\seq.encode.inter_keys[1] ),
    .RESET_B(net74),
    .Q(\seq.encode.keys_sync[1] ));
 sky130_fd_sc_hd__dfrtp_4 _7869_ (.CLK(net113),
    .D(\inputcont.u1.ff_intermediate[0] ),
    .RESET_B(net74),
    .Q(\inputcont.INTERNAL_SYNCED_I[0] ));
 sky130_fd_sc_hd__dfrtp_4 _7870_ (.CLK(net111),
    .D(\inputcont.u1.ff_intermediate[1] ),
    .RESET_B(net72),
    .Q(\inputcont.INTERNAL_SYNCED_I[1] ));
 sky130_fd_sc_hd__dfrtp_4 _7871_ (.CLK(net108),
    .D(\inputcont.u1.ff_intermediate[2] ),
    .RESET_B(net69),
    .Q(\inputcont.INTERNAL_SYNCED_I[2] ));
 sky130_fd_sc_hd__dfrtp_4 _7872_ (.CLK(net111),
    .D(\inputcont.u1.ff_intermediate[3] ),
    .RESET_B(net72),
    .Q(\inputcont.INTERNAL_SYNCED_I[3] ));
 sky130_fd_sc_hd__dfrtp_4 _7873_ (.CLK(net107),
    .D(\inputcont.u1.ff_intermediate[4] ),
    .RESET_B(net68),
    .Q(\inputcont.INTERNAL_SYNCED_I[4] ));
 sky130_fd_sc_hd__dfrtp_4 _7874_ (.CLK(net108),
    .D(\inputcont.u1.ff_intermediate[5] ),
    .RESET_B(net69),
    .Q(\inputcont.INTERNAL_SYNCED_I[5] ));
 sky130_fd_sc_hd__dfrtp_4 _7875_ (.CLK(net110),
    .D(\inputcont.u1.ff_intermediate[6] ),
    .RESET_B(net71),
    .Q(\inputcont.INTERNAL_SYNCED_I[6] ));
 sky130_fd_sc_hd__dfrtp_4 _7876_ (.CLK(net113),
    .D(\inputcont.u1.ff_intermediate[7] ),
    .RESET_B(net74),
    .Q(\inputcont.INTERNAL_SYNCED_I[7] ));
 sky130_fd_sc_hd__dfrtp_1 _7877_ (.CLK(net111),
    .D(\seq.encode.inter_keys[10] ),
    .RESET_B(net72),
    .Q(\seq.encode.keys_sync[10] ));
 sky130_fd_sc_hd__dfrtp_1 _7878_ (.CLK(net114),
    .D(seq_play_on),
    .RESET_B(net75),
    .Q(\seq.encode.inter_keys[0] ));
 sky130_fd_sc_hd__dfrtp_1 _7879_ (.CLK(net130),
    .D(seq_power_on),
    .RESET_B(net91),
    .Q(\seq.encode.inter_keys[1] ));
 sky130_fd_sc_hd__dfrtp_2 _7880_ (.CLK(net130),
    .D(net4),
    .RESET_B(net91),
    .Q(\inputcont.u1.ff_intermediate[0] ));
 sky130_fd_sc_hd__dfrtp_4 _7881_ (.CLK(net118),
    .D(net10),
    .RESET_B(net79),
    .Q(\inputcont.u1.ff_intermediate[1] ));
 sky130_fd_sc_hd__dfrtp_1 _7882_ (.CLK(net108),
    .D(net11),
    .RESET_B(net69),
    .Q(\inputcont.u1.ff_intermediate[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7883_ (.CLK(net110),
    .D(net12),
    .RESET_B(net71),
    .Q(\inputcont.u1.ff_intermediate[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7884_ (.CLK(net109),
    .D(net13),
    .RESET_B(net70),
    .Q(\inputcont.u1.ff_intermediate[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7885_ (.CLK(net108),
    .D(net14),
    .RESET_B(net69),
    .Q(\inputcont.u1.ff_intermediate[5] ));
 sky130_fd_sc_hd__dfrtp_1 _7886_ (.CLK(net110),
    .D(net15),
    .RESET_B(net71),
    .Q(\inputcont.u1.ff_intermediate[6] ));
 sky130_fd_sc_hd__dfrtp_4 _7887_ (.CLK(net144),
    .D(net16),
    .RESET_B(net105),
    .Q(\inputcont.u1.ff_intermediate[7] ));
 sky130_fd_sc_hd__dfrtp_1 _7888_ (.CLK(net111),
    .D(tempo_select_on),
    .RESET_B(net72),
    .Q(\seq.encode.inter_keys[10] ));
 sky130_fd_sc_hd__dfrtp_4 _7889_ (.CLK(net113),
    .D(\seq.encode.next_sequencer_on ),
    .RESET_B(net74),
    .Q(\select1.sequencer_on ));
 sky130_fd_sc_hd__dfrtp_4 _7890_ (.CLK(net114),
    .D(\seq.encode.next_play ),
    .RESET_B(net75),
    .Q(\seq.encode.play ));
 sky130_fd_sc_hd__dfrtp_1 _7891_ (.CLK(net114),
    .D(\seq.encode.keys_sync[0] ),
    .RESET_B(net75),
    .Q(\seq.encode.keys_edge_det[0] ));
 sky130_fd_sc_hd__dfrtp_1 _7892_ (.CLK(net113),
    .D(\seq.encode.keys_sync[1] ),
    .RESET_B(net74),
    .Q(\seq.encode.keys_edge_det[1] ));
 sky130_fd_sc_hd__dfrtp_1 _7893_ (.CLK(net114),
    .D(\inputcont.INTERNAL_SYNCED_I[0] ),
    .RESET_B(net75),
    .Q(\seq.encode.keys_edge_det[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7894_ (.CLK(net114),
    .D(\inputcont.INTERNAL_SYNCED_I[1] ),
    .RESET_B(net75),
    .Q(\seq.encode.keys_edge_det[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7895_ (.CLK(net114),
    .D(\inputcont.INTERNAL_SYNCED_I[2] ),
    .RESET_B(net75),
    .Q(\seq.encode.keys_edge_det[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7896_ (.CLK(net114),
    .D(\inputcont.INTERNAL_SYNCED_I[3] ),
    .RESET_B(net75),
    .Q(\seq.encode.keys_edge_det[5] ));
 sky130_fd_sc_hd__dfrtp_1 _7897_ (.CLK(net107),
    .D(\inputcont.INTERNAL_SYNCED_I[4] ),
    .RESET_B(net68),
    .Q(\seq.encode.keys_edge_det[6] ));
 sky130_fd_sc_hd__dfrtp_1 _7898_ (.CLK(net107),
    .D(\inputcont.INTERNAL_SYNCED_I[5] ),
    .RESET_B(net68),
    .Q(\seq.encode.keys_edge_det[7] ));
 sky130_fd_sc_hd__dfrtp_1 _7899_ (.CLK(net107),
    .D(\inputcont.INTERNAL_SYNCED_I[6] ),
    .RESET_B(net68),
    .Q(\seq.encode.keys_edge_det[8] ));
 sky130_fd_sc_hd__dfrtp_1 _7900_ (.CLK(net107),
    .D(\inputcont.INTERNAL_SYNCED_I[7] ),
    .RESET_B(net68),
    .Q(\seq.encode.keys_edge_det[9] ));
 sky130_fd_sc_hd__dfrtp_1 _7901_ (.CLK(net111),
    .D(\seq.encode.keys_sync[10] ),
    .RESET_B(net72),
    .Q(\seq.encode.keys_edge_det[10] ));
 sky130_fd_sc_hd__dfrtp_1 _7902_ (.CLK(net140),
    .D(\sound1.sdiv.next_dived ),
    .RESET_B(net101),
    .Q(\sound1.sdiv.dived ));
 sky130_fd_sc_hd__dfrtp_4 _7903_ (.CLK(net115),
    .D(_0066_),
    .RESET_B(net76),
    .Q(\seq.beat[0] ));
 sky130_fd_sc_hd__dfrtp_4 _7904_ (.CLK(net115),
    .D(_0067_),
    .RESET_B(net76),
    .Q(\seq.beat[1] ));
 sky130_fd_sc_hd__dfrtp_4 _7905_ (.CLK(net115),
    .D(_0068_),
    .RESET_B(net76),
    .Q(\seq.beat[2] ));
 sky130_fd_sc_hd__dfrtp_4 _7906_ (.CLK(net115),
    .D(_0069_),
    .RESET_B(net76),
    .Q(\seq.beat[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7907_ (.CLK(net128),
    .D(_0070_),
    .RESET_B(net89),
    .Q(\sound1.count_m[0] ));
 sky130_fd_sc_hd__dfrtp_1 _7908_ (.CLK(net128),
    .D(_0071_),
    .RESET_B(net89),
    .Q(\sound1.count_m[1] ));
 sky130_fd_sc_hd__dfrtp_1 _7909_ (.CLK(net128),
    .D(_0072_),
    .RESET_B(net89),
    .Q(\sound1.count_m[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7910_ (.CLK(net128),
    .D(_0073_),
    .RESET_B(net89),
    .Q(\sound1.count_m[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7911_ (.CLK(net126),
    .D(_0074_),
    .RESET_B(net87),
    .Q(\sound1.count_m[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7912_ (.CLK(net127),
    .D(_0075_),
    .RESET_B(net88),
    .Q(\sound1.count_m[5] ));
 sky130_fd_sc_hd__dfrtp_1 _7913_ (.CLK(net127),
    .D(_0076_),
    .RESET_B(net88),
    .Q(\sound1.count_m[6] ));
 sky130_fd_sc_hd__dfrtp_1 _7914_ (.CLK(net127),
    .D(_0077_),
    .RESET_B(net88),
    .Q(\sound1.count_m[7] ));
 sky130_fd_sc_hd__dfrtp_1 _7915_ (.CLK(net126),
    .D(_0078_),
    .RESET_B(net87),
    .Q(\sound1.count_m[8] ));
 sky130_fd_sc_hd__dfrtp_1 _7916_ (.CLK(net126),
    .D(_0079_),
    .RESET_B(net87),
    .Q(\sound1.count_m[9] ));
 sky130_fd_sc_hd__dfrtp_1 _7917_ (.CLK(net126),
    .D(_0080_),
    .RESET_B(net87),
    .Q(\sound1.count_m[10] ));
 sky130_fd_sc_hd__dfrtp_1 _7918_ (.CLK(net126),
    .D(_0081_),
    .RESET_B(net87),
    .Q(\sound1.count_m[11] ));
 sky130_fd_sc_hd__dfrtp_1 _7919_ (.CLK(net126),
    .D(_0082_),
    .RESET_B(net87),
    .Q(\sound1.count_m[12] ));
 sky130_fd_sc_hd__dfrtp_1 _7920_ (.CLK(net126),
    .D(_0083_),
    .RESET_B(net87),
    .Q(\sound1.count_m[13] ));
 sky130_fd_sc_hd__dfrtp_1 _7921_ (.CLK(net126),
    .D(_0084_),
    .RESET_B(net87),
    .Q(\sound1.count_m[14] ));
 sky130_fd_sc_hd__dfrtp_1 _7922_ (.CLK(net126),
    .D(_0085_),
    .RESET_B(net87),
    .Q(\sound1.count_m[15] ));
 sky130_fd_sc_hd__dfrtp_1 _7923_ (.CLK(net127),
    .D(_0086_),
    .RESET_B(net88),
    .Q(\sound1.count_m[16] ));
 sky130_fd_sc_hd__dfrtp_1 _7924_ (.CLK(net127),
    .D(_0087_),
    .RESET_B(net88),
    .Q(\sound1.count_m[17] ));
 sky130_fd_sc_hd__dfrtp_1 _7925_ (.CLK(net127),
    .D(_0088_),
    .RESET_B(net88),
    .Q(\sound1.count_m[18] ));
 sky130_fd_sc_hd__dfrtp_4 _7926_ (.CLK(net128),
    .D(_0089_),
    .RESET_B(net89),
    .Q(\sound1.divisor_m[0] ));
 sky130_fd_sc_hd__dfrtp_4 _7927_ (.CLK(net129),
    .D(_0090_),
    .RESET_B(net90),
    .Q(\sound1.divisor_m[1] ));
 sky130_fd_sc_hd__dfrtp_2 _7928_ (.CLK(net128),
    .D(_0091_),
    .RESET_B(net89),
    .Q(\sound1.divisor_m[2] ));
 sky130_fd_sc_hd__dfrtp_4 _7929_ (.CLK(net129),
    .D(_0092_),
    .RESET_B(net90),
    .Q(\sound1.divisor_m[3] ));
 sky130_fd_sc_hd__dfrtp_2 _7930_ (.CLK(net128),
    .D(_0093_),
    .RESET_B(net89),
    .Q(\sound1.divisor_m[4] ));
 sky130_fd_sc_hd__dfrtp_2 _7931_ (.CLK(net127),
    .D(_0094_),
    .RESET_B(net88),
    .Q(\sound1.divisor_m[5] ));
 sky130_fd_sc_hd__dfrtp_2 _7932_ (.CLK(net127),
    .D(_0095_),
    .RESET_B(net88),
    .Q(\sound1.divisor_m[6] ));
 sky130_fd_sc_hd__dfrtp_2 _7933_ (.CLK(net127),
    .D(_0096_),
    .RESET_B(net88),
    .Q(\sound1.divisor_m[7] ));
 sky130_fd_sc_hd__dfrtp_2 _7934_ (.CLK(net127),
    .D(_0097_),
    .RESET_B(net88),
    .Q(\sound1.divisor_m[8] ));
 sky130_fd_sc_hd__dfrtp_4 _7935_ (.CLK(net125),
    .D(_0098_),
    .RESET_B(net86),
    .Q(\sound1.divisor_m[9] ));
 sky130_fd_sc_hd__dfrtp_1 _7936_ (.CLK(net127),
    .D(_0099_),
    .RESET_B(net88),
    .Q(\sound1.divisor_m[10] ));
 sky130_fd_sc_hd__dfrtp_2 _7937_ (.CLK(net126),
    .D(_0100_),
    .RESET_B(net87),
    .Q(\sound1.divisor_m[11] ));
 sky130_fd_sc_hd__dfrtp_2 _7938_ (.CLK(net127),
    .D(_0101_),
    .RESET_B(net88),
    .Q(\sound1.divisor_m[12] ));
 sky130_fd_sc_hd__dfrtp_2 _7939_ (.CLK(net125),
    .D(_0102_),
    .RESET_B(net86),
    .Q(\sound1.divisor_m[13] ));
 sky130_fd_sc_hd__dfrtp_1 _7940_ (.CLK(net126),
    .D(_0103_),
    .RESET_B(net87),
    .Q(\sound1.divisor_m[14] ));
 sky130_fd_sc_hd__dfrtp_1 _7941_ (.CLK(net126),
    .D(_0104_),
    .RESET_B(net87),
    .Q(\sound1.divisor_m[15] ));
 sky130_fd_sc_hd__dfrtp_2 _7942_ (.CLK(net126),
    .D(_0105_),
    .RESET_B(net87),
    .Q(\sound1.divisor_m[16] ));
 sky130_fd_sc_hd__dfrtp_4 _7943_ (.CLK(net125),
    .D(_0106_),
    .RESET_B(net86),
    .Q(\sound1.divisor_m[17] ));
 sky130_fd_sc_hd__dfrtp_4 _7944_ (.CLK(net125),
    .D(_0107_),
    .RESET_B(net86),
    .Q(\sound1.divisor_m[18] ));
 sky130_fd_sc_hd__dfrtp_1 _7945_ (.CLK(net128),
    .D(_0108_),
    .RESET_B(net89),
    .Q(\sound1.sdiv.A[0] ));
 sky130_fd_sc_hd__dfrtp_1 _7946_ (.CLK(net128),
    .D(_0109_),
    .RESET_B(net89),
    .Q(\sound1.sdiv.A[1] ));
 sky130_fd_sc_hd__dfrtp_1 _7947_ (.CLK(net131),
    .D(_0110_),
    .RESET_B(net92),
    .Q(\sound1.sdiv.A[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7948_ (.CLK(net131),
    .D(_0111_),
    .RESET_B(net92),
    .Q(\sound1.sdiv.A[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7949_ (.CLK(net131),
    .D(_0112_),
    .RESET_B(net92),
    .Q(\sound1.sdiv.A[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7950_ (.CLK(net130),
    .D(_0113_),
    .RESET_B(net91),
    .Q(\sound1.sdiv.A[5] ));
 sky130_fd_sc_hd__dfrtp_1 _7951_ (.CLK(net131),
    .D(_0114_),
    .RESET_B(net92),
    .Q(\sound1.sdiv.A[6] ));
 sky130_fd_sc_hd__dfrtp_1 _7952_ (.CLK(net130),
    .D(_0115_),
    .RESET_B(net91),
    .Q(\sound1.sdiv.A[7] ));
 sky130_fd_sc_hd__dfrtp_1 _7953_ (.CLK(net130),
    .D(_0116_),
    .RESET_B(net91),
    .Q(\sound1.sdiv.A[8] ));
 sky130_fd_sc_hd__dfrtp_1 _7954_ (.CLK(net130),
    .D(_0117_),
    .RESET_B(net91),
    .Q(\sound1.sdiv.A[9] ));
 sky130_fd_sc_hd__dfrtp_1 _7955_ (.CLK(net130),
    .D(_0118_),
    .RESET_B(net91),
    .Q(\sound1.sdiv.A[10] ));
 sky130_fd_sc_hd__dfrtp_1 _7956_ (.CLK(net130),
    .D(_0119_),
    .RESET_B(net91),
    .Q(\sound1.sdiv.A[11] ));
 sky130_fd_sc_hd__dfrtp_1 _7957_ (.CLK(net130),
    .D(_0120_),
    .RESET_B(net91),
    .Q(\sound1.sdiv.A[12] ));
 sky130_fd_sc_hd__dfrtp_1 _7958_ (.CLK(net130),
    .D(_0121_),
    .RESET_B(net91),
    .Q(\sound1.sdiv.A[13] ));
 sky130_fd_sc_hd__dfrtp_1 _7959_ (.CLK(net130),
    .D(_0122_),
    .RESET_B(net91),
    .Q(\sound1.sdiv.A[14] ));
 sky130_fd_sc_hd__dfrtp_1 _7960_ (.CLK(net130),
    .D(_0123_),
    .RESET_B(net91),
    .Q(\sound1.sdiv.A[15] ));
 sky130_fd_sc_hd__dfrtp_1 _7961_ (.CLK(net130),
    .D(_0124_),
    .RESET_B(net91),
    .Q(\sound1.sdiv.A[16] ));
 sky130_fd_sc_hd__dfrtp_1 _7962_ (.CLK(net130),
    .D(_0125_),
    .RESET_B(net91),
    .Q(\sound1.sdiv.A[17] ));
 sky130_fd_sc_hd__dfrtp_1 _7963_ (.CLK(net130),
    .D(_0126_),
    .RESET_B(net91),
    .Q(\sound1.sdiv.A[18] ));
 sky130_fd_sc_hd__dfrtp_1 _7964_ (.CLK(net130),
    .D(_0127_),
    .RESET_B(net91),
    .Q(\sound1.sdiv.A[19] ));
 sky130_fd_sc_hd__dfrtp_2 _7965_ (.CLK(net130),
    .D(_0128_),
    .RESET_B(net91),
    .Q(\sound1.sdiv.A[20] ));
 sky130_fd_sc_hd__dfrtp_1 _7966_ (.CLK(net134),
    .D(_0129_),
    .RESET_B(net95),
    .Q(\sound1.sdiv.A[21] ));
 sky130_fd_sc_hd__dfrtp_1 _7967_ (.CLK(net134),
    .D(_0130_),
    .RESET_B(net95),
    .Q(\sound1.sdiv.A[22] ));
 sky130_fd_sc_hd__dfrtp_1 _7968_ (.CLK(net130),
    .D(_0131_),
    .RESET_B(net91),
    .Q(\sound1.sdiv.A[23] ));
 sky130_fd_sc_hd__dfrtp_1 _7969_ (.CLK(net134),
    .D(_0132_),
    .RESET_B(net95),
    .Q(\sound1.sdiv.A[24] ));
 sky130_fd_sc_hd__dfrtp_1 _7970_ (.CLK(net131),
    .D(_0133_),
    .RESET_B(net92),
    .Q(\sound1.sdiv.A[25] ));
 sky130_fd_sc_hd__dfrtp_4 _7971_ (.CLK(net130),
    .D(_0134_),
    .RESET_B(net91),
    .Q(\sound1.sdiv.A[26] ));
 sky130_fd_sc_hd__dfrtp_1 _7972_ (.CLK(net131),
    .D(_0135_),
    .RESET_B(net92),
    .Q(\sound1.sdiv.C[0] ));
 sky130_fd_sc_hd__dfrtp_1 _7973_ (.CLK(net131),
    .D(_0136_),
    .RESET_B(net92),
    .Q(\sound1.sdiv.C[1] ));
 sky130_fd_sc_hd__dfrtp_2 _7974_ (.CLK(net131),
    .D(_0137_),
    .RESET_B(net92),
    .Q(\sound1.sdiv.C[2] ));
 sky130_fd_sc_hd__dfrtp_2 _7975_ (.CLK(net131),
    .D(_0138_),
    .RESET_B(net92),
    .Q(\sound1.sdiv.C[3] ));
 sky130_fd_sc_hd__dfrtp_1 _7976_ (.CLK(net131),
    .D(_0139_),
    .RESET_B(net92),
    .Q(\sound1.sdiv.C[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7977_ (.CLK(net131),
    .D(_0140_),
    .RESET_B(net92),
    .Q(\sound1.sdiv.C[5] ));
 sky130_fd_sc_hd__dfrtp_1 _7978_ (.CLK(net131),
    .D(\sound1.sdiv.next_start ),
    .RESET_B(net92),
    .Q(\sound1.sdiv.start ));
 sky130_fd_sc_hd__dfstp_2 _7979_ (.CLK(net125),
    .D(\sound1.osc.next_count[0] ),
    .SET_B(net86),
    .Q(\sound1.count[0] ));
 sky130_fd_sc_hd__dfrtp_4 _7980_ (.CLK(net125),
    .D(\sound1.osc.next_count[1] ),
    .RESET_B(net86),
    .Q(\sound1.count[1] ));
 sky130_fd_sc_hd__dfrtp_2 _7981_ (.CLK(net125),
    .D(\sound1.osc.next_count[2] ),
    .RESET_B(net86),
    .Q(\sound1.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _7982_ (.CLK(net125),
    .D(\sound1.osc.next_count[3] ),
    .RESET_B(net86),
    .Q(\sound1.count[3] ));
 sky130_fd_sc_hd__dfrtp_2 _7983_ (.CLK(net134),
    .D(\sound1.osc.next_count[4] ),
    .RESET_B(net95),
    .Q(\sound1.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _7984_ (.CLK(net134),
    .D(\sound1.osc.next_count[5] ),
    .RESET_B(net95),
    .Q(\sound1.count[5] ));
 sky130_fd_sc_hd__dfrtp_2 _7985_ (.CLK(net134),
    .D(\sound1.osc.next_count[6] ),
    .RESET_B(net95),
    .Q(\sound1.count[6] ));
 sky130_fd_sc_hd__dfrtp_2 _7986_ (.CLK(net125),
    .D(\sound1.osc.next_count[7] ),
    .RESET_B(net86),
    .Q(\sound1.count[7] ));
 sky130_fd_sc_hd__dfrtp_1 _7987_ (.CLK(net125),
    .D(\sound1.osc.next_count[8] ),
    .RESET_B(net86),
    .Q(\sound1.count[8] ));
 sky130_fd_sc_hd__dfrtp_2 _7988_ (.CLK(net125),
    .D(\sound1.osc.next_count[9] ),
    .RESET_B(net86),
    .Q(\sound1.count[9] ));
 sky130_fd_sc_hd__dfrtp_2 _7989_ (.CLK(net125),
    .D(\sound1.osc.next_count[10] ),
    .RESET_B(net86),
    .Q(\sound1.count[10] ));
 sky130_fd_sc_hd__dfrtp_2 _7990_ (.CLK(net125),
    .D(\sound1.osc.next_count[11] ),
    .RESET_B(net86),
    .Q(\sound1.count[11] ));
 sky130_fd_sc_hd__dfrtp_2 _7991_ (.CLK(net125),
    .D(\sound1.osc.next_count[12] ),
    .RESET_B(net86),
    .Q(\sound1.count[12] ));
 sky130_fd_sc_hd__dfrtp_4 _7992_ (.CLK(net125),
    .D(\sound1.osc.next_count[13] ),
    .RESET_B(net86),
    .Q(\sound1.count[13] ));
 sky130_fd_sc_hd__dfrtp_1 _7993_ (.CLK(net125),
    .D(\sound1.osc.next_count[14] ),
    .RESET_B(net86),
    .Q(\sound1.count[14] ));
 sky130_fd_sc_hd__dfrtp_2 _7994_ (.CLK(net125),
    .D(\sound1.osc.next_count[15] ),
    .RESET_B(net86),
    .Q(\sound1.count[15] ));
 sky130_fd_sc_hd__dfrtp_2 _7995_ (.CLK(net125),
    .D(\sound1.osc.next_count[16] ),
    .RESET_B(net86),
    .Q(\sound1.count[16] ));
 sky130_fd_sc_hd__dfrtp_1 _7996_ (.CLK(net125),
    .D(\sound1.osc.next_count[17] ),
    .RESET_B(net86),
    .Q(\sound1.count[17] ));
 sky130_fd_sc_hd__dfrtp_2 _7997_ (.CLK(net134),
    .D(\sound1.osc.next_count[18] ),
    .RESET_B(net95),
    .Q(\sound1.count[18] ));
 sky130_fd_sc_hd__dfrtp_1 _7998_ (.CLK(net137),
    .D(\sound2.sdiv.next_dived ),
    .RESET_B(net98),
    .Q(\sound2.sdiv.dived ));
 sky130_fd_sc_hd__dfrtp_2 _7999_ (.CLK(net140),
    .D(_0141_),
    .RESET_B(net101),
    .Q(\sound1.sdiv.Q[0] ));
 sky130_fd_sc_hd__dfrtp_1 _8000_ (.CLK(net140),
    .D(_0142_),
    .RESET_B(net101),
    .Q(\sound1.sdiv.Q[1] ));
 sky130_fd_sc_hd__dfrtp_1 _8001_ (.CLK(net135),
    .D(_0143_),
    .RESET_B(net96),
    .Q(\sound1.sdiv.Q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _8002_ (.CLK(net135),
    .D(_0144_),
    .RESET_B(net96),
    .Q(\sound1.sdiv.Q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _8003_ (.CLK(net135),
    .D(_0145_),
    .RESET_B(net96),
    .Q(\sound1.sdiv.Q[4] ));
 sky130_fd_sc_hd__dfrtp_2 _8004_ (.CLK(net136),
    .D(_0146_),
    .RESET_B(net97),
    .Q(\sound1.sdiv.Q[5] ));
 sky130_fd_sc_hd__dfrtp_2 _8005_ (.CLK(net135),
    .D(_0147_),
    .RESET_B(net96),
    .Q(\sound1.sdiv.Q[6] ));
 sky130_fd_sc_hd__dfrtp_2 _8006_ (.CLK(net135),
    .D(_0148_),
    .RESET_B(net96),
    .Q(\sound1.sdiv.Q[7] ));
 sky130_fd_sc_hd__dfrtp_2 _8007_ (.CLK(net128),
    .D(_0149_),
    .RESET_B(net89),
    .Q(\sound1.sdiv.Q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _8008_ (.CLK(net128),
    .D(_0150_),
    .RESET_B(net89),
    .Q(\sound1.sdiv.Q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _8009_ (.CLK(net128),
    .D(_0151_),
    .RESET_B(net89),
    .Q(\sound1.sdiv.Q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _8010_ (.CLK(net128),
    .D(_0152_),
    .RESET_B(net89),
    .Q(\sound1.sdiv.Q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _8011_ (.CLK(net127),
    .D(_0153_),
    .RESET_B(net88),
    .Q(\sound1.sdiv.Q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _8012_ (.CLK(net127),
    .D(_0154_),
    .RESET_B(net88),
    .Q(\sound1.sdiv.Q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _8013_ (.CLK(net127),
    .D(_0155_),
    .RESET_B(net88),
    .Q(\sound1.sdiv.Q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _8014_ (.CLK(net127),
    .D(_0156_),
    .RESET_B(net88),
    .Q(\sound1.sdiv.Q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _8015_ (.CLK(net126),
    .D(_0157_),
    .RESET_B(net87),
    .Q(\sound1.sdiv.Q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _8016_ (.CLK(net126),
    .D(_0158_),
    .RESET_B(net87),
    .Q(\sound1.sdiv.Q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _8017_ (.CLK(net126),
    .D(_0159_),
    .RESET_B(net87),
    .Q(\sound1.sdiv.Q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _8018_ (.CLK(net126),
    .D(_0160_),
    .RESET_B(net87),
    .Q(\sound1.sdiv.Q[19] ));
 sky130_fd_sc_hd__dfrtp_1 _8019_ (.CLK(net126),
    .D(_0161_),
    .RESET_B(net87),
    .Q(\sound1.sdiv.Q[20] ));
 sky130_fd_sc_hd__dfrtp_1 _8020_ (.CLK(net126),
    .D(_0162_),
    .RESET_B(net87),
    .Q(\sound1.sdiv.Q[21] ));
 sky130_fd_sc_hd__dfrtp_1 _8021_ (.CLK(net126),
    .D(_0163_),
    .RESET_B(net87),
    .Q(\sound1.sdiv.Q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _8022_ (.CLK(net125),
    .D(_0164_),
    .RESET_B(net86),
    .Q(\sound1.sdiv.Q[23] ));
 sky130_fd_sc_hd__dfrtp_1 _8023_ (.CLK(net134),
    .D(_0165_),
    .RESET_B(net95),
    .Q(\sound1.sdiv.Q[24] ));
 sky130_fd_sc_hd__dfrtp_1 _8024_ (.CLK(net127),
    .D(_0166_),
    .RESET_B(net88),
    .Q(\sound1.sdiv.Q[25] ));
 sky130_fd_sc_hd__dfrtp_1 _8025_ (.CLK(net127),
    .D(_0167_),
    .RESET_B(net88),
    .Q(\sound1.sdiv.Q[26] ));
 sky130_fd_sc_hd__dfrtp_1 _8026_ (.CLK(net128),
    .D(_0168_),
    .RESET_B(net89),
    .Q(\sound1.sdiv.Q[27] ));
 sky130_fd_sc_hd__dfrtp_1 _8027_ (.CLK(net120),
    .D(_0169_),
    .RESET_B(net81),
    .Q(\sound2.count_m[0] ));
 sky130_fd_sc_hd__dfrtp_1 _8028_ (.CLK(net120),
    .D(_0170_),
    .RESET_B(net81),
    .Q(\sound2.count_m[1] ));
 sky130_fd_sc_hd__dfrtp_1 _8029_ (.CLK(net111),
    .D(_0171_),
    .RESET_B(net72),
    .Q(\sound2.count_m[2] ));
 sky130_fd_sc_hd__dfrtp_1 _8030_ (.CLK(net111),
    .D(_0172_),
    .RESET_B(net72),
    .Q(\sound2.count_m[3] ));
 sky130_fd_sc_hd__dfrtp_1 _8031_ (.CLK(net111),
    .D(_0173_),
    .RESET_B(net72),
    .Q(\sound2.count_m[4] ));
 sky130_fd_sc_hd__dfrtp_1 _8032_ (.CLK(net111),
    .D(_0174_),
    .RESET_B(net72),
    .Q(\sound2.count_m[5] ));
 sky130_fd_sc_hd__dfrtp_1 _8033_ (.CLK(net109),
    .D(_0175_),
    .RESET_B(net70),
    .Q(\sound2.count_m[6] ));
 sky130_fd_sc_hd__dfrtp_1 _8034_ (.CLK(net109),
    .D(_0176_),
    .RESET_B(net70),
    .Q(\sound2.count_m[7] ));
 sky130_fd_sc_hd__dfrtp_1 _8035_ (.CLK(net109),
    .D(_0177_),
    .RESET_B(net70),
    .Q(\sound2.count_m[8] ));
 sky130_fd_sc_hd__dfrtp_1 _8036_ (.CLK(net109),
    .D(_0178_),
    .RESET_B(net70),
    .Q(\sound2.count_m[9] ));
 sky130_fd_sc_hd__dfrtp_1 _8037_ (.CLK(net109),
    .D(_0179_),
    .RESET_B(net70),
    .Q(\sound2.count_m[10] ));
 sky130_fd_sc_hd__dfrtp_1 _8038_ (.CLK(net109),
    .D(_0180_),
    .RESET_B(net70),
    .Q(\sound2.count_m[11] ));
 sky130_fd_sc_hd__dfrtp_1 _8039_ (.CLK(net109),
    .D(_0181_),
    .RESET_B(net70),
    .Q(\sound2.count_m[12] ));
 sky130_fd_sc_hd__dfrtp_1 _8040_ (.CLK(net109),
    .D(_0182_),
    .RESET_B(net70),
    .Q(\sound2.count_m[13] ));
 sky130_fd_sc_hd__dfrtp_1 _8041_ (.CLK(net109),
    .D(_0183_),
    .RESET_B(net70),
    .Q(\sound2.count_m[14] ));
 sky130_fd_sc_hd__dfrtp_1 _8042_ (.CLK(net116),
    .D(_0184_),
    .RESET_B(net77),
    .Q(\sound2.count_m[15] ));
 sky130_fd_sc_hd__dfrtp_1 _8043_ (.CLK(net117),
    .D(_0185_),
    .RESET_B(net78),
    .Q(\sound2.count_m[16] ));
 sky130_fd_sc_hd__dfrtp_1 _8044_ (.CLK(net117),
    .D(_0186_),
    .RESET_B(net78),
    .Q(\sound2.count_m[17] ));
 sky130_fd_sc_hd__dfrtp_1 _8045_ (.CLK(net120),
    .D(_0187_),
    .RESET_B(net81),
    .Q(\sound2.count_m[18] ));
 sky130_fd_sc_hd__dfrtp_4 _8046_ (.CLK(net111),
    .D(_0188_),
    .RESET_B(net72),
    .Q(\sound2.divisor_m[0] ));
 sky130_fd_sc_hd__dfrtp_4 _8047_ (.CLK(net111),
    .D(_0189_),
    .RESET_B(net72),
    .Q(\sound2.divisor_m[1] ));
 sky130_fd_sc_hd__dfrtp_4 _8048_ (.CLK(net112),
    .D(_0190_),
    .RESET_B(net73),
    .Q(\sound2.divisor_m[2] ));
 sky130_fd_sc_hd__dfrtp_4 _8049_ (.CLK(net112),
    .D(_0191_),
    .RESET_B(net73),
    .Q(\sound2.divisor_m[3] ));
 sky130_fd_sc_hd__dfrtp_4 _8050_ (.CLK(net112),
    .D(_0192_),
    .RESET_B(net73),
    .Q(\sound2.divisor_m[4] ));
 sky130_fd_sc_hd__dfrtp_2 _8051_ (.CLK(net112),
    .D(_0193_),
    .RESET_B(net73),
    .Q(\sound2.divisor_m[5] ));
 sky130_fd_sc_hd__dfrtp_2 _8052_ (.CLK(net117),
    .D(_0194_),
    .RESET_B(net78),
    .Q(\sound2.divisor_m[6] ));
 sky130_fd_sc_hd__dfrtp_2 _8053_ (.CLK(net116),
    .D(_0195_),
    .RESET_B(net77),
    .Q(\sound2.divisor_m[7] ));
 sky130_fd_sc_hd__dfrtp_2 _8054_ (.CLK(net116),
    .D(_0196_),
    .RESET_B(net77),
    .Q(\sound2.divisor_m[8] ));
 sky130_fd_sc_hd__dfrtp_2 _8055_ (.CLK(net109),
    .D(_0197_),
    .RESET_B(net70),
    .Q(\sound2.divisor_m[9] ));
 sky130_fd_sc_hd__dfrtp_2 _8056_ (.CLK(net109),
    .D(_0198_),
    .RESET_B(net70),
    .Q(\sound2.divisor_m[10] ));
 sky130_fd_sc_hd__dfrtp_2 _8057_ (.CLK(net116),
    .D(_0199_),
    .RESET_B(net77),
    .Q(\sound2.divisor_m[11] ));
 sky130_fd_sc_hd__dfrtp_1 _8058_ (.CLK(net109),
    .D(_0200_),
    .RESET_B(net70),
    .Q(\sound2.divisor_m[12] ));
 sky130_fd_sc_hd__dfrtp_1 _8059_ (.CLK(net116),
    .D(_0201_),
    .RESET_B(net77),
    .Q(\sound2.divisor_m[13] ));
 sky130_fd_sc_hd__dfrtp_2 _8060_ (.CLK(net116),
    .D(_0202_),
    .RESET_B(net77),
    .Q(\sound2.divisor_m[14] ));
 sky130_fd_sc_hd__dfrtp_2 _8061_ (.CLK(net116),
    .D(_0203_),
    .RESET_B(net77),
    .Q(\sound2.divisor_m[15] ));
 sky130_fd_sc_hd__dfrtp_1 _8062_ (.CLK(net116),
    .D(_0204_),
    .RESET_B(net77),
    .Q(\sound2.divisor_m[16] ));
 sky130_fd_sc_hd__dfrtp_2 _8063_ (.CLK(net117),
    .D(_0205_),
    .RESET_B(net78),
    .Q(\sound2.divisor_m[17] ));
 sky130_fd_sc_hd__dfrtp_1 _8064_ (.CLK(net117),
    .D(_0206_),
    .RESET_B(net78),
    .Q(\sound2.divisor_m[18] ));
 sky130_fd_sc_hd__dfrtp_1 _8065_ (.CLK(net117),
    .D(_0207_),
    .RESET_B(net78),
    .Q(\sound2.sdiv.A[0] ));
 sky130_fd_sc_hd__dfrtp_1 _8066_ (.CLK(net117),
    .D(_0208_),
    .RESET_B(net78),
    .Q(\sound2.sdiv.A[1] ));
 sky130_fd_sc_hd__dfrtp_1 _8067_ (.CLK(net117),
    .D(_0209_),
    .RESET_B(net78),
    .Q(\sound2.sdiv.A[2] ));
 sky130_fd_sc_hd__dfrtp_1 _8068_ (.CLK(net117),
    .D(_0210_),
    .RESET_B(net78),
    .Q(\sound2.sdiv.A[3] ));
 sky130_fd_sc_hd__dfrtp_1 _8069_ (.CLK(net117),
    .D(_0211_),
    .RESET_B(net78),
    .Q(\sound2.sdiv.A[4] ));
 sky130_fd_sc_hd__dfrtp_1 _8070_ (.CLK(net117),
    .D(_0212_),
    .RESET_B(net78),
    .Q(\sound2.sdiv.A[5] ));
 sky130_fd_sc_hd__dfrtp_1 _8071_ (.CLK(net116),
    .D(_0213_),
    .RESET_B(net77),
    .Q(\sound2.sdiv.A[6] ));
 sky130_fd_sc_hd__dfrtp_1 _8072_ (.CLK(net116),
    .D(_0214_),
    .RESET_B(net77),
    .Q(\sound2.sdiv.A[7] ));
 sky130_fd_sc_hd__dfrtp_1 _8073_ (.CLK(net116),
    .D(_0215_),
    .RESET_B(net77),
    .Q(\sound2.sdiv.A[8] ));
 sky130_fd_sc_hd__dfrtp_1 _8074_ (.CLK(net116),
    .D(_0216_),
    .RESET_B(net77),
    .Q(\sound2.sdiv.A[9] ));
 sky130_fd_sc_hd__dfrtp_1 _8075_ (.CLK(net116),
    .D(_0217_),
    .RESET_B(net77),
    .Q(\sound2.sdiv.A[10] ));
 sky130_fd_sc_hd__dfrtp_1 _8076_ (.CLK(net116),
    .D(_0218_),
    .RESET_B(net77),
    .Q(\sound2.sdiv.A[11] ));
 sky130_fd_sc_hd__dfrtp_1 _8077_ (.CLK(net116),
    .D(_0219_),
    .RESET_B(net77),
    .Q(\sound2.sdiv.A[12] ));
 sky130_fd_sc_hd__dfrtp_1 _8078_ (.CLK(net116),
    .D(_0220_),
    .RESET_B(net77),
    .Q(\sound2.sdiv.A[13] ));
 sky130_fd_sc_hd__dfrtp_1 _8079_ (.CLK(net116),
    .D(_0221_),
    .RESET_B(net77),
    .Q(\sound2.sdiv.A[14] ));
 sky130_fd_sc_hd__dfrtp_1 _8080_ (.CLK(net116),
    .D(_0222_),
    .RESET_B(net77),
    .Q(\sound2.sdiv.A[15] ));
 sky130_fd_sc_hd__dfrtp_1 _8081_ (.CLK(net116),
    .D(_0223_),
    .RESET_B(net77),
    .Q(\sound2.sdiv.A[16] ));
 sky130_fd_sc_hd__dfrtp_1 _8082_ (.CLK(net119),
    .D(_0224_),
    .RESET_B(net80),
    .Q(\sound2.sdiv.A[17] ));
 sky130_fd_sc_hd__dfrtp_1 _8083_ (.CLK(net119),
    .D(_0225_),
    .RESET_B(net80),
    .Q(\sound2.sdiv.A[18] ));
 sky130_fd_sc_hd__dfrtp_1 _8084_ (.CLK(net118),
    .D(_0226_),
    .RESET_B(net79),
    .Q(\sound2.sdiv.A[19] ));
 sky130_fd_sc_hd__dfrtp_1 _8085_ (.CLK(net118),
    .D(_0227_),
    .RESET_B(net79),
    .Q(\sound2.sdiv.A[20] ));
 sky130_fd_sc_hd__dfrtp_1 _8086_ (.CLK(net119),
    .D(_0228_),
    .RESET_B(net80),
    .Q(\sound2.sdiv.A[21] ));
 sky130_fd_sc_hd__dfrtp_1 _8087_ (.CLK(net117),
    .D(_0229_),
    .RESET_B(net78),
    .Q(\sound2.sdiv.A[22] ));
 sky130_fd_sc_hd__dfrtp_1 _8088_ (.CLK(net118),
    .D(_0230_),
    .RESET_B(net79),
    .Q(\sound2.sdiv.A[23] ));
 sky130_fd_sc_hd__dfrtp_1 _8089_ (.CLK(net118),
    .D(_0231_),
    .RESET_B(net79),
    .Q(\sound2.sdiv.A[24] ));
 sky130_fd_sc_hd__dfrtp_1 _8090_ (.CLK(net118),
    .D(_0232_),
    .RESET_B(net79),
    .Q(\sound2.sdiv.A[25] ));
 sky130_fd_sc_hd__dfrtp_4 _8091_ (.CLK(net117),
    .D(_0233_),
    .RESET_B(net78),
    .Q(\sound2.sdiv.A[26] ));
 sky130_fd_sc_hd__dfrtp_1 _8092_ (.CLK(net117),
    .D(_0234_),
    .RESET_B(net78),
    .Q(\sound2.sdiv.C[0] ));
 sky130_fd_sc_hd__dfrtp_1 _8093_ (.CLK(net117),
    .D(_0235_),
    .RESET_B(net78),
    .Q(\sound2.sdiv.C[1] ));
 sky130_fd_sc_hd__dfrtp_2 _8094_ (.CLK(net119),
    .D(_0236_),
    .RESET_B(net80),
    .Q(\sound2.sdiv.C[2] ));
 sky130_fd_sc_hd__dfrtp_2 _8095_ (.CLK(net119),
    .D(_0237_),
    .RESET_B(net80),
    .Q(\sound2.sdiv.C[3] ));
 sky130_fd_sc_hd__dfrtp_1 _8096_ (.CLK(net118),
    .D(_0238_),
    .RESET_B(net79),
    .Q(\sound2.sdiv.C[4] ));
 sky130_fd_sc_hd__dfrtp_1 _8097_ (.CLK(net118),
    .D(_0239_),
    .RESET_B(net79),
    .Q(\sound2.sdiv.C[5] ));
 sky130_fd_sc_hd__dfrtp_1 _8098_ (.CLK(net136),
    .D(\sound2.sdiv.next_start ),
    .RESET_B(net97),
    .Q(\sound2.sdiv.start ));
 sky130_fd_sc_hd__dfstp_1 _8099_ (.CLK(net111),
    .D(\sound2.osc.next_count[0] ),
    .SET_B(net72),
    .Q(\sound2.count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _8100_ (.CLK(net111),
    .D(\sound2.osc.next_count[1] ),
    .RESET_B(net72),
    .Q(\sound2.count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _8101_ (.CLK(net111),
    .D(\sound2.osc.next_count[2] ),
    .RESET_B(net72),
    .Q(\sound2.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _8102_ (.CLK(net111),
    .D(\sound2.osc.next_count[3] ),
    .RESET_B(net72),
    .Q(\sound2.count[3] ));
 sky130_fd_sc_hd__dfrtp_2 _8103_ (.CLK(net111),
    .D(\sound2.osc.next_count[4] ),
    .RESET_B(net72),
    .Q(\sound2.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _8104_ (.CLK(net111),
    .D(\sound2.osc.next_count[5] ),
    .RESET_B(net72),
    .Q(\sound2.count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _8105_ (.CLK(net111),
    .D(\sound2.osc.next_count[6] ),
    .RESET_B(net72),
    .Q(\sound2.count[6] ));
 sky130_fd_sc_hd__dfrtp_1 _8106_ (.CLK(net111),
    .D(\sound2.osc.next_count[7] ),
    .RESET_B(net72),
    .Q(\sound2.count[7] ));
 sky130_fd_sc_hd__dfrtp_2 _8107_ (.CLK(net110),
    .D(\sound2.osc.next_count[8] ),
    .RESET_B(net71),
    .Q(\sound2.count[8] ));
 sky130_fd_sc_hd__dfrtp_1 _8108_ (.CLK(net110),
    .D(\sound2.osc.next_count[9] ),
    .RESET_B(net71),
    .Q(\sound2.count[9] ));
 sky130_fd_sc_hd__dfrtp_2 _8109_ (.CLK(net110),
    .D(\sound2.osc.next_count[10] ),
    .RESET_B(net71),
    .Q(\sound2.count[10] ));
 sky130_fd_sc_hd__dfrtp_2 _8110_ (.CLK(net110),
    .D(\sound2.osc.next_count[11] ),
    .RESET_B(net71),
    .Q(\sound2.count[11] ));
 sky130_fd_sc_hd__dfrtp_2 _8111_ (.CLK(net110),
    .D(\sound2.osc.next_count[12] ),
    .RESET_B(net71),
    .Q(\sound2.count[12] ));
 sky130_fd_sc_hd__dfrtp_4 _8112_ (.CLK(net110),
    .D(\sound2.osc.next_count[13] ),
    .RESET_B(net71),
    .Q(\sound2.count[13] ));
 sky130_fd_sc_hd__dfrtp_2 _8113_ (.CLK(net110),
    .D(\sound2.osc.next_count[14] ),
    .RESET_B(net71),
    .Q(\sound2.count[14] ));
 sky130_fd_sc_hd__dfrtp_2 _8114_ (.CLK(net112),
    .D(\sound2.osc.next_count[15] ),
    .RESET_B(net73),
    .Q(\sound2.count[15] ));
 sky130_fd_sc_hd__dfrtp_2 _8115_ (.CLK(net112),
    .D(\sound2.osc.next_count[16] ),
    .RESET_B(net73),
    .Q(\sound2.count[16] ));
 sky130_fd_sc_hd__dfrtp_2 _8116_ (.CLK(net112),
    .D(\sound2.osc.next_count[17] ),
    .RESET_B(net73),
    .Q(\sound2.count[17] ));
 sky130_fd_sc_hd__dfrtp_1 _8117_ (.CLK(net112),
    .D(\sound2.osc.next_count[18] ),
    .RESET_B(net73),
    .Q(\sound2.count[18] ));
 sky130_fd_sc_hd__dfrtp_1 _8118_ (.CLK(net140),
    .D(\sound3.sdiv.next_dived ),
    .RESET_B(net101),
    .Q(\sound3.sdiv.dived ));
 sky130_fd_sc_hd__dfrtp_2 _8119_ (.CLK(net136),
    .D(_0240_),
    .RESET_B(net97),
    .Q(\sound2.sdiv.Q[0] ));
 sky130_fd_sc_hd__dfrtp_2 _8120_ (.CLK(net136),
    .D(_0241_),
    .RESET_B(net97),
    .Q(\sound2.sdiv.Q[1] ));
 sky130_fd_sc_hd__dfrtp_2 _8121_ (.CLK(net136),
    .D(_0242_),
    .RESET_B(net97),
    .Q(\sound2.sdiv.Q[2] ));
 sky130_fd_sc_hd__dfrtp_1 _8122_ (.CLK(net136),
    .D(_0243_),
    .RESET_B(net97),
    .Q(\sound2.sdiv.Q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _8123_ (.CLK(net136),
    .D(_0244_),
    .RESET_B(net97),
    .Q(\sound2.sdiv.Q[4] ));
 sky130_fd_sc_hd__dfrtp_2 _8124_ (.CLK(net136),
    .D(_0245_),
    .RESET_B(net97),
    .Q(\sound2.sdiv.Q[5] ));
 sky130_fd_sc_hd__dfrtp_2 _8125_ (.CLK(net136),
    .D(_0246_),
    .RESET_B(net97),
    .Q(\sound2.sdiv.Q[6] ));
 sky130_fd_sc_hd__dfrtp_4 _8126_ (.CLK(net136),
    .D(_0247_),
    .RESET_B(net97),
    .Q(\sound2.sdiv.Q[7] ));
 sky130_fd_sc_hd__dfrtp_2 _8127_ (.CLK(net120),
    .D(_0248_),
    .RESET_B(net81),
    .Q(\sound2.sdiv.Q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _8128_ (.CLK(net120),
    .D(_0249_),
    .RESET_B(net81),
    .Q(\sound2.sdiv.Q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _8129_ (.CLK(net112),
    .D(_0250_),
    .RESET_B(net73),
    .Q(\sound2.sdiv.Q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _8130_ (.CLK(net112),
    .D(_0251_),
    .RESET_B(net73),
    .Q(\sound2.sdiv.Q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _8131_ (.CLK(net112),
    .D(_0252_),
    .RESET_B(net73),
    .Q(\sound2.sdiv.Q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _8132_ (.CLK(net112),
    .D(_0253_),
    .RESET_B(net73),
    .Q(\sound2.sdiv.Q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _8133_ (.CLK(net109),
    .D(_0254_),
    .RESET_B(net70),
    .Q(\sound2.sdiv.Q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _8134_ (.CLK(net109),
    .D(_0255_),
    .RESET_B(net70),
    .Q(\sound2.sdiv.Q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _8135_ (.CLK(net110),
    .D(_0256_),
    .RESET_B(net71),
    .Q(\sound2.sdiv.Q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _8136_ (.CLK(net110),
    .D(_0257_),
    .RESET_B(net71),
    .Q(\sound2.sdiv.Q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _8137_ (.CLK(net109),
    .D(_0258_),
    .RESET_B(net70),
    .Q(\sound2.sdiv.Q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _8138_ (.CLK(net109),
    .D(_0259_),
    .RESET_B(net70),
    .Q(\sound2.sdiv.Q[19] ));
 sky130_fd_sc_hd__dfrtp_1 _8139_ (.CLK(net109),
    .D(_0260_),
    .RESET_B(net70),
    .Q(\sound2.sdiv.Q[20] ));
 sky130_fd_sc_hd__dfrtp_1 _8140_ (.CLK(net109),
    .D(_0261_),
    .RESET_B(net70),
    .Q(\sound2.sdiv.Q[21] ));
 sky130_fd_sc_hd__dfrtp_1 _8141_ (.CLK(net109),
    .D(_0262_),
    .RESET_B(net70),
    .Q(\sound2.sdiv.Q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _8142_ (.CLK(net116),
    .D(_0263_),
    .RESET_B(net77),
    .Q(\sound2.sdiv.Q[23] ));
 sky130_fd_sc_hd__dfrtp_1 _8143_ (.CLK(net117),
    .D(_0264_),
    .RESET_B(net78),
    .Q(\sound2.sdiv.Q[24] ));
 sky130_fd_sc_hd__dfrtp_1 _8144_ (.CLK(net117),
    .D(_0265_),
    .RESET_B(net78),
    .Q(\sound2.sdiv.Q[25] ));
 sky130_fd_sc_hd__dfrtp_1 _8145_ (.CLK(net117),
    .D(_0266_),
    .RESET_B(net78),
    .Q(\sound2.sdiv.Q[26] ));
 sky130_fd_sc_hd__dfrtp_1 _8146_ (.CLK(net117),
    .D(_0267_),
    .RESET_B(net78),
    .Q(\sound2.sdiv.Q[27] ));
 sky130_fd_sc_hd__dfrtp_1 _8147_ (.CLK(net140),
    .D(_0268_),
    .RESET_B(net101),
    .Q(\sound3.count_m[0] ));
 sky130_fd_sc_hd__dfrtp_1 _8148_ (.CLK(net140),
    .D(_0269_),
    .RESET_B(net101),
    .Q(\sound3.count_m[1] ));
 sky130_fd_sc_hd__dfrtp_1 _8149_ (.CLK(net135),
    .D(_0270_),
    .RESET_B(net96),
    .Q(\sound3.count_m[2] ));
 sky130_fd_sc_hd__dfrtp_1 _8150_ (.CLK(net131),
    .D(_0271_),
    .RESET_B(net92),
    .Q(\sound3.count_m[3] ));
 sky130_fd_sc_hd__dfrtp_1 _8151_ (.CLK(net131),
    .D(_0272_),
    .RESET_B(net92),
    .Q(\sound3.count_m[4] ));
 sky130_fd_sc_hd__dfrtp_1 _8152_ (.CLK(net131),
    .D(_0273_),
    .RESET_B(net92),
    .Q(\sound3.count_m[5] ));
 sky130_fd_sc_hd__dfrtp_1 _8153_ (.CLK(net132),
    .D(_0274_),
    .RESET_B(net93),
    .Q(\sound3.count_m[6] ));
 sky130_fd_sc_hd__dfrtp_1 _8154_ (.CLK(net132),
    .D(_0275_),
    .RESET_B(net93),
    .Q(\sound3.count_m[7] ));
 sky130_fd_sc_hd__dfrtp_1 _8155_ (.CLK(net131),
    .D(_0276_),
    .RESET_B(net92),
    .Q(\sound3.count_m[8] ));
 sky130_fd_sc_hd__dfrtp_1 _8156_ (.CLK(net132),
    .D(_0277_),
    .RESET_B(net93),
    .Q(\sound3.count_m[9] ));
 sky130_fd_sc_hd__dfrtp_1 _8157_ (.CLK(net132),
    .D(_0278_),
    .RESET_B(net93),
    .Q(\sound3.count_m[10] ));
 sky130_fd_sc_hd__dfrtp_1 _8158_ (.CLK(net132),
    .D(_0279_),
    .RESET_B(net93),
    .Q(\sound3.count_m[11] ));
 sky130_fd_sc_hd__dfrtp_1 _8159_ (.CLK(net132),
    .D(_0280_),
    .RESET_B(net93),
    .Q(\sound3.count_m[12] ));
 sky130_fd_sc_hd__dfrtp_1 _8160_ (.CLK(net132),
    .D(_0281_),
    .RESET_B(net93),
    .Q(\sound3.count_m[13] ));
 sky130_fd_sc_hd__dfrtp_1 _8161_ (.CLK(net132),
    .D(_0282_),
    .RESET_B(net93),
    .Q(\sound3.count_m[14] ));
 sky130_fd_sc_hd__dfrtp_1 _8162_ (.CLK(net140),
    .D(_0283_),
    .RESET_B(net101),
    .Q(\sound3.count_m[15] ));
 sky130_fd_sc_hd__dfrtp_1 _8163_ (.CLK(net140),
    .D(_0284_),
    .RESET_B(net101),
    .Q(\sound3.count_m[16] ));
 sky130_fd_sc_hd__dfrtp_1 _8164_ (.CLK(net135),
    .D(_0285_),
    .RESET_B(net96),
    .Q(\sound3.count_m[17] ));
 sky130_fd_sc_hd__dfrtp_1 _8165_ (.CLK(net140),
    .D(_0286_),
    .RESET_B(net101),
    .Q(\sound3.count_m[18] ));
 sky130_fd_sc_hd__dfrtp_4 _8166_ (.CLK(net135),
    .D(_0287_),
    .RESET_B(net96),
    .Q(\sound3.divisor_m[0] ));
 sky130_fd_sc_hd__dfrtp_4 _8167_ (.CLK(net140),
    .D(_0288_),
    .RESET_B(net101),
    .Q(\sound3.divisor_m[1] ));
 sky130_fd_sc_hd__dfrtp_2 _8168_ (.CLK(net140),
    .D(_0289_),
    .RESET_B(net101),
    .Q(\sound3.divisor_m[2] ));
 sky130_fd_sc_hd__dfrtp_2 _8169_ (.CLK(net140),
    .D(_0290_),
    .RESET_B(net101),
    .Q(\sound3.divisor_m[3] ));
 sky130_fd_sc_hd__dfrtp_4 _8170_ (.CLK(net135),
    .D(_0291_),
    .RESET_B(net96),
    .Q(\sound3.divisor_m[4] ));
 sky130_fd_sc_hd__dfrtp_2 _8171_ (.CLK(net135),
    .D(_0292_),
    .RESET_B(net96),
    .Q(\sound3.divisor_m[5] ));
 sky130_fd_sc_hd__dfrtp_4 _8172_ (.CLK(net135),
    .D(_0293_),
    .RESET_B(net96),
    .Q(\sound3.divisor_m[6] ));
 sky130_fd_sc_hd__dfrtp_4 _8173_ (.CLK(net132),
    .D(_0294_),
    .RESET_B(net93),
    .Q(\sound3.divisor_m[7] ));
 sky130_fd_sc_hd__dfrtp_2 _8174_ (.CLK(net132),
    .D(_0295_),
    .RESET_B(net93),
    .Q(\sound3.divisor_m[8] ));
 sky130_fd_sc_hd__dfrtp_2 _8175_ (.CLK(net133),
    .D(_0296_),
    .RESET_B(net94),
    .Q(\sound3.divisor_m[9] ));
 sky130_fd_sc_hd__dfrtp_2 _8176_ (.CLK(net133),
    .D(_0297_),
    .RESET_B(net94),
    .Q(\sound3.divisor_m[10] ));
 sky130_fd_sc_hd__dfrtp_2 _8177_ (.CLK(net133),
    .D(_0298_),
    .RESET_B(net94),
    .Q(\sound3.divisor_m[11] ));
 sky130_fd_sc_hd__dfrtp_2 _8178_ (.CLK(net133),
    .D(_0299_),
    .RESET_B(net94),
    .Q(\sound3.divisor_m[12] ));
 sky130_fd_sc_hd__dfrtp_2 _8179_ (.CLK(net133),
    .D(_0300_),
    .RESET_B(net94),
    .Q(\sound3.divisor_m[13] ));
 sky130_fd_sc_hd__dfrtp_2 _8180_ (.CLK(net140),
    .D(_0301_),
    .RESET_B(net101),
    .Q(\sound3.divisor_m[14] ));
 sky130_fd_sc_hd__dfrtp_2 _8181_ (.CLK(net142),
    .D(_0302_),
    .RESET_B(net103),
    .Q(\sound3.divisor_m[15] ));
 sky130_fd_sc_hd__dfrtp_2 _8182_ (.CLK(net140),
    .D(_0303_),
    .RESET_B(net101),
    .Q(\sound3.divisor_m[16] ));
 sky130_fd_sc_hd__dfrtp_4 _8183_ (.CLK(net135),
    .D(_0304_),
    .RESET_B(net96),
    .Q(\sound3.divisor_m[17] ));
 sky130_fd_sc_hd__dfrtp_2 _8184_ (.CLK(net140),
    .D(_0305_),
    .RESET_B(net101),
    .Q(\sound3.divisor_m[18] ));
 sky130_fd_sc_hd__dfrtp_1 _8185_ (.CLK(net140),
    .D(_0306_),
    .RESET_B(net101),
    .Q(\sound3.sdiv.A[0] ));
 sky130_fd_sc_hd__dfrtp_1 _8186_ (.CLK(net141),
    .D(_0307_),
    .RESET_B(net102),
    .Q(\sound3.sdiv.A[1] ));
 sky130_fd_sc_hd__dfrtp_1 _8187_ (.CLK(net142),
    .D(_0308_),
    .RESET_B(net103),
    .Q(\sound3.sdiv.A[2] ));
 sky130_fd_sc_hd__dfrtp_1 _8188_ (.CLK(net142),
    .D(_0309_),
    .RESET_B(net103),
    .Q(\sound3.sdiv.A[3] ));
 sky130_fd_sc_hd__dfrtp_1 _8189_ (.CLK(net142),
    .D(_0310_),
    .RESET_B(net103),
    .Q(\sound3.sdiv.A[4] ));
 sky130_fd_sc_hd__dfrtp_1 _8190_ (.CLK(net142),
    .D(_0311_),
    .RESET_B(net103),
    .Q(\sound3.sdiv.A[5] ));
 sky130_fd_sc_hd__dfrtp_1 _8191_ (.CLK(net142),
    .D(_0312_),
    .RESET_B(net103),
    .Q(\sound3.sdiv.A[6] ));
 sky130_fd_sc_hd__dfrtp_1 _8192_ (.CLK(net142),
    .D(_0313_),
    .RESET_B(net103),
    .Q(\sound3.sdiv.A[7] ));
 sky130_fd_sc_hd__dfrtp_1 _8193_ (.CLK(net133),
    .D(_0314_),
    .RESET_B(net94),
    .Q(\sound3.sdiv.A[8] ));
 sky130_fd_sc_hd__dfrtp_1 _8194_ (.CLK(net133),
    .D(_0315_),
    .RESET_B(net94),
    .Q(\sound3.sdiv.A[9] ));
 sky130_fd_sc_hd__dfrtp_1 _8195_ (.CLK(net133),
    .D(_0316_),
    .RESET_B(net94),
    .Q(\sound3.sdiv.A[10] ));
 sky130_fd_sc_hd__dfrtp_1 _8196_ (.CLK(net133),
    .D(_0317_),
    .RESET_B(net94),
    .Q(\sound3.sdiv.A[11] ));
 sky130_fd_sc_hd__dfrtp_1 _8197_ (.CLK(net133),
    .D(_0318_),
    .RESET_B(net94),
    .Q(\sound3.sdiv.A[12] ));
 sky130_fd_sc_hd__dfrtp_1 _8198_ (.CLK(net133),
    .D(_0319_),
    .RESET_B(net94),
    .Q(\sound3.sdiv.A[13] ));
 sky130_fd_sc_hd__dfrtp_1 _8199_ (.CLK(net142),
    .D(_0320_),
    .RESET_B(net103),
    .Q(\sound3.sdiv.A[14] ));
 sky130_fd_sc_hd__dfrtp_1 _8200_ (.CLK(net142),
    .D(_0321_),
    .RESET_B(net103),
    .Q(\sound3.sdiv.A[15] ));
 sky130_fd_sc_hd__dfrtp_1 _8201_ (.CLK(net142),
    .D(_0322_),
    .RESET_B(net103),
    .Q(\sound3.sdiv.A[16] ));
 sky130_fd_sc_hd__dfrtp_1 _8202_ (.CLK(net142),
    .D(_0323_),
    .RESET_B(net103),
    .Q(\sound3.sdiv.A[17] ));
 sky130_fd_sc_hd__dfrtp_2 _8203_ (.CLK(net142),
    .D(_0324_),
    .RESET_B(net103),
    .Q(\sound3.sdiv.A[18] ));
 sky130_fd_sc_hd__dfrtp_2 _8204_ (.CLK(net142),
    .D(_0325_),
    .RESET_B(net103),
    .Q(\sound3.sdiv.A[19] ));
 sky130_fd_sc_hd__dfrtp_2 _8205_ (.CLK(net142),
    .D(_0326_),
    .RESET_B(net103),
    .Q(\sound3.sdiv.A[20] ));
 sky130_fd_sc_hd__dfrtp_1 _8206_ (.CLK(net144),
    .D(_0327_),
    .RESET_B(net105),
    .Q(\sound3.sdiv.A[21] ));
 sky130_fd_sc_hd__dfrtp_1 _8207_ (.CLK(net142),
    .D(_0328_),
    .RESET_B(net103),
    .Q(\sound3.sdiv.A[22] ));
 sky130_fd_sc_hd__dfrtp_1 _8208_ (.CLK(net144),
    .D(_0329_),
    .RESET_B(net105),
    .Q(\sound3.sdiv.A[23] ));
 sky130_fd_sc_hd__dfrtp_1 _8209_ (.CLK(net144),
    .D(_0330_),
    .RESET_B(net105),
    .Q(\sound3.sdiv.A[24] ));
 sky130_fd_sc_hd__dfrtp_1 _8210_ (.CLK(net144),
    .D(_0331_),
    .RESET_B(net105),
    .Q(\sound3.sdiv.A[25] ));
 sky130_fd_sc_hd__dfrtp_4 _8211_ (.CLK(net142),
    .D(_0332_),
    .RESET_B(net103),
    .Q(\sound3.sdiv.A[26] ));
 sky130_fd_sc_hd__dfrtp_1 _8212_ (.CLK(net142),
    .D(_0333_),
    .RESET_B(net103),
    .Q(\sound3.sdiv.C[0] ));
 sky130_fd_sc_hd__dfrtp_1 _8213_ (.CLK(net145),
    .D(_0334_),
    .RESET_B(net106),
    .Q(\sound3.sdiv.C[1] ));
 sky130_fd_sc_hd__dfrtp_2 _8214_ (.CLK(net145),
    .D(_0335_),
    .RESET_B(net106),
    .Q(\sound3.sdiv.C[2] ));
 sky130_fd_sc_hd__dfrtp_2 _8215_ (.CLK(net144),
    .D(_0336_),
    .RESET_B(net105),
    .Q(\sound3.sdiv.C[3] ));
 sky130_fd_sc_hd__dfrtp_1 _8216_ (.CLK(net141),
    .D(_0337_),
    .RESET_B(net102),
    .Q(\sound3.sdiv.C[4] ));
 sky130_fd_sc_hd__dfrtp_1 _8217_ (.CLK(net144),
    .D(_0338_),
    .RESET_B(net105),
    .Q(\sound3.sdiv.C[5] ));
 sky130_fd_sc_hd__dfrtp_1 _8218_ (.CLK(net141),
    .D(\sound3.sdiv.next_start ),
    .RESET_B(net102),
    .Q(\sound3.sdiv.start ));
 sky130_fd_sc_hd__dfstp_2 _8219_ (.CLK(net135),
    .D(\sound3.osc.next_count[0] ),
    .SET_B(net96),
    .Q(\sound3.count[0] ));
 sky130_fd_sc_hd__dfrtp_4 _8220_ (.CLK(net135),
    .D(\sound3.osc.next_count[1] ),
    .RESET_B(net96),
    .Q(\sound3.count[1] ));
 sky130_fd_sc_hd__dfrtp_2 _8221_ (.CLK(net128),
    .D(\sound3.osc.next_count[2] ),
    .RESET_B(net89),
    .Q(\sound3.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _8222_ (.CLK(net128),
    .D(\sound3.osc.next_count[3] ),
    .RESET_B(net89),
    .Q(\sound3.count[3] ));
 sky130_fd_sc_hd__dfrtp_4 _8223_ (.CLK(net129),
    .D(\sound3.osc.next_count[4] ),
    .RESET_B(net90),
    .Q(\sound3.count[4] ));
 sky130_fd_sc_hd__dfrtp_2 _8224_ (.CLK(net129),
    .D(\sound3.osc.next_count[5] ),
    .RESET_B(net90),
    .Q(\sound3.count[5] ));
 sky130_fd_sc_hd__dfrtp_2 _8225_ (.CLK(net129),
    .D(\sound3.osc.next_count[6] ),
    .RESET_B(net90),
    .Q(\sound3.count[6] ));
 sky130_fd_sc_hd__dfrtp_2 _8226_ (.CLK(net128),
    .D(\sound3.osc.next_count[7] ),
    .RESET_B(net89),
    .Q(\sound3.count[7] ));
 sky130_fd_sc_hd__dfrtp_2 _8227_ (.CLK(net129),
    .D(\sound3.osc.next_count[8] ),
    .RESET_B(net90),
    .Q(\sound3.count[8] ));
 sky130_fd_sc_hd__dfrtp_2 _8228_ (.CLK(net128),
    .D(\sound3.osc.next_count[9] ),
    .RESET_B(net89),
    .Q(\sound3.count[9] ));
 sky130_fd_sc_hd__dfrtp_2 _8229_ (.CLK(net128),
    .D(\sound3.osc.next_count[10] ),
    .RESET_B(net89),
    .Q(\sound3.count[10] ));
 sky130_fd_sc_hd__dfrtp_1 _8230_ (.CLK(net129),
    .D(\sound3.osc.next_count[11] ),
    .RESET_B(net90),
    .Q(\sound3.count[11] ));
 sky130_fd_sc_hd__dfrtp_2 _8231_ (.CLK(net129),
    .D(\sound3.osc.next_count[12] ),
    .RESET_B(net90),
    .Q(\sound3.count[12] ));
 sky130_fd_sc_hd__dfrtp_2 _8232_ (.CLK(net129),
    .D(\sound3.osc.next_count[13] ),
    .RESET_B(net90),
    .Q(\sound3.count[13] ));
 sky130_fd_sc_hd__dfrtp_1 _8233_ (.CLK(net129),
    .D(\sound3.osc.next_count[14] ),
    .RESET_B(net90),
    .Q(\sound3.count[14] ));
 sky130_fd_sc_hd__dfrtp_2 _8234_ (.CLK(net135),
    .D(\sound3.osc.next_count[15] ),
    .RESET_B(net96),
    .Q(\sound3.count[15] ));
 sky130_fd_sc_hd__dfrtp_2 _8235_ (.CLK(net135),
    .D(\sound3.osc.next_count[16] ),
    .RESET_B(net96),
    .Q(\sound3.count[16] ));
 sky130_fd_sc_hd__dfrtp_1 _8236_ (.CLK(net135),
    .D(\sound3.osc.next_count[17] ),
    .RESET_B(net96),
    .Q(\sound3.count[17] ));
 sky130_fd_sc_hd__dfrtp_1 _8237_ (.CLK(net135),
    .D(\sound3.osc.next_count[18] ),
    .RESET_B(net96),
    .Q(\sound3.count[18] ));
 sky130_fd_sc_hd__dfrtp_1 _8238_ (.CLK(net137),
    .D(\sound4.sdiv.next_dived ),
    .RESET_B(net98),
    .Q(\sound4.sdiv.dived ));
 sky130_fd_sc_hd__dfrtp_1 _8239_ (.CLK(net143),
    .D(_0339_),
    .RESET_B(net104),
    .Q(\sound3.sdiv.Q[0] ));
 sky130_fd_sc_hd__dfrtp_2 _8240_ (.CLK(net143),
    .D(_0340_),
    .RESET_B(net104),
    .Q(\sound3.sdiv.Q[1] ));
 sky130_fd_sc_hd__dfrtp_2 _8241_ (.CLK(net143),
    .D(_0341_),
    .RESET_B(net104),
    .Q(\sound3.sdiv.Q[2] ));
 sky130_fd_sc_hd__dfrtp_2 _8242_ (.CLK(net143),
    .D(_0342_),
    .RESET_B(net104),
    .Q(\sound3.sdiv.Q[3] ));
 sky130_fd_sc_hd__dfrtp_1 _8243_ (.CLK(net141),
    .D(_0343_),
    .RESET_B(net102),
    .Q(\sound3.sdiv.Q[4] ));
 sky130_fd_sc_hd__dfrtp_2 _8244_ (.CLK(net141),
    .D(_0344_),
    .RESET_B(net102),
    .Q(\sound3.sdiv.Q[5] ));
 sky130_fd_sc_hd__dfrtp_2 _8245_ (.CLK(net141),
    .D(_0345_),
    .RESET_B(net102),
    .Q(\sound3.sdiv.Q[6] ));
 sky130_fd_sc_hd__dfrtp_1 _8246_ (.CLK(net141),
    .D(_0346_),
    .RESET_B(net102),
    .Q(\sound3.sdiv.Q[7] ));
 sky130_fd_sc_hd__dfrtp_1 _8247_ (.CLK(net141),
    .D(_0347_),
    .RESET_B(net102),
    .Q(\sound3.sdiv.Q[8] ));
 sky130_fd_sc_hd__dfrtp_1 _8248_ (.CLK(net135),
    .D(_0348_),
    .RESET_B(net96),
    .Q(\sound3.sdiv.Q[9] ));
 sky130_fd_sc_hd__dfrtp_1 _8249_ (.CLK(net135),
    .D(_0349_),
    .RESET_B(net96),
    .Q(\sound3.sdiv.Q[10] ));
 sky130_fd_sc_hd__dfrtp_1 _8250_ (.CLK(net129),
    .D(_0350_),
    .RESET_B(net90),
    .Q(\sound3.sdiv.Q[11] ));
 sky130_fd_sc_hd__dfrtp_1 _8251_ (.CLK(net132),
    .D(_0351_),
    .RESET_B(net93),
    .Q(\sound3.sdiv.Q[12] ));
 sky130_fd_sc_hd__dfrtp_1 _8252_ (.CLK(net132),
    .D(_0352_),
    .RESET_B(net93),
    .Q(\sound3.sdiv.Q[13] ));
 sky130_fd_sc_hd__dfrtp_1 _8253_ (.CLK(net131),
    .D(_0353_),
    .RESET_B(net92),
    .Q(\sound3.sdiv.Q[14] ));
 sky130_fd_sc_hd__dfrtp_1 _8254_ (.CLK(net131),
    .D(_0354_),
    .RESET_B(net92),
    .Q(\sound3.sdiv.Q[15] ));
 sky130_fd_sc_hd__dfrtp_1 _8255_ (.CLK(net131),
    .D(_0355_),
    .RESET_B(net92),
    .Q(\sound3.sdiv.Q[16] ));
 sky130_fd_sc_hd__dfrtp_1 _8256_ (.CLK(net131),
    .D(_0356_),
    .RESET_B(net92),
    .Q(\sound3.sdiv.Q[17] ));
 sky130_fd_sc_hd__dfrtp_1 _8257_ (.CLK(net132),
    .D(_0357_),
    .RESET_B(net93),
    .Q(\sound3.sdiv.Q[18] ));
 sky130_fd_sc_hd__dfrtp_1 _8258_ (.CLK(net132),
    .D(_0358_),
    .RESET_B(net93),
    .Q(\sound3.sdiv.Q[19] ));
 sky130_fd_sc_hd__dfrtp_1 _8259_ (.CLK(net132),
    .D(_0359_),
    .RESET_B(net93),
    .Q(\sound3.sdiv.Q[20] ));
 sky130_fd_sc_hd__dfrtp_1 _8260_ (.CLK(net132),
    .D(_0360_),
    .RESET_B(net93),
    .Q(\sound3.sdiv.Q[21] ));
 sky130_fd_sc_hd__dfrtp_1 _8261_ (.CLK(net140),
    .D(_0361_),
    .RESET_B(net101),
    .Q(\sound3.sdiv.Q[22] ));
 sky130_fd_sc_hd__dfrtp_1 _8262_ (.CLK(net140),
    .D(_0362_),
    .RESET_B(net101),
    .Q(\sound3.sdiv.Q[23] ));
 sky130_fd_sc_hd__dfrtp_1 _8263_ (.CLK(net140),
    .D(_0363_),
    .RESET_B(net101),
    .Q(\sound3.sdiv.Q[24] ));
 sky130_fd_sc_hd__dfrtp_1 _8264_ (.CLK(net140),
    .D(_0364_),
    .RESET_B(net101),
    .Q(\sound3.sdiv.Q[25] ));
 sky130_fd_sc_hd__dfrtp_1 _8265_ (.CLK(net141),
    .D(_0365_),
    .RESET_B(net102),
    .Q(\sound3.sdiv.Q[26] ));
 sky130_fd_sc_hd__dfrtp_1 _8266_ (.CLK(net141),
    .D(_0366_),
    .RESET_B(net102),
    .Q(\sound3.sdiv.Q[27] ));
 sky130_fd_sc_hd__dfrtp_1 _8267_ (.CLK(net123),
    .D(_0367_),
    .RESET_B(net84),
    .Q(\sound4.count_m[0] ));
 sky130_fd_sc_hd__dfrtp_1 _8268_ (.CLK(net123),
    .D(_0368_),
    .RESET_B(net84),
    .Q(\sound4.count_m[1] ));
 sky130_fd_sc_hd__dfrtp_1 _8269_ (.CLK(net123),
    .D(_0369_),
    .RESET_B(net84),
    .Q(\sound4.count_m[2] ));
 sky130_fd_sc_hd__dfrtp_1 _8270_ (.CLK(net123),
    .D(_0370_),
    .RESET_B(net84),
    .Q(\sound4.count_m[3] ));
 sky130_fd_sc_hd__dfrtp_1 _8271_ (.CLK(net123),
    .D(_0371_),
    .RESET_B(net84),
    .Q(\sound4.count_m[4] ));
 sky130_fd_sc_hd__dfrtp_1 _8272_ (.CLK(net123),
    .D(_0372_),
    .RESET_B(net84),
    .Q(\sound4.count_m[5] ));
 sky130_fd_sc_hd__dfrtp_1 _8273_ (.CLK(net122),
    .D(_0373_),
    .RESET_B(net83),
    .Q(\sound4.count_m[6] ));
 sky130_fd_sc_hd__dfrtp_1 _8274_ (.CLK(net122),
    .D(_0374_),
    .RESET_B(net83),
    .Q(\sound4.count_m[7] ));
 sky130_fd_sc_hd__dfrtp_1 _8275_ (.CLK(net120),
    .D(_0375_),
    .RESET_B(net81),
    .Q(\sound4.count_m[8] ));
 sky130_fd_sc_hd__dfrtp_1 _8276_ (.CLK(net122),
    .D(_0376_),
    .RESET_B(net83),
    .Q(\sound4.count_m[9] ));
 sky130_fd_sc_hd__dfrtp_1 _8277_ (.CLK(net118),
    .D(_0377_),
    .RESET_B(net79),
    .Q(\sound4.count_m[10] ));
 sky130_fd_sc_hd__dfrtp_1 _8278_ (.CLK(net118),
    .D(_0378_),
    .RESET_B(net79),
    .Q(\sound4.count_m[11] ));
 sky130_fd_sc_hd__dfrtp_1 _8279_ (.CLK(net122),
    .D(_0379_),
    .RESET_B(net83),
    .Q(\sound4.count_m[12] ));
 sky130_fd_sc_hd__dfrtp_1 _8280_ (.CLK(net122),
    .D(_0380_),
    .RESET_B(net83),
    .Q(\sound4.count_m[13] ));
 sky130_fd_sc_hd__dfrtp_1 _8281_ (.CLK(net122),
    .D(_0381_),
    .RESET_B(net83),
    .Q(\sound4.count_m[14] ));
 sky130_fd_sc_hd__dfrtp_1 _8282_ (.CLK(net122),
    .D(_0382_),
    .RESET_B(net83),
    .Q(\sound4.count_m[15] ));
 sky130_fd_sc_hd__dfrtp_1 _8283_ (.CLK(net123),
    .D(_0383_),
    .RESET_B(net84),
    .Q(\sound4.count_m[16] ));
 sky130_fd_sc_hd__dfrtp_1 _8284_ (.CLK(net123),
    .D(_0384_),
    .RESET_B(net84),
    .Q(\sound4.count_m[17] ));
 sky130_fd_sc_hd__dfrtp_1 _8285_ (.CLK(net123),
    .D(_0385_),
    .RESET_B(net84),
    .Q(\sound4.count_m[18] ));
 sky130_fd_sc_hd__dfrtp_4 _8286_ (.CLK(net121),
    .D(_0386_),
    .RESET_B(net82),
    .Q(\sound4.divisor_m[0] ));
 sky130_fd_sc_hd__dfrtp_4 _8287_ (.CLK(net123),
    .D(_0387_),
    .RESET_B(net84),
    .Q(\sound4.divisor_m[1] ));
 sky130_fd_sc_hd__dfrtp_4 _8288_ (.CLK(net121),
    .D(_0388_),
    .RESET_B(net82),
    .Q(\sound4.divisor_m[2] ));
 sky130_fd_sc_hd__dfrtp_2 _8289_ (.CLK(net121),
    .D(_0389_),
    .RESET_B(net82),
    .Q(\sound4.divisor_m[3] ));
 sky130_fd_sc_hd__dfrtp_4 _8290_ (.CLK(net121),
    .D(_0390_),
    .RESET_B(net82),
    .Q(\sound4.divisor_m[4] ));
 sky130_fd_sc_hd__dfrtp_2 _8291_ (.CLK(net123),
    .D(_0391_),
    .RESET_B(net84),
    .Q(\sound4.divisor_m[5] ));
 sky130_fd_sc_hd__dfrtp_2 _8292_ (.CLK(net121),
    .D(_0392_),
    .RESET_B(net82),
    .Q(\sound4.divisor_m[6] ));
 sky130_fd_sc_hd__dfrtp_2 _8293_ (.CLK(net122),
    .D(_0393_),
    .RESET_B(net83),
    .Q(\sound4.divisor_m[7] ));
 sky130_fd_sc_hd__dfrtp_1 _8294_ (.CLK(net123),
    .D(_0394_),
    .RESET_B(net84),
    .Q(\sound4.divisor_m[8] ));
 sky130_fd_sc_hd__dfrtp_2 _8295_ (.CLK(net122),
    .D(_0395_),
    .RESET_B(net83),
    .Q(\sound4.divisor_m[9] ));
 sky130_fd_sc_hd__dfrtp_4 _8296_ (.CLK(net122),
    .D(_0396_),
    .RESET_B(net83),
    .Q(\sound4.divisor_m[10] ));
 sky130_fd_sc_hd__dfrtp_1 _8297_ (.CLK(net118),
    .D(_0397_),
    .RESET_B(net79),
    .Q(\sound4.divisor_m[11] ));
 sky130_fd_sc_hd__dfrtp_2 _8298_ (.CLK(net118),
    .D(_0398_),
    .RESET_B(net79),
    .Q(\sound4.divisor_m[12] ));
 sky130_fd_sc_hd__dfrtp_4 _8299_ (.CLK(net122),
    .D(_0399_),
    .RESET_B(net83),
    .Q(\sound4.divisor_m[13] ));
 sky130_fd_sc_hd__dfrtp_2 _8300_ (.CLK(net122),
    .D(_0400_),
    .RESET_B(net83),
    .Q(\sound4.divisor_m[14] ));
 sky130_fd_sc_hd__dfrtp_2 _8301_ (.CLK(net122),
    .D(_0401_),
    .RESET_B(net83),
    .Q(\sound4.divisor_m[15] ));
 sky130_fd_sc_hd__dfrtp_2 _8302_ (.CLK(net122),
    .D(_0402_),
    .RESET_B(net83),
    .Q(\sound4.divisor_m[16] ));
 sky130_fd_sc_hd__dfrtp_4 _8303_ (.CLK(net121),
    .D(_0403_),
    .RESET_B(net82),
    .Q(\sound4.divisor_m[17] ));
 sky130_fd_sc_hd__dfrtp_4 _8304_ (.CLK(net121),
    .D(_0404_),
    .RESET_B(net82),
    .Q(\sound4.divisor_m[18] ));
 sky130_fd_sc_hd__dfrtp_1 _8305_ (.CLK(net137),
    .D(_0405_),
    .RESET_B(net98),
    .Q(\sound4.sdiv.A[0] ));
 sky130_fd_sc_hd__dfrtp_1 _8306_ (.CLK(net138),
    .D(_0406_),
    .RESET_B(net99),
    .Q(\sound4.sdiv.A[1] ));
 sky130_fd_sc_hd__dfrtp_1 _8307_ (.CLK(net123),
    .D(_0407_),
    .RESET_B(net84),
    .Q(\sound4.sdiv.A[2] ));
 sky130_fd_sc_hd__dfrtp_1 _8308_ (.CLK(net123),
    .D(_0408_),
    .RESET_B(net84),
    .Q(\sound4.sdiv.A[3] ));
 sky130_fd_sc_hd__dfrtp_1 _8309_ (.CLK(net123),
    .D(_0409_),
    .RESET_B(net84),
    .Q(\sound4.sdiv.A[4] ));
 sky130_fd_sc_hd__dfrtp_1 _8310_ (.CLK(net123),
    .D(_0410_),
    .RESET_B(net84),
    .Q(\sound4.sdiv.A[5] ));
 sky130_fd_sc_hd__dfrtp_1 _8311_ (.CLK(net123),
    .D(_0411_),
    .RESET_B(net84),
    .Q(\sound4.sdiv.A[6] ));
 sky130_fd_sc_hd__dfrtp_1 _8312_ (.CLK(net123),
    .D(_0412_),
    .RESET_B(net84),
    .Q(\sound4.sdiv.A[7] ));
 sky130_fd_sc_hd__dfrtp_1 _8313_ (.CLK(net122),
    .D(_0413_),
    .RESET_B(net83),
    .Q(\sound4.sdiv.A[8] ));
 sky130_fd_sc_hd__dfrtp_1 _8314_ (.CLK(net124),
    .D(_0414_),
    .RESET_B(net85),
    .Q(\sound4.sdiv.A[9] ));
 sky130_fd_sc_hd__dfrtp_1 _8315_ (.CLK(net124),
    .D(_0415_),
    .RESET_B(net85),
    .Q(\sound4.sdiv.A[10] ));
 sky130_fd_sc_hd__dfrtp_1 _8316_ (.CLK(net118),
    .D(_0416_),
    .RESET_B(net79),
    .Q(\sound4.sdiv.A[11] ));
 sky130_fd_sc_hd__dfrtp_1 _8317_ (.CLK(net124),
    .D(_0417_),
    .RESET_B(net85),
    .Q(\sound4.sdiv.A[12] ));
 sky130_fd_sc_hd__dfrtp_1 _8318_ (.CLK(net124),
    .D(_0418_),
    .RESET_B(net85),
    .Q(\sound4.sdiv.A[13] ));
 sky130_fd_sc_hd__dfrtp_1 _8319_ (.CLK(net124),
    .D(_0419_),
    .RESET_B(net85),
    .Q(\sound4.sdiv.A[14] ));
 sky130_fd_sc_hd__dfrtp_1 _8320_ (.CLK(net124),
    .D(_0420_),
    .RESET_B(net85),
    .Q(\sound4.sdiv.A[15] ));
 sky130_fd_sc_hd__dfrtp_1 _8321_ (.CLK(net124),
    .D(_0421_),
    .RESET_B(net85),
    .Q(\sound4.sdiv.A[16] ));
 sky130_fd_sc_hd__dfrtp_1 _8322_ (.CLK(net123),
    .D(_0422_),
    .RESET_B(net84),
    .Q(\sound4.sdiv.A[17] ));
 sky130_fd_sc_hd__dfrtp_1 _8323_ (.CLK(net123),
    .D(_0423_),
    .RESET_B(net84),
    .Q(\sound4.sdiv.A[18] ));
 sky130_fd_sc_hd__dfrtp_4 _8324_ (.CLK(net124),
    .D(_0424_),
    .RESET_B(net85),
    .Q(\sound4.sdiv.A[19] ));
 sky130_fd_sc_hd__dfrtp_2 _8325_ (.CLK(net124),
    .D(_0425_),
    .RESET_B(net85),
    .Q(\sound4.sdiv.A[20] ));
 sky130_fd_sc_hd__dfrtp_2 _8326_ (.CLK(net138),
    .D(_0426_),
    .RESET_B(net99),
    .Q(\sound4.sdiv.A[21] ));
 sky130_fd_sc_hd__dfrtp_2 _8327_ (.CLK(net138),
    .D(_0427_),
    .RESET_B(net99),
    .Q(\sound4.sdiv.A[22] ));
 sky130_fd_sc_hd__dfrtp_1 _8328_ (.CLK(net138),
    .D(_0428_),
    .RESET_B(net99),
    .Q(\sound4.sdiv.A[23] ));
 sky130_fd_sc_hd__dfrtp_1 _8329_ (.CLK(net124),
    .D(_0429_),
    .RESET_B(net85),
    .Q(\sound4.sdiv.A[24] ));
 sky130_fd_sc_hd__dfrtp_1 _8330_ (.CLK(net124),
    .D(_0430_),
    .RESET_B(net85),
    .Q(\sound4.sdiv.A[25] ));
 sky130_fd_sc_hd__dfrtp_4 _8331_ (.CLK(net124),
    .D(_0431_),
    .RESET_B(net85),
    .Q(\sound4.sdiv.A[26] ));
 sky130_fd_sc_hd__dfrtp_1 _8332_ (.CLK(net138),
    .D(_0432_),
    .RESET_B(net99),
    .Q(\sound4.sdiv.C[0] ));
 sky130_fd_sc_hd__dfrtp_1 _8333_ (.CLK(net138),
    .D(_0433_),
    .RESET_B(net99),
    .Q(\sound4.sdiv.C[1] ));
 sky130_fd_sc_hd__dfrtp_2 _8334_ (.CLK(net138),
    .D(_0434_),
    .RESET_B(net99),
    .Q(\sound4.sdiv.C[2] ));
 sky130_fd_sc_hd__dfrtp_2 _8335_ (.CLK(net137),
    .D(_0435_),
    .RESET_B(net98),
    .Q(\sound4.sdiv.C[3] ));
 sky130_fd_sc_hd__dfrtp_1 _8336_ (.CLK(net137),
    .D(_0436_),
    .RESET_B(net98),
    .Q(\sound4.sdiv.C[4] ));
 sky130_fd_sc_hd__dfrtp_1 _8337_ (.CLK(net138),
    .D(_0437_),
    .RESET_B(net99),
    .Q(\sound4.sdiv.C[5] ));
 sky130_fd_sc_hd__dfrtp_2 _8338_ (.CLK(net139),
    .D(_0438_),
    .RESET_B(net100),
    .Q(\wave_comb.u1.M[0] ));
 sky130_fd_sc_hd__dfrtp_2 _8339_ (.CLK(net138),
    .D(_0439_),
    .RESET_B(net99),
    .Q(\wave_comb.u1.M[1] ));
 sky130_fd_sc_hd__dfrtp_1 _8340_ (.CLK(net145),
    .D(_0440_),
    .RESET_B(net106),
    .Q(\wave_comb.u1.M[2] ));
 sky130_fd_sc_hd__dfrtp_1 _8341_ (.CLK(net138),
    .D(\sound4.sdiv.next_start ),
    .RESET_B(net99),
    .Q(\sound4.sdiv.start ));
 sky130_fd_sc_hd__dfstp_2 _8342_ (.CLK(net121),
    .D(\sound4.osc.next_count[0] ),
    .SET_B(net82),
    .Q(\sound4.count[0] ));
 sky130_fd_sc_hd__dfrtp_4 _8343_ (.CLK(net121),
    .D(\sound4.osc.next_count[1] ),
    .RESET_B(net82),
    .Q(\sound4.count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _8344_ (.CLK(net121),
    .D(\sound4.osc.next_count[2] ),
    .RESET_B(net82),
    .Q(\sound4.count[2] ));
 sky130_fd_sc_hd__dfrtp_2 _8345_ (.CLK(net121),
    .D(\sound4.osc.next_count[3] ),
    .RESET_B(net82),
    .Q(\sound4.count[3] ));
 sky130_fd_sc_hd__dfrtp_2 _8346_ (.CLK(net120),
    .D(\sound4.osc.next_count[4] ),
    .RESET_B(net81),
    .Q(\sound4.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _8347_ (.CLK(net121),
    .D(\sound4.osc.next_count[5] ),
    .RESET_B(net82),
    .Q(\sound4.count[5] ));
 sky130_fd_sc_hd__dfrtp_2 _8348_ (.CLK(net120),
    .D(\sound4.osc.next_count[6] ),
    .RESET_B(net81),
    .Q(\sound4.count[6] ));
 sky130_fd_sc_hd__dfrtp_2 _8349_ (.CLK(net120),
    .D(\sound4.osc.next_count[7] ),
    .RESET_B(net81),
    .Q(\sound4.count[7] ));
 sky130_fd_sc_hd__dfrtp_1 _8350_ (.CLK(net120),
    .D(\sound4.osc.next_count[8] ),
    .RESET_B(net81),
    .Q(\sound4.count[8] ));
 sky130_fd_sc_hd__dfrtp_2 _8351_ (.CLK(net120),
    .D(\sound4.osc.next_count[9] ),
    .RESET_B(net81),
    .Q(\sound4.count[9] ));
 sky130_fd_sc_hd__dfrtp_2 _8352_ (.CLK(net119),
    .D(\sound4.osc.next_count[10] ),
    .RESET_B(net80),
    .Q(\sound4.count[10] ));
 sky130_fd_sc_hd__dfrtp_2 _8353_ (.CLK(net119),
    .D(\sound4.osc.next_count[11] ),
    .RESET_B(net80),
    .Q(\sound4.count[11] ));
 sky130_fd_sc_hd__dfrtp_2 _8354_ (.CLK(net120),
    .D(\sound4.osc.next_count[12] ),
    .RESET_B(net81),
    .Q(\sound4.count[12] ));
 sky130_fd_sc_hd__dfrtp_2 _8355_ (.CLK(net120),
    .D(\sound4.osc.next_count[13] ),
    .RESET_B(net81),
    .Q(\sound4.count[13] ));
 sky130_fd_sc_hd__dfrtp_1 _8356_ (.CLK(net120),
    .D(\sound4.osc.next_count[14] ),
    .RESET_B(net81),
    .Q(\sound4.count[14] ));
 sky130_fd_sc_hd__dfrtp_2 _8357_ (.CLK(net121),
    .D(\sound4.osc.next_count[15] ),
    .RESET_B(net82),
    .Q(\sound4.count[15] ));
 sky130_fd_sc_hd__dfrtp_4 _8358_ (.CLK(net136),
    .D(\sound4.osc.next_count[16] ),
    .RESET_B(net97),
    .Q(\sound4.count[16] ));
 sky130_fd_sc_hd__dfrtp_4 _8359_ (.CLK(net136),
    .D(\sound4.osc.next_count[17] ),
    .RESET_B(net97),
    .Q(\sound4.count[17] ));
 sky130_fd_sc_hd__dfrtp_1 _8360_ (.CLK(net136),
    .D(\sound4.osc.next_count[18] ),
    .RESET_B(net97),
    .Q(\sound4.count[18] ));
 sky130_fd_sc_hd__dfrtp_1 _8361_ (.CLK(net145),
    .D(\wave.next_state[0] ),
    .RESET_B(net106),
    .Q(\wave.mode[0] ));
 sky130_fd_sc_hd__dfrtp_2 _8362_ (.CLK(net145),
    .D(\wave.next_state[1] ),
    .RESET_B(net106),
    .Q(\wave.mode[1] ));
 sky130_fd_sc_hd__dfrtp_1 _8363_ (.CLK(net118),
    .D(\rate_clk.next_count[0] ),
    .RESET_B(net79),
    .Q(\rate_clk.count[0] ));
 sky130_fd_sc_hd__dfrtp_1 _8364_ (.CLK(net118),
    .D(\rate_clk.next_count[1] ),
    .RESET_B(net79),
    .Q(\rate_clk.count[1] ));
 sky130_fd_sc_hd__dfrtp_1 _8365_ (.CLK(net118),
    .D(\rate_clk.next_count[2] ),
    .RESET_B(net79),
    .Q(\rate_clk.count[2] ));
 sky130_fd_sc_hd__dfrtp_1 _8366_ (.CLK(net119),
    .D(\rate_clk.next_count[3] ),
    .RESET_B(net80),
    .Q(\rate_clk.count[3] ));
 sky130_fd_sc_hd__dfrtp_1 _8367_ (.CLK(net119),
    .D(\rate_clk.next_count[4] ),
    .RESET_B(net80),
    .Q(\rate_clk.count[4] ));
 sky130_fd_sc_hd__dfrtp_1 _8368_ (.CLK(net119),
    .D(\rate_clk.next_count[5] ),
    .RESET_B(net80),
    .Q(\rate_clk.count[5] ));
 sky130_fd_sc_hd__dfrtp_1 _8369_ (.CLK(net119),
    .D(\rate_clk.next_count[6] ),
    .RESET_B(net80),
    .Q(\rate_clk.count[6] ));
 sky130_fd_sc_hd__dfrtp_4 _8370_ (.CLK(net119),
    .D(\rate_clk.next_count[7] ),
    .RESET_B(net80),
    .Q(\rate_clk.count[7] ));
 sky130_fd_sc_hd__dfrtp_1 _8371_ (.CLK(net144),
    .D(\wave_comb.u1.next_dived ),
    .RESET_B(net105),
    .Q(\wave_comb.u1.dived ));
 sky130_fd_sc_hd__buf_8 fanout100 (.A(net106),
    .X(net100));
 sky130_fd_sc_hd__buf_8 fanout101 (.A(net106),
    .X(net101));
 sky130_fd_sc_hd__clkbuf_4 fanout102 (.A(net106),
    .X(net102));
 sky130_fd_sc_hd__buf_8 fanout103 (.A(net106),
    .X(net103));
 sky130_fd_sc_hd__buf_6 fanout104 (.A(net105),
    .X(net104));
 sky130_fd_sc_hd__buf_8 fanout105 (.A(net106),
    .X(net105));
 sky130_fd_sc_hd__buf_8 fanout106 (.A(net3),
    .X(net106));
 sky130_fd_sc_hd__buf_4 fanout107 (.A(net115),
    .X(net107));
 sky130_fd_sc_hd__buf_4 fanout108 (.A(net115),
    .X(net108));
 sky130_fd_sc_hd__buf_4 fanout109 (.A(net110),
    .X(net109));
 sky130_fd_sc_hd__buf_4 fanout110 (.A(net115),
    .X(net110));
 sky130_fd_sc_hd__buf_4 fanout111 (.A(net115),
    .X(net111));
 sky130_fd_sc_hd__clkbuf_4 fanout112 (.A(net115),
    .X(net112));
 sky130_fd_sc_hd__buf_4 fanout113 (.A(net114),
    .X(net113));
 sky130_fd_sc_hd__buf_4 fanout114 (.A(net115),
    .X(net114));
 sky130_fd_sc_hd__clkbuf_4 fanout115 (.A(net2),
    .X(net115));
 sky130_fd_sc_hd__buf_4 fanout116 (.A(net119),
    .X(net116));
 sky130_fd_sc_hd__buf_4 fanout117 (.A(net119),
    .X(net117));
 sky130_fd_sc_hd__clkbuf_8 fanout118 (.A(net119),
    .X(net118));
 sky130_fd_sc_hd__buf_4 fanout119 (.A(net2),
    .X(net119));
 sky130_fd_sc_hd__buf_4 fanout120 (.A(net2),
    .X(net120));
 sky130_fd_sc_hd__clkbuf_4 fanout121 (.A(net2),
    .X(net121));
 sky130_fd_sc_hd__buf_4 fanout122 (.A(net124),
    .X(net122));
 sky130_fd_sc_hd__clkbuf_8 fanout123 (.A(net124),
    .X(net123));
 sky130_fd_sc_hd__buf_4 fanout124 (.A(net2),
    .X(net124));
 sky130_fd_sc_hd__buf_4 fanout125 (.A(net134),
    .X(net125));
 sky130_fd_sc_hd__buf_4 fanout126 (.A(net134),
    .X(net126));
 sky130_fd_sc_hd__buf_4 fanout127 (.A(net134),
    .X(net127));
 sky130_fd_sc_hd__buf_4 fanout128 (.A(net129),
    .X(net128));
 sky130_fd_sc_hd__clkbuf_4 fanout129 (.A(net134),
    .X(net129));
 sky130_fd_sc_hd__clkbuf_8 fanout130 (.A(net134),
    .X(net130));
 sky130_fd_sc_hd__buf_4 fanout131 (.A(net133),
    .X(net131));
 sky130_fd_sc_hd__clkbuf_4 fanout132 (.A(net133),
    .X(net132));
 sky130_fd_sc_hd__clkbuf_4 fanout133 (.A(net134),
    .X(net133));
 sky130_fd_sc_hd__clkbuf_8 fanout134 (.A(net2),
    .X(net134));
 sky130_fd_sc_hd__buf_4 fanout135 (.A(net136),
    .X(net135));
 sky130_fd_sc_hd__buf_4 fanout136 (.A(net145),
    .X(net136));
 sky130_fd_sc_hd__buf_4 fanout137 (.A(net145),
    .X(net137));
 sky130_fd_sc_hd__buf_2 fanout138 (.A(net145),
    .X(net138));
 sky130_fd_sc_hd__buf_4 fanout139 (.A(net145),
    .X(net139));
 sky130_fd_sc_hd__buf_4 fanout140 (.A(net145),
    .X(net140));
 sky130_fd_sc_hd__buf_2 fanout141 (.A(net145),
    .X(net141));
 sky130_fd_sc_hd__buf_4 fanout142 (.A(net145),
    .X(net142));
 sky130_fd_sc_hd__buf_4 fanout143 (.A(net144),
    .X(net143));
 sky130_fd_sc_hd__clkbuf_8 fanout144 (.A(net145),
    .X(net144));
 sky130_fd_sc_hd__clkbuf_8 fanout145 (.A(net2),
    .X(net145));
 sky130_fd_sc_hd__buf_8 fanout68 (.A(net76),
    .X(net68));
 sky130_fd_sc_hd__buf_8 fanout69 (.A(net76),
    .X(net69));
 sky130_fd_sc_hd__buf_6 fanout70 (.A(net71),
    .X(net70));
 sky130_fd_sc_hd__buf_6 fanout71 (.A(net76),
    .X(net71));
 sky130_fd_sc_hd__buf_8 fanout72 (.A(net76),
    .X(net72));
 sky130_fd_sc_hd__buf_4 fanout73 (.A(net76),
    .X(net73));
 sky130_fd_sc_hd__buf_6 fanout74 (.A(net75),
    .X(net74));
 sky130_fd_sc_hd__buf_8 fanout75 (.A(net76),
    .X(net75));
 sky130_fd_sc_hd__buf_6 fanout76 (.A(net3),
    .X(net76));
 sky130_fd_sc_hd__buf_8 fanout77 (.A(net80),
    .X(net77));
 sky130_fd_sc_hd__buf_8 fanout78 (.A(net80),
    .X(net78));
 sky130_fd_sc_hd__buf_8 fanout79 (.A(net80),
    .X(net79));
 sky130_fd_sc_hd__buf_8 fanout80 (.A(net3),
    .X(net80));
 sky130_fd_sc_hd__buf_8 fanout81 (.A(net3),
    .X(net81));
 sky130_fd_sc_hd__clkbuf_8 fanout82 (.A(net3),
    .X(net82));
 sky130_fd_sc_hd__buf_8 fanout83 (.A(net85),
    .X(net83));
 sky130_fd_sc_hd__buf_8 fanout84 (.A(net85),
    .X(net84));
 sky130_fd_sc_hd__buf_6 fanout85 (.A(net3),
    .X(net85));
 sky130_fd_sc_hd__buf_8 fanout86 (.A(net95),
    .X(net86));
 sky130_fd_sc_hd__buf_6 fanout87 (.A(net95),
    .X(net87));
 sky130_fd_sc_hd__buf_6 fanout88 (.A(net95),
    .X(net88));
 sky130_fd_sc_hd__buf_6 fanout89 (.A(net90),
    .X(net89));
 sky130_fd_sc_hd__buf_4 fanout90 (.A(net95),
    .X(net90));
 sky130_fd_sc_hd__buf_8 fanout91 (.A(net95),
    .X(net91));
 sky130_fd_sc_hd__buf_8 fanout92 (.A(net94),
    .X(net92));
 sky130_fd_sc_hd__clkbuf_8 fanout93 (.A(net94),
    .X(net93));
 sky130_fd_sc_hd__clkbuf_8 fanout94 (.A(net95),
    .X(net94));
 sky130_fd_sc_hd__buf_8 fanout95 (.A(net3),
    .X(net95));
 sky130_fd_sc_hd__buf_6 fanout96 (.A(net97),
    .X(net96));
 sky130_fd_sc_hd__clkbuf_8 fanout97 (.A(net106),
    .X(net97));
 sky130_fd_sc_hd__buf_6 fanout98 (.A(net106),
    .X(net98));
 sky130_fd_sc_hd__buf_4 fanout99 (.A(net106),
    .X(net99));
 sky130_fd_sc_hd__buf_8 input1 (.A(cs),
    .X(net1));
 sky130_fd_sc_hd__clkbuf_1 input10 (.A(piano_keys[1]),
    .X(net10));
 sky130_fd_sc_hd__clkbuf_1 input11 (.A(piano_keys[2]),
    .X(net11));
 sky130_fd_sc_hd__clkbuf_1 input12 (.A(piano_keys[3]),
    .X(net12));
 sky130_fd_sc_hd__clkbuf_1 input13 (.A(piano_keys[4]),
    .X(net13));
 sky130_fd_sc_hd__clkbuf_1 input14 (.A(piano_keys[5]),
    .X(net14));
 sky130_fd_sc_hd__buf_1 input15 (.A(piano_keys[6]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_1 input16 (.A(piano_keys[7]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_1 input17 (.A(piano_keys[8]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_1 input18 (.A(piano_keys[9]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_1 input19 (.A(seq_play),
    .X(net19));
 sky130_fd_sc_hd__clkbuf_8 input2 (.A(hwclk),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_1 input20 (.A(seq_power),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(tempo_select),
    .X(net21));
 sky130_fd_sc_hd__buf_6 input3 (.A(n_rst),
    .X(net3));
 sky130_fd_sc_hd__clkbuf_1 input4 (.A(piano_keys[0]),
    .X(net4));
 sky130_fd_sc_hd__buf_1 input5 (.A(piano_keys[10]),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_1 input6 (.A(piano_keys[11]),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_1 input7 (.A(piano_keys[12]),
    .X(net7));
 sky130_fd_sc_hd__clkbuf_1 input8 (.A(piano_keys[13]),
    .X(net8));
 sky130_fd_sc_hd__clkbuf_1 input9 (.A(piano_keys[14]),
    .X(net9));
 sky130_fd_sc_hd__clkbuf_2 max_cap1 (.A(_0562_),
    .X(net147));
 sky130_fd_sc_hd__clkbuf_1 max_cap53 (.A(net54),
    .X(net53));
 sky130_fd_sc_hd__buf_2 max_cap56 (.A(_0542_),
    .X(net56));
 sky130_fd_sc_hd__buf_4 max_cap58 (.A(net35),
    .X(net58));
 sky130_fd_sc_hd__clkbuf_1 max_cap59 (.A(net60),
    .X(net59));
 sky130_fd_sc_hd__buf_8 max_cap63 (.A(_1040_),
    .X(net63));
 sky130_fd_sc_hd__buf_6 max_cap64 (.A(_0684_),
    .X(net64));
 sky130_fd_sc_hd__clkbuf_2 max_cap65 (.A(_0565_),
    .X(net65));
 sky130_fd_sc_hd__clkbuf_2 max_cap66 (.A(_0559_),
    .X(net66));
 sky130_fd_sc_hd__dlymetal6s2s_1 max_cap67 (.A(_0483_),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_4 output22 (.A(net22),
    .X(beat_led[0]));
 sky130_fd_sc_hd__clkbuf_4 output23 (.A(net23),
    .X(beat_led[1]));
 sky130_fd_sc_hd__clkbuf_4 output24 (.A(net24),
    .X(beat_led[2]));
 sky130_fd_sc_hd__clkbuf_4 output25 (.A(net25),
    .X(beat_led[3]));
 sky130_fd_sc_hd__buf_2 output26 (.A(net26),
    .X(beat_led[4]));
 sky130_fd_sc_hd__clkbuf_4 output27 (.A(net27),
    .X(beat_led[5]));
 sky130_fd_sc_hd__clkbuf_4 output28 (.A(net28),
    .X(beat_led[6]));
 sky130_fd_sc_hd__clkbuf_4 output29 (.A(net29),
    .X(beat_led[7]));
 sky130_fd_sc_hd__buf_2 output30 (.A(net30),
    .X(mode_out[0]));
 sky130_fd_sc_hd__buf_2 output31 (.A(net31),
    .X(mode_out[1]));
 sky130_fd_sc_hd__clkbuf_4 output32 (.A(net32),
    .X(multi[0]));
 sky130_fd_sc_hd__clkbuf_4 output33 (.A(net33),
    .X(multi[1]));
 sky130_fd_sc_hd__buf_2 output34 (.A(net34),
    .X(multi[2]));
 sky130_fd_sc_hd__clkbuf_4 output35 (.A(net58),
    .X(note1[0]));
 sky130_fd_sc_hd__clkbuf_4 output36 (.A(net36),
    .X(note1[1]));
 sky130_fd_sc_hd__clkbuf_4 output37 (.A(net37),
    .X(note1[2]));
 sky130_fd_sc_hd__clkbuf_4 output38 (.A(net38),
    .X(note1[3]));
 sky130_fd_sc_hd__clkbuf_4 output39 (.A(net39),
    .X(note2[0]));
 sky130_fd_sc_hd__clkbuf_4 output40 (.A(net40),
    .X(note2[1]));
 sky130_fd_sc_hd__buf_2 output41 (.A(net41),
    .X(note2[2]));
 sky130_fd_sc_hd__clkbuf_4 output42 (.A(net42),
    .X(note2[3]));
 sky130_fd_sc_hd__clkbuf_4 output43 (.A(net43),
    .X(note3[0]));
 sky130_fd_sc_hd__clkbuf_4 output44 (.A(net44),
    .X(note3[1]));
 sky130_fd_sc_hd__buf_2 output45 (.A(net45),
    .X(note3[2]));
 sky130_fd_sc_hd__buf_2 output46 (.A(net46),
    .X(note3[3]));
 sky130_fd_sc_hd__buf_2 output47 (.A(net47),
    .X(note4[0]));
 sky130_fd_sc_hd__clkbuf_4 output48 (.A(net48),
    .X(note4[1]));
 sky130_fd_sc_hd__clkbuf_4 output49 (.A(net49),
    .X(note4[2]));
 sky130_fd_sc_hd__clkbuf_4 output50 (.A(net50),
    .X(note4[3]));
 sky130_fd_sc_hd__clkbuf_4 output51 (.A(net51),
    .X(pwm_o));
 sky130_fd_sc_hd__clkbuf_4 output52 (.A(net52),
    .X(seq_led_on));
 sky130_fd_sc_hd__conb_1 sass_synth_146 (.LO(net146));
 sky130_fd_sc_hd__buf_1 wire54 (.A(_2797_),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_1 wire55 (.A(_3086_),
    .X(net55));
 sky130_fd_sc_hd__buf_1 wire57 (.A(_0537_),
    .X(net57));
 sky130_fd_sc_hd__clkbuf_1 wire60 (.A(_2541_),
    .X(net60));
 sky130_fd_sc_hd__clkbuf_1 wire61 (.A(net62),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_1 wire62 (.A(_2344_),
    .X(net62));
 assign multi[3] = net146;
endmodule

