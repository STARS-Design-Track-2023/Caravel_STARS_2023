* NGSPICE file created from top_asic.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_1 abstract view
.subckt sky130_fd_sc_hd__a311oi_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkdlybuf4s25_1 abstract view
.subckt sky130_fd_sc_hd__clkdlybuf4s25_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_4 abstract view
.subckt sky130_fd_sc_hd__inv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_2 abstract view
.subckt sky130_fd_sc_hd__nand4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_1 abstract view
.subckt sky130_fd_sc_hd__a221oi_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_1 abstract view
.subckt sky130_fd_sc_hd__nand2b_1 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_6 abstract view
.subckt sky130_fd_sc_hd__inv_6 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32oi_1 abstract view
.subckt sky130_fd_sc_hd__a32oi_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_1 abstract view
.subckt sky130_fd_sc_hd__nor2b_1 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

.subckt top_asic clk mode_out[0] mode_out[1] pb[0] pb[10] pb[11] pb[12] pb[13] pb[14]
+ pb[1] pb[2] pb[3] pb[4] pb[5] pb[6] pb[7] pb[8] pb[9] reset sigout vccd1 vssd1
XANTENNA__09523__A2 _04048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06883_ genblk1\[6\].osc.clkdiv_C.cnt\[11\] _01484_ _01728_ _01734_ _01736_ vssd1
+ vssd1 vccd1 vccd1 _01737_ sky130_fd_sc_hd__a2111o_1
X_09671_ _00006_ _04151_ net1174 vssd1 vssd1 vccd1 vccd1 _04153_ sky130_fd_sc_hd__a21oi_1
X_08622_ _03251_ _03308_ _03327_ vssd1 vssd1 vccd1 vccd1 _03329_ sky130_fd_sc_hd__nor3_1
X_08553_ genblk2\[6\].wave_shpr.div.fin_quo\[0\] genblk2\[6\].wave_shpr.div.fin_quo\[1\]
+ _02734_ _02261_ vssd1 vssd1 vccd1 vccd1 _03260_ sky130_fd_sc_hd__a31o_1
XANTENNA_fanout162_A net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07504_ net18 net17 vssd1 vssd1 vccd1 vccd1 _02225_ sky130_fd_sc_hd__nor2b_2
XANTENNA__11094__A1 _05055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08484_ _03188_ _03189_ _03190_ _02885_ vssd1 vssd1 vccd1 vccd1 _03191_ sky130_fd_sc_hd__a31o_1
XFILLER_0_92_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07435_ _02173_ vssd1 vssd1 vccd1 vccd1 _00011_ sky130_fd_sc_hd__buf_1
XFILLER_0_9_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11789__B genblk1\[9\].osc.clkdiv_C.cnt\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07366_ _02091_ _02120_ _02121_ vssd1 vssd1 vccd1 vccd1 _02122_ sky130_fd_sc_hd__and3_1
X_09105_ genblk2\[0\].wave_shpr.div.acc\[10\] genblk2\[0\].wave_shpr.div.b1\[10\]
+ vssd1 vssd1 vccd1 vccd1 _03753_ sky130_fd_sc_hd__or2b_1
XFILLER_0_73_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06317_ genblk1\[0\].osc.clkdiv_C.cnt\[3\] _01274_ vssd1 vssd1 vccd1 vccd1 _01276_
+ sky130_fd_sc_hd__and2_1
XANTENNA__10185__S _04507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07297_ _02062_ vssd1 vssd1 vccd1 vccd1 genblk1\[10\].osc.clkdiv_C.next_cnt\[16\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09036_ _03702_ _01432_ vssd1 vssd1 vccd1 vccd1 _03705_ sky130_fd_sc_hd__nand2_8
XFILLER_0_130_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06248_ _01209_ vssd1 vssd1 vccd1 vccd1 _01210_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_115_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold340 genblk2\[0\].wave_shpr.div.quo\[2\] vssd1 vssd1 vccd1 vccd1 net558 sky130_fd_sc_hd__dlygate4sd3_1
X_06179_ net765 vssd1 vssd1 vccd1 vccd1 _01151_ sky130_fd_sc_hd__inv_2
XANTENNA__10913__S _04848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold351 genblk2\[0\].wave_shpr.div.quo\[10\] vssd1 vssd1 vccd1 vccd1 net569 sky130_fd_sc_hd__dlygate4sd3_1
Xhold362 genblk2\[2\].wave_shpr.div.acc\[18\] vssd1 vssd1 vccd1 vccd1 net580 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold373 genblk2\[4\].wave_shpr.div.acc\[19\] vssd1 vssd1 vccd1 vccd1 net591 sky130_fd_sc_hd__dlygate4sd3_1
Xhold384 genblk2\[4\].wave_shpr.div.quo\[11\] vssd1 vssd1 vccd1 vccd1 net602 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07222__B1 _02002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09275__A _03804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold395 genblk2\[7\].wave_shpr.div.quo\[14\] vssd1 vssd1 vccd1 vccd1 net613 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08610__C _02789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09938_ genblk2\[2\].wave_shpr.div.acc\[21\] _04342_ _04343_ vssd1 vssd1 vccd1 vccd1
+ _04344_ sky130_fd_sc_hd__a21bo_1
XANTENNA_fanout75_A net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09514__A2 _04043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09869_ genblk2\[2\].wave_shpr.div.acc\[4\] _04291_ _04214_ vssd1 vssd1 vccd1 vccd1
+ _04292_ sky130_fd_sc_hd__mux2_1
Xhold1040 genblk2\[6\].wave_shpr.div.b1\[6\] vssd1 vssd1 vccd1 vccd1 net1258 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1051 genblk1\[11\].osc.clkdiv_C.cnt\[10\] vssd1 vssd1 vccd1 vccd1 net1269 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1062 genblk2\[8\].wave_shpr.div.b1\[8\] vssd1 vssd1 vccd1 vccd1 net1280 sky130_fd_sc_hd__dlygate4sd3_1
X_11900_ genblk2\[0\].wave_shpr.div.i\[1\] genblk2\[0\].wave_shpr.div.i\[0\] genblk2\[0\].wave_shpr.div.i\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05725_ sky130_fd_sc_hd__a21o_1
Xhold1073 genblk2\[0\].wave_shpr.div.b1\[14\] vssd1 vssd1 vccd1 vccd1 net1291 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12880_ clknet_leaf_119_clk _00211_ net146 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.quo\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1084 genblk2\[10\].wave_shpr.div.b1\[17\] vssd1 vssd1 vccd1 vccd1 net1302 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1095 genblk2\[9\].wave_shpr.div.quo\[1\] vssd1 vssd1 vccd1 vccd1 net1313 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11831_ _05590_ _05562_ vssd1 vssd1 vccd1 vccd1 _05675_ sky130_fd_sc_hd__or2b_1
XTAP_2545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11762_ _05464_ genblk1\[9\].osc.clkdiv_C.cnt\[3\] vssd1 vssd1 vccd1 vccd1 _05630_
+ sky130_fd_sc_hd__and2_1
XTAP_1855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13501_ clknet_leaf_86_clk net230 net180 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.quo\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10713_ _02183_ vssd1 vssd1 vccd1 vccd1 _04886_ sky130_fd_sc_hd__clkbuf_4
XTAP_1877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11693_ _05565_ _05583_ _05584_ vssd1 vssd1 vccd1 vccd1 _05585_ sky130_fd_sc_hd__a21o_1
XFILLER_0_138_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13432_ clknet_leaf_82_clk _00751_ net201 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.acc\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12034__B1 _05816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_536 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10644_ _03704_ net747 _04647_ vssd1 vssd1 vccd1 vccd1 _00539_ sky130_fd_sc_hd__a21o_1
XANTENNA__07896__C _02365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_895 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10575_ _04769_ _04801_ _04802_ vssd1 vssd1 vccd1 vccd1 _04803_ sky130_fd_sc_hd__a21o_1
X_13363_ clknet_leaf_3_clk _00682_ net53 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.i\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09450__A1 genblk2\[1\].wave_shpr.div.quo\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12314_ _03942_ vssd1 vssd1 vccd1 vccd1 _06014_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_106_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13294_ clknet_leaf_87_clk _00615_ net179 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.b1\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_12245_ genblk2\[11\].wave_shpr.div.fin_quo\[0\] _05982_ _00005_ vssd1 vssd1 vccd1
+ vccd1 _05983_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10899__A1 _03687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12176_ genblk2\[10\].wave_shpr.div.i\[1\] genblk2\[10\].wave_shpr.div.i\[0\] vssd1
+ vssd1 vccd1 vccd1 _05918_ sky130_fd_sc_hd__nand2_1
X_11127_ _05181_ _05185_ _05186_ vssd1 vssd1 vccd1 vccd1 _05187_ sky130_fd_sc_hd__a21o_1
XANTENNA__07417__B _02153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11058_ _04967_ _05013_ vssd1 vssd1 vccd1 vccd1 _05133_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_3_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10009_ genblk2\[3\].wave_shpr.div.b1\[13\] genblk2\[3\].wave_shpr.div.acc\[13\]
+ vssd1 vssd1 vccd1 vccd1 _04405_ sky130_fd_sc_hd__and2b_1
XFILLER_0_64_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10520__B1 _04655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07220_ _01365_ _01189_ vssd1 vssd1 vccd1 vccd1 _02002_ sky130_fd_sc_hd__or2_4
XFILLER_0_116_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12025__B1 _05817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07151_ _01928_ net34 _01944_ _01945_ _01950_ vssd1 vssd1 vccd1 vccd1 _01951_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_42_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09079__B _01210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07082_ genblk1\[8\].osc.clkdiv_C.cnt\[5\] genblk1\[8\].osc.clkdiv_C.cnt\[4\] _01892_
+ vssd1 vssd1 vccd1 vccd1 _01895_ sky130_fd_sc_hd__and3_1
XANTENNA__06255__B2 genblk1\[0\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_42_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10339__B1 _03717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12193__B_N genblk2\[11\].wave_shpr.div.b1\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout105 net106 vssd1 vssd1 vccd1 vccd1 net105 sky130_fd_sc_hd__clkbuf_4
Xfanout116 net118 vssd1 vssd1 vccd1 vccd1 net116 sky130_fd_sc_hd__clkbuf_4
Xfanout127 net16 vssd1 vssd1 vccd1 vccd1 net127 sky130_fd_sc_hd__clkbuf_4
Xfanout138 net145 vssd1 vssd1 vccd1 vccd1 net138 sky130_fd_sc_hd__clkbuf_4
Xfanout149 net150 vssd1 vssd1 vccd1 vccd1 net149 sky130_fd_sc_hd__clkbuf_2
X_07984_ genblk2\[7\].wave_shpr.div.fin_quo\[6\] vssd1 vssd1 vccd1 vccd1 _02691_ sky130_fd_sc_hd__inv_2
XANTENNA__06231__B _01192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09723_ genblk2\[2\].wave_shpr.div.b1\[15\] genblk2\[2\].wave_shpr.div.acc\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04203_ sky130_fd_sc_hd__and2b_1
XANTENNA__09823__A _04069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06935_ net1180 _01775_ _01778_ vssd1 vssd1 vccd1 vccd1 genblk1\[6\].osc.clkdiv_C.next_cnt\[10\]
+ sky130_fd_sc_hd__o21a_1
XANTENNA__11303__A2 _05279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09654_ genblk2\[1\].wave_shpr.div.acc\[22\] _04139_ genblk2\[1\].wave_shpr.div.acc\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04142_ sky130_fd_sc_hd__o21bai_1
XANTENNA__09542__B genblk1\[1\].osc.clkdiv_C.cnt\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06866_ net1115 _01719_ _01722_ vssd1 vssd1 vccd1 vccd1 genblk1\[5\].osc.clkdiv_C.next_cnt\[15\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_96_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06885__C _01439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08605_ genblk2\[3\].wave_shpr.div.fin_quo\[2\] _02467_ vssd1 vssd1 vccd1 vccd1 _03312_
+ sky130_fd_sc_hd__nand2_1
X_06797_ genblk1\[5\].osc.clkdiv_C.cnt\[7\] vssd1 vssd1 vccd1 vccd1 _01669_ sky130_fd_sc_hd__inv_2
X_09585_ genblk2\[1\].wave_shpr.div.b1\[6\] genblk2\[1\].wave_shpr.div.acc\[6\] vssd1
+ vssd1 vccd1 vccd1 _04090_ sky130_fd_sc_hd__xor2_1
XFILLER_0_145_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08536_ _03240_ _03242_ vssd1 vssd1 vccd1 vccd1 _03243_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10814__A1 _04855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08467_ _03048_ _03049_ _03050_ vssd1 vssd1 vccd1 vccd1 _03174_ sky130_fd_sc_hd__a21oi_2
XANTENNA__07997__B _01360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07418_ _02160_ vssd1 vssd1 vccd1 vccd1 _00007_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08398_ genblk1\[2\].osc.clkdiv_C.cnt\[15\] _01349_ vssd1 vssd1 vccd1 vccd1 _03105_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_46_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_93_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07349_ genblk1\[11\].osc.clkdiv_C.cnt\[5\] genblk1\[11\].osc.clkdiv_C.cnt\[4\] _02101_
+ vssd1 vssd1 vccd1 vccd1 _02108_ sky130_fd_sc_hd__and3_1
X_10360_ _04648_ vssd1 vssd1 vccd1 vccd1 _00456_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06125__C _01096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11790__A2 _02203_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09019_ genblk2\[9\].wave_shpr.div.i\[1\] genblk2\[9\].wave_shpr.div.i\[0\] genblk2\[9\].wave_shpr.div.i\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03691_ sky130_fd_sc_hd__a21o_1
X_10291_ _04572_ _04601_ _04602_ vssd1 vssd1 vccd1 vccd1 _04603_ sky130_fd_sc_hd__a21o_1
X_12030_ genblk2\[10\].wave_shpr.div.quo\[8\] _05813_ _05817_ net320 vssd1 vssd1 vccd1
+ vccd1 _00957_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold170 _00388_ vssd1 vssd1 vccd1 vccd1 net388 sky130_fd_sc_hd__dlygate4sd3_1
Xhold181 PWM.counter\[7\] vssd1 vssd1 vccd1 vccd1 net399 sky130_fd_sc_hd__dlygate4sd3_1
Xhold192 genblk2\[0\].wave_shpr.div.quo\[17\] vssd1 vssd1 vccd1 vccd1 net410 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11542__A2 _05441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_31_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12932_ clknet_leaf_31_clk _00261_ net103 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.i\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12863_ clknet_leaf_129_clk _00194_ net66 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.b1\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_46_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11814_ _05582_ _05566_ vssd1 vssd1 vccd1 vccd1 _05662_ sky130_fd_sc_hd__or2b_1
XTAP_2364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12794_ clknet_leaf_93_clk _00127_ net148 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.quo\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11745_ net746 _05623_ _05624_ _05613_ vssd1 vssd1 vccd1 vccd1 _00865_ sky130_fd_sc_hd__a22o_1
XTAP_1674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08474__A2 _02308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11676_ genblk2\[9\].wave_shpr.div.acc\[4\] genblk2\[9\].wave_shpr.div.b1\[4\] vssd1
+ vssd1 vccd1 vccd1 _05568_ sky130_fd_sc_hd__or2b_1
XFILLER_0_154_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13415_ clknet_leaf_120_clk net488 net141 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.quo\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10627_ _04840_ vssd1 vssd1 vccd1 vccd1 _00531_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_104_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06237__A1 genblk1\[0\].osc.clkdiv_C.cnt\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13346_ clknet_leaf_6_clk _00667_ net49 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.acc\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10558_ _04780_ _04784_ _04785_ vssd1 vssd1 vccd1 vccd1 _04786_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13277_ clknet_leaf_12_clk _00598_ net54 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.i\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__12334__A _03689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10489_ _04614_ _04566_ vssd1 vssd1 vccd1 vccd1 _04732_ sky130_fd_sc_hd__nor2_1
X_12228_ _05930_ _05964_ _05965_ vssd1 vssd1 vccd1 vccd1 _05966_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_119_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07147__B _01946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12159_ genblk2\[10\].wave_shpr.div.acc\[21\] _05904_ vssd1 vssd1 vccd1 vccd1 _05907_
+ sky130_fd_sc_hd__xor2_1
X_06720_ _01600_ _01606_ _01607_ vssd1 vssd1 vccd1 vccd1 _01608_ sky130_fd_sc_hd__and3_1
XANTENNA__07163__A genblk1\[9\].osc.clkdiv_C.cnt\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06651_ net1193 _01543_ _01546_ vssd1 vssd1 vccd1 vccd1 genblk1\[3\].osc.clkdiv_C.next_cnt\[12\]
+ sky130_fd_sc_hd__o21a_1
X_09370_ net821 _03841_ _03839_ _03939_ vssd1 vssd1 vccd1 vccd1 _00175_ sky130_fd_sc_hd__a22o_1
X_06582_ _01489_ vssd1 vssd1 vccd1 vccd1 _01490_ sky130_fd_sc_hd__buf_8
XFILLER_0_59_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08321_ _02310_ _03027_ _02314_ vssd1 vssd1 vccd1 vccd1 _03028_ sky130_fd_sc_hd__o21a_1
XFILLER_0_129_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10728__S _04821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09662__A1 _04042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08252_ _02738_ vssd1 vssd1 vccd1 vccd1 _02959_ sky130_fd_sc_hd__inv_2
XFILLER_0_46_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07610__B _01211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07673__B1 _02013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06507__A _01200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07203_ genblk1\[9\].osc.clkdiv_C.cnt\[16\] _01985_ vssd1 vssd1 vccd1 vccd1 _01987_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_131_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08183_ _02850_ _02888_ _02889_ vssd1 vssd1 vccd1 vccd1 _02890_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_145_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_12_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_12_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA_fanout125_A net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07134_ genblk1\[9\].osc.clkdiv_C.cnt\[4\] _01311_ _01923_ genblk1\[9\].osc.clkdiv_C.cnt\[11\]
+ vssd1 vssd1 vccd1 vccd1 _01934_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__09818__A _04250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11559__S _05417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07065_ genblk1\[8\].osc.clkdiv_C.cnt\[0\] _01211_ _01882_ vssd1 vssd1 vccd1 vccd1
+ _01883_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_113_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07967_ genblk1\[7\].osc.clkdiv_C.cnt\[12\] _01214_ _02673_ vssd1 vssd1 vccd1 vccd1
+ _02674_ sky130_fd_sc_hd__a21bo_1
XANTENNA__06896__B _01439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09706_ _04167_ _04184_ _04185_ vssd1 vssd1 vccd1 vccd1 _04186_ sky130_fd_sc_hd__a21o_1
X_06918_ _01761_ _01767_ vssd1 vssd1 vccd1 vccd1 genblk1\[6\].osc.clkdiv_C.next_cnt\[4\]
+ sky130_fd_sc_hd__nor2_1
X_07898_ genblk1\[8\].osc.clkdiv_C.cnt\[14\] _01309_ _01576_ genblk1\[8\].osc.clkdiv_C.cnt\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02605_ sky130_fd_sc_hd__a2bb2o_1
X_09637_ _04006_ _04129_ vssd1 vssd1 vccd1 vccd1 _04130_ sky130_fd_sc_hd__or2_1
XFILLER_0_69_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06849_ _01693_ _01710_ _01711_ vssd1 vssd1 vccd1 vccd1 genblk1\[5\].osc.clkdiv_C.next_cnt\[9\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_97_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07900__A1 genblk1\[8\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09568_ _03974_ _03969_ vssd1 vssd1 vccd1 vccd1 _04077_ sky130_fd_sc_hd__or2b_1
XFILLER_0_78_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout38_A net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08519_ _02216_ _02552_ genblk2\[11\].wave_shpr.div.fin_quo\[0\] vssd1 vssd1 vccd1
+ vccd1 _03226_ sky130_fd_sc_hd__and3_1
X_09499_ _04040_ vssd1 vssd1 vccd1 vccd1 _00203_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_92_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11530_ _05450_ genblk1\[8\].osc.clkdiv_C.cnt\[9\] vssd1 vssd1 vccd1 vccd1 _05462_
+ sky130_fd_sc_hd__and2_1
XANTENNA__11460__A1 _01819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06417__A _01360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11461_ _05427_ vssd1 vssd1 vccd1 vccd1 _00778_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06136__B net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13200_ clknet_leaf_115_clk _00523_ net134 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.fin_quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10412_ _04672_ genblk1\[4\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 _04675_
+ sky130_fd_sc_hd__and2_1
X_11392_ genblk2\[8\].wave_shpr.div.acc\[7\] genblk2\[8\].wave_shpr.div.b1\[7\] vssd1
+ vssd1 vccd1 vccd1 _05368_ sky130_fd_sc_hd__or2b_1
XFILLER_0_61_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13131_ clknet_leaf_4_clk _00456_ net46 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.b1\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10343_ _04638_ vssd1 vssd1 vccd1 vccd1 _00449_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10274_ _04431_ genblk2\[4\].wave_shpr.div.acc\[1\] _04585_ vssd1 vssd1 vccd1 vccd1
+ _04586_ sky130_fd_sc_hd__a21o_1
X_13062_ clknet_leaf_29_clk net635 net95 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.quo\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11515__A2 _05448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07719__B2 genblk1\[1\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12013_ _03726_ _05810_ _03735_ vssd1 vssd1 vccd1 vccd1 _00947_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_136_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12915_ clknet_leaf_36_clk _00246_ net105 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.acc\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12846_ clknet_leaf_68_clk _00177_ net211 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.i\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07711__A net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12777_ clknet_leaf_43_clk _00110_ net124 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.b1\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_83_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11233__A _05245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11728_ genblk2\[9\].wave_shpr.div.fin_quo\[3\] genblk2\[9\].wave_shpr.div.quo\[2\]
+ _00023_ vssd1 vssd1 vccd1 vccd1 _05617_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11659_ _03690_ _05551_ _05552_ vssd1 vssd1 vccd1 vccd1 _00851_ sky130_fd_sc_hd__nor3_1
XFILLER_0_126_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11203__A1 _03726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold906 genblk2\[11\].wave_shpr.div.i\[1\] vssd1 vssd1 vccd1 vccd1 net1124 sky130_fd_sc_hd__dlygate4sd3_1
Xhold917 genblk2\[10\].wave_shpr.div.acc\[19\] vssd1 vssd1 vccd1 vccd1 net1135 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_386 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13329_ clknet_leaf_25_clk _00650_ net91 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.quo\[23\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold928 genblk1\[6\].osc.clkdiv_C.cnt\[13\] vssd1 vssd1 vccd1 vccd1 net1146 sky130_fd_sc_hd__dlygate4sd3_1
Xhold939 PWM.final_sample_in\[6\] vssd1 vssd1 vccd1 vccd1 net1157 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12064__A _03833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08870_ sig_norm.b1\[2\] vssd1 vssd1 vccd1 vccd1 _03576_ sky130_fd_sc_hd__inv_2
X_07821_ genblk2\[1\].wave_shpr.div.fin_quo\[4\] _02521_ _02523_ _02527_ vssd1 vssd1
+ vccd1 vccd1 _02528_ sky130_fd_sc_hd__a22o_1
XANTENNA__06394__B1 _01337_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07605__B net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07752_ genblk1\[1\].osc.clkdiv_C.cnt\[16\] _01577_ genblk1\[1\].osc.clkdiv_C.cnt\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02459_ sky130_fd_sc_hd__a21oi_4
X_06703_ genblk1\[4\].osc.clkdiv_C.cnt\[9\] _01592_ vssd1 vssd1 vccd1 vccd1 _01593_
+ sky130_fd_sc_hd__nand2_1
X_07683_ _01174_ genblk1\[10\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 _02390_
+ sky130_fd_sc_hd__nand2_1
X_09422_ genblk2\[1\].wave_shpr.div.b1\[8\] genblk2\[1\].wave_shpr.div.acc\[8\] vssd1
+ vssd1 vccd1 vccd1 _03986_ sky130_fd_sc_hd__and2b_1
X_06634_ genblk1\[3\].osc.clkdiv_C.cnt\[6\] _01533_ vssd1 vssd1 vccd1 vccd1 _01536_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09353_ net1175 _03903_ _03910_ _03928_ vssd1 vssd1 vccd1 vccd1 _00169_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06565_ _01451_ _01476_ vssd1 vssd1 vccd1 vccd1 _01477_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08304_ _02969_ _03003_ vssd1 vssd1 vccd1 vccd1 _03011_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11442__A1 _05417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_631 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09284_ genblk2\[0\].wave_shpr.div.acc\[3\] _03875_ _03804_ vssd1 vssd1 vccd1 vccd1
+ _03876_ sky130_fd_sc_hd__mux2_1
X_06496_ genblk1\[2\].osc.clkdiv_C.cnt\[14\] genblk1\[2\].osc.clkdiv_C.cnt\[1\] _01327_
+ vssd1 vssd1 vccd1 vccd1 _01422_ sky130_fd_sc_hd__and3_1
XFILLER_0_118_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08235_ _02592_ _02940_ _02941_ _02467_ genblk2\[3\].wave_shpr.div.fin_quo\[6\] vssd1
+ vssd1 vccd1 vccd1 _02942_ sky130_fd_sc_hd__a32o_1
XFILLER_0_15_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08166_ genblk1\[3\].osc.clkdiv_C.cnt\[8\] _01423_ vssd1 vssd1 vccd1 vccd1 _02873_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_43_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_43_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11745__A2 _05623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11289__S _05222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07117_ _01918_ vssd1 vssd1 vccd1 vccd1 genblk1\[8\].osc.clkdiv_C.next_cnt\[16\]
+ sky130_fd_sc_hd__clkbuf_1
X_08097_ _02800_ _02801_ _02802_ _02803_ vssd1 vssd1 vccd1 vccd1 _02804_ sky130_fd_sc_hd__or4b_1
XFILLER_0_101_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_868 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10953__B1 _05055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07048_ _01174_ _01182_ _01336_ vssd1 vssd1 vccd1 vccd1 _01866_ sky130_fd_sc_hd__a21oi_2
XANTENNA__09571__B1 _04047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08999_ _03679_ vssd1 vssd1 vccd1 vccd1 _00064_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10961_ net620 _05062_ _05064_ genblk2\[6\].wave_shpr.div.quo\[12\] _05065_ vssd1
+ vssd1 vccd1 vccd1 _00640_ sky130_fd_sc_hd__a221o_1
XFILLER_0_97_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12700_ clknet_leaf_89_clk genblk1\[8\].osc.clkdiv_C.next_cnt\[13\] net172 vssd1
+ vssd1 vccd1 vccd1 genblk1\[8\].osc.clkdiv_C.cnt\[13\] sky130_fd_sc_hd__dfrtp_2
X_13680_ clknet_leaf_63_clk _00993_ net190 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.acc\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10484__A2 _04715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10892_ genblk2\[6\].wave_shpr.div.fin_quo\[6\] genblk2\[6\].wave_shpr.div.quo\[5\]
+ _00017_ vssd1 vssd1 vccd1 vccd1 _05030_ sky130_fd_sc_hd__mux2_1
XANTENNA__07531__A _01155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12631_ clknet_leaf_18_clk genblk1\[4\].osc.clkdiv_C.next_cnt\[16\] net112 vssd1
+ vssd1 vccd1 vccd1 genblk1\[4\].osc.clkdiv_C.cnt\[16\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_155_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10236__A2 _04457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12562_ clknet_leaf_30_clk genblk1\[1\].osc.clkdiv_C.next_cnt\[1\] net96 vssd1 vssd1
+ vccd1 vccd1 genblk1\[1\].osc.clkdiv_C.cnt\[1\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__06147__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11513_ genblk2\[8\].wave_shpr.div.quo\[10\] _05448_ _05449_ net329 _05452_ vssd1
+ vssd1 vccd1 vccd1 _00805_ sky130_fd_sc_hd__a221o_1
X_12493_ clknet_leaf_107_clk _00055_ net152 vssd1 vssd1 vccd1 vccd1 sig_norm.quo\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11444_ genblk2\[8\].wave_shpr.div.fin_quo\[1\] net1331 _00021_ vssd1 vssd1 vccd1
+ vccd1 _05419_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11375_ _05353_ vssd1 vssd1 vccd1 vccd1 _05354_ sky130_fd_sc_hd__inv_2
XFILLER_0_150_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10944__B1 _05056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13114_ clknet_leaf_115_clk _00439_ net135 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.fin_quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10326_ genblk2\[4\].wave_shpr.div.fin_quo\[7\] net1263 _00013_ vssd1 vssd1 vccd1
+ vccd1 _04631_ sky130_fd_sc_hd__mux2_1
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13045_ clknet_leaf_128_clk _00372_ net67 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.b1\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10257_ genblk2\[4\].wave_shpr.div.acc\[13\] genblk2\[4\].wave_shpr.div.b1\[13\]
+ vssd1 vssd1 vccd1 vccd1 _04569_ sky130_fd_sc_hd__or2b_1
XFILLER_0_147_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10188_ _04403_ _04366_ vssd1 vssd1 vccd1 vccd1 _04519_ sky130_fd_sc_hd__or2b_1
XANTENNA__10132__A _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_47 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10475__A2 _04715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_807 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12829_ clknet_leaf_64_clk _00162_ net189 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.acc\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12059__A _03833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07160__B genblk1\[9\].osc.clkdiv_C.cnt\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06350_ _01268_ _01296_ vssd1 vssd1 vccd1 vccd1 _01297_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_286 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06281_ genblk1\[0\].osc.clkdiv_C.cnt\[16\] _01242_ vssd1 vssd1 vccd1 vccd1 _01243_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_4_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08020_ _02700_ _02702_ _02701_ _02726_ vssd1 vssd1 vccd1 vccd1 _02727_ sky130_fd_sc_hd__and4_1
XFILLER_0_115_848 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold703 genblk2\[6\].wave_shpr.div.acc\[14\] vssd1 vssd1 vccd1 vccd1 net921 sky130_fd_sc_hd__dlygate4sd3_1
Xhold714 genblk2\[8\].wave_shpr.div.acc\[6\] vssd1 vssd1 vccd1 vccd1 net932 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold725 _00413_ vssd1 vssd1 vccd1 vccd1 net943 sky130_fd_sc_hd__dlygate4sd3_1
Xhold736 genblk2\[10\].wave_shpr.div.acc\[8\] vssd1 vssd1 vccd1 vccd1 net954 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold747 genblk2\[1\].wave_shpr.div.acc\[3\] vssd1 vssd1 vccd1 vccd1 net965 sky130_fd_sc_hd__dlygate4sd3_1
Xhold758 genblk2\[3\].wave_shpr.div.acc\[2\] vssd1 vssd1 vccd1 vccd1 net976 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06377__A_N _01188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09971_ genblk2\[3\].wave_shpr.div.acc\[11\] genblk2\[3\].wave_shpr.div.b1\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04367_ sky130_fd_sc_hd__or2b_1
XFILLER_0_40_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold769 genblk2\[9\].wave_shpr.div.acc\[17\] vssd1 vssd1 vccd1 vccd1 net987 sky130_fd_sc_hd__dlygate4sd3_1
X_08922_ net678 _03588_ vssd1 vssd1 vccd1 vccd1 _03620_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09553__B1 _04046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08853_ _03501_ _03502_ _03500_ _03503_ vssd1 vssd1 vccd1 vccd1 _03560_ sky130_fd_sc_hd__a211o_1
XFILLER_0_34_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07804_ genblk2\[0\].wave_shpr.div.fin_quo\[0\] genblk2\[0\].wave_shpr.div.fin_quo\[1\]
+ genblk2\[0\].wave_shpr.div.fin_quo\[2\] vssd1 vssd1 vccd1 vccd1 _02511_ sky130_fd_sc_hd__or3_1
X_08784_ _03474_ _03479_ _03490_ vssd1 vssd1 vccd1 vccd1 _03491_ sky130_fd_sc_hd__a21o_1
XANTENNA__09831__A _04069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07735_ genblk1\[1\].osc.clkdiv_C.cnt\[5\] _02433_ _01305_ genblk1\[1\].osc.clkdiv_C.cnt\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02442_ sky130_fd_sc_hd__o22a_1
XANTENNA__09856__A1 _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11572__S _05417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09550__B genblk1\[1\].osc.clkdiv_C.cnt\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07666_ _02368_ _02372_ genblk1\[10\].osc.clkdiv_C.cnt\[7\] _01190_ vssd1 vssd1 vccd1
+ vccd1 _02373_ sky130_fd_sc_hd__a2bb2o_1
X_09405_ genblk2\[1\].wave_shpr.div.acc\[2\] genblk2\[1\].wave_shpr.div.b1\[2\] vssd1
+ vssd1 vccd1 vccd1 _03969_ sky130_fd_sc_hd__or2b_1
X_06617_ _01522_ vssd1 vssd1 vccd1 vccd1 _01524_ sky130_fd_sc_hd__inv_2
XFILLER_0_153_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07597_ _02265_ genblk2\[9\].wave_shpr.div.fin_quo\[5\] _02303_ vssd1 vssd1 vccd1
+ vccd1 _02304_ sky130_fd_sc_hd__or3b_1
XFILLER_0_48_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09336_ genblk2\[0\].wave_shpr.div.acc\[15\] _03915_ _03889_ vssd1 vssd1 vccd1 vccd1
+ _03916_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06548_ _01452_ _01464_ _01465_ vssd1 vssd1 vccd1 vccd1 genblk1\[2\].osc.clkdiv_C.next_cnt\[8\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_118_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10916__S _05042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09267_ _03838_ vssd1 vssd1 vccd1 vccd1 _03863_ sky130_fd_sc_hd__inv_2
X_06479_ genblk1\[1\].osc.clkdiv_C.cnt\[16\] _01405_ vssd1 vssd1 vccd1 vccd1 _01407_
+ sky130_fd_sc_hd__and2_1
X_08218_ _02900_ _02922_ vssd1 vssd1 vccd1 vccd1 _02925_ sky130_fd_sc_hd__and2b_1
XFILLER_0_133_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09198_ _02005_ vssd1 vssd1 vccd1 vccd1 _03827_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08149_ genblk1\[3\].osc.clkdiv_C.cnt\[2\] _01513_ vssd1 vssd1 vccd1 vccd1 _02856_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_120_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10926__B1 _04647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11160_ genblk2\[7\].wave_shpr.div.acc\[23\] genblk2\[7\].wave_shpr.div.acc\[25\]
+ genblk2\[7\].wave_shpr.div.acc\[24\] genblk2\[7\].wave_shpr.div.acc\[26\] vssd1
+ vssd1 vccd1 vccd1 _05220_ sky130_fd_sc_hd__or4_2
X_10111_ net634 _04461_ _04462_ genblk2\[3\].wave_shpr.div.quo\[13\] _04466_ vssd1
+ vssd1 vccd1 vccd1 _00389_ sky130_fd_sc_hd__a221o_1
X_11091_ _05155_ vssd1 vssd1 vccd1 vccd1 _00680_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_101_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10042_ _04430_ vssd1 vssd1 vccd1 vccd1 _00356_ sky130_fd_sc_hd__clkbuf_1
Xhold30 _00975_ vssd1 vssd1 vccd1 vccd1 net248 sky130_fd_sc_hd__dlygate4sd3_1
Xhold41 genblk2\[2\].wave_shpr.div.quo\[24\] vssd1 vssd1 vccd1 vccd1 net259 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 _00130_ vssd1 vssd1 vccd1 vccd1 net270 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold63 genblk2\[4\].wave_shpr.div.i\[4\] vssd1 vssd1 vccd1 vccd1 net281 sky130_fd_sc_hd__dlygate4sd3_1
Xhold74 genblk2\[1\].wave_shpr.div.quo\[6\] vssd1 vssd1 vccd1 vccd1 net292 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold85 _00721_ vssd1 vssd1 vccd1 vccd1 net303 sky130_fd_sc_hd__dlygate4sd3_1
Xhold96 _00647_ vssd1 vssd1 vccd1 vccd1 net314 sky130_fd_sc_hd__dlygate4sd3_1
X_11993_ _05801_ vssd1 vssd1 vccd1 vccd1 _00936_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13732_ clknet_leaf_45_clk _01043_ net121 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.quo\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10944_ genblk2\[6\].wave_shpr.div.quo\[5\] _05052_ _05056_ net720 vssd1 vssd1 vccd1
+ vccd1 _00632_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13663_ clknet_leaf_44_clk _00976_ net121 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.acc\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10875_ genblk2\[6\].wave_shpr.div.acc\[19\] _05018_ vssd1 vssd1 vccd1 vccd1 _05019_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_38_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12614_ clknet_leaf_23_clk genblk1\[3\].osc.clkdiv_C.next_cnt\[17\] net109 vssd1
+ vssd1 vccd1 vccd1 genblk1\[3\].osc.clkdiv_C.cnt\[17\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13594_ clknet_leaf_72_clk _00909_ net216 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.acc\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12545_ clknet_leaf_60_clk genblk1\[0\].osc.clkdiv_C.next_cnt\[2\] net187 vssd1 vssd1
+ vccd1 vccd1 genblk1\[0\].osc.clkdiv_C.cnt\[2\] sky130_fd_sc_hd__dfrtp_4
Xclkbuf_leaf_132_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_132_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__10090__B1 _04456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12476_ clknet_leaf_106_clk _00038_ net151 vssd1 vssd1 vccd1 vccd1 sig_norm.acc\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_5 _04242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11427_ _05361_ _05401_ _05402_ vssd1 vssd1 vccd1 vccd1 _05403_ sky130_fd_sc_hd__a21o_1
XFILLER_0_105_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09783__B1 _04241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11358_ genblk2\[7\].wave_shpr.div.acc\[23\] _05219_ vssd1 vssd1 vccd1 vccd1 _05342_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10309_ genblk2\[4\].wave_shpr.div.acc\[23\] _04620_ vssd1 vssd1 vccd1 vccd1 _04621_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11289_ genblk2\[7\].wave_shpr.div.acc\[5\] _05290_ _05222_ vssd1 vssd1 vccd1 vccd1
+ _05291_ sky130_fd_sc_hd__mux2_1
XANTENNA__12342__A _03689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13028_ clknet_leaf_113_clk _00355_ net131 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.fin_quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10696__A2 _02183_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08966__S _01155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07520_ _02230_ PWM.final_sample_in\[5\] PWM.final_sample_in\[4\] _01163_ _02239_
+ vssd1 vssd1 vccd1 vccd1 _02240_ sky130_fd_sc_hd__o221a_1
X_07451_ genblk2\[6\].wave_shpr.div.i\[2\] genblk2\[6\].wave_shpr.div.i\[3\] genblk2\[6\].wave_shpr.div.i\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02185_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_146_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06402_ genblk1\[1\].osc.clkdiv_C.cnt\[1\] _01340_ _01197_ _01341_ _01345_ vssd1
+ vssd1 vccd1 vccd1 _01346_ sky130_fd_sc_hd__a221o_1
X_07382_ _02091_ _02131_ _02133_ vssd1 vssd1 vccd1 vccd1 _02134_ sky130_fd_sc_hd__and3_1
X_09121_ genblk2\[0\].wave_shpr.div.b1\[3\] genblk2\[0\].wave_shpr.div.acc\[3\] vssd1
+ vssd1 vccd1 vccd1 _03769_ sky130_fd_sc_hd__and2b_1
X_06333_ genblk1\[0\].osc.clkdiv_C.cnt\[9\] _01284_ vssd1 vssd1 vccd1 vccd1 _01286_
+ sky130_fd_sc_hd__and2_1
XANTENNA__10736__S _04821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_123_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_123_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__08274__B1 _02525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06264_ _01225_ vssd1 vssd1 vccd1 vccd1 _01226_ sky130_fd_sc_hd__buf_6
X_09052_ _03689_ _01242_ vssd1 vssd1 vccd1 vccd1 _03716_ sky130_fd_sc_hd__nand2_2
XFILLER_0_44_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06515__A _01440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_621 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08003_ genblk1\[6\].osc.clkdiv_C.cnt\[12\] _01666_ _02709_ vssd1 vssd1 vccd1 vccd1
+ _02710_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_5_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06195_ net996 _01159_ vssd1 vssd1 vccd1 vccd1 _01162_ sky130_fd_sc_hd__nor2_1
Xhold500 genblk1\[1\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 net718 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold511 genblk2\[5\].wave_shpr.div.quo\[4\] vssd1 vssd1 vccd1 vccd1 net729 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold522 genblk2\[10\].wave_shpr.div.quo\[0\] vssd1 vssd1 vccd1 vccd1 net740 sky130_fd_sc_hd__buf_1
Xhold533 genblk2\[8\].wave_shpr.div.quo\[5\] vssd1 vssd1 vccd1 vccd1 net751 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold544 genblk2\[11\].wave_shpr.div.acc\[9\] vssd1 vssd1 vccd1 vccd1 net762 sky130_fd_sc_hd__dlygate4sd3_1
Xhold555 _00579_ vssd1 vssd1 vccd1 vccd1 net773 sky130_fd_sc_hd__dlygate4sd3_1
Xhold566 genblk2\[4\].wave_shpr.div.acc\[15\] vssd1 vssd1 vccd1 vccd1 net784 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold577 genblk2\[8\].wave_shpr.div.quo\[4\] vssd1 vssd1 vccd1 vccd1 net795 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold588 genblk2\[6\].wave_shpr.div.acc\[9\] vssd1 vssd1 vccd1 vccd1 net806 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09954_ genblk2\[2\].wave_shpr.div.i\[1\] genblk2\[2\].wave_shpr.div.i\[0\] vssd1
+ vssd1 vccd1 vccd1 _04354_ sky130_fd_sc_hd__nand2_1
Xhold599 genblk2\[9\].wave_shpr.div.i\[4\] vssd1 vssd1 vccd1 vccd1 net817 sky130_fd_sc_hd__dlygate4sd3_1
X_08905_ _03596_ _03607_ _02248_ vssd1 vssd1 vccd1 vccd1 _03608_ sky130_fd_sc_hd__a21oi_1
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09885_ _04188_ _04303_ vssd1 vssd1 vccd1 vccd1 _04304_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10136__A1 _03819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08836_ _02509_ _02572_ _02518_ vssd1 vssd1 vccd1 vccd1 _03543_ sky130_fd_sc_hd__o21ai_1
XTAP_2705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08767_ _02798_ _03466_ _03468_ _03473_ vssd1 vssd1 vccd1 vccd1 _03474_ sky130_fd_sc_hd__a31o_1
XTAP_2716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11636__A1 _05449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07718_ _01360_ _01302_ vssd1 vssd1 vccd1 vccd1 _02425_ sky130_fd_sc_hd__nand2_4
XTAP_2749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08698_ _03403_ _03357_ _03173_ _03402_ vssd1 vssd1 vccd1 vccd1 _03405_ sky130_fd_sc_hd__o211ai_4
XFILLER_0_67_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07649_ genblk2\[11\].wave_shpr.div.fin_quo\[5\] _02355_ vssd1 vssd1 vccd1 vccd1
+ _02356_ sky130_fd_sc_hd__nor2_1
X_10660_ net729 _04853_ _04857_ net745 vssd1 vssd1 vccd1 vccd1 _00547_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09319_ net889 _03870_ _03877_ _03902_ vssd1 vssd1 vccd1 vccd1 _00161_ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10591_ genblk2\[5\].wave_shpr.div.acc\[23\] genblk2\[5\].wave_shpr.div.acc\[25\]
+ genblk2\[5\].wave_shpr.div.acc\[24\] genblk2\[5\].wave_shpr.div.acc\[26\] vssd1
+ vssd1 vccd1 vccd1 _04819_ sky130_fd_sc_hd__or4_2
Xclkbuf_leaf_114_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_114_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_118_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12330_ _03689_ genblk1\[11\].osc.clkdiv_C.cnt\[10\] vssd1 vssd1 vccd1 vccd1 _06023_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_51_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06291__A2 _01240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12261_ genblk2\[1\].wave_shpr.div.b1\[0\] _01329_ _05802_ vssd1 vssd1 vccd1 vccd1
+ _05991_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11212_ _05245_ vssd1 vssd1 vccd1 vccd1 _05246_ sky130_fd_sc_hd__clkbuf_4
X_12192_ genblk2\[11\].wave_shpr.div.acc\[12\] genblk2\[11\].wave_shpr.div.b1\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05930_ sky130_fd_sc_hd__or2b_1
XANTENNA__08640__A _02216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11143_ genblk2\[7\].wave_shpr.div.b1\[11\] genblk2\[7\].wave_shpr.div.acc\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05203_ sky130_fd_sc_hd__and2b_1
XFILLER_0_101_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09517__B1 _04047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11074_ net1001 _05119_ _05126_ _05144_ vssd1 vssd1 vccd1 vccd1 _00674_ sky130_fd_sc_hd__a22o_1
XFILLER_0_37_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10025_ _02170_ genblk2\[3\].wave_shpr.div.busy _02172_ vssd1 vssd1 vccd1 vccd1 _04421_
+ sky130_fd_sc_hd__and3_2
XANTENNA__09471__A _01418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10410__A _04058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11976_ genblk2\[10\].wave_shpr.div.fin_quo\[5\] genblk2\[10\].wave_shpr.div.quo\[4\]
+ _00003_ vssd1 vssd1 vccd1 vccd1 _05793_ sky130_fd_sc_hd__mux2_1
X_13715_ clknet_leaf_21_clk _01026_ net97 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.b1\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10927_ genblk2\[7\].wave_shpr.div.b1\[15\] _01365_ _05042_ vssd1 vssd1 vccd1 vccd1
+ _05048_ sky130_fd_sc_hd__mux2_1
X_13646_ clknet_leaf_48_clk _00959_ net114 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.quo\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10858_ genblk2\[6\].wave_shpr.div.b1\[10\] genblk2\[6\].wave_shpr.div.acc\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05002_ sky130_fd_sc_hd__and2b_1
XFILLER_0_128_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07059__A1 genblk1\[8\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07059__B2 genblk1\[8\].osc.clkdiv_C.cnt\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_105_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_105_clk
+ sky130_fd_sc_hd__clkbuf_16
X_13577_ clknet_leaf_76_clk _00892_ net207 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.acc\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10789_ net1345 _04941_ vssd1 vssd1 vccd1 vccd1 _04944_ sky130_fd_sc_hd__nand2_1
XPHY_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11241__A _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12528_ clknet_leaf_43_clk _00080_ net124 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.b1\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12459_ clknet_leaf_104_clk _00032_ net153 vssd1 vssd1 vccd1 vccd1 PWM.final_sample_in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09220__A2 _03836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09508__B1 _04011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07166__A genblk1\[9\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07782__A2 _01241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06951_ genblk1\[6\].osc.clkdiv_C.cnt\[16\] _01787_ vssd1 vssd1 vccd1 vccd1 _01789_
+ sky130_fd_sc_hd__or2_1
XANTENNA__11315__B1 _05283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10669__A2 _04858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09670_ _04045_ _04150_ _04152_ _04048_ net757 vssd1 vssd1 vccd1 vccd1 _00262_ sky130_fd_sc_hd__a32o_1
X_06882_ genblk1\[6\].osc.clkdiv_C.cnt\[9\] _01732_ _01735_ genblk1\[6\].osc.clkdiv_C.cnt\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01736_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__13338__RESET_B net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08621_ _03251_ _03308_ _03327_ vssd1 vssd1 vccd1 vccd1 _03328_ sky130_fd_sc_hd__o21a_1
X_08552_ genblk2\[6\].wave_shpr.div.fin_quo\[0\] _02734_ genblk2\[6\].wave_shpr.div.fin_quo\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03259_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07503_ _02223_ vssd1 vssd1 vccd1 vccd1 _02224_ sky130_fd_sc_hd__clkbuf_4
X_08483_ genblk2\[3\].wave_shpr.div.fin_quo\[2\] vssd1 vssd1 vccd1 vccd1 _03190_ sky130_fd_sc_hd__inv_2
XFILLER_0_92_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07434_ _02171_ genblk2\[3\].wave_shpr.div.busy _02172_ vssd1 vssd1 vccd1 vccd1 _02173_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_91_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08247__B1 _02223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07365_ genblk1\[11\].osc.clkdiv_C.cnt\[7\] genblk1\[11\].osc.clkdiv_C.cnt\[6\] _02108_
+ genblk1\[11\].osc.clkdiv_C.cnt\[8\] vssd1 vssd1 vccd1 vccd1 _02121_ sky130_fd_sc_hd__a31o_1
XFILLER_0_45_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09104_ genblk2\[0\].wave_shpr.div.acc\[11\] genblk2\[0\].wave_shpr.div.b1\[11\]
+ vssd1 vssd1 vccd1 vccd1 _03752_ sky130_fd_sc_hd__or2b_1
XFILLER_0_17_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06316_ _01269_ _01274_ _01275_ vssd1 vssd1 vccd1 vccd1 genblk1\[0\].osc.clkdiv_C.next_cnt\[2\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_33_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07296_ _02028_ _02060_ _02061_ vssd1 vssd1 vccd1 vccd1 _02062_ sky130_fd_sc_hd__and3_1
XFILLER_0_115_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09035_ _02171_ vssd1 vssd1 vccd1 vccd1 _03704_ sky130_fd_sc_hd__buf_6
X_06247_ _01208_ vssd1 vssd1 vccd1 vccd1 _01209_ sky130_fd_sc_hd__buf_4
XANTENNA__09556__A _03707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold330 genblk2\[7\].wave_shpr.div.quo\[16\] vssd1 vssd1 vccd1 vccd1 net548 sky130_fd_sc_hd__dlygate4sd3_1
X_06178_ _01144_ _01145_ _01147_ _01149_ vssd1 vssd1 vccd1 vccd1 _01150_ sky130_fd_sc_hd__or4bb_4
Xhold341 _00126_ vssd1 vssd1 vccd1 vccd1 net559 sky130_fd_sc_hd__dlygate4sd3_1
Xhold352 _00134_ vssd1 vssd1 vccd1 vccd1 net570 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11297__S _05222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold363 _00335_ vssd1 vssd1 vccd1 vccd1 net581 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold374 genblk1\[0\].osc.clkdiv_C.cnt\[7\] vssd1 vssd1 vccd1 vccd1 net592 sky130_fd_sc_hd__dlygate4sd3_1
Xhold385 _00470_ vssd1 vssd1 vccd1 vccd1 net603 sky130_fd_sc_hd__dlygate4sd3_1
Xhold396 genblk2\[3\].wave_shpr.div.b1\[9\] vssd1 vssd1 vccd1 vccd1 net614 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07773__A2 _01556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09937_ genblk2\[2\].wave_shpr.div.acc\[21\] genblk2\[2\].wave_shpr.div.acc\[20\]
+ _04210_ net22 vssd1 vssd1 vccd1 vccd1 _04343_ sky130_fd_sc_hd__or4_1
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09868_ _04290_ _04180_ vssd1 vssd1 vccd1 vccd1 _04291_ sky130_fd_sc_hd__xnor2_1
Xhold1030 genblk2\[6\].wave_shpr.div.b1\[12\] vssd1 vssd1 vccd1 vccd1 net1248 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1041 genblk2\[9\].wave_shpr.div.fin_quo\[7\] vssd1 vssd1 vccd1 vccd1 net1259
+ sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout68_A net85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1052 genblk2\[1\].wave_shpr.div.b1\[14\] vssd1 vssd1 vccd1 vccd1 net1270 sky130_fd_sc_hd__dlygate4sd3_1
X_08819_ _03461_ _03463_ vssd1 vssd1 vccd1 vccd1 _03526_ sky130_fd_sc_hd__nor2_1
Xhold1063 genblk2\[4\].wave_shpr.div.b1\[13\] vssd1 vssd1 vccd1 vccd1 net1281 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1074 genblk2\[10\].wave_shpr.div.b1\[11\] vssd1 vssd1 vccd1 vccd1 net1292 sky130_fd_sc_hd__dlygate4sd3_1
X_09799_ _04250_ vssd1 vssd1 vccd1 vccd1 _04252_ sky130_fd_sc_hd__clkbuf_4
XTAP_2502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1085 genblk2\[5\].wave_shpr.div.b1\[9\] vssd1 vssd1 vccd1 vccd1 net1303 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1096 genblk2\[0\].wave_shpr.div.quo\[2\] vssd1 vssd1 vccd1 vccd1 net1314 sky130_fd_sc_hd__dlygate4sd3_1
X_11830_ net974 _05652_ _05653_ _05674_ vssd1 vssd1 vccd1 vccd1 _00900_ sky130_fd_sc_hd__a22o_1
XTAP_2535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11085__A2 _05057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11761_ _03693_ vssd1 vssd1 vccd1 vccd1 _05629_ sky130_fd_sc_hd__clkbuf_4
XTAP_1845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13500_ clknet_leaf_87_clk _00817_ net179 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.quo\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10712_ net910 _04853_ _04857_ _04885_ vssd1 vssd1 vccd1 vccd1 _00571_ sky130_fd_sc_hd__a22o_1
XTAP_1867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11692_ genblk2\[9\].wave_shpr.div.b1\[6\] genblk2\[9\].wave_shpr.div.acc\[6\] vssd1
+ vssd1 vccd1 vccd1 _05584_ sky130_fd_sc_hd__and2b_1
XANTENNA__08635__A genblk2\[8\].wave_shpr.div.fin_quo\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_138_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13431_ clknet_leaf_82_clk _00750_ net201 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.acc\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10643_ _04849_ vssd1 vssd1 vccd1 vccd1 _00538_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12034__B2 genblk2\[10\].wave_shpr.div.quo\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_548 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10045__B1 _03717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13362_ clknet_leaf_6_clk _00681_ net47 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.i\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10574_ genblk2\[5\].wave_shpr.div.b1\[11\] genblk2\[5\].wave_shpr.div.acc\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04802_ sky130_fd_sc_hd__and2b_1
XFILLER_0_91_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10596__A1 genblk2\[5\].wave_shpr.div.quo\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_5_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12313_ genblk2\[11\].wave_shpr.div.quo\[11\] _03947_ _03944_ net467 _06013_ vssd1
+ vssd1 vccd1 vccd1 _01044_ sky130_fd_sc_hd__a221o_1
XFILLER_0_121_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13293_ clknet_leaf_87_clk _00614_ net179 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.b1\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12337__A2 _03942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12244_ _05981_ vssd1 vssd1 vccd1 vccd1 _05982_ sky130_fd_sc_hd__buf_4
XFILLER_0_121_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12175_ genblk2\[10\].wave_shpr.div.i\[1\] genblk2\[10\].wave_shpr.div.i\[0\] vssd1
+ vssd1 vccd1 vccd1 _05917_ sky130_fd_sc_hd__or2_1
XANTENNA__10405__A _04477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11000__S _05023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11126_ genblk2\[7\].wave_shpr.div.b1\[2\] genblk2\[7\].wave_shpr.div.acc\[2\] vssd1
+ vssd1 vccd1 vccd1 _05186_ sky130_fd_sc_hd__and2b_1
X_11057_ net1093 _05119_ _05126_ _05132_ vssd1 vssd1 vccd1 vccd1 _00669_ sky130_fd_sc_hd__a22o_1
X_10008_ _04366_ _04402_ _04403_ vssd1 vssd1 vccd1 vccd1 _04404_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_86_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11959_ _05731_ _05779_ _05780_ vssd1 vssd1 vccd1 vccd1 _05781_ sky130_fd_sc_hd__a21o_1
XANTENNA__08477__B1 _02222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13629_ clknet_leaf_38_clk _00942_ net116 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.b1\[11\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_27_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07150_ genblk1\[9\].osc.clkdiv_C.cnt\[12\] _01799_ _01948_ _01949_ vssd1 vssd1 vccd1
+ vccd1 _01950_ sky130_fd_sc_hd__o211a_1
XFILLER_0_70_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11784__B1 _03693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07081_ net1162 _01892_ _01894_ vssd1 vssd1 vccd1 vccd1 genblk1\[8\].osc.clkdiv_C.next_cnt\[4\]
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__06255__A2 _01211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10339__A1 _03732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12006__S _05802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout106 net107 vssd1 vssd1 vccd1 vccd1 net106 sky130_fd_sc_hd__buf_2
XANTENNA__06512__B _01437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout117 net118 vssd1 vssd1 vccd1 vccd1 net117 sky130_fd_sc_hd__clkbuf_2
Xfanout128 net129 vssd1 vssd1 vccd1 vccd1 net128 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11551__A3 _05417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07983_ _02683_ _02689_ vssd1 vssd1 vccd1 vccd1 _02690_ sky130_fd_sc_hd__nand2_1
Xfanout139 net140 vssd1 vssd1 vccd1 vccd1 net139 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06963__B1 _01238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09722_ _04159_ _04200_ _04201_ vssd1 vssd1 vccd1 vccd1 _04202_ sky130_fd_sc_hd__a21o_1
X_06934_ net28 _01777_ vssd1 vssd1 vccd1 vccd1 _01778_ sky130_fd_sc_hd__nor2_1
X_09653_ genblk2\[1\].wave_shpr.div.acc\[22\] _04139_ genblk2\[1\].wave_shpr.div.acc\[23\]
+ vssd1 vssd1 vccd1 vccd1 _04141_ sky130_fd_sc_hd__or3b_1
X_06865_ net27 _01721_ vssd1 vssd1 vccd1 vccd1 _01722_ sky130_fd_sc_hd__nor2_1
X_08604_ _02261_ _03309_ _03310_ vssd1 vssd1 vccd1 vccd1 _03311_ sky130_fd_sc_hd__or3b_1
X_09584_ net1260 _04076_ _04080_ _04089_ vssd1 vssd1 vccd1 vccd1 _00239_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06796_ genblk1\[5\].osc.clkdiv_C.cnt\[13\] _01666_ _01667_ genblk1\[5\].osc.clkdiv_C.cnt\[11\]
+ vssd1 vssd1 vccd1 vccd1 _01668_ sky130_fd_sc_hd__a2bb2o_1
XTAP_1108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08535_ _02314_ _03241_ vssd1 vssd1 vccd1 vccd1 _03242_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10985__A _05074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08466_ _03170_ _03171_ _03172_ vssd1 vssd1 vccd1 vccd1 _03173_ sky130_fd_sc_hd__nand3_4
XFILLER_0_77_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07140__B1 _01328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07417_ _02157_ _02153_ genblk2\[1\].wave_shpr.div.busy vssd1 vssd1 vccd1 vccd1 _02160_
+ sky130_fd_sc_hd__and3b_2
XFILLER_0_107_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08397_ genblk1\[2\].osc.clkdiv_C.cnt\[14\] _01209_ _02425_ genblk1\[2\].osc.clkdiv_C.cnt\[13\]
+ vssd1 vssd1 vccd1 vccd1 _03104_ sky130_fd_sc_hd__a22o_1
X_07348_ _02107_ vssd1 vssd1 vccd1 vccd1 genblk1\[11\].osc.clkdiv_C.next_cnt\[4\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07279_ genblk1\[10\].osc.clkdiv_C.cnt\[10\] _02048_ _02050_ _02028_ vssd1 vssd1
+ vccd1 vccd1 genblk1\[10\].osc.clkdiv_C.next_cnt\[10\] sky130_fd_sc_hd__o211a_1
XFILLER_0_21_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10924__S _05042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_492 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09286__A _03838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07994__A2 _01732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07132__A2_N _01578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09018_ genblk2\[9\].wave_shpr.div.busy net1039 genblk2\[9\].wave_shpr.div.i\[0\]
+ _03688_ _03690_ vssd1 vssd1 vccd1 vccd1 _00072_ sky130_fd_sc_hd__a311oi_1
XFILLER_0_60_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10290_ genblk2\[4\].wave_shpr.div.b1\[10\] genblk2\[4\].wave_shpr.div.acc\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04602_ sky130_fd_sc_hd__and2b_1
XFILLER_0_130_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09196__A1 _03712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold160 genblk2\[5\].wave_shpr.div.quo\[16\] vssd1 vssd1 vccd1 vccd1 net378 sky130_fd_sc_hd__dlygate4sd3_1
Xhold171 genblk2\[8\].wave_shpr.div.b1\[2\] vssd1 vssd1 vccd1 vccd1 net389 sky130_fd_sc_hd__dlygate4sd3_1
Xhold182 genblk2\[7\].wave_shpr.div.quo\[18\] vssd1 vssd1 vccd1 vccd1 net400 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06422__B _01249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold193 _00141_ vssd1 vssd1 vccd1 vccd1 net411 sky130_fd_sc_hd__dlygate4sd3_1
X_12931_ clknet_leaf_31_clk _00260_ net102 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.i\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_12862_ clknet_leaf_126_clk _00193_ net61 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.b1\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_34_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11813_ net999 _05652_ _05653_ _05661_ vssd1 vssd1 vccd1 vccd1 _00896_ sky130_fd_sc_hd__a22o_1
XANTENNA__08459__B1 _02261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12793_ clknet_leaf_93_clk net559 net148 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11744_ _03693_ vssd1 vssd1 vccd1 vccd1 _05624_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_139_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11675_ genblk2\[9\].wave_shpr.div.b1\[4\] genblk2\[9\].wave_shpr.div.acc\[4\] vssd1
+ vssd1 vccd1 vccd1 _05567_ sky130_fd_sc_hd__or2b_1
XFILLER_0_36_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09959__B1 _04253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13414_ clknet_leaf_120_clk _00733_ net141 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.quo\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10626_ net1258 net37 _04834_ vssd1 vssd1 vccd1 vccd1 _04840_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13345_ clknet_leaf_6_clk _00666_ net49 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.acc\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06237__A2 _01197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10557_ genblk2\[5\].wave_shpr.div.b1\[2\] genblk2\[5\].wave_shpr.div.acc\[2\] vssd1
+ vssd1 vccd1 vccd1 _04785_ sky130_fd_sc_hd__and2b_1
XFILLER_0_59_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13276_ clknet_leaf_12_clk _00597_ net54 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.i\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_110_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10488_ net881 _04715_ _04722_ _04731_ vssd1 vssd1 vccd1 vccd1 _00501_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11518__B1 _05449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12227_ genblk2\[11\].wave_shpr.div.b1\[12\] genblk2\[11\].wave_shpr.div.acc\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05965_ sky130_fd_sc_hd__and2b_1
XANTENNA__08934__A1 _01099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12158_ net1087 _05876_ _05883_ _05906_ vssd1 vssd1 vccd1 vccd1 _00996_ sky130_fd_sc_hd__a22o_1
X_11109_ genblk2\[7\].wave_shpr.div.acc\[12\] genblk2\[7\].wave_shpr.div.b1\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05169_ sky130_fd_sc_hd__or2b_1
X_12089_ _05754_ _05743_ vssd1 vssd1 vccd1 vccd1 _05854_ sky130_fd_sc_hd__nor2_1
X_06650_ _01523_ _01545_ vssd1 vssd1 vccd1 vccd1 _01546_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06581_ _01187_ vssd1 vssd1 vccd1 vccd1 _01489_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_86_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08320_ _03025_ _03026_ genblk2\[9\].wave_shpr.div.fin_quo\[4\] _02362_ vssd1 vssd1
+ vccd1 vccd1 _03027_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_86_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07122__B1 _01328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_702 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08251_ _02946_ _02951_ _02957_ vssd1 vssd1 vccd1 vccd1 _02958_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06507__B _01432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07202_ genblk1\[9\].osc.clkdiv_C.cnt\[15\] _01983_ _01986_ vssd1 vssd1 vccd1 vccd1
+ genblk1\[9\].osc.clkdiv_C.next_cnt\[15\] sky130_fd_sc_hd__o21a_1
X_08182_ _02850_ _02888_ _02224_ vssd1 vssd1 vccd1 vccd1 _02889_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11757__B1 _03694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07133_ genblk1\[9\].osc.clkdiv_C.cnt\[7\] _01513_ _01929_ _01931_ _01932_ vssd1
+ vssd1 vccd1 vccd1 _01933_ sky130_fd_sc_hd__a221o_1
XANTENNA__11221__A2 _05246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout118_A net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07064_ _01874_ _01876_ _01877_ _01881_ vssd1 vssd1 vccd1 vccd1 _01882_ sky130_fd_sc_hd__or4b_1
XFILLER_0_113_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09178__A1 _01342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08386__C1 _01441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07966_ genblk1\[7\].osc.clkdiv_C.cnt\[12\] _01214_ _01675_ genblk1\[7\].osc.clkdiv_C.cnt\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02673_ sky130_fd_sc_hd__o22a_1
X_09705_ genblk2\[2\].wave_shpr.div.b1\[6\] genblk2\[2\].wave_shpr.div.acc\[6\] vssd1
+ vssd1 vccd1 vccd1 _04185_ sky130_fd_sc_hd__and2b_1
XANTENNA__09045__S _03708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06917_ genblk1\[6\].osc.clkdiv_C.cnt\[4\] _01765_ vssd1 vssd1 vccd1 vccd1 _01767_
+ sky130_fd_sc_hd__xnor2_1
X_07897_ _02603_ vssd1 vssd1 vccd1 vccd1 _02604_ sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_94_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_94_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_97_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08153__A2 _01500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09636_ genblk2\[1\].wave_shpr.div.acc\[25\] genblk2\[1\].wave_shpr.div.acc\[26\]
+ _04009_ vssd1 vssd1 vccd1 vccd1 _04129_ sky130_fd_sc_hd__nor3_2
X_06848_ genblk1\[5\].osc.clkdiv_C.cnt\[9\] _01708_ vssd1 vssd1 vccd1 vccd1 _01711_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__07900__A2 _01172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09567_ _04042_ vssd1 vssd1 vccd1 vccd1 _04076_ sky130_fd_sc_hd__clkbuf_4
X_06779_ genblk1\[4\].osc.clkdiv_C.cnt\[16\] _01652_ vssd1 vssd1 vccd1 vccd1 _01653_
+ sky130_fd_sc_hd__or2_1
X_08518_ _03136_ _03224_ vssd1 vssd1 vccd1 vccd1 _03225_ sky130_fd_sc_hd__nor2_1
X_09498_ net1282 _01327_ _04039_ vssd1 vssd1 vccd1 vccd1 _04040_ sky130_fd_sc_hd__mux2_1
XFILLER_0_81_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_154_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08449_ genblk2\[8\].wave_shpr.div.fin_quo\[3\] net30 _02639_ _02316_ vssd1 vssd1
+ vccd1 vccd1 _03156_ sky130_fd_sc_hd__a31o_1
XFILLER_0_81_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_93_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07664__B2 _01182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11460_ genblk2\[9\].wave_shpr.div.b1\[1\] _01819_ _05237_ vssd1 vssd1 vccd1 vccd1
+ _05427_ sky130_fd_sc_hd__mux2_1
XANTENNA__11748__B1 _05624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10411_ net665 _04651_ _04663_ genblk2\[4\].wave_shpr.div.quo\[21\] _04674_ vssd1
+ vssd1 vccd1 vccd1 _00481_ sky130_fd_sc_hd__a221o_1
XFILLER_0_150_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11391_ genblk2\[8\].wave_shpr.div.acc\[8\] genblk2\[8\].wave_shpr.div.b1\[8\] vssd1
+ vssd1 vccd1 vccd1 _05367_ sky130_fd_sc_hd__or2b_1
XFILLER_0_104_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13130_ clknet_leaf_3_clk _00455_ net46 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.b1\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07967__A2 _01214_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07529__A _01099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10342_ genblk2\[5\].wave_shpr.div.b1\[8\] _01326_ _04637_ vssd1 vssd1 vccd1 vccd1
+ _04638_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13061_ clknet_leaf_29_clk net388 net95 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.quo\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10273_ genblk2\[4\].wave_shpr.div.b1\[0\] _04583_ _04584_ vssd1 vssd1 vccd1 vccd1
+ _04585_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12173__A0 _05815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13094__RESET_B net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07719__A2 _01309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12012_ net1086 vssd1 vssd1 vccd1 vccd1 _05810_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_85_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_85_clk sky130_fd_sc_hd__clkbuf_16
X_12914_ clknet_leaf_36_clk net367 net106 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.acc\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xmax_cap6 _01692_ vssd1 vssd1 vccd1 vccd1 net1355 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12845_ clknet_leaf_68_clk _00176_ net194 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.i\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_2151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_152_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10239__A0 _04455_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11514__A _04676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07711__B net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12776_ clknet_leaf_43_clk _00109_ net124 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.b1\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11727_ _05616_ vssd1 vssd1 vccd1 vccd1 _00855_ sky130_fd_sc_hd__clkbuf_1
XTAP_1494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11658_ genblk2\[8\].wave_shpr.div.i\[3\] _02197_ _05549_ vssd1 vssd1 vccd1 vccd1
+ _05552_ sky130_fd_sc_hd__and3_1
XFILLER_0_9_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10609_ _04829_ vssd1 vssd1 vccd1 vccd1 _00524_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11203__A2 _01869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11589_ genblk2\[8\].wave_shpr.div.acc\[9\] _05502_ _05493_ vssd1 vssd1 vccd1 vccd1
+ _05503_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_44 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold907 genblk2\[11\].wave_shpr.div.acc\[16\] vssd1 vssd1 vccd1 vccd1 net1125 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07439__A _02147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13328_ clknet_leaf_25_clk _00649_ net86 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.quo\[22\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold918 genblk1\[9\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 net1136 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08080__A1 _01200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold929 genblk2\[8\].wave_shpr.div.b1\[12\] vssd1 vssd1 vccd1 vccd1 net1147 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13259_ clknet_leaf_2_clk _00582_ net43 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.acc\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07820_ _02526_ vssd1 vssd1 vccd1 vccd1 _02527_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__06489__S _01210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06394__B2 genblk1\[1\].osc.clkdiv_C.cnt\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07751_ _02428_ _02450_ _02452_ _02457_ vssd1 vssd1 vccd1 vccd1 _02458_ sky130_fd_sc_hd__a31o_4
XANTENNA_clkbuf_leaf_92_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_76_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_76_clk sky130_fd_sc_hd__clkbuf_16
X_06702_ _01171_ _01591_ vssd1 vssd1 vccd1 vccd1 _01592_ sky130_fd_sc_hd__nand2_4
XFILLER_0_126_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06146__A1 net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07682_ genblk1\[10\].osc.clkdiv_C.cnt\[13\] _01246_ _02386_ vssd1 vssd1 vccd1 vccd1
+ _02389_ sky130_fd_sc_hd__a21oi_1
X_09421_ _03964_ _03983_ _03984_ vssd1 vssd1 vccd1 vccd1 _03985_ sky130_fd_sc_hd__a21o_1
X_06633_ genblk1\[3\].osc.clkdiv_C.cnt\[6\] _01533_ vssd1 vssd1 vccd1 vccd1 _01535_
+ sky130_fd_sc_hd__and2_1
XANTENNA__06697__A2 _01436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_47_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09352_ genblk2\[0\].wave_shpr.div.acc\[19\] _03924_ _03927_ vssd1 vssd1 vccd1 vccd1
+ _03928_ sky130_fd_sc_hd__a21o_1
XFILLER_0_75_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06564_ genblk1\[2\].osc.clkdiv_C.cnt\[14\] _01474_ vssd1 vssd1 vccd1 vccd1 _01476_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_75_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08303_ _03007_ _03005_ vssd1 vssd1 vccd1 vccd1 _03010_ sky130_fd_sc_hd__xnor2_1
X_09283_ _03768_ _03874_ vssd1 vssd1 vccd1 vccd1 _03875_ sky130_fd_sc_hd__xnor2_1
X_06495_ genblk1\[2\].osc.clkdiv_C.cnt\[14\] genblk1\[2\].osc.clkdiv_C.cnt\[1\] _01327_
+ vssd1 vssd1 vccd1 vccd1 _01421_ sky130_fd_sc_hd__nor3_1
XFILLER_0_145_643 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08234_ _02885_ _02887_ genblk2\[3\].wave_shpr.div.fin_quo\[5\] vssd1 vssd1 vccd1
+ vccd1 _02941_ sky130_fd_sc_hd__o21bai_1
XANTENNA__09829__A _04069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_30_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10474__S _04704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_598 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08165_ genblk1\[3\].osc.clkdiv_C.cnt\[10\] _01508_ vssd1 vssd1 vccd1 vccd1 _02872_
+ sky130_fd_sc_hd__or2_1
XANTENNA__09548__B genblk1\[1\].osc.clkdiv_C.cnt\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07116_ _01886_ _01916_ _01917_ vssd1 vssd1 vccd1 vccd1 _01918_ sky130_fd_sc_hd__and3b_1
X_08096_ _01174_ genblk1\[4\].osc.clkdiv_C.cnt\[15\] _01359_ vssd1 vssd1 vccd1 vccd1
+ _02803_ sky130_fd_sc_hd__or3_1
XANTENNA__06253__A _01213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07047_ _01336_ _01223_ vssd1 vssd1 vccd1 vccd1 _01865_ sky130_fd_sc_hd__or2_2
XANTENNA_clkbuf_leaf_45_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08998_ net1103 sig_norm.quo\[0\] _01154_ vssd1 vssd1 vccd1 vccd1 _03679_ sky130_fd_sc_hd__mux2_1
XANTENNA__06700__B _01589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07949_ _01172_ _02011_ vssd1 vssd1 vccd1 vccd1 _02656_ sky130_fd_sc_hd__nand2_2
Xclkbuf_leaf_67_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_67_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__08126__A2 _01340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_103_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10960_ _05059_ genblk1\[6\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 _05065_
+ sky130_fd_sc_hd__and2_1
XANTENNA_fanout50_A net85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09619_ net1019 _04109_ _04113_ _04116_ vssd1 vssd1 vccd1 vccd1 _00247_ sky130_fd_sc_hd__a22o_1
X_10891_ _05029_ vssd1 vssd1 vccd1 vccd1 _00606_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12630_ clknet_leaf_18_clk genblk1\[4\].osc.clkdiv_C.next_cnt\[15\] net82 vssd1 vssd1
+ vccd1 vccd1 genblk1\[4\].osc.clkdiv_C.cnt\[15\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_38_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_118_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12561_ clknet_leaf_29_clk genblk1\[1\].osc.clkdiv_C.next_cnt\[0\] net96 vssd1 vssd1
+ vccd1 vccd1 genblk1\[1\].osc.clkdiv_C.cnt\[0\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__10338__B1_N _03733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06147__B net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11512_ _05450_ genblk1\[8\].osc.clkdiv_C.cnt\[1\] vssd1 vssd1 vccd1 vccd1 _05452_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_25_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12492_ clknet_leaf_107_clk _00054_ net153 vssd1 vssd1 vccd1 vccd1 sig_norm.quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11443_ _05418_ vssd1 vssd1 vccd1 vccd1 _00769_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11374_ genblk2\[7\].wave_shpr.div.i\[1\] genblk2\[7\].wave_shpr.div.i\[0\] genblk2\[7\].wave_shpr.div.i\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05353_ sky130_fd_sc_hd__and3_1
XFILLER_0_22_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13113_ clknet_leaf_115_clk _00438_ net134 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.fin_quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10325_ _04630_ vssd1 vssd1 vccd1 vccd1 _00439_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_132_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13044_ clknet_leaf_128_clk _00371_ net67 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.b1\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10256_ genblk2\[4\].wave_shpr.div.acc\[14\] genblk2\[4\].wave_shpr.div.b1\[14\]
+ vssd1 vssd1 vccd1 vccd1 _04568_ sky130_fd_sc_hd__or2b_1
XANTENNA__11509__A _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12104__S _05865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10187_ _04451_ vssd1 vssd1 vccd1 vccd1 _04518_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_58_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_58_clk sky130_fd_sc_hd__clkbuf_16
Xclkbuf_4_11_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_11_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__07325__B1 _01925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08522__C1 _02364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06679__A2 _01363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10880__A0 genblk2\[6\].wave_shpr.div.fin_quo\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__07441__B _02153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12828_ clknet_leaf_62_clk _00161_ net190 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.acc\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_552 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07160__C genblk1\[9\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12759_ clknet_leaf_58_clk _00000_ net192 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.busy
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06280_ _01241_ vssd1 vssd1 vccd1 vccd1 _01242_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_127_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11188__A1 _01507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_696 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold704 genblk2\[8\].wave_shpr.div.acc\[9\] vssd1 vssd1 vccd1 vccd1 net922 sky130_fd_sc_hd__dlygate4sd3_1
Xhold715 genblk2\[0\].wave_shpr.div.acc\[22\] vssd1 vssd1 vccd1 vccd1 net933 sky130_fd_sc_hd__dlygate4sd3_1
Xhold726 genblk2\[10\].wave_shpr.div.acc\[15\] vssd1 vssd1 vccd1 vccd1 net944 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold737 genblk2\[11\].wave_shpr.div.acc\[22\] vssd1 vssd1 vccd1 vccd1 net955 sky130_fd_sc_hd__dlygate4sd3_1
Xhold748 genblk2\[3\].wave_shpr.div.acc\[8\] vssd1 vssd1 vccd1 vccd1 net966 sky130_fd_sc_hd__dlygate4sd3_1
X_09970_ genblk2\[3\].wave_shpr.div.acc\[12\] genblk2\[3\].wave_shpr.div.b1\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04366_ sky130_fd_sc_hd__or2b_1
XANTENNA__06603__A2 _01487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold759 genblk2\[10\].wave_shpr.div.acc\[5\] vssd1 vssd1 vccd1 vccd1 net977 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08921_ net678 _02260_ _03619_ _03574_ vssd1 vssd1 vccd1 vccd1 _00046_ sky130_fd_sc_hd__a22o_1
X_08852_ _03546_ _03551_ _03557_ _03558_ vssd1 vssd1 vccd1 vccd1 _03559_ sky130_fd_sc_hd__a211oi_2
XANTENNA__07564__B1 _01732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07803_ net31 vssd1 vssd1 vccd1 vccd1 _02510_ sky130_fd_sc_hd__buf_2
XFILLER_0_137_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08783_ _03478_ _03477_ vssd1 vssd1 vccd1 vccd1 _03490_ sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_49_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_49_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA_fanout185_A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07734_ _02435_ _02436_ vssd1 vssd1 vccd1 vccd1 _02441_ sky130_fd_sc_hd__nor2_1
X_07665_ _02369_ _02370_ _02371_ vssd1 vssd1 vccd1 vccd1 _02372_ sky130_fd_sc_hd__a21oi_1
X_09404_ genblk2\[1\].wave_shpr.div.acc\[3\] genblk2\[1\].wave_shpr.div.b1\[3\] vssd1
+ vssd1 vccd1 vccd1 _03968_ sky130_fd_sc_hd__or2b_1
X_06616_ net1101 _01523_ vssd1 vssd1 vccd1 vccd1 genblk1\[3\].osc.clkdiv_C.next_cnt\[0\]
+ sky130_fd_sc_hd__nor2_1
X_07596_ net32 vssd1 vssd1 vccd1 vccd1 _02303_ sky130_fd_sc_hd__buf_2
XANTENNA__06248__A _01209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09335_ _03792_ _03914_ vssd1 vssd1 vccd1 vccd1 _03915_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06547_ genblk1\[2\].osc.clkdiv_C.cnt\[7\] _01461_ genblk1\[2\].osc.clkdiv_C.cnt\[8\]
+ vssd1 vssd1 vccd1 vccd1 _01465_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_63_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09266_ net578 _03835_ _03838_ genblk2\[0\].wave_shpr.div.quo\[24\] _03862_ vssd1
+ vssd1 vccd1 vccd1 _00148_ sky130_fd_sc_hd__a221o_1
XFILLER_0_63_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06478_ genblk1\[1\].osc.clkdiv_C.cnt\[15\] _01403_ _01406_ vssd1 vssd1 vccd1 vccd1
+ genblk1\[1\].osc.clkdiv_C.next_cnt\[15\] sky130_fd_sc_hd__o21a_1
XFILLER_0_133_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08217_ _02899_ _02923_ vssd1 vssd1 vccd1 vccd1 _02924_ sky130_fd_sc_hd__or2b_1
XFILLER_0_132_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09197_ _03826_ vssd1 vssd1 vccd1 vccd1 _00115_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11179__A1 _03831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_90_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08044__A1 _01181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08148_ genblk1\[3\].osc.clkdiv_C.cnt\[1\] _01496_ _01513_ genblk1\[3\].osc.clkdiv_C.cnt\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02855_ sky130_fd_sc_hd__a22o_1
XANTENNA__10926__A1 _03704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08079_ genblk1\[5\].osc.clkdiv_C.cnt\[11\] _01355_ _02760_ _02782_ _02785_ vssd1
+ vssd1 vccd1 vccd1 _02786_ sky130_fd_sc_hd__o221a_1
XFILLER_0_30_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10110_ _04465_ genblk1\[3\].osc.clkdiv_C.cnt\[5\] vssd1 vssd1 vccd1 vccd1 _04466_
+ sky130_fd_sc_hd__and2_1
XANTENNA_fanout98_A net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11090_ _05054_ _05051_ genblk2\[6\].wave_shpr.div.i\[0\] vssd1 vssd1 vccd1 vccd1
+ _05155_ sky130_fd_sc_hd__mux2_1
X_10041_ genblk2\[3\].wave_shpr.div.fin_quo\[7\] genblk2\[3\].wave_shpr.div.quo\[6\]
+ _04422_ vssd1 vssd1 vccd1 vccd1 _04430_ sky130_fd_sc_hd__mux2_1
Xhold20 _00810_ vssd1 vssd1 vccd1 vccd1 net238 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 genblk2\[5\].wave_shpr.div.quo\[14\] vssd1 vssd1 vccd1 vccd1 net249 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 _00316_ vssd1 vssd1 vccd1 vccd1 net260 sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 genblk2\[6\].wave_shpr.div.quo\[3\] vssd1 vssd1 vccd1 vccd1 net271 sky130_fd_sc_hd__dlygate4sd3_1
Xhold64 genblk2\[2\].wave_shpr.div.i\[4\] vssd1 vssd1 vccd1 vccd1 net282 sky130_fd_sc_hd__dlygate4sd3_1
Xhold75 _00214_ vssd1 vssd1 vccd1 vccd1 net293 sky130_fd_sc_hd__dlygate4sd3_1
Xhold86 genblk2\[9\].wave_shpr.div.quo\[15\] vssd1 vssd1 vccd1 vccd1 net304 sky130_fd_sc_hd__dlygate4sd3_1
Xhold97 genblk2\[2\].wave_shpr.div.quo\[15\] vssd1 vssd1 vccd1 vccd1 net315 sky130_fd_sc_hd__dlygate4sd3_1
X_11992_ genblk2\[11\].wave_shpr.div.b1\[5\] _01855_ _05433_ vssd1 vssd1 vccd1 vccd1
+ _05801_ sky130_fd_sc_hd__mux2_1
XANTENNA__12300__B1 _06010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10943_ genblk2\[6\].wave_shpr.div.quo\[4\] _05052_ _05056_ net271 vssd1 vssd1 vccd1
+ vccd1 _00631_ sky130_fd_sc_hd__a22o_1
X_13731_ clknet_leaf_45_clk net356 net121 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.quo\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10874_ genblk2\[6\].wave_shpr.div.acc\[18\] _05017_ vssd1 vssd1 vccd1 vccd1 _05018_
+ sky130_fd_sc_hd__or2_1
X_13662_ clknet_leaf_45_clk net248 net121 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.acc\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06158__A net12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12613_ clknet_leaf_23_clk genblk1\[3\].osc.clkdiv_C.next_cnt\[16\] net94 vssd1 vssd1
+ vccd1 vccd1 genblk1\[3\].osc.clkdiv_C.cnt\[16\] sky130_fd_sc_hd__dfrtp_2
X_13593_ clknet_leaf_72_clk _00908_ net216 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.acc\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12544_ clknet_leaf_60_clk genblk1\[0\].osc.clkdiv_C.next_cnt\[1\] net192 vssd1 vssd1
+ vccd1 vccd1 genblk1\[0\].osc.clkdiv_C.cnt\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_93_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12475_ clknet_leaf_116_clk FSM.next_mode\[1\] net150 vssd1 vssd1 vccd1 vccd1 net18
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_151_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10408__A _04672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11426_ genblk2\[8\].wave_shpr.div.b1\[14\] genblk2\[8\].wave_shpr.div.acc\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05402_ sky130_fd_sc_hd__and2b_1
XFILLER_0_1_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_6 _04242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09232__B1 _03839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09783__A1 _03732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11357_ net873 _05251_ _05315_ _05341_ vssd1 vssd1 vccd1 vccd1 _00760_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_830 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10308_ genblk2\[4\].wave_shpr.div.acc\[22\] _04619_ vssd1 vssd1 vccd1 vccd1 _04620_
+ sky130_fd_sc_hd__or2_1
XANTENNA__07717__A net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11288_ _05289_ _05190_ vssd1 vssd1 vccd1 vccd1 _05290_ sky130_fd_sc_hd__xnor2_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13027_ clknet_leaf_113_clk _00354_ net131 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.fin_quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11239__A _05074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10239_ _04455_ _04451_ genblk2\[3\].wave_shpr.div.i\[0\] vssd1 vssd1 vccd1 vccd1
+ _04556_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07450_ _02184_ vssd1 vssd1 vccd1 vccd1 _00015_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_147_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06521__B2 _01436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06401_ _01342_ genblk1\[1\].osc.clkdiv_C.cnt\[8\] _01344_ genblk1\[1\].osc.clkdiv_C.cnt\[13\]
+ vssd1 vssd1 vccd1 vccd1 _01345_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07381_ _02132_ vssd1 vssd1 vccd1 vccd1 _02133_ sky130_fd_sc_hd__inv_2
XFILLER_0_146_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09120_ _03761_ genblk2\[0\].wave_shpr.div.acc\[2\] _03767_ vssd1 vssd1 vccd1 vccd1
+ _03768_ sky130_fd_sc_hd__a21o_1
X_06332_ _01269_ _01284_ _01285_ vssd1 vssd1 vccd1 vccd1 genblk1\[0\].osc.clkdiv_C.next_cnt\[8\]
+ sky130_fd_sc_hd__nor3_1
XANTENNA__09379__A _03942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09051_ _03702_ _01257_ vssd1 vssd1 vccd1 vccd1 _03715_ sky130_fd_sc_hd__nand2_1
X_06263_ _01175_ _01194_ vssd1 vssd1 vccd1 vccd1 _01225_ sky130_fd_sc_hd__nor2b_2
XFILLER_0_32_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08002_ genblk1\[6\].osc.clkdiv_C.cnt\[13\] _01675_ _01666_ genblk1\[6\].osc.clkdiv_C.cnt\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02709_ sky130_fd_sc_hd__o22a_1
XFILLER_0_130_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06194_ PWM.counter\[3\] _01159_ vssd1 vssd1 vccd1 vccd1 _01161_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_633 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold501 genblk2\[2\].wave_shpr.div.quo\[2\] vssd1 vssd1 vccd1 vccd1 net719 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09223__B1 _03840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold512 genblk2\[3\].wave_shpr.div.b1\[16\] vssd1 vssd1 vccd1 vccd1 net730 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09774__A1 _03831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold523 genblk2\[11\].wave_shpr.div.i\[2\] vssd1 vssd1 vccd1 vccd1 net741 sky130_fd_sc_hd__dlygate4sd3_1
Xhold534 genblk2\[1\].wave_shpr.div.acc\[0\] vssd1 vssd1 vccd1 vccd1 net752 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_13_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold545 genblk2\[4\].wave_shpr.div.acc\[26\] vssd1 vssd1 vccd1 vccd1 net763 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold556 genblk2\[1\].wave_shpr.div.acc\[16\] vssd1 vssd1 vccd1 vccd1 net774 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_111_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10384__A2 _04657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold567 genblk2\[11\].wave_shpr.div.acc\[11\] vssd1 vssd1 vccd1 vccd1 net785 sky130_fd_sc_hd__dlygate4sd3_1
Xhold578 genblk2\[3\].wave_shpr.div.acc\[9\] vssd1 vssd1 vccd1 vccd1 net796 sky130_fd_sc_hd__dlygate4sd3_1
X_09953_ genblk2\[2\].wave_shpr.div.i\[1\] genblk2\[2\].wave_shpr.div.i\[0\] vssd1
+ vssd1 vccd1 vccd1 _04353_ sky130_fd_sc_hd__or2_1
Xhold589 genblk2\[9\].wave_shpr.div.acc\[11\] vssd1 vssd1 vccd1 vccd1 net807 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08904_ _03584_ _03592_ vssd1 vssd1 vccd1 vccd1 _03607_ sky130_fd_sc_hd__xnor2_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09884_ _04189_ _04165_ vssd1 vssd1 vccd1 vccd1 _04303_ sky130_fd_sc_hd__or2b_1
XFILLER_0_148_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08835_ net8 _02744_ _03541_ vssd1 vssd1 vccd1 vccd1 _03542_ sky130_fd_sc_hd__and3_1
XANTENNA__10988__A _03719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11884__A2 _03696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08766_ _03470_ _03472_ vssd1 vssd1 vccd1 vccd1 _03473_ sky130_fd_sc_hd__and2_1
XTAP_2706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07717_ net7 _02364_ _02365_ vssd1 vssd1 vccd1 vccd1 _02424_ sky130_fd_sc_hd__nand3_2
XANTENNA__10199__S _04507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08697_ _03173_ _03402_ _03403_ _03357_ vssd1 vssd1 vccd1 vccd1 _03404_ sky130_fd_sc_hd__a211o_1
XFILLER_0_95_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07648_ genblk2\[11\].wave_shpr.div.fin_quo\[4\] _02354_ vssd1 vssd1 vccd1 vccd1
+ _02355_ sky130_fd_sc_hd__or2_1
XFILLER_0_95_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10927__S _05042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07579_ _02283_ _02284_ _02285_ vssd1 vssd1 vccd1 vccd1 _02286_ sky130_fd_sc_hd__or3b_1
X_09318_ genblk2\[0\].wave_shpr.div.acc\[11\] _03901_ _03889_ vssd1 vssd1 vccd1 vccd1
+ _03902_ sky130_fd_sc_hd__mux2_1
X_10590_ genblk2\[5\].wave_shpr.div.acc\[22\] _04817_ vssd1 vssd1 vccd1 vccd1 _04818_
+ sky130_fd_sc_hd__or2_2
XFILLER_0_75_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09249_ _03707_ vssd1 vssd1 vccd1 vccd1 _03853_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_145_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12260_ _05990_ vssd1 vssd1 vccd1 vccd1 _01014_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11211_ _02193_ vssd1 vssd1 vccd1 vccd1 _05245_ sky130_fd_sc_hd__clkbuf_4
X_12191_ genblk2\[11\].wave_shpr.div.acc\[13\] genblk2\[11\].wave_shpr.div.b1\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05929_ sky130_fd_sc_hd__or2b_1
XFILLER_0_120_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11142_ _05171_ _05200_ _05201_ vssd1 vssd1 vccd1 vccd1 _05202_ sky130_fd_sc_hd__a21o_1
XANTENNA__07240__A2 _02013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09517__A1 genblk2\[1\].wave_shpr.div.quo\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09517__B2 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11073_ genblk2\[6\].wave_shpr.div.acc\[20\] _05142_ vssd1 vssd1 vccd1 vccd1 _05144_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__10127__A2 _04451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10024_ _04419_ vssd1 vssd1 vccd1 vccd1 _04420_ sky130_fd_sc_hd__buf_4
XFILLER_0_98_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11975_ _05792_ vssd1 vssd1 vccd1 vccd1 _00927_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08087__B _02789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13714_ clknet_leaf_31_clk _01025_ net102 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.b1\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10926_ _03704_ net484 _04647_ vssd1 vssd1 vccd1 vccd1 _00623_ sky130_fd_sc_hd__a21o_1
XFILLER_0_85_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10857_ _04974_ _04999_ _05000_ vssd1 vssd1 vccd1 vccd1 _05001_ sky130_fd_sc_hd__a21o_1
X_13645_ clknet_leaf_48_clk net433 net114 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.quo\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10788_ genblk2\[5\].wave_shpr.div.acc\[20\] _04941_ vssd1 vssd1 vccd1 vccd1 _04943_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_54_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13576_ clknet_leaf_84_clk net1210 net202 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.acc\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XPHY_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12527_ clknet_leaf_67_clk _00079_ net193 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.b1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10138__A _04480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12458_ clknet_leaf_104_clk _00031_ net155 vssd1 vssd1 vccd1 vccd1 PWM.final_sample_in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11409_ _05370_ _05383_ _05384_ vssd1 vssd1 vccd1 vccd1 _05385_ sky130_fd_sc_hd__a21o_1
X_12389_ _05960_ _06063_ vssd1 vssd1 vccd1 vccd1 _06064_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07767__B1 _01208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09508__A1 genblk2\[1\].wave_shpr.div.quo\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06950_ genblk1\[6\].osc.clkdiv_C.cnt\[15\] _01785_ _01788_ vssd1 vssd1 vccd1 vccd1
+ genblk1\[6\].osc.clkdiv_C.next_cnt\[15\] sky130_fd_sc_hd__o21a_1
XANTENNA__09508__B2 _04045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06881_ _01189_ _01678_ vssd1 vssd1 vccd1 vccd1 _01735_ sky130_fd_sc_hd__or2_2
XFILLER_0_118_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_27_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08620_ _03313_ _03326_ vssd1 vssd1 vccd1 vccd1 _03327_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08551_ _03256_ _03257_ vssd1 vssd1 vccd1 vccd1 _03258_ sky130_fd_sc_hd__or2_2
X_07502_ _02222_ vssd1 vssd1 vccd1 vccd1 _02223_ sky130_fd_sc_hd__buf_4
XFILLER_0_77_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08482_ genblk2\[3\].wave_shpr.div.fin_quo\[1\] vssd1 vssd1 vccd1 vccd1 _03189_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07433_ genblk2\[3\].wave_shpr.div.i\[1\] _02166_ genblk2\[3\].wave_shpr.div.i\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02172_ sky130_fd_sc_hd__nor3b_1
XFILLER_0_58_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout148_A net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07364_ _02119_ vssd1 vssd1 vccd1 vccd1 _02120_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09103_ genblk2\[0\].wave_shpr.div.acc\[12\] genblk2\[0\].wave_shpr.div.b1\[12\]
+ vssd1 vssd1 vccd1 vccd1 _03751_ sky130_fd_sc_hd__or2b_1
X_06315_ genblk1\[0\].osc.clkdiv_C.cnt\[1\] genblk1\[0\].osc.clkdiv_C.cnt\[0\] genblk1\[0\].osc.clkdiv_C.cnt\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01275_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_352 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07295_ genblk1\[10\].osc.clkdiv_C.cnt\[16\] _02058_ vssd1 vssd1 vccd1 vccd1 _02061_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_385 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09034_ _03700_ _03703_ vssd1 vssd1 vccd1 vccd1 _00075_ sky130_fd_sc_hd__nor2_1
XFILLER_0_142_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09837__A _04269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06246_ _01207_ vssd1 vssd1 vccd1 vccd1 _01208_ sky130_fd_sc_hd__buf_4
XFILLER_0_115_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold320 genblk2\[3\].wave_shpr.div.quo\[9\] vssd1 vssd1 vccd1 vccd1 net538 sky130_fd_sc_hd__dlygate4sd3_1
X_06177_ _01140_ _01148_ vssd1 vssd1 vccd1 vccd1 _01149_ sky130_fd_sc_hd__or2_1
XFILLER_0_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold331 _00728_ vssd1 vssd1 vccd1 vccd1 net549 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold342 genblk2\[6\].wave_shpr.div.acc\[18\] vssd1 vssd1 vccd1 vccd1 net560 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09048__S _03708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold353 genblk2\[11\].wave_shpr.div.quo\[16\] vssd1 vssd1 vccd1 vccd1 net571 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold364 genblk2\[6\].wave_shpr.div.quo\[17\] vssd1 vssd1 vccd1 vccd1 net582 sky130_fd_sc_hd__dlygate4sd3_1
Xhold375 genblk2\[8\].wave_shpr.div.b1\[4\] vssd1 vssd1 vccd1 vccd1 net593 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold386 genblk2\[0\].wave_shpr.div.acc\[18\] vssd1 vssd1 vccd1 vccd1 net604 sky130_fd_sc_hd__dlygate4sd3_1
Xhold397 genblk2\[8\].wave_shpr.div.acc\[26\] vssd1 vssd1 vccd1 vccd1 net615 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07773__A3 _01564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09936_ genblk2\[2\].wave_shpr.div.acc\[20\] _04210_ net1351 vssd1 vssd1 vccd1 vccd1
+ _04342_ sky130_fd_sc_hd__or3_1
XANTENNA__09572__A _04046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09867_ _04181_ _04169_ vssd1 vssd1 vccd1 vccd1 _04290_ sky130_fd_sc_hd__or2b_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1020 genblk2\[0\].wave_shpr.div.b1\[3\] vssd1 vssd1 vccd1 vccd1 net1238 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1031 genblk2\[10\].wave_shpr.div.b1\[3\] vssd1 vssd1 vccd1 vccd1 net1249 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1042 genblk2\[1\].wave_shpr.div.acc\[6\] vssd1 vssd1 vccd1 vccd1 net1260 sky130_fd_sc_hd__dlygate4sd3_1
X_08818_ _03508_ _03519_ _03523_ _03524_ vssd1 vssd1 vccd1 vccd1 _03525_ sky130_fd_sc_hd__o31a_1
Xhold1053 genblk2\[2\].wave_shpr.div.b1\[13\] vssd1 vssd1 vccd1 vccd1 net1271 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1064 genblk2\[2\].wave_shpr.div.b1\[14\] vssd1 vssd1 vccd1 vccd1 net1282 sky130_fd_sc_hd__dlygate4sd3_1
X_09798_ net1054 _04248_ _04214_ _04251_ vssd1 vssd1 vccd1 vccd1 _00291_ sky130_fd_sc_hd__a22o_1
Xhold1075 genblk2\[7\].wave_shpr.div.b1\[5\] vssd1 vssd1 vccd1 vccd1 net1293 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1086 genblk2\[2\].wave_shpr.div.b1\[10\] vssd1 vssd1 vccd1 vccd1 net1304 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1097 genblk2\[5\].wave_shpr.div.quo\[5\] vssd1 vssd1 vccd1 vccd1 net1315 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08749_ genblk2\[8\].wave_shpr.div.fin_quo\[0\] _02309_ _02636_ vssd1 vssd1 vccd1
+ vccd1 _03456_ sky130_fd_sc_hd__a21oi_1
XTAP_2536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11760_ _02203_ vssd1 vssd1 vccd1 vccd1 _05628_ sky130_fd_sc_hd__clkbuf_4
XTAP_2569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08486__B2 _02592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07820__A _02526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10711_ genblk2\[5\].wave_shpr.div.acc\[1\] _04884_ _04821_ vssd1 vssd1 vccd1 vccd1
+ _04885_ sky130_fd_sc_hd__mux2_1
XTAP_1857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11691_ _05566_ _05581_ _05582_ vssd1 vssd1 vccd1 vccd1 _05583_ sky130_fd_sc_hd__a21o_1
XFILLER_0_36_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10642_ genblk2\[6\].wave_shpr.div.b1\[13\] _04645_ _04848_ vssd1 vssd1 vccd1 vccd1
+ _04849_ sky130_fd_sc_hd__mux2_1
X_13430_ clknet_leaf_82_clk net853 net201 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.acc\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12034__A2 _05818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10045__A1 _03714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13361_ clknet_leaf_6_clk _00680_ net47 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.i\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_106_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10573_ _04770_ _04799_ _04800_ vssd1 vssd1 vccd1 vccd1 _04801_ sky130_fd_sc_hd__a21o_1
XFILLER_0_51_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12312_ _05835_ genblk1\[11\].osc.clkdiv_C.cnt\[2\] vssd1 vssd1 vccd1 vccd1 _06013_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_23_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13292_ clknet_leaf_88_clk _00613_ net177 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.b1\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_32_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12243_ genblk2\[11\].wave_shpr.div.acc\[25\] genblk2\[11\].wave_shpr.div.acc\[24\]
+ genblk2\[11\].wave_shpr.div.acc\[26\] _05980_ vssd1 vssd1 vccd1 vccd1 _05981_ sky130_fd_sc_hd__or4_2
XFILLER_0_20_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12174_ _05916_ vssd1 vssd1 vccd1 vccd1 _01002_ sky130_fd_sc_hd__clkbuf_1
X_11125_ _05033_ genblk2\[7\].wave_shpr.div.acc\[1\] _05184_ vssd1 vssd1 vccd1 vccd1
+ _05185_ sky130_fd_sc_hd__a21o_1
X_11056_ genblk2\[6\].wave_shpr.div.acc\[15\] _05131_ _05105_ vssd1 vssd1 vccd1 vccd1
+ _05132_ sky130_fd_sc_hd__mux2_1
XFILLER_0_155_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10007_ genblk2\[3\].wave_shpr.div.b1\[12\] genblk2\[3\].wave_shpr.div.acc\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04403_ sky130_fd_sc_hd__and2b_1
XFILLER_0_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12112__S _05865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08098__A _01440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10520__A2 _04657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11958_ genblk2\[10\].wave_shpr.div.b1\[17\] genblk2\[10\].wave_shpr.div.acc\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05780_ sky130_fd_sc_hd__and2b_1
XFILLER_0_80_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09674__B1 _03819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07730__A _01188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10909_ net1202 _04432_ _04848_ vssd1 vssd1 vccd1 vccd1 _05039_ sky130_fd_sc_hd__mux2_1
X_11889_ genblk2\[9\].wave_shpr.div.acc\[24\] vssd1 vssd1 vccd1 vccd1 _05718_ sky130_fd_sc_hd__inv_2
X_13628_ clknet_leaf_65_clk _00941_ net197 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.b1\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12025__A2 _05813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13559_ clknet_leaf_85_clk _00874_ net184 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.quo\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_07080_ genblk1\[8\].osc.clkdiv_C.cnt\[4\] _01892_ _01886_ vssd1 vssd1 vccd1 vccd1
+ _01894_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_81_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_777 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout107 net127 vssd1 vssd1 vccd1 vccd1 net107 sky130_fd_sc_hd__buf_2
Xfanout118 net126 vssd1 vssd1 vccd1 vccd1 net118 sky130_fd_sc_hd__buf_2
XFILLER_0_10_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout129 net131 vssd1 vssd1 vccd1 vccd1 net129 sky130_fd_sc_hd__clkbuf_2
X_07982_ genblk2\[7\].wave_shpr.div.fin_quo\[4\] _02688_ vssd1 vssd1 vccd1 vccd1 _02689_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__06963__A1 _01229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09721_ genblk2\[2\].wave_shpr.div.b1\[14\] genblk2\[2\].wave_shpr.div.acc\[14\]
+ vssd1 vssd1 vccd1 vccd1 _04201_ sky130_fd_sc_hd__and2b_1
X_06933_ genblk1\[6\].osc.clkdiv_C.cnt\[10\] genblk1\[6\].osc.clkdiv_C.cnt\[9\] _01773_
+ vssd1 vssd1 vccd1 vccd1 _01777_ sky130_fd_sc_hd__and3_1
X_09652_ net803 _04048_ _04113_ _04140_ vssd1 vssd1 vccd1 vccd1 _00256_ sky130_fd_sc_hd__a22o_1
X_06864_ genblk1\[5\].osc.clkdiv_C.cnt\[15\] genblk1\[5\].osc.clkdiv_C.cnt\[14\] _01717_
+ vssd1 vssd1 vccd1 vccd1 _01721_ sky130_fd_sc_hd__and3_1
XANTENNA__10511__A2 _04657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08603_ _03188_ _02885_ _03189_ vssd1 vssd1 vccd1 vccd1 _03310_ sky130_fd_sc_hd__o21ai_1
X_09583_ genblk2\[1\].wave_shpr.div.acc\[5\] _04088_ _04011_ vssd1 vssd1 vccd1 vccd1
+ _04089_ sky130_fd_sc_hd__mux2_1
X_06795_ _01325_ _01254_ vssd1 vssd1 vccd1 vccd1 _01667_ sky130_fd_sc_hd__or2_2
X_08534_ genblk2\[9\].wave_shpr.div.fin_quo\[0\] _02526_ _02308_ genblk2\[9\].wave_shpr.div.fin_quo\[1\]
+ _02310_ vssd1 vssd1 vccd1 vccd1 _03241_ sky130_fd_sc_hd__a221o_1
XTAP_1109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08465_ _03153_ _03152_ vssd1 vssd1 vccd1 vccd1 _03172_ sky130_fd_sc_hd__xnor2_2
XANTENNA__07140__B2 genblk1\[9\].osc.clkdiv_C.cnt\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07416_ _02159_ vssd1 vssd1 vccd1 vccd1 _00006_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08396_ genblk1\[2\].osc.clkdiv_C.cnt\[15\] _01349_ _01209_ genblk1\[2\].osc.clkdiv_C.cnt\[14\]
+ vssd1 vssd1 vccd1 vccd1 _03103_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_70_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10027__A1 _04420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11224__B1 _05250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07347_ _02092_ _02105_ _02106_ vssd1 vssd1 vccd1 vccd1 _02107_ sky130_fd_sc_hd__and3_1
XFILLER_0_116_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09567__A _04042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07278_ genblk1\[10\].osc.clkdiv_C.cnt\[10\] _02048_ vssd1 vssd1 vccd1 vccd1 _02050_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_115_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09017_ _03689_ vssd1 vssd1 vccd1 vccd1 _03690_ sky130_fd_sc_hd__buf_8
XFILLER_0_131_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06229_ freq_div.state\[2\] vssd1 vssd1 vccd1 vccd1 _01191_ sky130_fd_sc_hd__buf_4
XFILLER_0_20_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06703__B _01592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold150 smpl_rt_clkdiv.clkDiv_inst.cnt\[3\] vssd1 vssd1 vccd1 vccd1 net368 sky130_fd_sc_hd__dlygate4sd3_1
Xhold161 genblk2\[0\].wave_shpr.div.quo\[7\] vssd1 vssd1 vccd1 vccd1 net379 sky130_fd_sc_hd__dlygate4sd3_1
Xhold172 genblk2\[9\].wave_shpr.div.b1\[15\] vssd1 vssd1 vccd1 vccd1 net390 sky130_fd_sc_hd__dlygate4sd3_1
Xhold183 genblk2\[3\].wave_shpr.div.quo\[7\] vssd1 vssd1 vccd1 vccd1 net401 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_0_6 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold194 genblk2\[11\].wave_shpr.div.quo\[24\] vssd1 vssd1 vccd1 vccd1 net412 sky130_fd_sc_hd__dlygate4sd3_1
X_09919_ _04329_ _04204_ vssd1 vssd1 vccd1 vccd1 _04330_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08156__B1 _01576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12930_ clknet_leaf_116_clk _00009_ net150 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.done
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12861_ clknet_leaf_129_clk _00192_ net64 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.b1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11812_ genblk2\[9\].wave_shpr.div.acc\[4\] _05660_ _05613_ vssd1 vssd1 vccd1 vccd1
+ _05661_ sky130_fd_sc_hd__mux2_1
XTAP_2344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12792_ clknet_leaf_91_clk _00125_ net148 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.quo\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11743_ _02203_ vssd1 vssd1 vccd1 vccd1 _05623_ sky130_fd_sc_hd__clkbuf_4
XTAP_2399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11674_ genblk2\[9\].wave_shpr.div.acc\[5\] genblk2\[9\].wave_shpr.div.b1\[5\] vssd1
+ vssd1 vccd1 vccd1 _05566_ sky130_fd_sc_hd__or2b_1
XANTENNA__07682__A2 _01246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09959__A1 _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11215__B1 _05222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13413_ clknet_leaf_120_clk net528 net142 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.quo\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10625_ _04839_ vssd1 vssd1 vccd1 vccd1 _00530_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__06890__B1 _01739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10556_ _04633_ genblk2\[5\].wave_shpr.div.acc\[1\] _04783_ vssd1 vssd1 vccd1 vccd1
+ _04784_ sky130_fd_sc_hd__a21o_1
X_13344_ clknet_leaf_7_clk _00665_ net49 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.acc\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10487_ genblk2\[4\].wave_shpr.div.acc\[15\] _04730_ _04704_ vssd1 vssd1 vccd1 vccd1
+ _04731_ sky130_fd_sc_hd__mux2_1
X_13275_ clknet_leaf_12_clk _00596_ net54 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.i\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_121_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12226_ _05931_ _05962_ _05963_ vssd1 vssd1 vccd1 vccd1 _05964_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12157_ _05904_ _05905_ vssd1 vssd1 vccd1 vccd1 _05906_ sky130_fd_sc_hd__or2_1
X_11108_ genblk2\[7\].wave_shpr.div.acc\[13\] genblk2\[7\].wave_shpr.div.b1\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05168_ sky130_fd_sc_hd__or2b_1
X_12088_ net868 _05844_ _05850_ _05853_ vssd1 vssd1 vccd1 vccd1 _00979_ sky130_fd_sc_hd__a22o_1
XANTENNA__08147__B1 _01519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11039_ net838 _05086_ _05093_ _05118_ vssd1 vssd1 vccd1 vccd1 _00665_ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06580_ genblk1\[3\].osc.clkdiv_C.cnt\[12\] _01344_ genblk1\[3\].osc.clkdiv_C.cnt\[13\]
+ vssd1 vssd1 vccd1 vccd1 _01488_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07122__B2 genblk1\[9\].osc.clkdiv_C.cnt\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08250_ _02955_ _02956_ _02604_ vssd1 vssd1 vccd1 vccd1 _02957_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07673__A2 _02001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07201_ _01952_ _01985_ vssd1 vssd1 vccd1 vccd1 _01986_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08181_ genblk2\[3\].wave_shpr.div.fin_quo\[5\] _02885_ _02887_ vssd1 vssd1 vccd1
+ vccd1 _02888_ sky130_fd_sc_hd__or3b_1
XFILLER_0_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07132_ genblk1\[9\].osc.clkdiv_C.cnt\[16\] _01578_ _01349_ genblk1\[9\].osc.clkdiv_C.cnt\[15\]
+ vssd1 vssd1 vccd1 vccd1 _01932_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_42_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09387__A _03726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07063_ _01441_ _01878_ genblk1\[8\].osc.clkdiv_C.cnt\[2\] _01880_ vssd1 vssd1 vccd1
+ vccd1 _01881_ sky130_fd_sc_hd__a31o_1
XFILLER_0_113_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10980__A2 _05051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07965_ genblk1\[7\].osc.clkdiv_C.cnt\[15\] _01577_ _01675_ genblk1\[7\].osc.clkdiv_C.cnt\[13\]
+ _02671_ vssd1 vssd1 vccd1 vccd1 _02672_ sky130_fd_sc_hd__a221o_1
X_09704_ _04168_ _04182_ _04183_ vssd1 vssd1 vccd1 vccd1 _04184_ sky130_fd_sc_hd__a21o_1
XANTENNA__10061__A _03701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06916_ _01761_ _01765_ _01766_ vssd1 vssd1 vccd1 vccd1 genblk1\[6\].osc.clkdiv_C.next_cnt\[3\]
+ sky130_fd_sc_hd__nor3_1
X_07896_ net14 net136 _02365_ vssd1 vssd1 vccd1 vccd1 _02603_ sky130_fd_sc_hd__and3_1
X_09635_ net664 _04109_ _04113_ _04128_ vssd1 vssd1 vccd1 vccd1 _00251_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_4_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06847_ genblk1\[5\].osc.clkdiv_C.cnt\[9\] _01708_ vssd1 vssd1 vccd1 vccd1 _01710_
+ sky130_fd_sc_hd__and2_1
X_06778_ _01650_ _01648_ vssd1 vssd1 vccd1 vccd1 _01652_ sky130_fd_sc_hd__nor2_1
X_09566_ net990 _04043_ _04047_ _04075_ vssd1 vssd1 vccd1 vccd1 _00235_ sky130_fd_sc_hd__a22o_1
X_08517_ _03219_ _03223_ vssd1 vssd1 vccd1 vccd1 _03224_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09497_ _03701_ vssd1 vssd1 vccd1 vccd1 _04039_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_81_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07113__A1 genblk1\[8\].osc.clkdiv_C.cnt\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08185__B _02539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08448_ _02638_ _02639_ genblk2\[8\].wave_shpr.div.fin_quo\[3\] vssd1 vssd1 vccd1
+ vccd1 _03155_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07664__A2 _02336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08379_ genblk1\[2\].osc.clkdiv_C.cnt\[6\] _01433_ vssd1 vssd1 vccd1 vccd1 _03086_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10410_ _04058_ _01644_ vssd1 vssd1 vccd1 vccd1 _04674_ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11390_ genblk2\[8\].wave_shpr.div.acc\[9\] genblk2\[8\].wave_shpr.div.b1\[9\] vssd1
+ vssd1 vccd1 vccd1 _05366_ sky130_fd_sc_hd__or2b_1
XANTENNA__09810__B1 _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10341_ _03701_ vssd1 vssd1 vccd1 vccd1 _04637_ sky130_fd_sc_hd__buf_4
XFILLER_0_131_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13060_ clknet_leaf_21_clk _00387_ net95 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.quo\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10272_ genblk2\[4\].wave_shpr.div.b1\[1\] genblk2\[4\].wave_shpr.div.acc\[1\] vssd1
+ vssd1 vccd1 vccd1 _04584_ sky130_fd_sc_hd__xor2_1
X_12011_ _03687_ net424 _03717_ vssd1 vssd1 vccd1 vccd1 _00946_ sky130_fd_sc_hd__a21bo_1
X_12913_ clknet_leaf_34_clk _00244_ net106 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.acc\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xmax_cap7 _01760_ vssd1 vssd1 vccd1 vccd1 net1356 sky130_fd_sc_hd__buf_1
XTAP_2130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12844_ clknet_leaf_116_clk _00007_ net150 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.done
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10239__A1 _04451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12775_ clknet_leaf_41_clk _00108_ net123 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.b1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07104__A1 genblk1\[8\].osc.clkdiv_C.cnt\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08095__B _01196_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06608__B _01210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11726_ genblk2\[9\].wave_shpr.div.fin_quo\[2\] net1313 _00023_ vssd1 vssd1 vccd1
+ vccd1 _05616_ sky130_fd_sc_hd__mux2_1
XTAP_1484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11657_ _00020_ _05549_ net1164 vssd1 vssd1 vccd1 vccd1 _05551_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_52_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10608_ genblk2\[5\].wave_shpr.div.fin_quo\[7\] net1344 _00015_ vssd1 vssd1 vccd1
+ vccd1 _04829_ sky130_fd_sc_hd__mux2_1
XFILLER_0_3_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09801__B1 _04252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11588_ _05391_ _05501_ vssd1 vssd1 vccd1 vccd1 _05502_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_51_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold908 sig_norm.quo\[1\] vssd1 vssd1 vccd1 vccd1 net1126 sky130_fd_sc_hd__dlygate4sd3_1
X_13327_ clknet_leaf_25_clk net568 net86 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.quo\[21\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold919 genblk2\[2\].wave_shpr.div.acc\[2\] vssd1 vssd1 vccd1 vccd1 net1137 sky130_fd_sc_hd__dlygate4sd3_1
X_10539_ genblk2\[5\].wave_shpr.div.acc\[13\] genblk2\[5\].wave_shpr.div.b1\[13\]
+ vssd1 vssd1 vccd1 vccd1 _04767_ sky130_fd_sc_hd__or2b_1
XFILLER_0_150_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13258_ clknet_leaf_2_clk _00581_ net51 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.acc\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12209_ genblk2\[11\].wave_shpr.div.b1\[3\] genblk2\[11\].wave_shpr.div.acc\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05947_ sky130_fd_sc_hd__and2b_1
X_13189_ clknet_leaf_122_clk _00512_ net78 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.i\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__06394__A2 _01210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07750_ _02428_ _02453_ _02452_ _02456_ vssd1 vssd1 vccd1 vccd1 _02457_ sky130_fd_sc_hd__a31o_1
X_06701_ _01173_ _01175_ _01191_ vssd1 vssd1 vccd1 vccd1 _01591_ sky130_fd_sc_hd__or3b_4
X_07681_ _02387_ vssd1 vssd1 vccd1 vccd1 _02388_ sky130_fd_sc_hd__inv_2
XFILLER_0_126_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06632_ _01523_ _01533_ _01534_ vssd1 vssd1 vccd1 vccd1 genblk1\[3\].osc.clkdiv_C.next_cnt\[5\]
+ sky130_fd_sc_hd__nor3_1
X_09420_ genblk2\[1\].wave_shpr.div.b1\[7\] genblk2\[1\].wave_shpr.div.acc\[7\] vssd1
+ vssd1 vccd1 vccd1 _03984_ sky130_fd_sc_hd__and2b_1
XFILLER_0_149_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09351_ _03800_ net23 vssd1 vssd1 vccd1 vccd1 _03927_ sky130_fd_sc_hd__nor2_1
X_06563_ net1166 _01472_ _01475_ vssd1 vssd1 vccd1 vccd1 genblk1\[2\].osc.clkdiv_C.next_cnt\[13\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_19_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09096__A1 _01490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08302_ _02602_ _02924_ _02927_ _03008_ vssd1 vssd1 vccd1 vccd1 _03009_ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09282_ _03769_ _03760_ vssd1 vssd1 vccd1 vccd1 _03874_ sky130_fd_sc_hd__or2b_1
XFILLER_0_145_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06494_ _01242_ _01223_ vssd1 vssd1 vccd1 vccd1 _01420_ sky130_fd_sc_hd__nor2_2
XFILLER_0_74_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08233_ _02887_ _02885_ genblk2\[3\].wave_shpr.div.fin_quo\[5\] vssd1 vssd1 vccd1
+ vccd1 _02940_ sky130_fd_sc_hd__or3b_1
XFILLER_0_144_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08164_ _01181_ genblk1\[3\].osc.clkdiv_C.cnt\[9\] _01182_ vssd1 vssd1 vccd1 vccd1
+ _02871_ sky130_fd_sc_hd__and3_1
XFILLER_0_133_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07115_ genblk1\[8\].osc.clkdiv_C.cnt\[16\] _01914_ vssd1 vssd1 vccd1 vccd1 _01917_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08095_ _01650_ _01196_ vssd1 vssd1 vccd1 vccd1 _02802_ sky130_fd_sc_hd__nor2_1
XFILLER_0_70_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06253__B _01214_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10953__A2 _05057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09845__A _04269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07046_ genblk1\[8\].osc.clkdiv_C.cnt\[13\] _01328_ vssd1 vssd1 vccd1 vccd1 _01864_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_11_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09056__S _03708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08997_ _03678_ vssd1 vssd1 vccd1 vccd1 _00063_ sky130_fd_sc_hd__clkbuf_1
X_07948_ genblk1\[7\].osc.clkdiv_C.cnt\[7\] _01947_ _02652_ _02653_ _02654_ vssd1
+ vssd1 vccd1 vccd1 _02655_ sky130_fd_sc_hd__o221a_1
X_07879_ _02548_ _02561_ _02585_ vssd1 vssd1 vccd1 vccd1 _02586_ sky130_fd_sc_hd__or3_2
XANTENNA__06970__A2_N _01805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09618_ genblk2\[1\].wave_shpr.div.acc\[13\] _04115_ _04095_ vssd1 vssd1 vccd1 vccd1
+ _04116_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout43_A net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10890_ genblk2\[6\].wave_shpr.div.fin_quo\[5\] net720 _00017_ vssd1 vssd1 vccd1
+ vccd1 _05029_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09549_ genblk2\[1\].wave_shpr.div.quo\[21\] _04052_ _04053_ net257 _04065_ vssd1
+ vssd1 vccd1 vccd1 _00228_ sky130_fd_sc_hd__a221o_1
XFILLER_0_93_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12560_ clknet_leaf_57_clk genblk1\[0\].osc.clkdiv_C.next_cnt\[17\] net181 vssd1
+ vssd1 vccd1 vccd1 genblk1\[0\].osc.clkdiv_C.cnt\[17\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_53_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11511_ net329 _05448_ _05449_ net450 _05451_ vssd1 vssd1 vccd1 vccd1 _00804_ sky130_fd_sc_hd__a221o_1
XFILLER_0_136_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12491_ clknet_leaf_107_clk _00053_ net158 vssd1 vssd1 vccd1 vccd1 sig_norm.quo\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11442_ genblk2\[8\].wave_shpr.div.fin_quo\[0\] _05417_ _00021_ vssd1 vssd1 vccd1
+ vccd1 _05418_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08598__B1 _02467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11373_ genblk2\[7\].wave_shpr.div.i\[1\] genblk2\[7\].wave_shpr.div.i\[0\] genblk2\[7\].wave_shpr.div.i\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05352_ sky130_fd_sc_hd__a21o_1
XANTENNA_hold976_A genblk1\[9\].osc.clkdiv_C.cnt\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10944__A2 _05052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13112_ clknet_leaf_115_clk _00437_ net134 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.fin_quo\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10324_ genblk2\[4\].wave_shpr.div.fin_quo\[6\] genblk2\[4\].wave_shpr.div.quo\[5\]
+ _00013_ vssd1 vssd1 vccd1 vccd1 _04630_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13043_ clknet_leaf_128_clk _00370_ net66 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.b1\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10255_ genblk2\[4\].wave_shpr.div.acc\[15\] genblk2\[4\].wave_shpr.div.b1\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04567_ sky130_fd_sc_hd__or2b_1
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09562__A2 _04011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10186_ net942 _04486_ _04490_ _04517_ vssd1 vssd1 vccd1 vccd1 _00413_ sky130_fd_sc_hd__a22o_1
XANTENNA__08522__B1 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12827_ clknet_leaf_62_clk _00160_ net190 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.acc\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10880__A1 _05023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12758_ clknet_leaf_52_clk genblk1\[11\].osc.clkdiv_C.next_cnt\[17\] net110 vssd1
+ vssd1 vccd1 vccd1 genblk1\[11\].osc.clkdiv_C.cnt\[17\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__07628__A2 _01256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10632__A1 _01923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11709_ _05557_ _05599_ _05600_ vssd1 vssd1 vccd1 vccd1 _05601_ sky130_fd_sc_hd__a21o_1
XFILLER_0_71_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12689_ clknet_leaf_53_clk genblk1\[8\].osc.clkdiv_C.next_cnt\[2\] net174 vssd1 vssd1
+ vccd1 vccd1 genblk1\[8\].osc.clkdiv_C.cnt\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_126_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold705 genblk2\[7\].wave_shpr.div.acc\[20\] vssd1 vssd1 vccd1 vccd1 net923 sky130_fd_sc_hd__dlygate4sd3_1
Xhold716 genblk2\[0\].wave_shpr.div.acc\[10\] vssd1 vssd1 vccd1 vccd1 net934 sky130_fd_sc_hd__dlygate4sd3_1
Xhold727 genblk2\[10\].wave_shpr.div.acc\[14\] vssd1 vssd1 vccd1 vccd1 net945 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold738 genblk2\[0\].wave_shpr.div.acc\[9\] vssd1 vssd1 vccd1 vccd1 net956 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold749 genblk2\[9\].wave_shpr.div.acc\[13\] vssd1 vssd1 vccd1 vccd1 net967 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08920_ _03588_ _03602_ _03618_ vssd1 vssd1 vccd1 vccd1 _03619_ sky130_fd_sc_hd__o21ai_1
X_08851_ _03555_ _03556_ _03552_ vssd1 vssd1 vccd1 vccd1 _03558_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09553__A2 _04042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07802_ _02221_ net31 vssd1 vssd1 vccd1 vccd1 _02509_ sky130_fd_sc_hd__nor2_2
X_08782_ _03487_ _03488_ vssd1 vssd1 vccd1 vccd1 _03489_ sky130_fd_sc_hd__nand2_1
XANTENNA__09604__S _04095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11648__A0 _05444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07733_ _02430_ _02431_ _02432_ _02434_ _02439_ vssd1 vssd1 vccd1 vccd1 _02440_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_1_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07664_ genblk1\[10\].osc.clkdiv_C.cnt\[6\] _02336_ _01794_ genblk1\[10\].osc.clkdiv_C.cnt\[5\]
+ _01182_ vssd1 vssd1 vccd1 vccd1 _02371_ sky130_fd_sc_hd__a32o_1
XFILLER_0_95_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09403_ genblk2\[1\].wave_shpr.div.acc\[4\] genblk2\[1\].wave_shpr.div.b1\[4\] vssd1
+ vssd1 vccd1 vccd1 _03967_ sky130_fd_sc_hd__and2b_1
X_06615_ _01522_ vssd1 vssd1 vccd1 vccd1 _01523_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07595_ _02266_ _02277_ _02301_ genblk1\[9\].osc.clkdiv_C.cnt\[17\] genblk1\[9\].osc.clkdiv_C.cnt\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02302_ sky130_fd_sc_hd__a311oi_4
XFILLER_0_87_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09334_ _03793_ _03748_ vssd1 vssd1 vccd1 vccd1 _03914_ sky130_fd_sc_hd__or2b_1
XFILLER_0_47_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06546_ genblk1\[2\].osc.clkdiv_C.cnt\[8\] genblk1\[2\].osc.clkdiv_C.cnt\[7\] _01461_
+ vssd1 vssd1 vccd1 vccd1 _01464_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07619__A2 _01595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06477_ net29 _01405_ vssd1 vssd1 vccd1 vccd1 _01406_ sky130_fd_sc_hd__nor2_1
X_09265_ _03853_ genblk1\[0\].osc.clkdiv_C.cnt\[16\] vssd1 vssd1 vccd1 vccd1 _03862_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_7_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08216_ _02900_ _02922_ vssd1 vssd1 vccd1 vccd1 _02923_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_118_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09196_ net1224 _03712_ _03822_ vssd1 vssd1 vccd1 vccd1 _03826_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08147_ genblk1\[3\].osc.clkdiv_C.cnt\[1\] _01496_ _01519_ genblk1\[3\].osc.clkdiv_C.cnt\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02854_ sky130_fd_sc_hd__o211a_1
XFILLER_0_132_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08078_ genblk1\[5\].osc.clkdiv_C.cnt\[10\] _01667_ _02757_ vssd1 vssd1 vccd1 vccd1
+ _02785_ sky130_fd_sc_hd__or3_1
XFILLER_0_101_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07029_ genblk1\[7\].osc.clkdiv_C.cnt\[16\] _01847_ vssd1 vssd1 vccd1 vccd1 _01849_
+ sky130_fd_sc_hd__or2_1
X_10040_ _04429_ vssd1 vssd1 vccd1 vccd1 _00355_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold10 modein.delay_octave_up_in\[0\] vssd1 vssd1 vccd1 vccd1 net228 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 genblk2\[11\].wave_shpr.div.quo\[20\] vssd1 vssd1 vccd1 vccd1 net239 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 _00558_ vssd1 vssd1 vccd1 vccd1 net250 sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 genblk2\[2\].wave_shpr.div.quo\[21\] vssd1 vssd1 vccd1 vccd1 net261 sky130_fd_sc_hd__dlygate4sd3_1
Xhold54 _00631_ vssd1 vssd1 vccd1 vccd1 net272 sky130_fd_sc_hd__dlygate4sd3_1
Xhold65 genblk2\[6\].wave_shpr.div.acc_next\[0\] vssd1 vssd1 vccd1 vccd1 net283 sky130_fd_sc_hd__dlygate4sd3_1
Xhold76 genblk2\[5\].wave_shpr.div.quo\[13\] vssd1 vssd1 vccd1 vccd1 net294 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11639__B1 _05417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold87 _00881_ vssd1 vssd1 vccd1 vccd1 net305 sky130_fd_sc_hd__dlygate4sd3_1
Xhold98 _00307_ vssd1 vssd1 vccd1 vccd1 net316 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11991_ _05800_ vssd1 vssd1 vccd1 vccd1 _00935_ sky130_fd_sc_hd__clkbuf_1
X_13730_ clknet_leaf_74_clk _01041_ net212 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.quo\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10942_ net271 _05052_ _05056_ net671 vssd1 vssd1 vccd1 vccd1 _00630_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13661_ clknet_leaf_47_clk _00974_ net120 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.acc_next\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10873_ _04966_ _05015_ _05016_ vssd1 vssd1 vccd1 vccd1 _05017_ sky130_fd_sc_hd__a21o_1
X_12612_ clknet_leaf_23_clk genblk1\[3\].osc.clkdiv_C.next_cnt\[15\] net94 vssd1 vssd1
+ vccd1 vccd1 genblk1\[3\].osc.clkdiv_C.cnt\[15\] sky130_fd_sc_hd__dfrtp_4
X_13592_ clknet_leaf_72_clk _00907_ net216 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.acc\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06818__B1 _01675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12543_ clknet_leaf_60_clk genblk1\[0\].osc.clkdiv_C.next_cnt\[0\] net187 vssd1 vssd1
+ vccd1 vccd1 genblk1\[0\].osc.clkdiv_C.cnt\[0\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__09480__A1 _04028_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10090__A2 _04452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12474_ clknet_leaf_116_clk FSM.next_mode\[0\] net150 vssd1 vssd1 vccd1 vccd1 net17
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA_clkbuf_leaf_91_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11425_ _05362_ _05399_ _05400_ vssd1 vssd1 vccd1 vccd1 _05401_ sky130_fd_sc_hd__a21o_1
XFILLER_0_151_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_7 _04242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11356_ genblk2\[7\].wave_shpr.div.acc\[22\] _05218_ _05340_ vssd1 vssd1 vccd1 vccd1
+ _05341_ sky130_fd_sc_hd__a21o_1
XFILLER_0_120_842 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10307_ genblk2\[4\].wave_shpr.div.acc\[21\] genblk2\[4\].wave_shpr.div.acc\[20\]
+ _04617_ _04618_ vssd1 vssd1 vccd1 vccd1 _04619_ sky130_fd_sc_hd__or4_1
XANTENNA__07717__B _02364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11287_ _05191_ _05176_ vssd1 vssd1 vccd1 vccd1 _05289_ sky130_fd_sc_hd__or2b_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13026_ clknet_leaf_113_clk _00353_ net134 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.fin_quo\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10238_ net375 _04457_ _04454_ _04555_ vssd1 vssd1 vccd1 vccd1 _00427_ sky130_fd_sc_hd__a22o_1
X_10169_ net966 _04486_ _04490_ _04504_ vssd1 vssd1 vccd1 vccd1 _00409_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06349__A genblk1\[0\].osc.clkdiv_C.cnt\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_44_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06400_ _01343_ vssd1 vssd1 vccd1 vccd1 _01344_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_29_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07380_ genblk1\[11\].osc.clkdiv_C.cnt\[12\] _02130_ vssd1 vssd1 vccd1 vccd1 _02132_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_128_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06331_ genblk1\[0\].osc.clkdiv_C.cnt\[7\] _01281_ genblk1\[0\].osc.clkdiv_C.cnt\[8\]
+ vssd1 vssd1 vccd1 vccd1 _01285_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_29_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09050_ _03708_ vssd1 vssd1 vccd1 vccd1 _03714_ sky130_fd_sc_hd__buf_8
XFILLER_0_32_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06262_ _01220_ _01221_ _01223_ vssd1 vssd1 vccd1 vccd1 _01224_ sky130_fd_sc_hd__a21oi_4
XANTENNA_clkbuf_leaf_59_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08001_ genblk1\[6\].osc.clkdiv_C.cnt\[15\] _01577_ _01675_ genblk1\[6\].osc.clkdiv_C.cnt\[13\]
+ _02707_ vssd1 vssd1 vccd1 vccd1 _02708_ sky130_fd_sc_hd__a221o_1
XFILLER_0_114_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06193_ _01159_ net832 vssd1 vssd1 vccd1 vccd1 PWM.next_counter\[2\] sky130_fd_sc_hd__nor2_1
XFILLER_0_53_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_102_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold502 genblk2\[6\].wave_shpr.div.quo\[4\] vssd1 vssd1 vccd1 vccd1 net720 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold513 genblk2\[11\].wave_shpr.div.quo\[5\] vssd1 vssd1 vccd1 vccd1 net731 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold524 genblk2\[6\].wave_shpr.div.quo\[5\] vssd1 vssd1 vccd1 vccd1 net742 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_399 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06812__A _01189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold535 _00234_ vssd1 vssd1 vccd1 vccd1 net753 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold546 genblk2\[1\].wave_shpr.div.quo\[0\] vssd1 vssd1 vccd1 vccd1 net764 sky130_fd_sc_hd__buf_1
XFILLER_0_40_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold557 genblk2\[0\].wave_shpr.div.i\[2\] vssd1 vssd1 vccd1 vccd1 net775 sky130_fd_sc_hd__dlygate4sd3_1
Xhold568 genblk2\[0\].wave_shpr.div.acc\[17\] vssd1 vssd1 vccd1 vccd1 net786 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09952_ _04352_ vssd1 vssd1 vccd1 vccd1 _00344_ sky130_fd_sc_hd__clkbuf_1
Xhold579 genblk2\[7\].wave_shpr.div.acc\[10\] vssd1 vssd1 vccd1 vccd1 net797 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08903_ _03574_ _03604_ _03606_ _01157_ net1065 vssd1 vssd1 vccd1 vccd1 _00041_ sky130_fd_sc_hd__a32o_1
XANTENNA_clkbuf_leaf_117_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09883_ net903 _04282_ _04289_ _04302_ vssd1 vssd1 vccd1 vccd1 _00325_ sky130_fd_sc_hd__a22o_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08834_ genblk2\[2\].wave_shpr.div.fin_quo\[0\] _02468_ _03114_ vssd1 vssd1 vccd1
+ vccd1 _03541_ sky130_fd_sc_hd__a21o_1
XTAP_884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08765_ _03471_ _03468_ vssd1 vssd1 vccd1 vccd1 _03472_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09561__C _04011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07716_ _02315_ _02421_ _02422_ vssd1 vssd1 vccd1 vccd1 _02423_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12294__B1 _03733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08696_ _03355_ _03353_ vssd1 vssd1 vccd1 vccd1 _03403_ sky130_fd_sc_hd__and2b_1
XFILLER_0_73_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07647_ genblk2\[11\].wave_shpr.div.fin_quo\[3\] _02353_ vssd1 vssd1 vccd1 vccd1
+ _02354_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07578_ genblk1\[9\].osc.clkdiv_C.cnt\[7\] _01234_ vssd1 vssd1 vccd1 vccd1 _02285_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_153_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09317_ _03784_ _03900_ vssd1 vssd1 vccd1 vccd1 _03901_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_91_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06529_ _01452_ _01453_ vssd1 vssd1 vccd1 vccd1 genblk1\[2\].osc.clkdiv_C.next_cnt\[1\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_118_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06706__B _01595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09248_ net410 _03845_ _03847_ net522 _03852_ vssd1 vssd1 vccd1 vccd1 _00140_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_4_10_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_10_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_121_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09179_ _03816_ vssd1 vssd1 vccd1 vccd1 _00107_ sky130_fd_sc_hd__clkbuf_1
X_11210_ _05244_ vssd1 vssd1 vccd1 vccd1 _00710_ sky130_fd_sc_hd__clkbuf_1
X_12190_ genblk2\[11\].wave_shpr.div.acc\[14\] genblk2\[11\].wave_shpr.div.b1\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05928_ sky130_fd_sc_hd__or2b_1
XFILLER_0_31_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11141_ genblk2\[7\].wave_shpr.div.b1\[10\] genblk2\[7\].wave_shpr.div.acc\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05201_ sky130_fd_sc_hd__and2b_1
XFILLER_0_101_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11072_ net1138 _05119_ _05126_ _05143_ vssd1 vssd1 vccd1 vccd1 _00673_ sky130_fd_sc_hd__a22o_1
XANTENNA__09517__A2 _04043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10023_ _04417_ _04418_ vssd1 vssd1 vccd1 vccd1 _04419_ sky130_fd_sc_hd__or2_1
XANTENNA__07553__A _01157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11974_ genblk2\[10\].wave_shpr.div.fin_quo\[4\] net1323 _00003_ vssd1 vssd1 vccd1
+ vccd1 _05792_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_317 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13713_ clknet_leaf_31_clk _01024_ net99 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.b1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10925_ _05047_ vssd1 vssd1 vccd1 vccd1 _00622_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__06503__A2 _01411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13644_ clknet_leaf_69_clk net321 net211 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.quo\[8\]
+ sky130_fd_sc_hd__dfrtp_4
X_10856_ genblk2\[6\].wave_shpr.div.b1\[9\] genblk2\[6\].wave_shpr.div.acc\[9\] vssd1
+ vssd1 vccd1 vccd1 _05000_ sky130_fd_sc_hd__and2b_1
XFILLER_0_85_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13575_ clknet_leaf_84_clk net307 net183 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.acc_next\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10787_ net982 _04918_ _04922_ _04942_ vssd1 vssd1 vccd1 vccd1 _00589_ sky130_fd_sc_hd__a22o_1
XANTENNA__10419__A _04654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12526_ clknet_leaf_66_clk _00078_ net197 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.b1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09205__A1 _03704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12457_ clknet_leaf_106_clk _00030_ net155 vssd1 vssd1 vccd1 vccd1 PWM.final_sample_in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11408_ genblk2\[8\].wave_shpr.div.b1\[5\] genblk2\[8\].wave_shpr.div.acc\[5\] vssd1
+ vssd1 vccd1 vccd1 _05384_ sky130_fd_sc_hd__and2b_1
XANTENNA__07728__A _01342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12388_ _05961_ _05932_ vssd1 vssd1 vccd1 vccd1 _06063_ sky130_fd_sc_hd__or2b_1
XANTENNA__07767__A1 genblk1\[0\].osc.clkdiv_C.cnt\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07767__B2 genblk1\[0\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11339_ _05214_ _05328_ vssd1 vssd1 vccd1 vccd1 _05329_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09508__A2 _04043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11315__A2 _05279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13009_ clknet_leaf_133_clk _00338_ net59 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.acc\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_06880_ _01729_ _01684_ _01730_ genblk1\[6\].osc.clkdiv_C.cnt\[4\] _01733_ vssd1
+ vssd1 vccd1 vccd1 _01734_ sky130_fd_sc_hd__a221o_1
X_08550_ _03245_ _03235_ vssd1 vssd1 vccd1 vccd1 _03257_ sky130_fd_sc_hd__xor2_1
XFILLER_0_77_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07501_ net17 net18 vssd1 vssd1 vccd1 vccd1 _02222_ sky130_fd_sc_hd__nand2b_4
X_08481_ genblk2\[3\].wave_shpr.div.fin_quo\[0\] vssd1 vssd1 vccd1 vccd1 _03188_ sky130_fd_sc_hd__inv_2
X_07432_ _02170_ vssd1 vssd1 vccd1 vccd1 _02171_ sky130_fd_sc_hd__buf_8
XANTENNA__12028__B1 _05817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_84 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07363_ genblk1\[11\].osc.clkdiv_C.cnt\[8\] genblk1\[11\].osc.clkdiv_C.cnt\[7\] _02112_
+ vssd1 vssd1 vccd1 vccd1 _02119_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09102_ genblk2\[0\].wave_shpr.div.acc\[13\] genblk2\[0\].wave_shpr.div.b1\[13\]
+ vssd1 vssd1 vccd1 vccd1 _03750_ sky130_fd_sc_hd__or2b_1
XFILLER_0_73_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06314_ genblk1\[0\].osc.clkdiv_C.cnt\[2\] genblk1\[0\].osc.clkdiv_C.cnt\[1\] genblk1\[0\].osc.clkdiv_C.cnt\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01274_ sky130_fd_sc_hd__and3_1
XFILLER_0_33_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07294_ genblk1\[10\].osc.clkdiv_C.cnt\[16\] _02058_ vssd1 vssd1 vccd1 vccd1 _02060_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_33_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06245_ freq_div.state\[0\] freq_div.state\[2\] freq_div.state\[1\] vssd1 vssd1 vccd1
+ vccd1 _01207_ sky130_fd_sc_hd__or3b_1
X_09033_ net817 _02202_ _03698_ _03702_ vssd1 vssd1 vccd1 vccd1 _03703_ sky130_fd_sc_hd__a31o_1
XFILLER_0_60_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout210_A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06176_ _01139_ _01133_ _01137_ vssd1 vssd1 vccd1 vccd1 _01148_ sky130_fd_sc_hd__and3_1
Xhold310 _00732_ vssd1 vssd1 vccd1 vccd1 net528 sky130_fd_sc_hd__dlygate4sd3_1
Xhold321 _00384_ vssd1 vssd1 vccd1 vccd1 net539 sky130_fd_sc_hd__dlygate4sd3_1
Xhold332 genblk2\[7\].wave_shpr.div.quo\[15\] vssd1 vssd1 vccd1 vccd1 net550 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold343 genblk2\[3\].wave_shpr.div.quo\[24\] vssd1 vssd1 vccd1 vccd1 net561 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold354 genblk2\[5\].wave_shpr.div.quo\[10\] vssd1 vssd1 vccd1 vccd1 net572 sky130_fd_sc_hd__dlygate4sd3_1
Xhold365 genblk2\[10\].wave_shpr.div.quo\[12\] vssd1 vssd1 vccd1 vccd1 net583 sky130_fd_sc_hd__dlygate4sd3_1
Xhold376 genblk2\[6\].wave_shpr.div.quo\[15\] vssd1 vssd1 vccd1 vccd1 net594 sky130_fd_sc_hd__dlygate4sd3_1
Xhold387 genblk2\[2\].wave_shpr.div.acc\[19\] vssd1 vssd1 vccd1 vccd1 net605 sky130_fd_sc_hd__dlygate4sd3_1
Xhold398 genblk2\[6\].wave_shpr.div.quo\[21\] vssd1 vssd1 vccd1 vccd1 net616 sky130_fd_sc_hd__dlygate4sd3_1
X_09935_ net1034 _04315_ _04322_ _04341_ vssd1 vssd1 vccd1 vccd1 _00338_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08707__B1 _02224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12911__RESET_B net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09866_ _04250_ vssd1 vssd1 vccd1 vccd1 _04289_ sky130_fd_sc_hd__clkbuf_4
Xhold1010 genblk2\[1\].wave_shpr.div.acc\[25\] vssd1 vssd1 vccd1 vccd1 net1228 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10514__B1 _04655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1021 genblk2\[9\].wave_shpr.div.b1\[17\] vssd1 vssd1 vccd1 vccd1 net1239 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09380__B1 _03947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08817_ _03518_ _03521_ _03517_ vssd1 vssd1 vccd1 vccd1 _03524_ sky130_fd_sc_hd__a21o_1
Xhold1032 genblk2\[7\].wave_shpr.div.b1\[3\] vssd1 vssd1 vccd1 vccd1 net1250 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1043 sig_norm.quo\[10\] vssd1 vssd1 vccd1 vccd1 net1261 sky130_fd_sc_hd__dlygate4sd3_1
X_09797_ _04250_ vssd1 vssd1 vccd1 vccd1 _04251_ sky130_fd_sc_hd__clkbuf_4
Xhold1054 genblk2\[1\].wave_shpr.div.b1\[5\] vssd1 vssd1 vccd1 vccd1 net1272 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1065 genblk2\[5\].wave_shpr.div.b1\[10\] vssd1 vssd1 vccd1 vccd1 net1283 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1076 genblk2\[9\].wave_shpr.div.b1\[2\] vssd1 vssd1 vccd1 vccd1 net1294 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1087 genblk2\[0\].wave_shpr.div.acc\[24\] vssd1 vssd1 vccd1 vccd1 net1305 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08748_ net14 _02744_ _02365_ vssd1 vssd1 vccd1 vccd1 _03455_ sky130_fd_sc_hd__nand3_1
Xhold1098 genblk2\[1\].wave_shpr.div.quo\[3\] vssd1 vssd1 vccd1 vccd1 net1316 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08486__A2 _02467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08679_ _02584_ _03385_ vssd1 vssd1 vccd1 vccd1 _03386_ sky130_fd_sc_hd__xnor2_2
XTAP_1825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10710_ _04783_ _04883_ vssd1 vssd1 vccd1 vccd1 _04884_ sky130_fd_sc_hd__nor2_1
XTAP_1847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11690_ genblk2\[9\].wave_shpr.div.b1\[5\] genblk2\[9\].wave_shpr.div.acc\[5\] vssd1
+ vssd1 vccd1 vccd1 _05582_ sky130_fd_sc_hd__and2b_1
XFILLER_0_95_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10641_ _03707_ vssd1 vssd1 vccd1 vccd1 _04848_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_107_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13360_ clknet_leaf_116_clk _00019_ net139 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.done
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10572_ genblk2\[5\].wave_shpr.div.b1\[10\] genblk2\[5\].wave_shpr.div.acc\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04800_ sky130_fd_sc_hd__and2b_1
XFILLER_0_118_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12311_ net467 _03947_ _03944_ net479 _06012_ vssd1 vssd1 vccd1 vccd1 _01043_ sky130_fd_sc_hd__a221o_1
XFILLER_0_134_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13291_ clknet_leaf_88_clk _00612_ net177 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.b1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12242_ genblk2\[11\].wave_shpr.div.acc\[23\] _05979_ vssd1 vssd1 vccd1 vccd1 _05980_
+ sky130_fd_sc_hd__or2_2
XANTENNA__06452__A genblk1\[1\].osc.clkdiv_C.cnt\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12173_ _05815_ _05812_ genblk2\[10\].wave_shpr.div.i\[0\] vssd1 vssd1 vccd1 vccd1
+ _05916_ sky130_fd_sc_hd__mux2_1
X_11124_ genblk2\[7\].wave_shpr.div.b1\[0\] _05182_ _05183_ vssd1 vssd1 vccd1 vccd1
+ _05184_ sky130_fd_sc_hd__a21oi_1
X_11055_ _05011_ _05130_ vssd1 vssd1 vccd1 vccd1 _05131_ sky130_fd_sc_hd__xnor2_1
X_10006_ _04367_ _04400_ _04401_ vssd1 vssd1 vccd1 vccd1 _04402_ sky130_fd_sc_hd__a21o_1
XANTENNA__11517__B genblk1\[8\].osc.clkdiv_C.cnt\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11009__S _05023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08098__B _01576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11957_ _05732_ _05777_ _05778_ vssd1 vssd1 vccd1 vccd1 _05779_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_98_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10908_ _05038_ vssd1 vssd1 vccd1 vccd1 _00614_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07730__B genblk1\[1\].osc.clkdiv_C.cnt\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11888_ _03694_ _05611_ _05717_ _03696_ net1026 vssd1 vssd1 vccd1 vccd1 _00915_ sky130_fd_sc_hd__a32o_1
XFILLER_0_39_372 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13627_ clknet_leaf_66_clk _00940_ net197 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.b1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10839_ genblk2\[6\].wave_shpr.div.acc\[0\] genblk2\[6\].wave_shpr.div.b1\[0\] vssd1
+ vssd1 vccd1 vccd1 _04983_ sky130_fd_sc_hd__and2b_1
XFILLER_0_82_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13558_ clknet_leaf_78_clk _00873_ net208 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.quo\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_89_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11784__A2 _02203_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12509_ clknet_leaf_84_clk _00071_ net202 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.i\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_140_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13489_ clknet_leaf_88_clk net470 net177 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.quo\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08401__A2 _01591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout108 net109 vssd1 vssd1 vccd1 vccd1 net108 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09673__A _03690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07981_ _02684_ _02687_ vssd1 vssd1 vccd1 vccd1 _02688_ sky130_fd_sc_hd__nand2_1
Xfanout119 net122 vssd1 vssd1 vccd1 vccd1 net119 sky130_fd_sc_hd__clkbuf_4
X_09720_ _04160_ _04198_ _04199_ vssd1 vssd1 vccd1 vccd1 _04200_ sky130_fd_sc_hd__a21o_1
X_06932_ _01761_ _01775_ _01776_ vssd1 vssd1 vccd1 vccd1 genblk1\[6\].osc.clkdiv_C.next_cnt\[9\]
+ sky130_fd_sc_hd__nor3_1
XANTENNA__10612__A _01738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07905__B _01870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09651_ genblk2\[1\].wave_shpr.div.acc\[22\] _04139_ vssd1 vssd1 vccd1 vccd1 _04140_
+ sky130_fd_sc_hd__xnor2_1
X_06863_ genblk1\[5\].osc.clkdiv_C.cnt\[14\] _01717_ _01720_ vssd1 vssd1 vccd1 vccd1
+ genblk1\[5\].osc.clkdiv_C.next_cnt\[14\] sky130_fd_sc_hd__o21a_1
X_08602_ _03188_ _03189_ _02885_ vssd1 vssd1 vccd1 vccd1 _03309_ sky130_fd_sc_hd__nor3_1
XFILLER_0_78_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09582_ _04087_ _03979_ vssd1 vssd1 vccd1 vccd1 _04088_ sky130_fd_sc_hd__xnor2_1
X_06794_ _01440_ _01171_ vssd1 vssd1 vccd1 vccd1 _01666_ sky130_fd_sc_hd__nand2_4
XFILLER_0_54_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07921__A genblk1\[8\].osc.clkdiv_C.cnt\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08533_ _03237_ _03239_ vssd1 vssd1 vccd1 vccd1 _03240_ sky130_fd_sc_hd__xnor2_1
XANTENNA__13599__RESET_B net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06693__A2_N _01313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08464_ _03163_ _03164_ _03169_ vssd1 vssd1 vccd1 vccd1 _03171_ sky130_fd_sc_hd__a21o_1
XFILLER_0_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07140__A2 _01334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07415_ _02155_ _02158_ vssd1 vssd1 vccd1 vccd1 _02159_ sky130_fd_sc_hd__nor2_1
X_08395_ genblk1\[2\].osc.clkdiv_C.cnt\[10\] _01420_ _03099_ _03100_ _03101_ vssd1
+ vssd1 vccd1 vccd1 _03102_ sky130_fd_sc_hd__o221a_1
XANTENNA__13181__RESET_B net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09848__A _03702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07346_ genblk1\[11\].osc.clkdiv_C.cnt\[4\] _02101_ vssd1 vssd1 vccd1 vccd1 _02106_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_73_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07277_ _02027_ _02048_ _02049_ vssd1 vssd1 vccd1 vccd1 genblk1\[10\].osc.clkdiv_C.next_cnt\[9\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_115_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09016_ _02155_ vssd1 vssd1 vccd1 vccd1 _03689_ sky130_fd_sc_hd__buf_4
XANTENNA__09059__S _03719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06228_ _01186_ _01189_ vssd1 vssd1 vccd1 vccd1 _01190_ sky130_fd_sc_hd__nor2_4
XFILLER_0_103_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06159_ _01114_ _01116_ vssd1 vssd1 vccd1 vccd1 _01131_ sky130_fd_sc_hd__nand2_1
Xhold140 genblk2\[11\].wave_shpr.div.quo\[7\] vssd1 vssd1 vccd1 vccd1 net358 sky130_fd_sc_hd__dlygate4sd3_1
Xhold151 genblk2\[2\].wave_shpr.div.b1\[15\] vssd1 vssd1 vccd1 vccd1 net369 sky130_fd_sc_hd__dlygate4sd3_1
Xhold162 smpl_rt_clkdiv.clkDiv_inst.cnt\[4\] vssd1 vssd1 vccd1 vccd1 net380 sky130_fd_sc_hd__dlygate4sd3_1
Xhold173 genblk2\[8\].wave_shpr.div.b1\[15\] vssd1 vssd1 vccd1 vccd1 net391 sky130_fd_sc_hd__dlygate4sd3_1
Xhold184 genblk2\[11\].wave_shpr.div.quo\[2\] vssd1 vssd1 vccd1 vccd1 net402 sky130_fd_sc_hd__dlygate4sd3_1
Xhold195 _01058_ vssd1 vssd1 vccd1 vccd1 net413 sky130_fd_sc_hd__dlygate4sd3_1
X_09918_ _04205_ _04157_ vssd1 vssd1 vccd1 vccd1 _04329_ sky130_fd_sc_hd__or2b_1
XANTENNA_fanout73_A net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09849_ genblk2\[2\].wave_shpr.div.acc\[0\] _00008_ _04275_ net914 _04276_ vssd1
+ vssd1 vccd1 vccd1 _00317_ sky130_fd_sc_hd__o221a_1
X_12860_ clknet_leaf_129_clk _00191_ net64 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.b1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08927__A _01099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11811_ _05569_ _05580_ vssd1 vssd1 vccd1 vccd1 _05660_ sky130_fd_sc_hd__xor2_1
XTAP_2334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12791_ clknet_leaf_91_clk _00124_ net146 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.quo\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11742_ _02248_ _01144_ _05622_ net1088 vssd1 vssd1 vccd1 vccd1 _00864_ sky130_fd_sc_hd__a22o_1
XFILLER_0_68_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11673_ genblk2\[9\].wave_shpr.div.acc\[6\] genblk2\[9\].wave_shpr.div.b1\[6\] vssd1
+ vssd1 vccd1 vccd1 _05565_ sky130_fd_sc_hd__or2b_1
XFILLER_0_154_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13412_ clknet_leaf_120_clk net232 net142 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.quo\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10624_ genblk2\[6\].wave_shpr.div.b1\[5\] _04838_ _04834_ vssd1 vssd1 vccd1 vccd1
+ _04839_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11215__B2 _05248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13343_ clknet_leaf_7_clk _00664_ net49 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.acc\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10555_ genblk2\[5\].wave_shpr.div.b1\[0\] _04781_ _04782_ vssd1 vssd1 vccd1 vccd1
+ _04783_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_91_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12184__A _03690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13274_ clknet_leaf_118_clk _00017_ net138 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.done
+ sky130_fd_sc_hd__dfrtp_1
X_10486_ _04611_ _04729_ vssd1 vssd1 vccd1 vccd1 _04730_ sky130_fd_sc_hd__xnor2_1
X_12225_ genblk2\[11\].wave_shpr.div.b1\[11\] genblk2\[11\].wave_shpr.div.acc\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05963_ sky130_fd_sc_hd__and2b_1
XFILLER_0_121_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12156_ genblk2\[10\].wave_shpr.div.acc\[19\] _05900_ genblk2\[10\].wave_shpr.div.acc\[20\]
+ vssd1 vssd1 vccd1 vccd1 _05905_ sky130_fd_sc_hd__o21a_1
X_11107_ genblk2\[7\].wave_shpr.div.acc\[14\] genblk2\[7\].wave_shpr.div.b1\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05167_ sky130_fd_sc_hd__or2b_1
XFILLER_0_75_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12087_ genblk2\[10\].wave_shpr.div.acc\[3\] _05852_ _05787_ vssd1 vssd1 vccd1 vccd1
+ _05853_ sky130_fd_sc_hd__mux2_1
X_11038_ genblk2\[6\].wave_shpr.div.acc\[11\] _05117_ _05105_ vssd1 vssd1 vccd1 vccd1
+ _05118_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12989_ clknet_leaf_132_clk _00318_ net64 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.acc\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07122__A2 _01334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07200_ genblk1\[9\].osc.clkdiv_C.cnt\[15\] genblk1\[9\].osc.clkdiv_C.cnt\[14\] _01981_
+ vssd1 vssd1 vccd1 vccd1 _01985_ sky130_fd_sc_hd__and3_1
XANTENNA__11206__A1 _03831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08180_ genblk2\[3\].wave_shpr.div.fin_quo\[4\] _02886_ vssd1 vssd1 vccd1 vccd1 _02887_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_161 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11757__A2 _03696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07131_ _01930_ _01250_ vssd1 vssd1 vccd1 vccd1 _01931_ sky130_fd_sc_hd__nand2_1
XFILLER_0_125_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07062_ genblk1\[8\].osc.clkdiv_C.cnt\[6\] _01249_ _01879_ _01490_ genblk1\[8\].osc.clkdiv_C.cnt\[7\]
+ vssd1 vssd1 vccd1 vccd1 _01880_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_70_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10717__B1 _04857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08386__A1 _01200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07916__A genblk1\[8\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07964_ _02670_ vssd1 vssd1 vccd1 vccd1 _02671_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09703_ genblk2\[2\].wave_shpr.div.b1\[5\] genblk2\[2\].wave_shpr.div.acc\[5\] vssd1
+ vssd1 vccd1 vccd1 _04183_ sky130_fd_sc_hd__and2b_1
XANTENNA__08138__B2 _02527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06915_ genblk1\[6\].osc.clkdiv_C.cnt\[3\] _01763_ vssd1 vssd1 vccd1 vccd1 _01766_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07895_ _02423_ _02601_ vssd1 vssd1 vccd1 vccd1 _02602_ sky130_fd_sc_hd__nand2_1
X_09634_ genblk2\[1\].wave_shpr.div.acc\[17\] _04127_ _04010_ vssd1 vssd1 vccd1 vccd1
+ _04128_ sky130_fd_sc_hd__mux2_1
XANTENNA__10496__A2 _04715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06846_ _01693_ _01708_ _01709_ vssd1 vssd1 vccd1 vccd1 genblk1\[5\].osc.clkdiv_C.next_cnt\[8\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_78_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09565_ genblk2\[1\].wave_shpr.div.acc\[1\] _04074_ _04011_ vssd1 vssd1 vccd1 vccd1
+ _04075_ sky130_fd_sc_hd__mux2_1
X_06777_ _01650_ _01648_ _01651_ _01600_ vssd1 vssd1 vccd1 vccd1 genblk1\[4\].osc.clkdiv_C.next_cnt\[15\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08516_ _03220_ _03221_ _03219_ _03222_ vssd1 vssd1 vccd1 vccd1 _03223_ sky130_fd_sc_hd__a211oi_2
X_09496_ _04038_ vssd1 vssd1 vccd1 vccd1 _00202_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_65_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08447_ _03152_ _03153_ vssd1 vssd1 vccd1 vccd1 _03154_ sky130_fd_sc_hd__or2b_1
XFILLER_0_135_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07664__A3 _01794_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08378_ _03071_ _03074_ _03084_ vssd1 vssd1 vccd1 vccd1 _03085_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_80_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11748__A2 _05623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07329_ genblk1\[11\].osc.clkdiv_C.cnt\[0\] _02092_ vssd1 vssd1 vccd1 vccd1 _02093_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_104_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10340_ _03714_ net1097 _04432_ _03727_ vssd1 vssd1 vccd1 vccd1 _00448_ sky130_fd_sc_hd__o22a_1
X_10271_ genblk2\[4\].wave_shpr.div.acc\[0\] vssd1 vssd1 vccd1 vccd1 _04583_ sky130_fd_sc_hd__inv_2
XANTENNA__10708__B1 _04858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12010_ _03732_ net384 _03733_ vssd1 vssd1 vccd1 vccd1 _00945_ sky130_fd_sc_hd__o21a_1
X_12912_ clknet_leaf_34_clk _00243_ net107 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.acc\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12843_ clknet_leaf_30_clk _00006_ net104 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.busy
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12774_ clknet_leaf_44_clk _00107_ net120 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.b1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11725_ _05615_ vssd1 vssd1 vccd1 vccd1 _00854_ sky130_fd_sc_hd__clkbuf_1
XTAP_1474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11656_ _05449_ _05548_ _05550_ _05448_ net726 vssd1 vssd1 vccd1 vccd1 _00850_ sky130_fd_sc_hd__a32o_1
Xfanout90 net91 vssd1 vssd1 vccd1 vccd1 net90 sky130_fd_sc_hd__clkbuf_4
X_10607_ _04828_ vssd1 vssd1 vccd1 vccd1 _00523_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11587_ _05392_ _05366_ vssd1 vssd1 vccd1 vccd1 _05501_ sky130_fd_sc_hd__or2b_1
XFILLER_0_3_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10947__B1 _05056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13326_ clknet_leaf_25_clk net314 net86 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.quo\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10538_ genblk2\[5\].wave_shpr.div.acc\[14\] genblk2\[5\].wave_shpr.div.b1\[14\]
+ vssd1 vssd1 vccd1 vccd1 _04766_ sky130_fd_sc_hd__or2b_1
XANTENNA__10411__A2 _04651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold909 genblk2\[11\].wave_shpr.div.acc\[2\] vssd1 vssd1 vccd1 vccd1 net1127 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13257_ clknet_leaf_3_clk _00580_ net46 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.acc\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09014__C1 _03687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10469_ _04603_ _04716_ vssd1 vssd1 vccd1 vccd1 _04717_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_110_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12208_ _05940_ genblk2\[11\].wave_shpr.div.acc\[2\] _05945_ vssd1 vssd1 vccd1 vccd1
+ _05946_ sky130_fd_sc_hd__a21o_1
X_13188_ clknet_leaf_118_clk _00015_ net139 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.done
+ sky130_fd_sc_hd__dfrtp_1
X_12139_ net870 _05876_ _05883_ _05892_ vssd1 vssd1 vccd1 vccd1 _00991_ sky130_fd_sc_hd__a22o_1
X_06700_ _01588_ _01589_ vssd1 vssd1 vccd1 vccd1 _01590_ sky130_fd_sc_hd__nor2_1
X_07680_ _01181_ genblk1\[10\].osc.clkdiv_C.cnt\[12\] vssd1 vssd1 vccd1 vccd1 _02387_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06631_ genblk1\[3\].osc.clkdiv_C.cnt\[4\] _01530_ genblk1\[3\].osc.clkdiv_C.cnt\[5\]
+ vssd1 vssd1 vccd1 vccd1 _01534_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_149_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09350_ net688 _03903_ _03910_ _03926_ vssd1 vssd1 vccd1 vccd1 _00168_ sky130_fd_sc_hd__a22o_1
X_06562_ _01451_ _01474_ vssd1 vssd1 vccd1 vccd1 _01475_ sky130_fd_sc_hd__nor2_1
X_08301_ _03005_ _03007_ vssd1 vssd1 vccd1 vccd1 _03008_ sky130_fd_sc_hd__or2b_1
X_09281_ net854 _03870_ _03840_ _03873_ vssd1 vssd1 vccd1 vccd1 _00152_ sky130_fd_sc_hd__a22o_1
XFILLER_0_142_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06493_ _01197_ _01417_ _01418_ genblk1\[2\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1
+ vccd1 _01419_ sky130_fd_sc_hd__o22a_1
XFILLER_0_117_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08232_ _02225_ _02885_ vssd1 vssd1 vccd1 vccd1 _02939_ sky130_fd_sc_hd__and2_2
XFILLER_0_142_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_824 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08163_ genblk1\[3\].osc.clkdiv_C.cnt\[13\] _01498_ _02869_ vssd1 vssd1 vccd1 vccd1
+ _02870_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_27_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_654 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10938__B1 _05023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07114_ genblk1\[8\].osc.clkdiv_C.cnt\[16\] _01914_ vssd1 vssd1 vccd1 vccd1 _01916_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_30_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08094_ genblk1\[4\].osc.clkdiv_C.cnt\[14\] _01359_ _01498_ genblk1\[4\].osc.clkdiv_C.cnt\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02801_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07045_ genblk1\[8\].osc.clkdiv_C.cnt\[8\] _01430_ vssd1 vssd1 vccd1 vccd1 _01863_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_141_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08996_ net1134 _03596_ _01154_ vssd1 vssd1 vccd1 vccd1 _03678_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07947_ genblk1\[7\].osc.clkdiv_C.cnt\[6\] _01574_ vssd1 vssd1 vccd1 vccd1 _02654_
+ sky130_fd_sc_hd__or2_1
X_07878_ _02562_ _02584_ vssd1 vssd1 vccd1 vccd1 _02585_ sky130_fd_sc_hd__nor2_1
XANTENNA__09072__S _03722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09617_ _03995_ _04114_ vssd1 vssd1 vccd1 vccd1 _04115_ sky130_fd_sc_hd__xnor2_1
X_06829_ genblk1\[5\].osc.clkdiv_C.cnt\[1\] genblk1\[5\].osc.clkdiv_C.cnt\[0\] genblk1\[5\].osc.clkdiv_C.cnt\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01699_ sky130_fd_sc_hd__a21oi_1
X_09548_ _04055_ genblk1\[1\].osc.clkdiv_C.cnt\[12\] vssd1 vssd1 vccd1 vccd1 _04065_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_66_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09479_ _01433_ vssd1 vssd1 vccd1 vccd1 _04028_ sky130_fd_sc_hd__inv_2
XANTENNA__08834__A2 _02468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11510_ _05450_ genblk1\[8\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 _05451_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_25_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12490_ clknet_leaf_109_clk _00052_ net158 vssd1 vssd1 vccd1 vccd1 sig_norm.quo\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11441_ _05416_ vssd1 vssd1 vccd1 vccd1 _05417_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_123_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12496__RESET_B net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_637 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11372_ _05248_ _05350_ _05351_ _05251_ net1113 vssd1 vssd1 vccd1 vccd1 _00765_ sky130_fd_sc_hd__a32o_1
X_13111_ clknet_leaf_115_clk _00436_ net134 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.fin_quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10323_ _04629_ vssd1 vssd1 vccd1 vccd1 _00438_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07898__A2_N _01309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13042_ clknet_leaf_128_clk _00369_ net67 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.b1\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10254_ _04449_ genblk2\[4\].wave_shpr.div.acc\[16\] vssd1 vssd1 vccd1 vccd1 _04566_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__06460__A genblk1\[1\].osc.clkdiv_C.cnt\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10185_ genblk2\[3\].wave_shpr.div.acc\[11\] _04516_ _04507_ vssd1 vssd1 vccd1 vccd1
+ _04517_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11017__S _05023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12826_ clknet_leaf_62_clk _00159_ net190 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.acc\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_output17_A net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12757_ clknet_leaf_52_clk genblk1\[11\].osc.clkdiv_C.next_cnt\[16\] net110 vssd1
+ vssd1 vccd1 vccd1 genblk1\[11\].osc.clkdiv_C.cnt\[16\] sky130_fd_sc_hd__dfrtp_4
Xclkbuf_leaf_135_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_135_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10093__B1 _04456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11708_ genblk2\[9\].wave_shpr.div.b1\[14\] genblk2\[9\].wave_shpr.div.acc\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05600_ sky130_fd_sc_hd__and2b_1
XFILLER_0_16_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12688_ clknet_leaf_53_clk genblk1\[8\].osc.clkdiv_C.next_cnt\[1\] net112 vssd1 vssd1
+ vccd1 vccd1 genblk1\[8\].osc.clkdiv_C.cnt\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_126_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_154_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11639_ net704 _05507_ _05417_ _05539_ vssd1 vssd1 vccd1 vccd1 _00844_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_3_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold706 genblk2\[7\].wave_shpr.div.acc\[17\] vssd1 vssd1 vccd1 vccd1 net924 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold717 genblk2\[9\].wave_shpr.div.acc\[20\] vssd1 vssd1 vccd1 vccd1 net935 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13309_ clknet_leaf_117_clk _00630_ net137 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold728 genblk2\[8\].wave_shpr.div.acc\[24\] vssd1 vssd1 vccd1 vccd1 net946 sky130_fd_sc_hd__dlygate4sd3_1
Xhold739 genblk2\[10\].wave_shpr.div.acc\[12\] vssd1 vssd1 vccd1 vccd1 net957 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08850_ _03552_ _03555_ _03556_ vssd1 vssd1 vccd1 vccd1 _03557_ sky130_fd_sc_hd__and3_1
XANTENNA__07564__A2 _01227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07801_ genblk1\[0\].osc.clkdiv_C.cnt\[16\] _01577_ _02501_ _02507_ genblk1\[0\].osc.clkdiv_C.cnt\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02508_ sky130_fd_sc_hd__a221oi_2
X_08781_ _02583_ _03486_ _02582_ vssd1 vssd1 vccd1 vccd1 _03488_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_46_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11648__A1 _05441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07732_ genblk1\[1\].osc.clkdiv_C.cnt\[5\] _02433_ _02435_ _02436_ _02438_ vssd1
+ vssd1 vccd1 vccd1 _02439_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_79_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07663_ _01360_ _01224_ _01241_ genblk1\[10\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1
+ vccd1 _02370_ sky130_fd_sc_hd__a211o_1
X_09402_ genblk2\[1\].wave_shpr.div.acc\[5\] genblk2\[1\].wave_shpr.div.b1\[5\] vssd1
+ vssd1 vccd1 vccd1 _03966_ sky130_fd_sc_hd__and2b_1
XFILLER_0_149_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06614_ genblk1\[3\].osc.clkdiv_C.cnt\[8\] _01483_ _01484_ genblk1\[3\].osc.clkdiv_C.cnt\[0\]
+ _01521_ vssd1 vssd1 vccd1 vccd1 _01522_ sky130_fd_sc_hd__o221a_1
XFILLER_0_48_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07594_ _02276_ _02296_ _02300_ vssd1 vssd1 vccd1 vccd1 _02301_ sky130_fd_sc_hd__or3_1
X_09333_ net840 _03903_ _03910_ _03913_ vssd1 vssd1 vccd1 vccd1 _00164_ sky130_fd_sc_hd__a22o_1
X_06545_ _01452_ _01463_ vssd1 vssd1 vccd1 vccd1 genblk1\[2\].osc.clkdiv_C.next_cnt\[7\]
+ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_126_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_126_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_62_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09264_ genblk2\[0\].wave_shpr.div.quo\[24\] _03835_ _03838_ net454 _03861_ vssd1
+ vssd1 vccd1 vccd1 _00147_ sky130_fd_sc_hd__a221o_1
XFILLER_0_118_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06476_ genblk1\[1\].osc.clkdiv_C.cnt\[15\] genblk1\[1\].osc.clkdiv_C.cnt\[14\] _01401_
+ vssd1 vssd1 vccd1 vccd1 _01405_ sky130_fd_sc_hd__and3_1
XFILLER_0_145_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08215_ _02918_ _02921_ vssd1 vssd1 vccd1 vccd1 _02922_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09195_ _03825_ vssd1 vssd1 vccd1 vccd1 _00114_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08146_ _02851_ _02852_ vssd1 vssd1 vccd1 vccd1 _02853_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08077_ _02755_ _02760_ _02781_ _02783_ vssd1 vssd1 vccd1 vccd1 _02784_ sky130_fd_sc_hd__or4_1
XFILLER_0_31_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07028_ genblk1\[7\].osc.clkdiv_C.cnt\[15\] _01846_ _01848_ vssd1 vssd1 vccd1 vccd1
+ genblk1\[7\].osc.clkdiv_C.next_cnt\[15\] sky130_fd_sc_hd__o21a_1
XANTENNA__06280__A _01241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold11 genblk2\[8\].wave_shpr.div.quo\[22\] vssd1 vssd1 vccd1 vccd1 net229 sky130_fd_sc_hd__dlygate4sd3_1
Xhold22 _01054_ vssd1 vssd1 vccd1 vccd1 net240 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 genblk2\[4\].wave_shpr.div.quo\[8\] vssd1 vssd1 vccd1 vccd1 net251 sky130_fd_sc_hd__buf_1
X_08979_ net372 _01157_ vssd1 vssd1 vccd1 vccd1 _03665_ sky130_fd_sc_hd__nand2_1
Xhold44 _00313_ vssd1 vssd1 vccd1 vccd1 net262 sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 genblk2\[0\].wave_shpr.div.i\[4\] vssd1 vssd1 vccd1 vccd1 net273 sky130_fd_sc_hd__dlygate4sd3_1
Xhold66 _00653_ vssd1 vssd1 vccd1 vccd1 net284 sky130_fd_sc_hd__dlygate4sd3_1
Xhold77 _00557_ vssd1 vssd1 vccd1 vccd1 net295 sky130_fd_sc_hd__dlygate4sd3_1
Xhold88 genblk2\[9\].wave_shpr.div.quo\[24\] vssd1 vssd1 vccd1 vccd1 net306 sky130_fd_sc_hd__dlygate4sd3_1
X_11990_ genblk2\[11\].wave_shpr.div.b1\[4\] _04230_ _05433_ vssd1 vssd1 vccd1 vccd1
+ _05800_ sky130_fd_sc_hd__mux2_1
Xhold99 genblk2\[7\].wave_shpr.div.quo\[6\] vssd1 vssd1 vccd1 vccd1 net317 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12300__A2 _06009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10941_ net671 _05052_ _05056_ net756 vssd1 vssd1 vccd1 vccd1 _00629_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13660_ clknet_leaf_47_clk net447 net120 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.quo\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10872_ genblk2\[6\].wave_shpr.div.b1\[17\] genblk2\[6\].wave_shpr.div.acc\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05016_ sky130_fd_sc_hd__and2b_1
XFILLER_0_85_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12611_ clknet_leaf_23_clk genblk1\[3\].osc.clkdiv_C.next_cnt\[14\] net94 vssd1 vssd1
+ vccd1 vccd1 genblk1\[3\].osc.clkdiv_C.cnt\[14\] sky130_fd_sc_hd__dfrtp_4
Xclkbuf_leaf_117_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_117_clk
+ sky130_fd_sc_hd__clkbuf_16
X_13591_ clknet_leaf_72_clk _00906_ net216 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.acc\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_66_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12542_ clknet_leaf_100_clk net287 net164 vssd1 vssd1 vccd1 vccd1 PWM.pwm_out sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12473_ clknet_leaf_32_clk smpl_rt_clkdiv.clkDiv_inst.next_cnt\[7\] net99 vssd1 vssd1
+ vccd1 vccd1 smpl_rt_clkdiv.clkDiv_inst.cnt\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09766__A _01302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11424_ genblk2\[8\].wave_shpr.div.b1\[13\] genblk2\[8\].wave_shpr.div.acc\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05400_ sky130_fd_sc_hd__and2b_1
XFILLER_0_22_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09232__A2 _03841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_8 _04242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11355_ _05219_ _05220_ vssd1 vssd1 vccd1 vccd1 _05340_ sky130_fd_sc_hd__and2b_1
XFILLER_0_120_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10306_ genblk2\[4\].wave_shpr.div.acc\[19\] genblk2\[4\].wave_shpr.div.acc\[18\]
+ vssd1 vssd1 vccd1 vccd1 _04618_ sky130_fd_sc_hd__or2_1
XFILLER_0_120_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11286_ net1030 _05279_ _05283_ _05288_ vssd1 vssd1 vccd1 vccd1 _00742_ sky130_fd_sc_hd__a22o_1
XANTENNA__07717__C _02365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13025_ clknet_leaf_113_clk _00352_ net134 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.fin_quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12011__B1_N _03717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10237_ genblk2\[3\].wave_shpr.div.acc\[25\] _04553_ vssd1 vssd1 vccd1 vccd1 _04555_
+ sky130_fd_sc_hd__xnor2_1
X_10168_ genblk2\[3\].wave_shpr.div.acc\[7\] _04503_ _04420_ vssd1 vssd1 vccd1 vccd1
+ _04504_ sky130_fd_sc_hd__mux2_1
X_10099_ _04269_ genblk1\[3\].osc.clkdiv_C.cnt\[1\] vssd1 vssd1 vccd1 vccd1 _04459_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_88_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12809_ clknet_leaf_60_clk _00142_ net187 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.quo\[19\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_108_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_108_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__08564__B _02521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06330_ genblk1\[0\].osc.clkdiv_C.cnt\[8\] genblk1\[0\].osc.clkdiv_C.cnt\[7\] _01281_
+ vssd1 vssd1 vccd1 vccd1 _01284_ sky130_fd_sc_hd__and3_1
XTAP_1090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06365__A _01171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06261_ _01222_ vssd1 vssd1 vccd1 vccd1 _01223_ sky130_fd_sc_hd__buf_4
X_08000_ _02706_ vssd1 vssd1 vccd1 vccd1 _02707_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06192_ net642 PWM.counter\[0\] net831 vssd1 vssd1 vccd1 vccd1 _01160_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_142_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09223__A2 _03836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_102_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold503 _00632_ vssd1 vssd1 vccd1 vccd1 net721 sky130_fd_sc_hd__dlygate4sd3_1
Xhold514 genblk2\[4\].wave_shpr.div.quo\[3\] vssd1 vssd1 vccd1 vccd1 net732 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08431__B1 _02222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold525 genblk2\[8\].wave_shpr.div.quo\[0\] vssd1 vssd1 vccd1 vccd1 net743 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07908__B _01870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold536 genblk2\[7\].wave_shpr.div.quo\[5\] vssd1 vssd1 vccd1 vccd1 net754 sky130_fd_sc_hd__dlygate4sd3_1
Xhold547 sig_norm.i\[2\] vssd1 vssd1 vccd1 vccd1 net765 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06812__B _01678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09951_ _04250_ _04247_ genblk2\[2\].wave_shpr.div.i\[0\] vssd1 vssd1 vccd1 vccd1
+ _04352_ sky130_fd_sc_hd__mux2_1
Xhold558 genblk2\[11\].wave_shpr.div.quo\[3\] vssd1 vssd1 vccd1 vccd1 net776 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold569 genblk2\[4\].wave_shpr.div.acc\[23\] vssd1 vssd1 vccd1 vccd1 net787 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08902_ _03583_ _03605_ _03596_ vssd1 vssd1 vccd1 vccd1 _03606_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_148_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09882_ genblk2\[2\].wave_shpr.div.acc\[7\] _04300_ _04301_ vssd1 vssd1 vccd1 vccd1
+ _04302_ sky130_fd_sc_hd__mux2_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08833_ _03538_ _03539_ vssd1 vssd1 vccd1 vccd1 _03540_ sky130_fd_sc_hd__nor2_1
XTAP_874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout190_A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08764_ _02798_ _03466_ vssd1 vssd1 vccd1 vccd1 _03471_ sky130_fd_sc_hd__nand2_1
XANTENNA__07643__B genblk1\[11\].osc.clkdiv_C.cnt\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07715_ _02367_ _02420_ vssd1 vssd1 vccd1 vccd1 _02422_ sky130_fd_sc_hd__nor2_1
XTAP_2719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12294__A1 _03732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08695_ _03170_ _03171_ _03172_ vssd1 vssd1 vccd1 vccd1 _03402_ sky130_fd_sc_hd__a21o_1
XFILLER_0_79_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07646_ genblk2\[11\].wave_shpr.div.fin_quo\[2\] _02352_ vssd1 vssd1 vccd1 vccd1
+ _02353_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07577_ genblk1\[9\].osc.clkdiv_C.cnt\[6\] _01512_ vssd1 vssd1 vccd1 vccd1 _02284_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_76_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09316_ _03785_ _03752_ vssd1 vssd1 vccd1 vccd1 _03900_ sky130_fd_sc_hd__or2b_1
XFILLER_0_48_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06528_ genblk1\[2\].osc.clkdiv_C.cnt\[1\] genblk1\[2\].osc.clkdiv_C.cnt\[0\] vssd1
+ vssd1 vccd1 vccd1 _01453_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_63_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_35_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09247_ _03725_ genblk1\[0\].osc.clkdiv_C.cnt\[8\] vssd1 vssd1 vccd1 vccd1 _03852_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_133_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06459_ genblk1\[1\].osc.clkdiv_C.cnt\[9\] _01392_ vssd1 vssd1 vccd1 vccd1 _01394_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_63_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09178_ net1171 _01342_ _03722_ vssd1 vssd1 vccd1 vccd1 _03816_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08129_ _02808_ _02815_ _02821_ _02835_ vssd1 vssd1 vccd1 vccd1 _02836_ sky130_fd_sc_hd__or4_2
XFILLER_0_114_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11140_ _05172_ _05198_ _05199_ vssd1 vssd1 vccd1 vccd1 _05200_ sky130_fd_sc_hd__a21o_1
XFILLER_0_113_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11071_ net622 _05139_ _05142_ vssd1 vssd1 vccd1 vccd1 _05143_ sky130_fd_sc_hd__a21o_1
X_10022_ genblk2\[3\].wave_shpr.div.acc\[23\] genblk2\[3\].wave_shpr.div.acc\[25\]
+ genblk2\[3\].wave_shpr.div.acc\[24\] genblk2\[3\].wave_shpr.div.acc\[26\] vssd1
+ vssd1 vccd1 vccd1 _04418_ sky130_fd_sc_hd__or4_2
XFILLER_0_99_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11973_ _05791_ vssd1 vssd1 vccd1 vccd1 _00926_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10924_ genblk2\[7\].wave_shpr.div.b1\[13\] _02374_ _05042_ vssd1 vssd1 vccd1 vccd1
+ _05047_ sky130_fd_sc_hd__mux2_1
X_13712_ clknet_leaf_31_clk _01023_ net100 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.b1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07161__B1 genblk1\[9\].osc.clkdiv_C.cnt\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10855_ _04975_ _04997_ _04998_ vssd1 vssd1 vccd1 vccd1 _04999_ sky130_fd_sc_hd__a21o_1
XFILLER_0_128_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13643_ clknet_leaf_68_clk _00956_ net211 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13574_ clknet_leaf_85_clk _00889_ net183 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.quo\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10786_ genblk2\[5\].wave_shpr.div.acc\[19\] _04816_ _04941_ vssd1 vssd1 vccd1 vccd1
+ _04942_ sky130_fd_sc_hd__a21bo_1
XPHY_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11796__B1 _03696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12525_ clknet_leaf_67_clk _00077_ net194 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.b1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08661__B1 _02525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12456_ clknet_leaf_20_clk net225 net108 vssd1 vssd1 vccd1 vccd1 modein.delay_octave_down_in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_304 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11407_ _05371_ _05381_ _05382_ vssd1 vssd1 vccd1 vccd1 _05383_ sky130_fd_sc_hd__a21o_1
XFILLER_0_105_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12387_ net816 _06039_ _06040_ _06062_ vssd1 vssd1 vccd1 vccd1 _01069_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07728__B genblk1\[1\].osc.clkdiv_C.cnt\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07767__A2 _01309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11338_ _05215_ _05164_ vssd1 vssd1 vccd1 vccd1 _05328_ sky130_fd_sc_hd__or2b_1
XFILLER_0_120_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11269_ _05248_ _05274_ _05275_ _05251_ net1070 vssd1 vssd1 vccd1 vccd1 _00738_ sky130_fd_sc_hd__a32o_1
X_13008_ clknet_leaf_133_clk _00337_ net59 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.acc\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07463__B _02153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07500_ _02220_ vssd1 vssd1 vccd1 vccd1 _02221_ sky130_fd_sc_hd__buf_4
X_08480_ _03182_ _03186_ vssd1 vssd1 vccd1 vccd1 _03187_ sky130_fd_sc_hd__xor2_1
XFILLER_0_89_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07431_ _02152_ vssd1 vssd1 vccd1 vccd1 _02170_ sky130_fd_sc_hd__buf_6
XANTENNA__12028__A1 genblk2\[10\].wave_shpr.div.quo\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06807__B _01678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07362_ _02118_ vssd1 vssd1 vccd1 vccd1 genblk1\[11\].osc.clkdiv_C.next_cnt\[7\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_128_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09101_ genblk2\[0\].wave_shpr.div.acc\[14\] genblk2\[0\].wave_shpr.div.b1\[14\]
+ vssd1 vssd1 vccd1 vccd1 _03749_ sky130_fd_sc_hd__or2b_1
XFILLER_0_84_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_72_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06313_ _01273_ vssd1 vssd1 vccd1 vccd1 genblk1\[0\].osc.clkdiv_C.next_cnt\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_150_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07293_ net1143 _02057_ _02059_ vssd1 vssd1 vccd1 vccd1 genblk1\[10\].osc.clkdiv_C.next_cnt\[15\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_127_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09032_ _03701_ vssd1 vssd1 vccd1 vccd1 _03702_ sky130_fd_sc_hd__buf_8
XFILLER_0_115_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06244_ genblk1\[0\].osc.clkdiv_C.cnt\[2\] _01190_ _01204_ _01205_ vssd1 vssd1 vccd1
+ vccd1 _01206_ sky130_fd_sc_hd__o211a_1
XFILLER_0_150_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_142_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold300 genblk2\[10\].wave_shpr.div.quo\[18\] vssd1 vssd1 vccd1 vccd1 net518 sky130_fd_sc_hd__dlygate4sd3_1
X_06175_ _01137_ _01146_ vssd1 vssd1 vccd1 vccd1 _01147_ sky130_fd_sc_hd__nand2_1
Xhold311 genblk2\[3\].wave_shpr.div.quo\[22\] vssd1 vssd1 vccd1 vccd1 net529 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold322 genblk2\[7\].wave_shpr.div.acc_next\[0\] vssd1 vssd1 vccd1 vccd1 net540 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold333 genblk2\[5\].wave_shpr.div.quo\[15\] vssd1 vssd1 vccd1 vccd1 net551 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13316__RESET_B net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold344 _00400_ vssd1 vssd1 vccd1 vccd1 net562 sky130_fd_sc_hd__dlygate4sd3_1
Xhold355 genblk2\[2\].wave_shpr.div.quo\[16\] vssd1 vssd1 vccd1 vccd1 net573 sky130_fd_sc_hd__dlygate4sd3_1
Xhold366 genblk2\[0\].wave_shpr.div.quo\[12\] vssd1 vssd1 vccd1 vccd1 net584 sky130_fd_sc_hd__dlygate4sd3_1
Xhold377 genblk2\[6\].wave_shpr.div.quo\[16\] vssd1 vssd1 vccd1 vccd1 net595 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold388 _00336_ vssd1 vssd1 vccd1 vccd1 net606 sky130_fd_sc_hd__dlygate4sd3_1
X_09934_ genblk2\[2\].wave_shpr.div.acc\[20\] _04339_ vssd1 vssd1 vccd1 vccd1 _04341_
+ sky130_fd_sc_hd__xor2_1
Xhold399 genblk2\[8\].wave_shpr.div.quo\[18\] vssd1 vssd1 vccd1 vccd1 net617 sky130_fd_sc_hd__dlygate4sd3_1
X_09865_ net975 _04282_ _04252_ _04288_ vssd1 vssd1 vccd1 vccd1 _00321_ sky130_fd_sc_hd__a22o_1
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1000 genblk2\[0\].wave_shpr.div.fin_quo\[7\] vssd1 vssd1 vccd1 vccd1 net1218
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1011 genblk1\[5\].osc.clkdiv_C.cnt\[13\] vssd1 vssd1 vccd1 vccd1 net1229 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1022 sig_norm.acc\[4\] vssd1 vssd1 vccd1 vccd1 net1240 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09380__A1 _03944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1033 genblk2\[10\].wave_shpr.div.b1\[13\] vssd1 vssd1 vccd1 vccd1 net1251 sky130_fd_sc_hd__dlygate4sd3_1
X_08816_ _03521_ _03522_ vssd1 vssd1 vccd1 vccd1 _03523_ sky130_fd_sc_hd__nand2_1
Xhold1044 genblk2\[4\].wave_shpr.div.b1\[14\] vssd1 vssd1 vccd1 vccd1 net1262 sky130_fd_sc_hd__dlygate4sd3_1
X_09796_ _04249_ vssd1 vssd1 vccd1 vccd1 _04250_ sky130_fd_sc_hd__buf_4
Xhold1055 genblk2\[10\].wave_shpr.div.b1\[4\] vssd1 vssd1 vccd1 vccd1 net1273 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1066 genblk2\[10\].wave_shpr.div.b1\[9\] vssd1 vssd1 vccd1 vccd1 net1284 sky130_fd_sc_hd__dlygate4sd3_1
X_08747_ _02742_ _03453_ _02745_ vssd1 vssd1 vccd1 vccd1 _03454_ sky130_fd_sc_hd__o21ai_2
XANTENNA_clkbuf_leaf_90_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1077 genblk2\[1\].wave_shpr.div.b1\[2\] vssd1 vssd1 vccd1 vccd1 net1295 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1088 _00173_ vssd1 vssd1 vccd1 vccd1 net1306 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1099 genblk2\[9\].wave_shpr.div.quo\[4\] vssd1 vssd1 vccd1 vccd1 net1317 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08678_ _02561_ _02562_ vssd1 vssd1 vccd1 vccd1 _03385_ sky130_fd_sc_hd__or2_1
XANTENNA__10135__B_N _04455_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07629_ _01174_ _01177_ vssd1 vssd1 vccd1 vccd1 _02336_ sky130_fd_sc_hd__nand2_4
XTAP_1859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10640_ _04847_ vssd1 vssd1 vccd1 vccd1 _00537_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10571_ _04771_ _04797_ _04798_ vssd1 vssd1 vccd1 vccd1 _04799_ sky130_fd_sc_hd__a21o_1
XFILLER_0_63_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12310_ _05835_ genblk1\[11\].osc.clkdiv_C.cnt\[1\] vssd1 vssd1 vccd1 vccd1 _06012_
+ sky130_fd_sc_hd__and2_1
X_13290_ clknet_leaf_88_clk _00611_ net177 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.b1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12241_ genblk2\[11\].wave_shpr.div.acc\[22\] genblk2\[11\].wave_shpr.div.acc\[21\]
+ genblk2\[11\].wave_shpr.div.acc\[20\] _05978_ vssd1 vssd1 vccd1 vccd1 _05979_ sky130_fd_sc_hd__or4_1
X_12172_ net1081 _05818_ _05816_ _05915_ vssd1 vssd1 vccd1 vccd1 _01001_ sky130_fd_sc_hd__a22o_1
XANTENNA__06957__B1 _01732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11123_ genblk2\[7\].wave_shpr.div.b1\[1\] genblk2\[7\].wave_shpr.div.acc\[1\] vssd1
+ vssd1 vccd1 vccd1 _05183_ sky130_fd_sc_hd__xor2_1
XANTENNA_clkbuf_leaf_43_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11054_ _05012_ _04968_ vssd1 vssd1 vccd1 vccd1 _05130_ sky130_fd_sc_hd__or2b_1
X_10005_ genblk2\[3\].wave_shpr.div.b1\[11\] genblk2\[3\].wave_shpr.div.acc\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04401_ sky130_fd_sc_hd__and2b_1
XANTENNA_clkbuf_leaf_58_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_101_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11956_ _03832_ genblk2\[10\].wave_shpr.div.acc\[16\] vssd1 vssd1 vccd1 vccd1 _05778_
+ sky130_fd_sc_hd__and2_1
XANTENNA__07134__B1 _01923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10907_ net1293 _05037_ _04848_ vssd1 vssd1 vccd1 vccd1 _05038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11887_ _05715_ _05716_ vssd1 vssd1 vccd1 vccd1 _05717_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13626_ clknet_leaf_67_clk _00939_ net195 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.b1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10838_ genblk2\[6\].wave_shpr.div.acc\[1\] genblk2\[6\].wave_shpr.div.b1\[1\] vssd1
+ vssd1 vccd1 vccd1 _04982_ sky130_fd_sc_hd__xor2_1
XFILLER_0_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_116_clk_A clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10769_ _04810_ _04765_ vssd1 vssd1 vccd1 vccd1 _04929_ sky130_fd_sc_hd__or2b_1
X_13557_ clknet_leaf_97_clk net268 net169 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12508_ clknet_leaf_103_clk _00070_ net156 vssd1 vssd1 vccd1 vccd1 PWM.final_in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13488_ clknet_leaf_88_clk net330 net177 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.quo\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10992__B2 _05052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12439_ genblk2\[11\].wave_shpr.div.acc\[24\] _03947_ _03944_ _06100_ vssd1 vssd1
+ vccd1 vccd1 _01083_ sky130_fd_sc_hd__a22o_1
XFILLER_0_140_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07980_ _02685_ _02686_ vssd1 vssd1 vccd1 vccd1 _02687_ sky130_fd_sc_hd__and2_1
Xfanout109 net127 vssd1 vssd1 vccd1 vccd1 net109 sky130_fd_sc_hd__buf_2
XFILLER_0_38_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06931_ genblk1\[6\].osc.clkdiv_C.cnt\[9\] _01773_ vssd1 vssd1 vccd1 vccd1 _01776_
+ sky130_fd_sc_hd__nor2_1
X_09650_ genblk2\[1\].wave_shpr.div.acc\[21\] _04007_ _04129_ vssd1 vssd1 vccd1 vccd1
+ _04139_ sky130_fd_sc_hd__or3_1
X_06862_ net27 _01719_ vssd1 vssd1 vccd1 vccd1 _01720_ sky130_fd_sc_hd__nor2_1
X_08601_ _03251_ _03252_ _03255_ vssd1 vssd1 vccd1 vccd1 _03308_ sky130_fd_sc_hd__and3b_1
X_09581_ _03980_ _03966_ vssd1 vssd1 vccd1 vccd1 _04087_ sky130_fd_sc_hd__nor2_1
X_06793_ genblk1\[5\].osc.clkdiv_C.cnt\[3\] _01592_ vssd1 vssd1 vccd1 vccd1 _01665_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08532_ _02416_ _03238_ net2 _02364_ vssd1 vssd1 vccd1 vccd1 _03239_ sky130_fd_sc_hd__o211a_1
XANTENNA__07921__B _01430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08463_ _03163_ _03164_ _03169_ vssd1 vssd1 vccd1 vccd1 _03170_ sky130_fd_sc_hd__nand3_2
XFILLER_0_49_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07414_ genblk2\[1\].wave_shpr.div.busy _02157_ vssd1 vssd1 vccd1 vccd1 _02158_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08394_ genblk1\[2\].osc.clkdiv_C.cnt\[11\] _01411_ vssd1 vssd1 vccd1 vccd1 _03101_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_57_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07345_ genblk1\[11\].osc.clkdiv_C.cnt\[4\] _02101_ vssd1 vssd1 vccd1 vccd1 _02105_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__11224__A2 _05246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_30_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_30_clk sky130_fd_sc_hd__clkbuf_16
X_07276_ genblk1\[10\].osc.clkdiv_C.cnt\[9\] _02046_ vssd1 vssd1 vccd1 vccd1 _02049_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09015_ genblk2\[9\].wave_shpr.div.i\[0\] _02202_ genblk2\[9\].wave_shpr.div.i\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03688_ sky130_fd_sc_hd__a21oi_1
X_06227_ _01174_ _01187_ _01188_ vssd1 vssd1 vccd1 vccd1 _01189_ sky130_fd_sc_hd__a21boi_4
XFILLER_0_115_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12185__B1 _03855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold130 genblk2\[9\].wave_shpr.div.acc\[26\] vssd1 vssd1 vccd1 vccd1 net348 sky130_fd_sc_hd__dlygate4sd3_1
Xhold141 smpl_rt_clkdiv.clkDiv_inst.cnt\[2\] vssd1 vssd1 vccd1 vccd1 net359 sky130_fd_sc_hd__dlygate4sd3_1
X_06158_ net12 vssd1 vssd1 vccd1 vccd1 _01130_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold152 genblk2\[7\].wave_shpr.div.quo\[11\] vssd1 vssd1 vccd1 vccd1 net370 sky130_fd_sc_hd__dlygate4sd3_1
Xhold163 genblk2\[7\].wave_shpr.div.acc\[26\] vssd1 vssd1 vccd1 vccd1 net381 sky130_fd_sc_hd__dlygate4sd3_1
Xhold174 genblk2\[5\].wave_shpr.div.acc\[26\] vssd1 vssd1 vccd1 vccd1 net392 sky130_fd_sc_hd__dlygate4sd3_1
Xhold185 _01036_ vssd1 vssd1 vccd1 vccd1 net403 sky130_fd_sc_hd__dlygate4sd3_1
Xhold196 genblk2\[1\].wave_shpr.div.quo\[4\] vssd1 vssd1 vccd1 vccd1 net414 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09917_ net845 _04315_ _04322_ _04328_ vssd1 vssd1 vccd1 vccd1 _00333_ sky130_fd_sc_hd__a22o_1
Xclkbuf_leaf_97_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_97_clk sky130_fd_sc_hd__clkbuf_16
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09848_ _03702_ _01416_ vssd1 vssd1 vccd1 vccd1 _04276_ sky130_fd_sc_hd__nand2_1
XANTENNA_fanout66_A net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09779_ _04239_ vssd1 vssd1 vccd1 vccd1 _00284_ sky130_fd_sc_hd__clkbuf_1
XTAP_2302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11810_ net886 _05652_ _05653_ _05659_ vssd1 vssd1 vccd1 vccd1 _00895_ sky130_fd_sc_hd__a22o_1
XTAP_2324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12790_ clknet_leaf_57_clk _00123_ net182 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.quo\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11741_ _02248_ _01145_ _05622_ net1073 vssd1 vssd1 vccd1 vccd1 _00863_ sky130_fd_sc_hd__a22o_1
XTAP_2368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11672_ genblk2\[9\].wave_shpr.div.acc\[7\] genblk2\[9\].wave_shpr.div.b1\[7\] vssd1
+ vssd1 vccd1 vccd1 _05564_ sky130_fd_sc_hd__or2b_1
XTAP_1689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13411_ clknet_leaf_91_clk _00730_ net144 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.quo\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10623_ _01747_ vssd1 vssd1 vccd1 vccd1 _04838_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11215__A2 _05246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06890__A2 _01519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_21_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_21_clk sky130_fd_sc_hd__clkbuf_16
X_13342_ clknet_leaf_7_clk _00663_ net49 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.acc\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10554_ genblk2\[5\].wave_shpr.div.b1\[1\] genblk2\[5\].wave_shpr.div.acc\[1\] vssd1
+ vssd1 vccd1 vccd1 _04782_ sky130_fd_sc_hd__xor2_1
XFILLER_0_63_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13273_ clknet_leaf_12_clk _00016_ net51 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.busy
+ sky130_fd_sc_hd__dfrtp_1
X_10485_ _04612_ _04567_ vssd1 vssd1 vccd1 vccd1 _04729_ sky130_fd_sc_hd__or2b_1
XFILLER_0_121_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12224_ _05932_ _05960_ _05961_ vssd1 vssd1 vccd1 vccd1 _05962_ sky130_fd_sc_hd__a21o_1
XFILLER_0_122_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12155_ _05783_ _05899_ vssd1 vssd1 vccd1 vccd1 _05904_ sky130_fd_sc_hd__nor2_1
XANTENNA__10713__A _02183_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11106_ genblk2\[7\].wave_shpr.div.acc\[15\] genblk2\[7\].wave_shpr.div.b1\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05166_ sky130_fd_sc_hd__or2b_1
X_12086_ _05751_ _05851_ vssd1 vssd1 vccd1 vccd1 _05852_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_leaf_88_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_88_clk sky130_fd_sc_hd__clkbuf_16
X_11037_ _05003_ _05116_ vssd1 vssd1 vccd1 vccd1 _05117_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_87_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12988_ clknet_leaf_124_clk net915 net71 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.acc\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_148_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11939_ _05741_ _05759_ _05760_ vssd1 vssd1 vccd1 vccd1 _05761_ sky130_fd_sc_hd__a21o_1
XFILLER_0_28_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10662__B1 _04857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10594__S _00015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13609_ clknet_leaf_58_clk _00922_ net194 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.i\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_12_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_12_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_131_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07130_ genblk1\[9\].osc.clkdiv_C.cnt\[9\] vssd1 vssd1 vccd1 vccd1 _01930_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07061_ genblk1\[8\].osc.clkdiv_C.cnt\[2\] vssd1 vssd1 vccd1 vccd1 _01879_ sky130_fd_sc_hd__inv_2
XFILLER_0_112_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07916__B _01487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07963_ _01200_ genblk1\[7\].osc.clkdiv_C.cnt\[15\] _01361_ _02668_ _02669_ vssd1
+ vssd1 vccd1 vccd1 _02670_ sky130_fd_sc_hd__o311a_1
Xclkbuf_leaf_79_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_79_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__08138__A2 _02309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09702_ _04169_ _04180_ _04181_ vssd1 vssd1 vccd1 vccd1 _04182_ sky130_fd_sc_hd__a21o_1
X_06914_ genblk1\[6\].osc.clkdiv_C.cnt\[3\] _01763_ vssd1 vssd1 vccd1 vccd1 _01765_
+ sky130_fd_sc_hd__and2_1
X_07894_ _02520_ net24 _02599_ _02600_ vssd1 vssd1 vccd1 vccd1 _02601_ sky130_fd_sc_hd__o31a_1
XFILLER_0_4_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07932__A genblk2\[8\].wave_shpr.div.fin_quo\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09633_ _04003_ _04126_ vssd1 vssd1 vccd1 vccd1 _04127_ sky130_fd_sc_hd__xnor2_1
X_06845_ genblk1\[5\].osc.clkdiv_C.cnt\[7\] _01705_ genblk1\[5\].osc.clkdiv_C.cnt\[8\]
+ vssd1 vssd1 vccd1 vccd1 _01709_ sky130_fd_sc_hd__a21oi_1
X_09564_ _03970_ _03971_ vssd1 vssd1 vccd1 vccd1 _04074_ sky130_fd_sc_hd__xor2_1
X_06776_ genblk1\[4\].osc.clkdiv_C.cnt\[15\] _01647_ vssd1 vssd1 vccd1 vccd1 _01651_
+ sky130_fd_sc_hd__or2_1
X_08515_ _03127_ _03218_ _03204_ _03217_ vssd1 vssd1 vccd1 vccd1 _03222_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_78_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09495_ net1271 net35 _04024_ vssd1 vssd1 vccd1 vccd1 _04038_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08446_ _03024_ _03028_ vssd1 vssd1 vccd1 vccd1 _03153_ sky130_fd_sc_hd__xor2_2
XFILLER_0_93_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08763__A net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08377_ _03073_ _03072_ vssd1 vssd1 vccd1 vccd1 _03084_ sky130_fd_sc_hd__and2b_1
XFILLER_0_80_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12285__A _03702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07328_ _02091_ vssd1 vssd1 vccd1 vccd1 _02092_ sky130_fd_sc_hd__buf_2
XANTENNA__09810__A2 _04253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07259_ genblk1\[10\].osc.clkdiv_C.cnt\[4\] _02034_ vssd1 vssd1 vccd1 vccd1 _02037_
+ sky130_fd_sc_hd__or2_1
XANTENNA__07821__B2 _02527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10270_ genblk2\[4\].wave_shpr.div.acc\[2\] genblk2\[4\].wave_shpr.div.b1\[2\] vssd1
+ vssd1 vccd1 vccd1 _04582_ sky130_fd_sc_hd__or2b_1
XANTENNA__10708__A1 _04855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12911_ clknet_leaf_34_clk _00242_ net107 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.acc\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12842_ clknet_leaf_65_clk _00175_ net197 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.acc\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12773_ clknet_leaf_47_clk _00106_ net119 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.b1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10644__B1 _04647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11724_ genblk2\[9\].wave_shpr.div.fin_quo\[1\] net1328 _00023_ vssd1 vssd1 vccd1
+ vccd1 _05615_ sky130_fd_sc_hd__mux2_1
XTAP_1464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11655_ _05549_ vssd1 vssd1 vccd1 vccd1 _05550_ sky130_fd_sc_hd__inv_2
XFILLER_0_138_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout80 net83 vssd1 vssd1 vccd1 vccd1 net80 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_154_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout91 net127 vssd1 vssd1 vccd1 vccd1 net91 sky130_fd_sc_hd__clkbuf_4
X_10606_ genblk2\[5\].wave_shpr.div.fin_quo\[6\] net1315 _00015_ vssd1 vssd1 vccd1
+ vccd1 _04828_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11586_ net922 _05447_ _05484_ _05500_ vssd1 vssd1 vccd1 vccd1 _00830_ sky130_fd_sc_hd__a22o_1
XANTENNA__09262__B1 _03838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09801__A2 _04248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10537_ genblk2\[5\].wave_shpr.div.acc\[15\] genblk2\[5\].wave_shpr.div.b1\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04765_ sky130_fd_sc_hd__or2b_1
X_13325_ clknet_leaf_26_clk _00646_ net87 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.quo\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10468_ _04604_ _04571_ vssd1 vssd1 vccd1 vccd1 _04716_ sky130_fd_sc_hd__or2b_1
X_13256_ clknet_leaf_3_clk net773 net51 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.acc\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12207_ _05940_ genblk2\[11\].wave_shpr.div.acc\[2\] _05944_ vssd1 vssd1 vccd1 vccd1
+ _05945_ sky130_fd_sc_hd__o21a_1
XANTENNA__12134__S _05865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13187_ clknet_leaf_11_clk _00014_ net56 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.busy
+ sky130_fd_sc_hd__dfrtp_1
X_10399_ _04477_ genblk1\[4\].osc.clkdiv_C.cnt\[8\] vssd1 vssd1 vccd1 vccd1 _04668_
+ sky130_fd_sc_hd__and2_1
XANTENNA__11372__A1 _05248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07576__B1 _01234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12138_ genblk2\[10\].wave_shpr.div.acc\[15\] _05891_ _05865_ vssd1 vssd1 vccd1 vccd1
+ _05892_ sky130_fd_sc_hd__mux2_1
X_12069_ net247 _05812_ _05815_ net446 _05839_ vssd1 vssd1 vccd1 vccd1 _00974_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_1_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_1_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_29_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11274__A _05245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06630_ genblk1\[3\].osc.clkdiv_C.cnt\[5\] genblk1\[3\].osc.clkdiv_C.cnt\[4\] _01530_
+ vssd1 vssd1 vccd1 vccd1 _01533_ sky130_fd_sc_hd__and3_1
XFILLER_0_126_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06368__A _01309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06561_ genblk1\[2\].osc.clkdiv_C.cnt\[13\] genblk1\[2\].osc.clkdiv_C.cnt\[12\] _01470_
+ vssd1 vssd1 vccd1 vccd1 _01474_ sky130_fd_sc_hd__and3_1
XFILLER_0_59_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08300_ _02927_ _03006_ vssd1 vssd1 vccd1 vccd1 _03007_ sky130_fd_sc_hd__and2_1
X_09280_ genblk2\[0\].wave_shpr.div.acc\[2\] _03872_ _03804_ vssd1 vssd1 vccd1 vccd1
+ _03873_ sky130_fd_sc_hd__mux2_1
X_06492_ _01229_ _01182_ vssd1 vssd1 vccd1 vccd1 _01418_ sky130_fd_sc_hd__nand2_2
XANTENNA__06303__A1 genblk1\[0\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08231_ _02937_ _02936_ vssd1 vssd1 vccd1 vccd1 _02938_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_74_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06815__B _01355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08162_ _02866_ _02867_ _02868_ vssd1 vssd1 vccd1 vccd1 _02869_ sky130_fd_sc_hd__and3_1
XFILLER_0_133_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10938__A1 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10938__B2 _05055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07113_ genblk1\[8\].osc.clkdiv_C.cnt\[15\] _01912_ _01915_ vssd1 vssd1 vccd1 vccd1
+ genblk1\[8\].osc.clkdiv_C.next_cnt\[15\] sky130_fd_sc_hd__o21a_1
XFILLER_0_15_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08093_ genblk1\[4\].osc.clkdiv_C.cnt\[14\] _01360_ vssd1 vssd1 vccd1 vccd1 _02800_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_141_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09618__S _04095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07044_ _01854_ _01856_ _01857_ _01861_ vssd1 vssd1 vccd1 vccd1 _01862_ sky130_fd_sc_hd__or4_1
XFILLER_0_100_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07567__B1 _01349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08995_ net428 _00024_ _03676_ _03677_ vssd1 vssd1 vccd1 vccd1 _00062_ sky130_fd_sc_hd__o22a_1
XFILLER_0_76_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07946_ genblk1\[7\].osc.clkdiv_C.cnt\[6\] _01574_ _01802_ genblk1\[7\].osc.clkdiv_C.cnt\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02653_ sky130_fd_sc_hd__a22o_1
X_07877_ _02571_ _02582_ _02583_ vssd1 vssd1 vccd1 vccd1 _02584_ sky130_fd_sc_hd__a21o_1
XANTENNA__08531__A2 _02525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09616_ _03996_ _03958_ vssd1 vssd1 vccd1 vccd1 _04114_ sky130_fd_sc_hd__or2b_1
X_06828_ genblk1\[5\].osc.clkdiv_C.cnt\[2\] genblk1\[5\].osc.clkdiv_C.cnt\[1\] genblk1\[5\].osc.clkdiv_C.cnt\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01698_ sky130_fd_sc_hd__and3_1
XANTENNA__06278__A _01238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06759_ _01637_ vssd1 vssd1 vccd1 vccd1 _01638_ sky130_fd_sc_hd__inv_2
X_09547_ net257 _04052_ _04053_ net417 _04064_ vssd1 vssd1 vccd1 vccd1 _00227_ sky130_fd_sc_hd__a221o_1
X_09478_ _04027_ vssd1 vssd1 vccd1 vccd1 _00195_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_109_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08429_ _03131_ _03132_ vssd1 vssd1 vccd1 vccd1 _03136_ sky130_fd_sc_hd__xor2_1
XFILLER_0_81_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11440_ _05415_ vssd1 vssd1 vccd1 vccd1 _05416_ sky130_fd_sc_hd__buf_2
XFILLER_0_135_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_123_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08598__A2 _02592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11371_ genblk2\[7\].wave_shpr.div.i\[1\] genblk2\[7\].wave_shpr.div.i\[0\] vssd1
+ vssd1 vccd1 vccd1 _05351_ sky130_fd_sc_hd__nand2_1
X_10322_ genblk2\[4\].wave_shpr.div.fin_quo\[5\] genblk2\[4\].wave_shpr.div.quo\[4\]
+ _00013_ vssd1 vssd1 vccd1 vccd1 _04629_ sky130_fd_sc_hd__mux2_1
X_13110_ clknet_leaf_114_clk _00435_ net133 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.fin_quo\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13041_ clknet_leaf_126_clk _00368_ net66 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.b1\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10253_ genblk2\[4\].wave_shpr.div.acc\[17\] genblk2\[4\].wave_shpr.div.b1\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04565_ sky130_fd_sc_hd__or2b_1
X_10184_ _04400_ _04515_ vssd1 vssd1 vccd1 vccd1 _04516_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12303__B1 _06010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07572__A genblk1\[9\].osc.clkdiv_C.cnt\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12825_ clknet_leaf_62_clk _00158_ net190 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.acc\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12756_ clknet_leaf_50_clk genblk1\[11\].osc.clkdiv_C.next_cnt\[15\] net110 vssd1
+ vssd1 vccd1 vccd1 genblk1\[11\].osc.clkdiv_C.cnt\[15\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11290__B1 _05283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11541__B genblk1\[8\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11707_ _05558_ _05597_ _05598_ vssd1 vssd1 vccd1 vccd1 _05599_ sky130_fd_sc_hd__a21o_1
XFILLER_0_127_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12687_ clknet_leaf_54_clk genblk1\[8\].osc.clkdiv_C.next_cnt\[0\] net174 vssd1 vssd1
+ vccd1 vccd1 genblk1\[8\].osc.clkdiv_C.cnt\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_115_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11638_ _05412_ _05538_ _05471_ vssd1 vssd1 vccd1 vccd1 _05539_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11569_ net898 _05447_ _05484_ _05487_ vssd1 vssd1 vccd1 vccd1 _00826_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold707 genblk2\[5\].wave_shpr.div.acc\[16\] vssd1 vssd1 vccd1 vccd1 net925 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13308_ clknet_leaf_117_clk _00629_ net137 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.quo\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold718 _00911_ vssd1 vssd1 vccd1 vccd1 net936 sky130_fd_sc_hd__dlygate4sd3_1
Xhold729 genblk2\[8\].wave_shpr.div.acc\[15\] vssd1 vssd1 vccd1 vccd1 net947 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13239_ clknet_leaf_10_clk _00562_ net57 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.quo\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06370__B _01313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09962__A _03690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07800_ _02475_ _02476_ _02478_ _02504_ _02506_ vssd1 vssd1 vccd1 vccd1 _02507_ sky130_fd_sc_hd__o221a_1
X_08780_ _02583_ _03486_ _02582_ vssd1 vssd1 vccd1 vccd1 _03487_ sky130_fd_sc_hd__or3b_1
X_07731_ genblk1\[1\].osc.clkdiv_C.cnt\[6\] _01360_ net37 _02437_ vssd1 vssd1 vccd1
+ vccd1 _02438_ sky130_fd_sc_hd__a31o_1
XANTENNA__07482__A _02147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07662_ genblk1\[10\].osc.clkdiv_C.cnt\[5\] _01182_ vssd1 vssd1 vccd1 vccd1 _02369_
+ sky130_fd_sc_hd__or2_1
X_06613_ _01485_ _01256_ _01511_ _01518_ _01520_ vssd1 vssd1 vccd1 vccd1 _01521_ sky130_fd_sc_hd__o2111a_1
X_09401_ genblk2\[1\].wave_shpr.div.b1\[6\] vssd1 vssd1 vccd1 vccd1 _03965_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07593_ _02270_ _02297_ _02299_ vssd1 vssd1 vccd1 vccd1 _02300_ sky130_fd_sc_hd__or3b_1
X_09332_ genblk2\[0\].wave_shpr.div.acc\[14\] _03912_ _03889_ vssd1 vssd1 vccd1 vccd1
+ _03913_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06544_ genblk1\[2\].osc.clkdiv_C.cnt\[7\] _01461_ vssd1 vssd1 vccd1 vccd1 _01463_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__12073__A2 _05787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09263_ _03853_ genblk1\[0\].osc.clkdiv_C.cnt\[15\] vssd1 vssd1 vccd1 vccd1 _03861_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_8_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06475_ genblk1\[1\].osc.clkdiv_C.cnt\[14\] _01401_ _01404_ vssd1 vssd1 vccd1 vccd1
+ genblk1\[1\].osc.clkdiv_C.next_cnt\[14\] sky130_fd_sc_hd__o21a_1
X_08214_ _02747_ _02919_ _02920_ vssd1 vssd1 vccd1 vccd1 _02921_ sky130_fd_sc_hd__nand3_1
XFILLER_0_8_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09194_ net1284 _01991_ _03822_ vssd1 vssd1 vccd1 vccd1 _03825_ sky130_fd_sc_hd__mux2_1
XANTENNA__09226__B1 _03840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08145_ _01201_ genblk1\[3\].osc.clkdiv_C.cnt\[15\] genblk1\[3\].osc.clkdiv_C.cnt\[14\]
+ _01362_ vssd1 vssd1 vccd1 vccd1 _02852_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_16_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_636 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07657__A net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08076_ genblk1\[5\].osc.clkdiv_C.cnt\[8\] _01678_ _02782_ vssd1 vssd1 vccd1 vccd1
+ _02783_ sky130_fd_sc_hd__a21bo_1
X_07027_ _01822_ _01847_ vssd1 vssd1 vccd1 vccd1 _01848_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10083__A _02170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10139__A2 _04420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold12 _00818_ vssd1 vssd1 vccd1 vccd1 net230 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 genblk2\[6\].wave_shpr.div.quo\[6\] vssd1 vssd1 vccd1 vccd1 net241 sky130_fd_sc_hd__dlygate4sd3_1
X_08978_ _03661_ _03663_ _02248_ vssd1 vssd1 vccd1 vccd1 _03664_ sky130_fd_sc_hd__mux2_1
Xhold34 _00468_ vssd1 vssd1 vccd1 vccd1 net252 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 genblk2\[8\].wave_shpr.div.quo\[17\] vssd1 vssd1 vccd1 vccd1 net263 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 genblk2\[8\].wave_shpr.div.acc_next\[0\] vssd1 vssd1 vccd1 vccd1 net274 sky130_fd_sc_hd__buf_1
Xhold67 genblk2\[1\].wave_shpr.div.i\[4\] vssd1 vssd1 vccd1 vccd1 net285 sky130_fd_sc_hd__dlygate4sd3_1
X_07929_ _02221_ net30 vssd1 vssd1 vccd1 vccd1 _02636_ sky130_fd_sc_hd__nor2_2
Xhold78 genblk2\[3\].wave_shpr.div.quo\[19\] vssd1 vssd1 vccd1 vccd1 net296 sky130_fd_sc_hd__dlygate4sd3_1
Xhold89 _00890_ vssd1 vssd1 vccd1 vccd1 net307 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10940_ net756 _05052_ _05056_ net792 vssd1 vssd1 vccd1 vccd1 _00628_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10871_ _04851_ genblk2\[6\].wave_shpr.div.acc\[16\] _05014_ vssd1 vssd1 vccd1 vccd1
+ _05015_ sky130_fd_sc_hd__a21o_1
XPHY_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12610_ clknet_leaf_22_clk genblk1\[3\].osc.clkdiv_C.next_cnt\[13\] net93 vssd1 vssd1
+ vccd1 vccd1 genblk1\[3\].osc.clkdiv_C.cnt\[13\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_94_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13590_ clknet_leaf_73_clk _00905_ net215 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.acc\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_93_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10075__A1 _01365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12541_ clknet_leaf_64_clk _00093_ net189 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.b1\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12472_ clknet_leaf_32_clk smpl_rt_clkdiv.clkDiv_inst.next_cnt\[6\] net99 vssd1 vssd1
+ vccd1 vccd1 smpl_rt_clkdiv.clkDiv_inst.cnt\[6\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__09768__A1 _01262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11423_ _05363_ _05397_ _05398_ vssd1 vssd1 vccd1 vccd1 _05399_ sky130_fd_sc_hd__a21o_1
XFILLER_0_151_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09766__B _03727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_9 _04242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11354_ net706 _05311_ _05315_ _05339_ vssd1 vssd1 vccd1 vccd1 _00759_ sky130_fd_sc_hd__a22o_1
XANTENNA__07243__A2 _01235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10305_ _04565_ _04615_ _04616_ vssd1 vssd1 vccd1 vccd1 _04617_ sky130_fd_sc_hd__a21o_1
X_11285_ net877 _05287_ _05222_ vssd1 vssd1 vccd1 vccd1 _05288_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10236_ net1021 _04457_ _04454_ _04554_ vssd1 vssd1 vccd1 vccd1 _00426_ sky130_fd_sc_hd__a22o_1
X_13024_ clknet_leaf_114_clk _00351_ net132 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.fin_quo\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09782__A _03702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10167_ _04392_ _04502_ vssd1 vssd1 vccd1 vccd1 _04503_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07951__B1 _01732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10098_ net538 _04457_ _04454_ genblk2\[3\].wave_shpr.div.quo\[8\] _04458_ vssd1
+ vssd1 vccd1 vccd1 _00384_ sky130_fd_sc_hd__a221o_1
XFILLER_0_89_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12808_ clknet_leaf_60_clk net411 net187 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.quo\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10066__A1 _04229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09022__A _03693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11263__B1 _05249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12739_ clknet_leaf_48_clk genblk1\[10\].osc.clkdiv_C.next_cnt\[16\] net114 vssd1
+ vssd1 vccd1 vccd1 genblk1\[10\].osc.clkdiv_C.cnt\[16\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_155_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_120_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06260_ freq_div.state\[0\] freq_div.state\[1\] freq_div.state\[2\] vssd1 vssd1 vccd1
+ vccd1 _01222_ sky130_fd_sc_hd__and3b_1
XFILLER_0_115_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06690__B1 _01578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06191_ PWM.counter\[1\] PWM.counter\[0\] PWM.counter\[2\] vssd1 vssd1 vccd1 vccd1
+ _01159_ sky130_fd_sc_hd__and3_1
Xhold504 genblk2\[8\].wave_shpr.div.b1\[14\] vssd1 vssd1 vccd1 vccd1 net722 sky130_fd_sc_hd__dlygate4sd3_1
Xhold515 _00463_ vssd1 vssd1 vccd1 vccd1 net733 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold526 _00796_ vssd1 vssd1 vccd1 vccd1 net744 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold537 genblk2\[1\].wave_shpr.div.quo\[2\] vssd1 vssd1 vccd1 vccd1 net755 sky130_fd_sc_hd__dlygate4sd3_1
Xhold548 _00028_ vssd1 vssd1 vccd1 vccd1 net766 sky130_fd_sc_hd__dlygate4sd3_1
Xhold559 genblk2\[4\].wave_shpr.div.acc\[25\] vssd1 vssd1 vccd1 vccd1 net777 sky130_fd_sc_hd__dlygate4sd3_1
X_09950_ net962 _04253_ _04251_ _04351_ vssd1 vssd1 vccd1 vccd1 _00343_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08901_ _03582_ _03577_ _03581_ vssd1 vssd1 vccd1 vccd1 _03605_ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_4_9_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09881_ _04213_ vssd1 vssd1 vccd1 vccd1 _04301_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_148_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08832_ _03531_ _03537_ _03536_ vssd1 vssd1 vccd1 vccd1 _03539_ sky130_fd_sc_hd__a21oi_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_148_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07942__B1 _01925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08763_ net9 _02744_ _03469_ vssd1 vssd1 vccd1 vccd1 _03470_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout183_A net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07714_ _02367_ _02420_ vssd1 vssd1 vccd1 vccd1 _02421_ sky130_fd_sc_hd__xor2_1
XTAP_2709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08694_ _03397_ _03400_ vssd1 vssd1 vccd1 vccd1 _03401_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07940__A net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07645_ genblk2\[11\].wave_shpr.div.fin_quo\[0\] genblk2\[11\].wave_shpr.div.fin_quo\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02352_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07576_ genblk1\[9\].osc.clkdiv_C.cnt\[6\] _01512_ _01234_ genblk1\[9\].osc.clkdiv_C.cnt\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02283_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_75_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10057__A1 _01329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09315_ net1004 _03870_ _03877_ _03899_ vssd1 vssd1 vccd1 vccd1 _00160_ sky130_fd_sc_hd__a22o_1
X_06527_ net1051 _01452_ vssd1 vssd1 vccd1 vccd1 genblk1\[2\].osc.clkdiv_C.next_cnt\[0\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_363 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06458_ _01373_ _01392_ _01393_ vssd1 vssd1 vccd1 vccd1 genblk1\[1\].osc.clkdiv_C.next_cnt\[8\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_118_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09246_ net522 _03845_ _03847_ net543 _03851_ vssd1 vssd1 vccd1 vccd1 _00139_ sky130_fd_sc_hd__a221o_1
XFILLER_0_90_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06681__B1 _01248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09177_ _03815_ vssd1 vssd1 vccd1 vccd1 _00106_ sky130_fd_sc_hd__clkbuf_1
X_06389_ _01179_ _01332_ _01225_ vssd1 vssd1 vccd1 vccd1 _01333_ sky130_fd_sc_hd__or3_1
X_08128_ _02826_ _02828_ _02832_ _02833_ _02834_ vssd1 vssd1 vccd1 vccd1 _02835_ sky130_fd_sc_hd__o311a_1
XFILLER_0_102_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08059_ genblk1\[5\].osc.clkdiv_C.cnt\[5\] _01238_ net36 genblk1\[5\].osc.clkdiv_C.cnt\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02766_ sky130_fd_sc_hd__o22a_1
XFILLER_0_101_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout96_A net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11070_ _05019_ net21 vssd1 vssd1 vccd1 vccd1 _05142_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10021_ genblk2\[3\].wave_shpr.div.acc\[22\] _04416_ vssd1 vssd1 vccd1 vccd1 _04417_
+ sky130_fd_sc_hd__or2_2
XFILLER_0_101_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11972_ genblk2\[10\].wave_shpr.div.fin_quo\[3\] genblk2\[10\].wave_shpr.div.quo\[2\]
+ _00003_ vssd1 vssd1 vccd1 vccd1 _05791_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_2_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13711_ clknet_leaf_31_clk _01022_ net100 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.b1\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10923_ _05046_ vssd1 vssd1 vccd1 vccd1 _00621_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07161__A1 genblk1\[9\].osc.clkdiv_C.cnt\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13642_ clknet_leaf_95_clk _00955_ net161 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.quo\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_10854_ genblk2\[6\].wave_shpr.div.b1\[8\] genblk2\[6\].wave_shpr.div.acc\[8\] vssd1
+ vssd1 vccd1 vccd1 _04998_ sky130_fd_sc_hd__and2b_1
XANTENNA__10048__A1 _01223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13573_ clknet_leaf_86_clk net227 net183 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.quo\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10785_ genblk2\[5\].wave_shpr.div.acc\[19\] _04938_ vssd1 vssd1 vccd1 vccd1 _04941_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_27_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06185__B _01097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11796__A1 _03694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09777__A _03701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12524_ clknet_leaf_59_clk _00076_ net193 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.b1\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06672__B1 _01498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12480__RESET_B net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12455_ clknet_leaf_33_clk net4 net101 vssd1 vssd1 vccd1 vccd1 modein.delay_octave_down_in\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_151_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11406_ genblk2\[8\].wave_shpr.div.b1\[4\] genblk2\[8\].wave_shpr.div.acc\[4\] vssd1
+ vssd1 vccd1 vccd1 _05382_ sky130_fd_sc_hd__and2b_1
XFILLER_0_34_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12386_ genblk2\[11\].wave_shpr.div.acc\[9\] _06061_ _06055_ vssd1 vssd1 vccd1 vccd1
+ _06062_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_316 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11337_ net924 _05311_ _05315_ _05327_ vssd1 vssd1 vccd1 vccd1 _00754_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11268_ genblk2\[7\].wave_shpr.div.b1\[0\] _05222_ genblk2\[7\].wave_shpr.div.acc\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05275_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13007_ clknet_leaf_138_clk net606 net40 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.acc\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11547__A _05444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12142__S _05865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10219_ net1055 _04518_ _04522_ _04542_ vssd1 vssd1 vccd1 vccd1 _00421_ sky130_fd_sc_hd__a22o_1
X_11199_ _05240_ vssd1 vssd1 vccd1 vccd1 _00703_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09017__A _03689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07760__A _02362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11484__B1 _03687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07430_ _02169_ vssd1 vssd1 vccd1 vccd1 _00010_ sky130_fd_sc_hd__inv_2
XANTENNA__12028__A2 _05813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07361_ _02091_ _02116_ _02117_ vssd1 vssd1 vccd1 vccd1 _02118_ sky130_fd_sc_hd__and3_1
XFILLER_0_45_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09100_ genblk2\[0\].wave_shpr.div.acc\[15\] genblk2\[0\].wave_shpr.div.b1\[15\]
+ vssd1 vssd1 vccd1 vccd1 _03748_ sky130_fd_sc_hd__or2b_1
X_06312_ _01270_ _01271_ _01272_ vssd1 vssd1 vccd1 vccd1 _01273_ sky130_fd_sc_hd__and3_1
XFILLER_0_84_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07292_ _02026_ _02058_ vssd1 vssd1 vccd1 vccd1 _02059_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09031_ _02155_ vssd1 vssd1 vccd1 vccd1 _03701_ sky130_fd_sc_hd__buf_8
XFILLER_0_14_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06243_ genblk1\[0\].osc.clkdiv_C.cnt\[17\] _01197_ _01198_ vssd1 vssd1 vccd1 vccd1
+ _01205_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_4_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_794 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06174_ _01134_ _01136_ vssd1 vssd1 vccd1 vccd1 _01146_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08404__A1 _01201_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold301 genblk2\[1\].wave_shpr.div.quo\[13\] vssd1 vssd1 vccd1 vccd1 net519 sky130_fd_sc_hd__dlygate4sd3_1
Xhold312 genblk2\[9\].wave_shpr.div.quo\[17\] vssd1 vssd1 vccd1 vccd1 net530 sky130_fd_sc_hd__dlygate4sd3_1
Xhold323 genblk2\[9\].wave_shpr.div.quo\[13\] vssd1 vssd1 vccd1 vccd1 net541 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold334 genblk2\[1\].wave_shpr.div.quo\[17\] vssd1 vssd1 vccd1 vccd1 net552 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold345 genblk2\[7\].wave_shpr.div.quo\[1\] vssd1 vssd1 vccd1 vccd1 net563 sky130_fd_sc_hd__dlygate4sd3_1
Xhold356 genblk2\[2\].wave_shpr.div.quo\[9\] vssd1 vssd1 vccd1 vccd1 net574 sky130_fd_sc_hd__dlygate4sd3_1
Xhold367 genblk2\[7\].wave_shpr.div.quo\[17\] vssd1 vssd1 vccd1 vccd1 net585 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09626__S _04095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold378 genblk2\[4\].wave_shpr.div.quo\[14\] vssd1 vssd1 vccd1 vccd1 net596 sky130_fd_sc_hd__dlygate4sd3_1
X_09933_ net648 _04315_ _04322_ _04340_ vssd1 vssd1 vccd1 vccd1 _00337_ sky130_fd_sc_hd__a22o_1
Xhold389 genblk2\[3\].wave_shpr.div.quo\[21\] vssd1 vssd1 vccd1 vccd1 net607 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08707__A2 net25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09864_ genblk2\[2\].wave_shpr.div.acc\[3\] _04287_ _04214_ vssd1 vssd1 vccd1 vccd1
+ _04288_ sky130_fd_sc_hd__mux2_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10514__A2 _04657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1001 _03812_ vssd1 vssd1 vccd1 vccd1 net1219 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07915__B1 _01487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1012 genblk2\[9\].wave_shpr.div.b1\[3\] vssd1 vssd1 vccd1 vccd1 net1230 sky130_fd_sc_hd__dlygate4sd3_1
X_08815_ _03516_ _03520_ _03445_ _03450_ vssd1 vssd1 vccd1 vccd1 _03522_ sky130_fd_sc_hd__a211o_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1023 genblk2\[10\].wave_shpr.div.acc\[6\] vssd1 vssd1 vccd1 vccd1 net1241 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09795_ _02152_ genblk2\[2\].wave_shpr.div.busy _02162_ vssd1 vssd1 vccd1 vccd1 _04249_
+ sky130_fd_sc_hd__and3_1
Xhold1034 genblk1\[7\].osc.clkdiv_C.cnt\[1\] vssd1 vssd1 vccd1 vccd1 net1252 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1045 genblk2\[4\].wave_shpr.div.quo\[6\] vssd1 vssd1 vccd1 vccd1 net1263 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1056 genblk2\[1\].wave_shpr.div.b1\[7\] vssd1 vssd1 vccd1 vccd1 net1274 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1067 genblk2\[3\].wave_shpr.div.b1\[12\] vssd1 vssd1 vccd1 vccd1 net1285 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08746_ _02217_ _02553_ genblk2\[6\].wave_shpr.div.fin_quo\[0\] vssd1 vssd1 vccd1
+ vccd1 _03453_ sky130_fd_sc_hd__and3_1
XTAP_2506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1078 genblk1\[9\].osc.clkdiv_C.cnt\[12\] vssd1 vssd1 vccd1 vccd1 net1296 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1089 PWM.counter\[4\] vssd1 vssd1 vccd1 vccd1 net1307 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08677_ _03298_ _03333_ _03381_ _03382_ vssd1 vssd1 vccd1 vccd1 _03384_ sky130_fd_sc_hd__a211oi_1
XTAP_1805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07628_ genblk1\[11\].osc.clkdiv_C.cnt\[12\] _01256_ _02333_ _02334_ vssd1 vssd1
+ vccd1 vccd1 _02335_ sky130_fd_sc_hd__a211o_1
XTAP_1849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07559_ _01200_ genblk1\[9\].osc.clkdiv_C.cnt\[14\] _01361_ genblk1\[9\].osc.clkdiv_C.cnt\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02266_ sky130_fd_sc_hd__a211o_1
X_10570_ genblk2\[5\].wave_shpr.div.b1\[9\] genblk2\[5\].wave_shpr.div.acc\[9\] vssd1
+ vssd1 vccd1 vccd1 _04798_ sky130_fd_sc_hd__and2b_1
XFILLER_0_63_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09229_ _03725_ genblk1\[0\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 _03842_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_134_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12240_ genblk2\[11\].wave_shpr.div.acc\[19\] _05977_ vssd1 vssd1 vccd1 vccd1 _05978_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_121_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06406__B1 genblk1\[1\].osc.clkdiv_C.cnt\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12171_ genblk2\[10\].wave_shpr.div.acc\[25\] _05785_ _05914_ vssd1 vssd1 vccd1 vccd1
+ _05915_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_32_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07845__A net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11122_ genblk2\[7\].wave_shpr.div.acc\[0\] vssd1 vssd1 vccd1 vccd1 _05182_ sky130_fd_sc_hd__inv_2
XANTENNA__10047__A2_N _04432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold890 genblk2\[4\].wave_shpr.div.i\[1\] vssd1 vssd1 vccd1 vccd1 net1108 sky130_fd_sc_hd__dlygate4sd3_1
X_11053_ net818 _05119_ _05126_ _05129_ vssd1 vssd1 vccd1 vccd1 _00668_ sky130_fd_sc_hd__a22o_1
XANTENNA_hold944_A genblk1\[8\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10505__A2 _04715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10004_ _04368_ _04398_ _04399_ vssd1 vssd1 vccd1 vccd1 _04400_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11955_ _05733_ _05775_ _05776_ vssd1 vssd1 vccd1 vccd1 _05777_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_99_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08331__B1 _02526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10906_ _01805_ vssd1 vssd1 vccd1 vccd1 _05037_ sky130_fd_sc_hd__inv_2
X_11886_ genblk2\[9\].wave_shpr.div.acc\[23\] _05610_ vssd1 vssd1 vccd1 vccd1 _05716_
+ sky130_fd_sc_hd__and2_1
XANTENNA__11218__B1 _05250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13625_ clknet_leaf_68_clk _00938_ net194 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.b1\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10837_ genblk2\[6\].wave_shpr.div.b1\[2\] vssd1 vssd1 vccd1 vccd1 _04981_ sky130_fd_sc_hd__inv_2
XANTENNA__12661__RESET_B net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13556_ clknet_leaf_101_clk _00871_ net164 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08634__A1 genblk2\[8\].wave_shpr.div.fin_quo\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10768_ net835 _04918_ _04922_ _04928_ vssd1 vssd1 vccd1 vccd1 _00584_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12507_ clknet_leaf_103_clk _00069_ net156 vssd1 vssd1 vccd1 vccd1 PWM.final_in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_13487_ clknet_leaf_89_clk _00804_ net177 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.quo\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10699_ _04869_ genblk1\[5\].osc.clkdiv_C.cnt\[15\] vssd1 vssd1 vccd1 vccd1 _04877_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_113_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12438_ genblk2\[11\].wave_shpr.div.acc\[23\] _05979_ _06099_ vssd1 vssd1 vccd1 vccd1
+ _06100_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12369_ genblk2\[11\].wave_shpr.div.acc\[5\] _06048_ _05982_ vssd1 vssd1 vccd1 vccd1
+ _06049_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06930_ genblk1\[6\].osc.clkdiv_C.cnt\[9\] _01773_ vssd1 vssd1 vccd1 vccd1 _01775_
+ sky130_fd_sc_hd__and2_1
X_06861_ genblk1\[5\].osc.clkdiv_C.cnt\[14\] _01717_ vssd1 vssd1 vccd1 vccd1 _01719_
+ sky130_fd_sc_hd__and2_1
X_08600_ _03304_ _03306_ _03302_ vssd1 vssd1 vccd1 vccd1 _03307_ sky130_fd_sc_hd__a21o_1
X_09580_ net825 _04076_ _04080_ _04086_ vssd1 vssd1 vccd1 vccd1 _00238_ sky130_fd_sc_hd__a22o_1
X_06792_ _01659_ _01661_ _01662_ _01663_ vssd1 vssd1 vccd1 vccd1 _01664_ sky130_fd_sc_hd__or4_1
X_08531_ genblk2\[10\].wave_shpr.div.fin_quo\[0\] _02525_ _02307_ genblk2\[10\].wave_shpr.div.fin_quo\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03238_ sky130_fd_sc_hd__a22o_1
XFILLER_0_49_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08462_ _02742_ _03167_ _03168_ _02745_ vssd1 vssd1 vccd1 vccd1 _03169_ sky130_fd_sc_hd__o31a_1
XANTENNA__07676__A2 _01190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07413_ genblk2\[1\].wave_shpr.div.i\[1\] _02156_ genblk2\[1\].wave_shpr.div.i\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02157_ sky130_fd_sc_hd__or3b_1
XFILLER_0_148_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08393_ genblk1\[2\].osc.clkdiv_C.cnt\[10\] _01420_ _01431_ genblk1\[2\].osc.clkdiv_C.cnt\[9\]
+ vssd1 vssd1 vccd1 vccd1 _03100_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_92_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout146_A net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07344_ _02104_ vssd1 vssd1 vccd1 vccd1 genblk1\[11\].osc.clkdiv_C.next_cnt\[3\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09210__A _02170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07275_ genblk1\[10\].osc.clkdiv_C.cnt\[9\] _02046_ vssd1 vssd1 vccd1 vccd1 _02048_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_72_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06226_ _01178_ vssd1 vssd1 vccd1 vccd1 _01188_ sky130_fd_sc_hd__buf_4
X_09014_ genblk2\[9\].wave_shpr.div.busy genblk2\[9\].wave_shpr.div.i\[0\] _03686_
+ _03687_ vssd1 vssd1 vccd1 vccd1 _00071_ sky130_fd_sc_hd__o211a_1
XFILLER_0_41_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold120 smpl_rt_clkdiv.clkDiv_inst.cnt\[0\] vssd1 vssd1 vccd1 vccd1 net338 sky130_fd_sc_hd__dlymetal6s2s_1
X_06157_ _01113_ _01117_ _01128_ vssd1 vssd1 vccd1 vccd1 _01129_ sky130_fd_sc_hd__a21oi_1
Xhold131 genblk2\[9\].wave_shpr.div.quo\[16\] vssd1 vssd1 vccd1 vccd1 net349 sky130_fd_sc_hd__dlygate4sd3_1
Xhold142 _01090_ vssd1 vssd1 vccd1 vccd1 net360 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold153 _00723_ vssd1 vssd1 vccd1 vccd1 net371 sky130_fd_sc_hd__dlygate4sd3_1
Xhold164 _00763_ vssd1 vssd1 vccd1 vccd1 net382 sky130_fd_sc_hd__dlygate4sd3_1
Xhold175 genblk2\[2\].wave_shpr.div.quo\[17\] vssd1 vssd1 vccd1 vccd1 net393 sky130_fd_sc_hd__dlygate4sd3_1
Xhold186 genblk2\[8\].wave_shpr.div.quo\[7\] vssd1 vssd1 vccd1 vccd1 net404 sky130_fd_sc_hd__dlygate4sd3_1
Xhold197 _00212_ vssd1 vssd1 vccd1 vccd1 net415 sky130_fd_sc_hd__dlygate4sd3_1
X_09916_ genblk2\[2\].wave_shpr.div.acc\[15\] _04327_ _04301_ vssd1 vssd1 vccd1 vccd1
+ _04328_ sky130_fd_sc_hd__mux2_1
X_09847_ _04250_ vssd1 vssd1 vccd1 vccd1 _04275_ sky130_fd_sc_hd__inv_2
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09778_ net1297 _01487_ _04238_ vssd1 vssd1 vccd1 vccd1 _04239_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout59_A net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11448__A0 genblk2\[8\].wave_shpr.div.fin_quo\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_2303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08729_ _03434_ _03435_ genblk2\[2\].wave_shpr.div.fin_quo\[5\] _02468_ vssd1 vssd1
+ vccd1 vccd1 _03436_ sky130_fd_sc_hd__a2bb2o_1
XTAP_2325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08313__B1 _02525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11999__A1 _03687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11740_ _01099_ _01149_ _05622_ net497 vssd1 vssd1 vccd1 vccd1 _00862_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_68_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11671_ genblk2\[9\].wave_shpr.div.acc\[8\] genblk2\[9\].wave_shpr.div.b1\[8\] vssd1
+ vssd1 vccd1 vccd1 _05563_ sky130_fd_sc_hd__or2b_1
X_13410_ clknet_leaf_90_clk _00729_ net144 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.quo\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_48_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10622_ _04837_ vssd1 vssd1 vccd1 vccd1 _00529_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13341_ clknet_leaf_7_clk _00662_ net49 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.acc\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10553_ genblk2\[5\].wave_shpr.div.acc\[0\] vssd1 vssd1 vccd1 vccd1 _04781_ sky130_fd_sc_hd__inv_2
XFILLER_0_106_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13272_ clknet_leaf_136_clk _00595_ net41 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.acc\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10484_ net784 _04715_ _04722_ _04728_ vssd1 vssd1 vccd1 vccd1 _00500_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_550 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12223_ genblk2\[11\].wave_shpr.div.b1\[10\] genblk2\[11\].wave_shpr.div.acc\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05961_ sky130_fd_sc_hd__and2b_1
XFILLER_0_32_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09041__A1 _03706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12154_ net705 _05876_ _05883_ _05903_ vssd1 vssd1 vccd1 vccd1 _00995_ sky130_fd_sc_hd__a22o_1
X_11105_ _05049_ genblk2\[7\].wave_shpr.div.acc\[16\] vssd1 vssd1 vccd1 vccd1 _05165_
+ sky130_fd_sc_hd__nor2_1
X_12085_ _05752_ _05744_ vssd1 vssd1 vccd1 vccd1 _05851_ sky130_fd_sc_hd__or2b_1
X_11036_ _05004_ _04972_ vssd1 vssd1 vccd1 vccd1 _05116_ sky130_fd_sc_hd__or2b_1
XANTENNA__08552__B1 genblk2\[6\].wave_shpr.div.fin_quo\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_99_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12987_ clknet_leaf_125_clk net260 net69 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.acc_next\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11938_ genblk2\[10\].wave_shpr.div.b1\[7\] genblk2\[10\].wave_shpr.div.acc\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05760_ sky130_fd_sc_hd__and2b_1
XFILLER_0_24_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11869_ _05608_ _05646_ vssd1 vssd1 vccd1 vccd1 _05704_ sky130_fd_sc_hd__or2_1
XFILLER_0_27_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13608_ clknet_leaf_58_clk _00921_ net194 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.i\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_145_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09804__B1 _04252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_450 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13539_ clknet_leaf_100_clk _00854_ net165 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.fin_quo\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_42_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06373__B _01240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07060_ genblk1\[8\].osc.clkdiv_C.cnt\[7\] vssd1 vssd1 vccd1 vccd1 _01878_ sky130_fd_sc_hd__inv_2
XFILLER_0_140_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_30 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07485__A _02209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07043__B1 _01858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09176__S _03722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07962_ genblk1\[7\].osc.clkdiv_C.cnt\[14\] _01361_ vssd1 vssd1 vccd1 vccd1 _02669_
+ sky130_fd_sc_hd__nand2_1
X_09701_ genblk2\[2\].wave_shpr.div.b1\[4\] genblk2\[2\].wave_shpr.div.acc\[4\] vssd1
+ vssd1 vccd1 vccd1 _04181_ sky130_fd_sc_hd__and2b_1
X_06913_ _01761_ _01763_ _01764_ vssd1 vssd1 vccd1 vccd1 genblk1\[6\].osc.clkdiv_C.next_cnt\[2\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_4_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07893_ _02529_ _02594_ _02518_ _02598_ vssd1 vssd1 vccd1 vccd1 _02600_ sky130_fd_sc_hd__a22o_1
X_09632_ _04004_ _03954_ vssd1 vssd1 vccd1 vccd1 _04126_ sky130_fd_sc_hd__or2b_1
XANTENNA__07932__B genblk2\[8\].wave_shpr.div.fin_quo\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_06844_ genblk1\[5\].osc.clkdiv_C.cnt\[8\] genblk1\[5\].osc.clkdiv_C.cnt\[7\] _01705_
+ vssd1 vssd1 vccd1 vccd1 _01708_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09563_ _04045_ _04072_ _04073_ _04048_ genblk2\[1\].wave_shpr.div.acc\[1\] vssd1
+ vssd1 vccd1 vccd1 _00234_ sky130_fd_sc_hd__a32o_1
X_06775_ genblk1\[4\].osc.clkdiv_C.cnt\[15\] vssd1 vssd1 vccd1 vccd1 _01650_ sky130_fd_sc_hd__inv_2
X_08514_ _03208_ _03215_ vssd1 vssd1 vccd1 vccd1 _03221_ sky130_fd_sc_hd__or2b_1
X_09494_ _04037_ vssd1 vssd1 vccd1 vccd1 _00201_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10102__B1 _04454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08445_ _03140_ _03150_ _03151_ vssd1 vssd1 vccd1 vccd1 _03152_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_77_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_42_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08376_ _03081_ _03082_ vssd1 vssd1 vccd1 vccd1 _03083_ sky130_fd_sc_hd__nand2_1
XFILLER_0_92_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06609__B1 _01513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07327_ _02069_ _02072_ _02073_ _02090_ vssd1 vssd1 vccd1 vccd1 _02091_ sky130_fd_sc_hd__or4_4
XFILLER_0_144_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07258_ genblk1\[10\].osc.clkdiv_C.cnt\[4\] _02034_ vssd1 vssd1 vccd1 vccd1 _02036_
+ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_57_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07821__A2 _02521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06209_ _01170_ vssd1 vssd1 vccd1 vccd1 _01171_ sky130_fd_sc_hd__buf_4
X_07189_ genblk1\[9\].osc.clkdiv_C.cnt\[11\] genblk1\[9\].osc.clkdiv_C.cnt\[10\] _01974_
+ vssd1 vssd1 vccd1 vccd1 _01978_ sky130_fd_sc_hd__and3_1
XFILLER_0_131_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_100_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07585__A1 genblk1\[9\].osc.clkdiv_C.cnt\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_115_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08534__B1 _02308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12910_ clknet_leaf_33_clk _00241_ net100 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.acc\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_12841_ clknet_leaf_64_clk _00174_ net196 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.acc\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12772_ clknet_leaf_47_clk _00105_ net121 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.b1\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11723_ _05614_ vssd1 vssd1 vccd1 vccd1 _00853_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10644__A1 _03704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11654_ genblk2\[8\].wave_shpr.div.i\[1\] genblk2\[8\].wave_shpr.div.i\[0\] genblk2\[8\].wave_shpr.div.i\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05549_ sky130_fd_sc_hd__and3_1
XFILLER_0_126_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout70 net75 vssd1 vssd1 vccd1 vccd1 net70 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_25_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout81 net83 vssd1 vssd1 vccd1 vccd1 net81 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_154_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10605_ _04827_ vssd1 vssd1 vccd1 vccd1 _00522_ sky130_fd_sc_hd__clkbuf_1
Xfanout92 net94 vssd1 vssd1 vccd1 vccd1 net92 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_64_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11585_ genblk2\[8\].wave_shpr.div.acc\[8\] _05499_ _05493_ vssd1 vssd1 vccd1 vccd1
+ _05500_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10947__A2 _05052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13324_ clknet_leaf_26_clk _00645_ net87 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.quo\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10536_ _04649_ genblk2\[5\].wave_shpr.div.acc\[16\] vssd1 vssd1 vccd1 vccd1 _04764_
+ sky130_fd_sc_hd__nor2_1
X_13255_ clknet_leaf_2_clk _00578_ net51 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.acc\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10467_ _04651_ vssd1 vssd1 vccd1 vccd1 _04715_ sky130_fd_sc_hd__clkbuf_4
X_12206_ _05941_ _05942_ _05943_ vssd1 vssd1 vccd1 vccd1 _05944_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_20_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13186_ clknet_leaf_112_clk _00511_ net129 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.acc\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10398_ net680 _04661_ _04663_ genblk2\[4\].wave_shpr.div.quo\[15\] _04667_ vssd1
+ vssd1 vccd1 vccd1 _00475_ sky130_fd_sc_hd__a221o_1
XFILLER_0_103_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12137_ _05775_ _05890_ vssd1 vssd1 vccd1 vccd1 _05891_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12068_ _05835_ genblk1\[10\].osc.clkdiv_C.cnt\[16\] vssd1 vssd1 vccd1 vccd1 _05839_
+ sky130_fd_sc_hd__and2_1
XANTENNA__11555__A _05417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11019_ _04996_ _04976_ vssd1 vssd1 vccd1 vccd1 _05103_ sky130_fd_sc_hd__or2b_1
XFILLER_0_149_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06368__B _01221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_531 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06560_ net1256 _01470_ _01473_ vssd1 vssd1 vccd1 vccd1 genblk1\[2\].osc.clkdiv_C.next_cnt\[12\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_59_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06491_ genblk1\[2\].osc.clkdiv_C.cnt\[16\] _01363_ _01416_ vssd1 vssd1 vccd1 vccd1
+ _01417_ sky130_fd_sc_hd__o21a_1
XFILLER_0_51_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06303__A2 _01256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08230_ _02798_ _02931_ vssd1 vssd1 vccd1 vccd1 _02937_ sky130_fd_sc_hd__nand2_1
XFILLER_0_51_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_117_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08161_ genblk1\[3\].osc.clkdiv_C.cnt\[13\] _01498_ vssd1 vssd1 vccd1 vccd1 _02868_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_43_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10938__A2 _05052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07112_ _01886_ _01914_ vssd1 vssd1 vccd1 vccd1 _01915_ sky130_fd_sc_hd__nor2_1
X_08092_ _02791_ _02796_ _02798_ vssd1 vssd1 vccd1 vccd1 _02799_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_70_464 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07043_ genblk1\[8\].osc.clkdiv_C.cnt\[5\] _01487_ _01858_ genblk1\[8\].osc.clkdiv_C.cnt\[6\]
+ _01860_ vssd1 vssd1 vccd1 vccd1 _01861_ sky130_fd_sc_hd__a221o_1
XFILLER_0_140_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout109_A net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11899__B1 _03841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07567__A1 genblk1\[9\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08994_ sig_norm.quo\[10\] _01099_ _01157_ vssd1 vssd1 vccd1 vccd1 _03677_ sky130_fd_sc_hd__a21o_1
X_07945_ genblk1\[7\].osc.clkdiv_C.cnt\[5\] _01802_ _01805_ genblk1\[7\].osc.clkdiv_C.cnt\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02652_ sky130_fd_sc_hd__o22a_1
XANTENNA__07662__B _01182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07876_ _02517_ _02570_ _02566_ vssd1 vssd1 vccd1 vccd1 _02583_ sky130_fd_sc_hd__and3_1
X_09615_ _04046_ vssd1 vssd1 vccd1 vccd1 _04113_ sky130_fd_sc_hd__buf_2
X_06827_ _01697_ vssd1 vssd1 vccd1 vccd1 genblk1\[5\].osc.clkdiv_C.next_cnt\[1\] sky130_fd_sc_hd__clkbuf_1
X_09546_ _04055_ genblk1\[1\].osc.clkdiv_C.cnt\[11\] vssd1 vssd1 vccd1 vccd1 _04064_
+ sky130_fd_sc_hd__and2_1
X_06758_ genblk1\[4\].osc.clkdiv_C.cnt\[11\] genblk1\[4\].osc.clkdiv_C.cnt\[10\] _01631_
+ vssd1 vssd1 vccd1 vccd1 _01637_ sky130_fd_sc_hd__and3_1
XANTENNA__10626__A1 net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09477_ genblk2\[2\].wave_shpr.div.b1\[6\] _01437_ _04024_ vssd1 vssd1 vccd1 vccd1
+ _04027_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06689_ genblk1\[4\].osc.clkdiv_C.cnt\[12\] _01574_ _01578_ genblk1\[4\].osc.clkdiv_C.cnt\[16\]
+ vssd1 vssd1 vccd1 vccd1 _01579_ sky130_fd_sc_hd__a2bb2o_1
X_08428_ _03129_ _03133_ _03010_ vssd1 vssd1 vccd1 vccd1 _03135_ sky130_fd_sc_hd__o21a_1
XFILLER_0_93_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06294__A _01255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08359_ _03060_ _03065_ vssd1 vssd1 vccd1 vccd1 _03066_ sky130_fd_sc_hd__xor2_1
XANTENNA__08047__A2 _01666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11370_ genblk2\[7\].wave_shpr.div.i\[1\] genblk2\[7\].wave_shpr.div.i\[0\] vssd1
+ vssd1 vccd1 vccd1 _05350_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07053__A1_N genblk1\[8\].osc.clkdiv_C.cnt\[12\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10321_ _04628_ vssd1 vssd1 vccd1 vccd1 _00437_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13040_ clknet_leaf_126_clk _00367_ net61 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.b1\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10252_ net333 _04563_ _04564_ vssd1 vssd1 vccd1 vccd1 _00432_ sky130_fd_sc_hd__a21oi_1
X_10183_ _04401_ _04367_ vssd1 vssd1 vccd1 vccd1 _04515_ sky130_fd_sc_hd__or2b_1
X_12824_ clknet_leaf_62_clk _00157_ net189 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.acc\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12067__B1 _05815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12755_ clknet_leaf_52_clk genblk1\[11\].osc.clkdiv_C.next_cnt\[14\] net110 vssd1
+ vssd1 vccd1 vccd1 genblk1\[11\].osc.clkdiv_C.cnt\[14\] sky130_fd_sc_hd__dfrtp_1
XTAP_1251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10093__A2 _04452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11706_ genblk2\[9\].wave_shpr.div.b1\[13\] genblk2\[9\].wave_shpr.div.acc\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05598_ sky130_fd_sc_hd__and2b_1
XFILLER_0_126_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12686_ clknet_leaf_119_clk genblk1\[7\].osc.clkdiv_C.next_cnt\[17\] net141 vssd1
+ vssd1 vccd1 vccd1 genblk1\[7\].osc.clkdiv_C.cnt\[17\] sky130_fd_sc_hd__dfrtp_1
X_11637_ genblk2\[8\].wave_shpr.div.acc\[22\] _05411_ vssd1 vssd1 vccd1 vccd1 _05538_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_126_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11568_ genblk2\[8\].wave_shpr.div.acc\[4\] _05486_ _05417_ vssd1 vssd1 vccd1 vccd1
+ _05487_ sky130_fd_sc_hd__mux2_1
XFILLER_0_141_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08994__B1 _01157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold708 genblk2\[4\].wave_shpr.div.acc\[17\] vssd1 vssd1 vccd1 vccd1 net926 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13307_ clknet_leaf_122_clk _00628_ net137 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.quo\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold719 genblk2\[4\].wave_shpr.div.acc\[2\] vssd1 vssd1 vccd1 vccd1 net937 sky130_fd_sc_hd__dlygate4sd3_1
X_10519_ genblk2\[4\].wave_shpr.div.acc\[25\] _04751_ vssd1 vssd1 vccd1 vccd1 _04753_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07747__B _01172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11499_ net709 _05442_ _05446_ net871 vssd1 vssd1 vccd1 vccd1 _00797_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13238_ clknet_leaf_11_clk net236 net57 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.quo\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_862 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13169_ clknet_leaf_127_clk _00494_ net66 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.acc\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09454__S _00007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_137_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07730_ _01188_ genblk1\[1\].osc.clkdiv_C.cnt\[7\] vssd1 vssd1 vccd1 vccd1 _02437_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_137_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07661_ genblk1\[10\].osc.clkdiv_C.cnt\[7\] _01190_ _01235_ genblk1\[10\].osc.clkdiv_C.cnt\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02368_ sky130_fd_sc_hd__o22ai_1
XANTENNA__06524__A2 _01231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07721__A1 genblk1\[1\].osc.clkdiv_C.cnt\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09400_ genblk2\[1\].wave_shpr.div.acc\[7\] genblk2\[1\].wave_shpr.div.b1\[7\] vssd1
+ vssd1 vccd1 vccd1 _03964_ sky130_fd_sc_hd__or2b_1
X_06612_ genblk1\[3\].osc.clkdiv_C.cnt\[1\] _01519_ vssd1 vssd1 vccd1 vccd1 _01520_
+ sky130_fd_sc_hd__xor2_1
XANTENNA__08594__A net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07592_ _02298_ _02269_ _02272_ _02267_ vssd1 vssd1 vccd1 vccd1 _02299_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_88_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09331_ _03790_ _03911_ vssd1 vssd1 vccd1 vccd1 _03912_ sky130_fd_sc_hd__xnor2_1
X_06543_ _01452_ _01461_ _01462_ vssd1 vssd1 vccd1 vccd1 genblk1\[2\].osc.clkdiv_C.next_cnt\[6\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_5_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09262_ net454 _03835_ _03838_ net476 _03860_ vssd1 vssd1 vccd1 vccd1 _00146_ sky130_fd_sc_hd__a221o_1
X_06474_ net29 _01403_ vssd1 vssd1 vccd1 vccd1 _01404_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08213_ _02917_ _02916_ vssd1 vssd1 vccd1 vccd1 _02920_ sky130_fd_sc_hd__xnor2_1
X_09193_ _03824_ vssd1 vssd1 vccd1 vccd1 _00113_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09226__B2 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_488 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08144_ genblk1\[3\].osc.clkdiv_C.cnt\[15\] _01576_ vssd1 vssd1 vccd1 vccd1 _02851_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08075_ genblk1\[5\].osc.clkdiv_C.cnt\[8\] _01678_ _01726_ genblk1\[5\].osc.clkdiv_C.cnt\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02782_ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07026_ genblk1\[7\].osc.clkdiv_C.cnt\[15\] _01846_ vssd1 vssd1 vccd1 vccd1 _01847_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_87_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold13 genblk2\[7\].wave_shpr.div.quo\[19\] vssd1 vssd1 vccd1 vccd1 net231 sky130_fd_sc_hd__dlygate4sd3_1
X_08977_ _03519_ _03662_ vssd1 vssd1 vccd1 vccd1 _03663_ sky130_fd_sc_hd__xnor2_1
Xhold24 _00634_ vssd1 vssd1 vccd1 vccd1 net242 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 genblk2\[5\].wave_shpr.div.quo\[5\] vssd1 vssd1 vccd1 vccd1 net253 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 _00813_ vssd1 vssd1 vccd1 vccd1 net264 sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 genblk2\[2\].wave_shpr.div.quo\[7\] vssd1 vssd1 vccd1 vccd1 net275 sky130_fd_sc_hd__dlygate4sd3_1
X_07928_ _02632_ _02633_ _02634_ genblk1\[8\].osc.clkdiv_C.cnt\[17\] genblk1\[8\].osc.clkdiv_C.cnt\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02635_ sky130_fd_sc_hd__a311oi_2
Xhold68 PWM.final_sample_in\[7\] vssd1 vssd1 vccd1 vccd1 net286 sky130_fd_sc_hd__dlygate4sd3_1
Xhold79 _00395_ vssd1 vssd1 vccd1 vccd1 net297 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06289__A _01246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07859_ _02563_ _02564_ _02565_ _02509_ vssd1 vssd1 vccd1 vccd1 _02566_ sky130_fd_sc_hd__a211o_1
XFILLER_0_98_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10870_ _04967_ _05013_ vssd1 vssd1 vccd1 vccd1 _05014_ sky130_fd_sc_hd__and2b_1
XFILLER_0_79_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09529_ net537 _04052_ _04053_ net645 _04054_ vssd1 vssd1 vccd1 vccd1 _00219_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12540_ clknet_leaf_62_clk _00092_ net189 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.b1\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_47_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12471_ clknet_leaf_31_clk smpl_rt_clkdiv.clkDiv_inst.next_cnt\[5\] net100 vssd1
+ vssd1 vccd1 vccd1 smpl_rt_clkdiv.clkDiv_inst.cnt\[5\] sky130_fd_sc_hd__dfrtp_1
X_11422_ genblk2\[8\].wave_shpr.div.b1\[12\] genblk2\[8\].wave_shpr.div.acc\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05398_ sky130_fd_sc_hd__and2b_1
XANTENNA__07228__B1 _01227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07779__A1 _01181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11353_ _05218_ _05273_ _05336_ genblk2\[7\].wave_shpr.div.acc\[21\] vssd1 vssd1
+ vccd1 vccd1 _05339_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_104_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_105_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10304_ genblk2\[4\].wave_shpr.div.b1\[17\] genblk2\[4\].wave_shpr.div.acc\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04616_ sky130_fd_sc_hd__and2b_1
X_11284_ _05179_ _05189_ vssd1 vssd1 vccd1 vccd1 _05287_ sky130_fd_sc_hd__xor2_1
XANTENNA__08728__B1 _02224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13023_ clknet_leaf_113_clk _00350_ net128 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.fin_quo\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_10235_ _04552_ _04549_ _04553_ vssd1 vssd1 vccd1 vccd1 _04554_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09782__B _01490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10166_ _04393_ _04371_ vssd1 vssd1 vccd1 vccd1 _04502_ sky130_fd_sc_hd__or2b_1
XANTENNA__08398__B _01349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10097_ _04269_ genblk1\[3\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 _04458_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_88_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12807_ clknet_leaf_59_clk _00140_ net187 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.quo\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10999_ _04985_ _05087_ vssd1 vssd1 vccd1 vccd1 _05088_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_84_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12738_ clknet_leaf_38_clk genblk1\[10\].osc.clkdiv_C.next_cnt\[15\] net114 vssd1
+ vssd1 vccd1 vccd1 genblk1\[10\].osc.clkdiv_C.cnt\[15\] sky130_fd_sc_hd__dfrtp_2
XTAP_1081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_45_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12669_ clknet_leaf_90_clk genblk1\[7\].osc.clkdiv_C.next_cnt\[0\] net173 vssd1 vssd1
+ vccd1 vccd1 genblk1\[7\].osc.clkdiv_C.cnt\[0\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_115_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06190_ net642 net361 vssd1 vssd1 vccd1 vccd1 PWM.next_counter\[1\] sky130_fd_sc_hd__xor2_1
XFILLER_0_13_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold505 genblk2\[10\].wave_shpr.div.quo\[4\] vssd1 vssd1 vccd1 vccd1 net723 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07477__B _02153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08431__A2 net32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold516 genblk2\[4\].wave_shpr.div.i\[2\] vssd1 vssd1 vccd1 vccd1 net734 sky130_fd_sc_hd__dlygate4sd3_1
Xhold527 genblk2\[5\].wave_shpr.div.quo\[3\] vssd1 vssd1 vccd1 vccd1 net745 sky130_fd_sc_hd__dlygate4sd3_1
Xhold538 genblk2\[6\].wave_shpr.div.quo\[1\] vssd1 vssd1 vccd1 vccd1 net756 sky130_fd_sc_hd__dlygate4sd3_1
Xhold549 genblk2\[11\].wave_shpr.div.quo\[4\] vssd1 vssd1 vccd1 vccd1 net767 sky130_fd_sc_hd__buf_1
XFILLER_0_110_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08900_ sig_norm.acc\[2\] _03596_ vssd1 vssd1 vccd1 vccd1 _03604_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09880_ _04186_ _04299_ vssd1 vssd1 vccd1 vccd1 _04300_ sky130_fd_sc_hd__xnor2_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07493__A modein.delay_in\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08831_ _03531_ _03536_ _03537_ vssd1 vssd1 vccd1 vccd1 _03538_ sky130_fd_sc_hd__and3_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12279__A0 _01308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08762_ genblk2\[3\].wave_shpr.div.fin_quo\[0\] _02539_ _02939_ vssd1 vssd1 vccd1
+ vccd1 _03469_ sky130_fd_sc_hd__a21o_1
X_07713_ _02414_ _02417_ _02419_ vssd1 vssd1 vccd1 vccd1 _02420_ sky130_fd_sc_hd__a21bo_1
X_08693_ _03398_ _03399_ vssd1 vssd1 vccd1 vccd1 _03400_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout176_A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11743__A _02203_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07940__B _02364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07644_ _02350_ vssd1 vssd1 vccd1 vccd1 _02351_ sky130_fd_sc_hd__buf_2
XFILLER_0_76_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07575_ genblk1\[9\].osc.clkdiv_C.cnt\[4\] _01925_ _02280_ _02281_ vssd1 vssd1 vccd1
+ vccd1 _02282_ sky130_fd_sc_hd__a211o_1
X_09314_ genblk2\[0\].wave_shpr.div.acc\[10\] _03898_ _03889_ vssd1 vssd1 vccd1 vccd1
+ _03899_ sky130_fd_sc_hd__mux2_1
X_06526_ _01451_ vssd1 vssd1 vccd1 vccd1 _01452_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_8_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_898 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09245_ _03725_ genblk1\[0\].osc.clkdiv_C.cnt\[7\] vssd1 vssd1 vccd1 vccd1 _03851_
+ sky130_fd_sc_hd__and2_1
X_06457_ genblk1\[1\].osc.clkdiv_C.cnt\[7\] _01387_ genblk1\[1\].osc.clkdiv_C.cnt\[8\]
+ vssd1 vssd1 vccd1 vccd1 _01393_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09176_ genblk2\[10\].wave_shpr.div.b1\[1\] _01368_ _03722_ vssd1 vssd1 vccd1 vccd1
+ _03815_ sky130_fd_sc_hd__mux2_1
X_06388_ _01194_ _01176_ vssd1 vssd1 vccd1 vccd1 _01332_ sky130_fd_sc_hd__and2b_1
XFILLER_0_71_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08127_ _02830_ _02827_ _02831_ _02829_ vssd1 vssd1 vccd1 vccd1 _02834_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_133_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08058_ genblk1\[5\].osc.clkdiv_C.cnt\[6\] _01172_ _01180_ _02764_ vssd1 vssd1 vccd1
+ vccd1 _02765_ sky130_fd_sc_hd__a31o_1
XFILLER_0_141_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07009_ _01823_ _01835_ _01836_ vssd1 vssd1 vccd1 vccd1 genblk1\[7\].osc.clkdiv_C.next_cnt\[8\]
+ sky130_fd_sc_hd__nor3_1
X_10020_ genblk2\[3\].wave_shpr.div.acc\[21\] genblk2\[3\].wave_shpr.div.acc\[20\]
+ genblk2\[3\].wave_shpr.div.acc\[19\] _04415_ vssd1 vssd1 vccd1 vccd1 _04416_ sky130_fd_sc_hd__or4_1
X_11971_ _05790_ vssd1 vssd1 vccd1 vccd1 _00925_ sky130_fd_sc_hd__clkbuf_1
X_13710_ clknet_leaf_31_clk _01021_ net103 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.b1\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10922_ net1301 _01811_ _05042_ vssd1 vssd1 vccd1 vccd1 _05046_ sky130_fd_sc_hd__mux2_1
XANTENNA__07161__A2 genblk1\[9\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13641_ clknet_leaf_94_clk _00954_ net160 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10853_ _04976_ _04995_ _04996_ vssd1 vssd1 vccd1 vccd1 _04997_ sky130_fd_sc_hd__a21o_1
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13572_ clknet_leaf_85_clk _00887_ net184 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.quo\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10784_ net896 _04918_ _04922_ _04940_ vssd1 vssd1 vccd1 vccd1 _00588_ sky130_fd_sc_hd__a22o_1
XPHY_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11799__S _05613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12523_ clknet_leaf_103_clk PWM.next_counter\[7\] net157 vssd1 vssd1 vccd1 vccd1
+ PWM.counter\[7\] sky130_fd_sc_hd__dfrtp_1
XPHY_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08661__A2 _02789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12454_ clknet_leaf_39_clk net228 net115 vssd1 vssd1 vccd1 vccd1 modein.delay_octave_up_in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11405_ _05372_ _05379_ _05380_ vssd1 vssd1 vccd1 vccd1 _05381_ sky130_fd_sc_hd__a21o_1
XFILLER_0_78_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12385_ _05958_ _06060_ vssd1 vssd1 vccd1 vccd1 _06061_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09071__C1 _03728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11336_ genblk2\[7\].wave_shpr.div.acc\[16\] _05326_ _05300_ vssd1 vssd1 vccd1 vccd1
+ _05327_ sky130_fd_sc_hd__mux2_1
X_11267_ _05273_ _05182_ genblk2\[7\].wave_shpr.div.b1\[0\] vssd1 vssd1 vccd1 vccd1
+ _05274_ sky130_fd_sc_hd__or3b_1
XFILLER_0_120_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09374__A0 _03941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13006_ clknet_leaf_133_clk net581 net40 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.acc\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10218_ net904 _04415_ _04541_ vssd1 vssd1 vccd1 vccd1 _04542_ sky130_fd_sc_hd__a21bo_1
X_11198_ genblk2\[8\].wave_shpr.div.b1\[10\] _05239_ _05237_ vssd1 vssd1 vccd1 vccd1
+ _05240_ sky130_fd_sc_hd__mux2_1
X_10149_ net1057 _04486_ _04456_ _04489_ vssd1 vssd1 vccd1 vccd1 _00404_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07688__B1 _02011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07360_ genblk1\[11\].osc.clkdiv_C.cnt\[7\] _02112_ vssd1 vssd1 vccd1 vccd1 _02117_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_85_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06311_ genblk1\[0\].osc.clkdiv_C.cnt\[1\] genblk1\[0\].osc.clkdiv_C.cnt\[0\] vssd1
+ vssd1 vccd1 vccd1 _01272_ sky130_fd_sc_hd__nand2_1
XFILLER_0_155_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07291_ genblk1\[10\].osc.clkdiv_C.cnt\[15\] _02057_ vssd1 vssd1 vccd1 vccd1 _02058_
+ sky130_fd_sc_hd__and2_1
X_09030_ genblk2\[9\].wave_shpr.div.busy _03698_ net817 vssd1 vssd1 vccd1 vccd1 _03700_
+ sky130_fd_sc_hd__a21oi_1
X_06242_ genblk1\[0\].osc.clkdiv_C.cnt\[9\] _01193_ _01199_ _01202_ _01203_ vssd1
+ vssd1 vccd1 vccd1 _01204_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_150_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_143_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06392__A _01179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06173_ _01141_ _01143_ vssd1 vssd1 vccd1 vccd1 _01145_ sky130_fd_sc_hd__xor2_1
XFILLER_0_142_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold302 genblk2\[2\].wave_shpr.div.quo\[23\] vssd1 vssd1 vccd1 vccd1 net520 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold313 genblk2\[4\].wave_shpr.div.quo\[17\] vssd1 vssd1 vccd1 vccd1 net531 sky130_fd_sc_hd__dlygate4sd3_1
Xhold324 genblk2\[7\].wave_shpr.div.quo\[21\] vssd1 vssd1 vccd1 vccd1 net542 sky130_fd_sc_hd__dlygate4sd3_1
Xhold335 genblk2\[2\].wave_shpr.div.quo\[12\] vssd1 vssd1 vccd1 vccd1 net553 sky130_fd_sc_hd__dlygate4sd3_1
Xhold346 _00713_ vssd1 vssd1 vccd1 vccd1 net564 sky130_fd_sc_hd__dlygate4sd3_1
Xhold357 genblk2\[8\].wave_shpr.div.quo\[21\] vssd1 vssd1 vccd1 vccd1 net575 sky130_fd_sc_hd__dlygate4sd3_1
X_09932_ net605 _04336_ _04339_ vssd1 vssd1 vccd1 vccd1 _04340_ sky130_fd_sc_hd__a21o_1
XANTENNA__11738__A _02248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold368 genblk2\[9\].wave_shpr.div.quo\[4\] vssd1 vssd1 vccd1 vccd1 net586 sky130_fd_sc_hd__dlygate4sd3_1
Xhold379 _00474_ vssd1 vssd1 vccd1 vccd1 net597 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09863_ _04178_ _04286_ vssd1 vssd1 vccd1 vccd1 _04287_ sky130_fd_sc_hd__xnor2_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07915__A1 genblk1\[8\].osc.clkdiv_C.cnt\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08814_ _03445_ _03450_ _03516_ _03520_ vssd1 vssd1 vccd1 vccd1 _03521_ sky130_fd_sc_hd__o211ai_2
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07915__B2 genblk1\[8\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1002 genblk1\[11\].osc.clkdiv_C.cnt\[17\] vssd1 vssd1 vccd1 vccd1 net1220 sky130_fd_sc_hd__clkbuf_2
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1013 genblk2\[9\].wave_shpr.div.b1\[10\] vssd1 vssd1 vccd1 vccd1 net1231 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09794_ _04247_ vssd1 vssd1 vccd1 vccd1 _04248_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1024 genblk2\[11\].wave_shpr.div.b1\[6\] vssd1 vssd1 vccd1 vccd1 net1242 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1035 genblk2\[7\].wave_shpr.div.b1\[10\] vssd1 vssd1 vccd1 vccd1 net1253 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1046 _04631_ vssd1 vssd1 vccd1 vccd1 net1264 sky130_fd_sc_hd__dlygate4sd3_1
X_08745_ _03256_ _03257_ vssd1 vssd1 vccd1 vccd1 _03452_ sky130_fd_sc_hd__nand2_1
Xhold1057 genblk2\[11\].wave_shpr.div.b1\[7\] vssd1 vssd1 vccd1 vccd1 net1275 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1068 genblk2\[7\].wave_shpr.div.b1\[9\] vssd1 vssd1 vccd1 vccd1 net1286 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1079 genblk2\[3\].wave_shpr.div.b1\[11\] vssd1 vssd1 vccd1 vccd1 net1297 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11475__A1 net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08676_ _03298_ _03333_ _03381_ _03382_ vssd1 vssd1 vccd1 vccd1 _03383_ sky130_fd_sc_hd__a211o_1
XFILLER_0_67_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07627_ genblk1\[11\].osc.clkdiv_C.cnt\[13\] _01209_ _01256_ genblk1\[11\].osc.clkdiv_C.cnt\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02334_ sky130_fd_sc_hd__o22ai_1
XTAP_1839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07558_ genblk2\[9\].wave_shpr.div.fin_quo\[4\] _02264_ vssd1 vssd1 vccd1 vccd1 _02265_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_36_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06509_ _01416_ _01365_ _01326_ genblk1\[2\].osc.clkdiv_C.cnt\[11\] genblk1\[2\].osc.clkdiv_C.cnt\[16\]
+ vssd1 vssd1 vccd1 vccd1 _01435_ sky130_fd_sc_hd__a221o_1
XFILLER_0_90_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07489_ _02147_ _02212_ vssd1 vssd1 vccd1 vccd1 _02213_ sky130_fd_sc_hd__nor2_1
XANTENNA__10986__B1 _05054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09228_ _03835_ vssd1 vssd1 vccd1 vccd1 _03841_ sky130_fd_sc_hd__clkbuf_4
X_09159_ genblk2\[0\].wave_shpr.div.fin_quo\[1\] genblk2\[0\].wave_shpr.div.quo\[0\]
+ _00001_ vssd1 vssd1 vccd1 vccd1 _03806_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06406__A1 _01201_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12170_ _05785_ genblk2\[10\].wave_shpr.div.acc\[25\] genblk2\[10\].wave_shpr.div.acc\[26\]
+ vssd1 vssd1 vccd1 vccd1 _05914_ sky130_fd_sc_hd__or3b_1
XFILLER_0_102_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06957__A2 _01227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11121_ genblk2\[7\].wave_shpr.div.acc\[2\] genblk2\[7\].wave_shpr.div.b1\[2\] vssd1
+ vssd1 vccd1 vccd1 _05181_ sky130_fd_sc_hd__or2b_1
XFILLER_0_7_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold880 genblk2\[8\].wave_shpr.div.i\[1\] vssd1 vssd1 vccd1 vccd1 net1098 sky130_fd_sc_hd__dlygate4sd3_1
Xhold891 genblk2\[1\].wave_shpr.div.acc\[21\] vssd1 vssd1 vccd1 vccd1 net1109 sky130_fd_sc_hd__dlygate4sd3_1
X_11052_ genblk2\[6\].wave_shpr.div.acc\[14\] _05128_ _05105_ vssd1 vssd1 vccd1 vccd1
+ _05129_ sky130_fd_sc_hd__mux2_1
XANTENNA__11163__A0 genblk2\[7\].wave_shpr.div.fin_quo\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10003_ genblk2\[3\].wave_shpr.div.b1\[10\] genblk2\[3\].wave_shpr.div.acc\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04399_ sky130_fd_sc_hd__and2b_1
XFILLER_0_99_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_4_13_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11466__A1 _02433_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11954_ genblk2\[10\].wave_shpr.div.b1\[15\] genblk2\[10\].wave_shpr.div.acc\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05776_ sky130_fd_sc_hd__and2b_1
XFILLER_0_59_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10905_ _05036_ vssd1 vssd1 vccd1 vccd1 _00613_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11885_ genblk2\[9\].wave_shpr.div.acc\[23\] _05610_ vssd1 vssd1 vccd1 vccd1 _05715_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13624_ clknet_leaf_68_clk _00937_ net194 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.b1\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10836_ genblk2\[6\].wave_shpr.div.acc\[3\] genblk2\[6\].wave_shpr.div.b1\[3\] vssd1
+ vssd1 vccd1 vccd1 _04980_ sky130_fd_sc_hd__or2b_1
XFILLER_0_39_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13555_ clknet_leaf_101_clk net587 net164 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10767_ genblk2\[5\].wave_shpr.div.acc\[14\] _04927_ _04907_ vssd1 vssd1 vccd1 vccd1
+ _04928_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08634__A2 genblk2\[8\].wave_shpr.div.fin_quo\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_137_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12506_ clknet_leaf_104_clk _00068_ net154 vssd1 vssd1 vccd1 vccd1 PWM.final_in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13486_ clknet_leaf_79_clk net405 net206 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.quo\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10698_ net459 _02183_ _04856_ net471 _04876_ vssd1 vssd1 vccd1 vccd1 _00566_ sky130_fd_sc_hd__a221o_1
XFILLER_0_35_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12437_ _05980_ _06088_ vssd1 vssd1 vccd1 vccd1 _06099_ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12368_ _06047_ _05950_ vssd1 vssd1 vccd1 vccd1 _06048_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11319_ genblk2\[7\].wave_shpr.div.acc\[12\] _05313_ _05300_ vssd1 vssd1 vccd1 vccd1
+ _05314_ sky130_fd_sc_hd__mux2_1
X_12299_ net430 _06009_ _06010_ _05982_ vssd1 vssd1 vccd1 vccd1 _01033_ sky130_fd_sc_hd__a22o_1
X_06860_ net1229 _01715_ _01718_ vssd1 vssd1 vccd1 vccd1 genblk1\[5\].osc.clkdiv_C.next_cnt\[13\]
+ sky130_fd_sc_hd__o21a_1
XANTENNA__09462__S _00007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06791_ genblk1\[5\].osc.clkdiv_C.cnt\[16\] _01578_ vssd1 vssd1 vccd1 vccd1 _01663_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08530_ _03141_ _03236_ net3 net163 vssd1 vssd1 vccd1 vccd1 _03237_ sky130_fd_sc_hd__o211a_1
XFILLER_0_54_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08461_ _02217_ _02553_ genblk2\[6\].wave_shpr.div.fin_quo\[4\] vssd1 vssd1 vccd1
+ vccd1 _03168_ sky130_fd_sc_hd__and3_1
XFILLER_0_148_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07412_ genblk2\[1\].wave_shpr.div.i\[2\] genblk2\[1\].wave_shpr.div.i\[3\] genblk2\[1\].wave_shpr.div.i\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02156_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_46_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08392_ genblk1\[2\].osc.clkdiv_C.cnt\[9\] _01431_ _03096_ _03097_ _03098_ vssd1
+ vssd1 vccd1 vccd1 _03099_ sky130_fd_sc_hd__o221a_1
XFILLER_0_85_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07343_ _02092_ _02102_ _02103_ vssd1 vssd1 vccd1 vccd1 _02104_ sky130_fd_sc_hd__and3_1
XFILLER_0_45_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07274_ _02027_ _02046_ _02047_ vssd1 vssd1 vccd1 vccd1 genblk1\[10\].osc.clkdiv_C.next_cnt\[8\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_61_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_72_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09013_ _02171_ vssd1 vssd1 vccd1 vccd1 _03687_ sky130_fd_sc_hd__buf_6
XFILLER_0_14_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06225_ _01176_ vssd1 vssd1 vccd1 vccd1 _01187_ sky130_fd_sc_hd__buf_4
XFILLER_0_5_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_214 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold110 genblk2\[7\].wave_shpr.div.i\[4\] vssd1 vssd1 vccd1 vccd1 net328 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08389__B2 _02011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06156_ _01126_ _01127_ vssd1 vssd1 vccd1 vccd1 _01128_ sky130_fd_sc_hd__or2_1
Xhold121 genblk2\[2\].wave_shpr.div.quo\[18\] vssd1 vssd1 vccd1 vccd1 net339 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold132 _00882_ vssd1 vssd1 vccd1 vccd1 net350 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_1_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold143 PWM.counter\[0\] vssd1 vssd1 vccd1 vccd1 net361 sky130_fd_sc_hd__buf_1
Xhold154 sig_norm.quo\[8\] vssd1 vssd1 vccd1 vccd1 net372 sky130_fd_sc_hd__dlygate4sd3_1
Xhold165 genblk2\[10\].wave_shpr.div.quo\[20\] vssd1 vssd1 vccd1 vccd1 net383 sky130_fd_sc_hd__dlygate4sd3_1
Xhold176 genblk2\[0\].wave_shpr.div.b1\[6\] vssd1 vssd1 vccd1 vccd1 net394 sky130_fd_sc_hd__dlygate4sd3_1
Xhold187 _00803_ vssd1 vssd1 vccd1 vccd1 net405 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold198 genblk2\[9\].wave_shpr.div.quo\[21\] vssd1 vssd1 vccd1 vccd1 net416 sky130_fd_sc_hd__dlygate4sd3_1
X_09915_ _04202_ _04326_ vssd1 vssd1 vccd1 vccd1 _04327_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10499__A2 _04715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09846_ genblk2\[2\].wave_shpr.div.acc_next\[0\] _04247_ _04250_ net259 _04274_ vssd1
+ vssd1 vccd1 vccd1 _00316_ sky130_fd_sc_hd__a221o_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09777_ _03701_ vssd1 vssd1 vccd1 vccd1 _04238_ sky130_fd_sc_hd__buf_4
X_06989_ genblk1\[7\].osc.clkdiv_C.cnt\[1\] genblk1\[7\].osc.clkdiv_C.cnt\[0\] vssd1
+ vssd1 vccd1 vccd1 _01824_ sky130_fd_sc_hd__xnor2_1
X_08728_ genblk2\[2\].wave_shpr.div.fin_quo\[4\] _03113_ _03117_ _02224_ vssd1 vssd1
+ vccd1 vccd1 _03435_ sky130_fd_sc_hd__a31o_1
XTAP_2304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08659_ _02939_ _03365_ _02943_ vssd1 vssd1 vccd1 vccd1 _03366_ sky130_fd_sc_hd__o21ai_1
XTAP_2359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11670_ genblk2\[9\].wave_shpr.div.acc\[9\] genblk2\[9\].wave_shpr.div.b1\[9\] vssd1
+ vssd1 vccd1 vccd1 _05562_ sky130_fd_sc_hd__or2b_1
XTAP_1669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10621_ genblk2\[6\].wave_shpr.div.b1\[4\] _04836_ _04834_ vssd1 vssd1 vccd1 vccd1
+ _04837_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13340_ clknet_leaf_7_clk _00661_ net49 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.acc\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10552_ genblk2\[5\].wave_shpr.div.acc\[2\] genblk2\[5\].wave_shpr.div.b1\[2\] vssd1
+ vssd1 vccd1 vccd1 _04780_ sky130_fd_sc_hd__or2b_1
XFILLER_0_91_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13271_ clknet_leaf_137_clk _00594_ net41 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.acc\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10483_ genblk2\[4\].wave_shpr.div.acc\[14\] _04727_ _04704_ vssd1 vssd1 vccd1 vccd1
+ _04728_ sky130_fd_sc_hd__mux2_1
XFILLER_0_134_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12222_ _05933_ _05958_ _05959_ vssd1 vssd1 vccd1 vccd1 _05960_ sky130_fd_sc_hd__a21o_1
XFILLER_0_106_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12153_ genblk2\[10\].wave_shpr.div.acc\[19\] _05900_ vssd1 vssd1 vccd1 vccd1 _05903_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11104_ genblk2\[7\].wave_shpr.div.acc\[17\] genblk2\[7\].wave_shpr.div.b1\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05164_ sky130_fd_sc_hd__or2b_1
X_12084_ _05815_ vssd1 vssd1 vccd1 vccd1 _05850_ sky130_fd_sc_hd__clkbuf_4
X_11035_ net900 _05086_ _05093_ _05115_ vssd1 vssd1 vccd1 vccd1 _00664_ sky130_fd_sc_hd__a22o_1
XANTENNA__08001__B1 _01675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08552__A1 genblk2\[6\].wave_shpr.div.fin_quo\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_12986_ clknet_leaf_13_clk _00315_ net69 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.quo\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12100__A2 _05844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11937_ _03821_ genblk2\[10\].wave_shpr.div.acc\[6\] _05758_ vssd1 vssd1 vccd1 vccd1
+ _05759_ sky130_fd_sc_hd__a21o_1
XFILLER_0_86_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10662__A2 _04853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11868_ net669 _05684_ _05685_ _05703_ vssd1 vssd1 vccd1 vccd1 _00909_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10819_ genblk2\[5\].wave_shpr.div.busy _04962_ net855 vssd1 vssd1 vccd1 vccd1 _04964_
+ sky130_fd_sc_hd__a21oi_1
X_13607_ clknet_leaf_68_clk _00920_ net194 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.i\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11799_ genblk2\[9\].wave_shpr.div.acc\[1\] _05650_ _05613_ vssd1 vssd1 vccd1 vccd1
+ _05651_ sky130_fd_sc_hd__mux2_1
XFILLER_0_144_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13538_ clknet_leaf_100_clk _00853_ net165 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.fin_quo\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_40_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13469_ clknet_leaf_85_clk _00786_ net204 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.b1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_445 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07043__A1 genblk1\[8\].osc.clkdiv_C.cnt\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10192__A _04455_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07043__B2 genblk1\[8\].osc.clkdiv_C.cnt\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07961_ genblk1\[7\].osc.clkdiv_C.cnt\[14\] _01360_ vssd1 vssd1 vccd1 vccd1 _02668_
+ sky130_fd_sc_hd__or2_1
X_09700_ _04170_ _04178_ _04179_ vssd1 vssd1 vccd1 vccd1 _04180_ sky130_fd_sc_hd__a21o_1
X_06912_ genblk1\[6\].osc.clkdiv_C.cnt\[1\] net837 genblk1\[6\].osc.clkdiv_C.cnt\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01764_ sky130_fd_sc_hd__a21oi_1
X_07892_ _02529_ _02594_ _02518_ _02598_ vssd1 vssd1 vccd1 vccd1 _02599_ sky130_fd_sc_hd__and4_1
XANTENNA__09192__S _03822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08543__A1 _02225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09631_ net973 _04109_ _04113_ _04125_ vssd1 vssd1 vccd1 vccd1 _00250_ sky130_fd_sc_hd__a22o_1
XFILLER_0_4_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06843_ net1072 _01705_ _01707_ vssd1 vssd1 vccd1 vccd1 genblk1\[5\].osc.clkdiv_C.next_cnt\[7\]
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__07932__C genblk2\[8\].wave_shpr.div.fin_quo\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09562_ genblk2\[1\].wave_shpr.div.b1\[0\] _04011_ net752 vssd1 vssd1 vccd1 vccd1
+ _04073_ sky130_fd_sc_hd__a21o_1
X_06774_ _01649_ vssd1 vssd1 vccd1 vccd1 genblk1\[4\].osc.clkdiv_C.next_cnt\[14\]
+ sky130_fd_sc_hd__clkbuf_1
X_08513_ _03210_ _03214_ vssd1 vssd1 vccd1 vccd1 _03220_ sky130_fd_sc_hd__or2b_1
XFILLER_0_77_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09493_ net1277 _04036_ _04024_ vssd1 vssd1 vccd1 vccd1 _04037_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08444_ _03145_ _03149_ vssd1 vssd1 vccd1 vccd1 _03151_ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08059__B1 net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08375_ _02600_ _03080_ net24 _02520_ vssd1 vssd1 vccd1 vccd1 _03082_ sky130_fd_sc_hd__a211o_1
XANTENNA__10367__A _02152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07326_ _02074_ _02084_ _02088_ _02089_ vssd1 vssd1 vccd1 vccd1 _02090_ sky130_fd_sc_hd__nand4_1
XFILLER_0_34_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07257_ _02027_ _02034_ _02035_ vssd1 vssd1 vccd1 vccd1 genblk1\[10\].osc.clkdiv_C.next_cnt\[3\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_116_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06208_ freq_div.state\[1\] freq_div.state\[2\] freq_div.state\[0\] vssd1 vssd1 vccd1
+ vccd1 _01170_ sky130_fd_sc_hd__or3b_1
XFILLER_0_131_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07188_ genblk1\[9\].osc.clkdiv_C.cnt\[10\] _01974_ genblk1\[9\].osc.clkdiv_C.cnt\[11\]
+ vssd1 vssd1 vccd1 vccd1 _01977_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06139_ _01107_ _01110_ vssd1 vssd1 vccd1 vccd1 _01111_ sky130_fd_sc_hd__xor2_1
XFILLER_0_112_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07585__A2 _01311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09829_ _04069_ genblk1\[2\].osc.clkdiv_C.cnt\[9\] vssd1 vssd1 vccd1 vccd1 _04265_
+ sky130_fd_sc_hd__and2_1
X_12840_ clknet_leaf_65_clk net1306 net197 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.acc\[24\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_2101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12771_ clknet_leaf_93_clk _00104_ net148 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.fin_quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11722_ genblk2\[9\].wave_shpr.div.fin_quo\[0\] _05613_ _00023_ vssd1 vssd1 vccd1
+ vccd1 _05614_ sky130_fd_sc_hd__mux2_1
XFILLER_0_56_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11653_ genblk2\[8\].wave_shpr.div.i\[1\] genblk2\[8\].wave_shpr.div.i\[0\] genblk2\[8\].wave_shpr.div.i\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05548_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout60 net63 vssd1 vssd1 vccd1 vccd1 net60 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_126_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout71 net72 vssd1 vssd1 vccd1 vccd1 net71 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_153_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10604_ genblk2\[5\].wave_shpr.div.fin_quo\[5\] net1330 _00015_ vssd1 vssd1 vccd1
+ vccd1 _04827_ sky130_fd_sc_hd__mux2_1
XANTENNA__09798__B1 _04214_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout82 net83 vssd1 vssd1 vccd1 vccd1 net82 sky130_fd_sc_hd__clkbuf_2
X_11584_ _05389_ _05498_ vssd1 vssd1 vccd1 vccd1 _05499_ sky130_fd_sc_hd__xnor2_1
Xfanout93 net94 vssd1 vssd1 vccd1 vccd1 net93 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_92_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_326 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13323_ clknet_leaf_26_clk _00644_ net87 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.quo\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10535_ genblk2\[5\].wave_shpr.div.acc\[17\] genblk2\[5\].wave_shpr.div.b1\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04763_ sky130_fd_sc_hd__or2b_1
XFILLER_0_135_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13254_ clknet_leaf_2_clk _00577_ net43 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.acc\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10466_ net1008 _04683_ _04690_ _04714_ vssd1 vssd1 vccd1 vccd1 _00496_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12205_ genblk2\[11\].wave_shpr.div.b1\[1\] genblk2\[11\].wave_shpr.div.acc\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05943_ sky130_fd_sc_hd__or2b_1
X_13185_ clknet_leaf_112_clk _00510_ net128 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.acc\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10397_ _04477_ genblk1\[4\].osc.clkdiv_C.cnt\[7\] vssd1 vssd1 vccd1 vccd1 _04667_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_103_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12136_ _05776_ _05733_ vssd1 vssd1 vccd1 vccd1 _05890_ sky130_fd_sc_hd__or2b_1
XANTENNA__13081__RESET_B net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12067_ net446 _05812_ _05815_ genblk2\[10\].wave_shpr.div.quo\[23\] _05838_ vssd1
+ vssd1 vccd1 vccd1 _00973_ sky130_fd_sc_hd__a221o_1
X_11018_ net826 _05086_ _05093_ _05102_ vssd1 vssd1 vccd1 vccd1 _00660_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_138_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_138_clk
+ sky130_fd_sc_hd__clkbuf_16
X_12969_ clknet_leaf_111_clk _00298_ net128 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06490_ genblk1\[2\].osc.clkdiv_C.cnt\[17\] vssd1 vssd1 vccd1 vccd1 _01416_ sky130_fd_sc_hd__inv_2
XTAP_2690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10187__A _04451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06384__B _01327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_602 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08160_ _01489_ genblk1\[3\].osc.clkdiv_C.cnt\[12\] vssd1 vssd1 vccd1 vccd1 _02867_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_55_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07111_ genblk1\[8\].osc.clkdiv_C.cnt\[15\] genblk1\[8\].osc.clkdiv_C.cnt\[14\] _01910_
+ vssd1 vssd1 vccd1 vccd1 _01914_ sky130_fd_sc_hd__and3_1
XFILLER_0_132_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08091_ _02797_ vssd1 vssd1 vccd1 vccd1 _02798_ sky130_fd_sc_hd__buf_2
XFILLER_0_141_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10915__A _03707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07042_ genblk1\[8\].osc.clkdiv_C.cnt\[1\] _01436_ _01855_ _01859_ genblk1\[8\].osc.clkdiv_C.cnt\[10\]
+ vssd1 vssd1 vccd1 vccd1 _01860_ sky130_fd_sc_hd__a32o_1
XFILLER_0_141_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11899__A1 _03839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_1_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08993_ _03572_ _03675_ vssd1 vssd1 vccd1 vccd1 _03676_ sky130_fd_sc_hd__nor2_1
XFILLER_0_76_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07944_ genblk1\[7\].osc.clkdiv_C.cnt\[8\] _01920_ _01514_ genblk1\[7\].osc.clkdiv_C.cnt\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02651_ sky130_fd_sc_hd__o22a_1
XANTENNA__07319__A2 _01242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07875_ _02575_ _02580_ _02581_ vssd1 vssd1 vccd1 vccd1 _02582_ sky130_fd_sc_hd__a21o_1
XANTENNA__11520__B1 _05449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09614_ net865 _04109_ _04080_ _04112_ vssd1 vssd1 vccd1 vccd1 _00246_ sky130_fd_sc_hd__a22o_1
X_06826_ _01694_ _01695_ _01696_ vssd1 vssd1 vccd1 vccd1 _01697_ sky130_fd_sc_hd__and3_1
X_09545_ net417 _04052_ _04053_ net426 _04063_ vssd1 vssd1 vccd1 vccd1 _00226_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_129_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_129_clk
+ sky130_fd_sc_hd__clkbuf_16
X_06757_ genblk1\[4\].osc.clkdiv_C.cnt\[10\] genblk1\[4\].osc.clkdiv_C.cnt\[9\] _01627_
+ genblk1\[4\].osc.clkdiv_C.cnt\[11\] vssd1 vssd1 vccd1 vccd1 _01636_ sky130_fd_sc_hd__a31o_1
XFILLER_0_116_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09476_ _04026_ vssd1 vssd1 vccd1 vccd1 _00194_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__06575__A _01196_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06688_ _01577_ vssd1 vssd1 vccd1 vccd1 _01578_ sky130_fd_sc_hd__buf_4
XFILLER_0_136_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08427_ _03010_ _03129_ _03133_ vssd1 vssd1 vccd1 vccd1 _03134_ sky130_fd_sc_hd__nor3_1
XFILLER_0_136_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10097__A _04269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08358_ _02846_ _03064_ vssd1 vssd1 vccd1 vccd1 _03065_ sky130_fd_sc_hd__and2_1
XFILLER_0_73_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07309_ genblk1\[11\].osc.clkdiv_C.cnt\[7\] _01430_ vssd1 vssd1 vccd1 vccd1 _02073_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_132_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_668 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08289_ _02993_ _02994_ _02995_ vssd1 vssd1 vccd1 vccd1 _02996_ sky130_fd_sc_hd__and3_1
XFILLER_0_150_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10320_ genblk2\[4\].wave_shpr.div.fin_quo\[4\] net1333 _00013_ vssd1 vssd1 vccd1
+ vccd1 _04628_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12000__A1 _03706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10251_ net333 _04563_ _03855_ vssd1 vssd1 vccd1 vccd1 _04564_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_104_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08014__B _01367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10182_ net791 _04486_ _04490_ _04514_ vssd1 vssd1 vccd1 vccd1 _00412_ sky130_fd_sc_hd__a22o_1
XANTENNA__12303__A2 _06009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06518__B1 _01439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07572__C _01437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11511__B1 _05449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11484__A1_N _03727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09180__A1 _01356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12823_ clknet_leaf_62_clk _00156_ net189 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.acc\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12474__RESET_B net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10078__B1 _03736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06485__A _01241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12754_ clknet_leaf_51_clk genblk1\[11\].osc.clkdiv_C.next_cnt\[13\] net110 vssd1
+ vssd1 vccd1 vccd1 genblk1\[11\].osc.clkdiv_C.cnt\[13\] sky130_fd_sc_hd__dfrtp_2
XTAP_1252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11705_ _05559_ _05595_ _05596_ vssd1 vssd1 vccd1 vccd1 _05597_ sky130_fd_sc_hd__a21o_1
X_12685_ clknet_leaf_119_clk genblk1\[7\].osc.clkdiv_C.next_cnt\[16\] net141 vssd1
+ vssd1 vccd1 vccd1 genblk1\[7\].osc.clkdiv_C.cnt\[16\] sky130_fd_sc_hd__dfrtp_2
XTAP_1285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11290__A2 _05279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_112_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11636_ _05449_ _05536_ _05537_ _05448_ net456 vssd1 vssd1 vccd1 vccd1 _00843_ sky130_fd_sc_hd__a32o_1
XFILLER_0_142_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_624 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11567_ _05485_ _05381_ vssd1 vssd1 vccd1 vccd1 _05486_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10518_ net777 _04657_ _04655_ _04752_ vssd1 vssd1 vccd1 vccd1 _00510_ sky130_fd_sc_hd__a22o_1
X_13306_ clknet_leaf_3_clk _00627_ net51 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.quo\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold709 genblk2\[5\].wave_shpr.div.acc\[8\] vssd1 vssd1 vccd1 vccd1 net927 sky130_fd_sc_hd__dlygate4sd3_1
X_11498_ genblk2\[8\].wave_shpr.div.quo\[1\] _05442_ _05446_ net743 vssd1 vssd1 vccd1
+ vccd1 _00796_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13237_ clknet_leaf_10_clk _00560_ net57 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.quo\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13262__RESET_B net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10449_ net971 _04683_ _04690_ _04701_ vssd1 vssd1 vccd1 vccd1 _00492_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09735__S _00009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13168_ clknet_leaf_127_clk _00493_ net66 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.acc\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11750__B1 _05624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06889__A2_N _01519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12119_ _05768_ _05737_ vssd1 vssd1 vccd1 vccd1 _05877_ sky130_fd_sc_hd__or2b_1
XANTENNA_clkbuf_leaf_41_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13099_ clknet_leaf_137_clk _00426_ net42 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.acc\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09036__A _03702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06509__B1 _01326_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11502__B1 _05446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07660_ _02359_ _02360_ _02363_ _02366_ vssd1 vssd1 vccd1 vccd1 _02367_ sky130_fd_sc_hd__a31o_1
XANTENNA_clkbuf_leaf_56_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06611_ _01186_ _01354_ _01171_ vssd1 vssd1 vccd1 vccd1 _01519_ sky130_fd_sc_hd__o21a_2
XANTENNA__07721__A2 _02425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07591_ _01928_ _01801_ vssd1 vssd1 vccd1 vccd1 _02298_ sky130_fd_sc_hd__nor2_1
XANTENNA__08594__B _02364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09330_ _03791_ _03749_ vssd1 vssd1 vccd1 vccd1 _03911_ sky130_fd_sc_hd__or2b_1
X_06542_ genblk1\[2\].osc.clkdiv_C.cnt\[6\] _01459_ vssd1 vssd1 vccd1 vccd1 _01462_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09261_ _03853_ genblk1\[0\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 _03860_
+ sky130_fd_sc_hd__and2_1
X_06473_ genblk1\[1\].osc.clkdiv_C.cnt\[14\] _01401_ vssd1 vssd1 vccd1 vccd1 _01403_
+ sky130_fd_sc_hd__and2_1
XANTENNA__08682__B1 _02224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08212_ _02697_ _02698_ _02746_ vssd1 vssd1 vccd1 vccd1 _02919_ sky130_fd_sc_hd__a21o_1
XFILLER_0_117_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09192_ net1244 _02002_ _03822_ vssd1 vssd1 vccd1 vccd1 _03824_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09226__A2 _03836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_114_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08143_ genblk2\[3\].wave_shpr.div.fin_quo\[6\] vssd1 vssd1 vccd1 vccd1 _02850_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07237__A1 _01242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08434__B1 _02221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07237__B2 _01197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08074_ _02763_ _02765_ _02769_ _02778_ _02780_ vssd1 vssd1 vccd1 vccd1 _02781_ sky130_fd_sc_hd__o41a_1
XFILLER_0_113_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07025_ _01822_ _01845_ _01846_ vssd1 vssd1 vccd1 vccd1 genblk1\[7\].osc.clkdiv_C.next_cnt\[14\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_12_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_129_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_101_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_87_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10380__A _04651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold14 _00731_ vssd1 vssd1 vccd1 vccd1 net232 sky130_fd_sc_hd__dlygate4sd3_1
X_08976_ _03656_ _03523_ _03521_ vssd1 vssd1 vccd1 vccd1 _03662_ sky130_fd_sc_hd__o21a_1
Xhold25 genblk2\[9\].wave_shpr.div.quo\[12\] vssd1 vssd1 vccd1 vccd1 net243 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 _00549_ vssd1 vssd1 vccd1 vccd1 net254 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07960__A2 _01514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold47 genblk2\[0\].wave_shpr.div.quo\[21\] vssd1 vssd1 vccd1 vccd1 net265 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 _00299_ vssd1 vssd1 vccd1 vccd1 net276 sky130_fd_sc_hd__dlygate4sd3_1
X_07927_ _01200_ genblk1\[8\].osc.clkdiv_C.cnt\[14\] _01362_ genblk1\[8\].osc.clkdiv_C.cnt\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02634_ sky130_fd_sc_hd__a211o_1
Xhold69 PWM.next_pwm_out vssd1 vssd1 vccd1 vccd1 net287 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06289__B _01250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07858_ _02216_ _02552_ genblk2\[0\].wave_shpr.div.fin_quo\[2\] vssd1 vssd1 vccd1
+ vccd1 _02565_ sky130_fd_sc_hd__and3_1
X_06809_ _01676_ _01677_ _01679_ _01680_ vssd1 vssd1 vccd1 vccd1 _01681_ sky130_fd_sc_hd__or4b_1
X_07789_ genblk1\[0\].osc.clkdiv_C.cnt\[11\] _01263_ vssd1 vssd1 vccd1 vccd1 _02496_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_78_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09528_ _03853_ genblk1\[1\].osc.clkdiv_C.cnt\[3\] vssd1 vssd1 vccd1 vccd1 _04054_
+ sky130_fd_sc_hd__and2_1
XPHY_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09459_ _04017_ vssd1 vssd1 vccd1 vccd1 _00186_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12470_ clknet_leaf_33_clk smpl_rt_clkdiv.clkDiv_inst.next_cnt\[4\] net100 vssd1
+ vssd1 vccd1 vccd1 smpl_rt_clkdiv.clkDiv_inst.cnt\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13773__RESET_B net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11421_ _05364_ _05395_ _05396_ vssd1 vssd1 vccd1 vccd1 _05397_ sky130_fd_sc_hd__a21o_1
XANTENNA__10232__B1 _04457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11352_ net679 _05311_ _05315_ _05338_ vssd1 vssd1 vccd1 vccd1 _00758_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10303_ _04566_ _04613_ _04614_ vssd1 vssd1 vccd1 vccd1 _04615_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_120_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_132_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11283_ net877 _05279_ _05283_ _05286_ vssd1 vssd1 vccd1 vccd1 _00741_ sky130_fd_sc_hd__a22o_1
XFILLER_0_104_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_hold967_A genblk1\[8\].osc.clkdiv_C.cnt\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13022_ clknet_leaf_128_clk _00349_ net67 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.fin_quo\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_10234_ genblk2\[3\].wave_shpr.div.acc\[24\] _04480_ _04549_ vssd1 vssd1 vccd1 vccd1
+ _04553_ sky130_fd_sc_hd__or3b_1
X_10165_ net890 _04486_ _04490_ _04501_ vssd1 vssd1 vccd1 vccd1 _00408_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07951__A2 _01556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10096_ _04451_ vssd1 vssd1 vccd1 vccd1 _04457_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12806_ clknet_leaf_59_clk _00139_ net187 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.quo\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10998_ genblk2\[6\].wave_shpr.div.b1\[2\] genblk2\[6\].wave_shpr.div.acc\[2\] vssd1
+ vssd1 vccd1 vccd1 _05087_ sky130_fd_sc_hd__xor2_1
XFILLER_0_128_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11263__A2 _05245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12737_ clknet_leaf_37_clk genblk1\[10\].osc.clkdiv_C.next_cnt\[14\] net114 vssd1
+ vssd1 vccd1 vccd1 genblk1\[10\].osc.clkdiv_C.cnt\[14\] sky130_fd_sc_hd__dfrtp_2
XTAP_1082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12668_ clknet_leaf_24_clk genblk1\[6\].osc.clkdiv_C.next_cnt\[17\] net92 vssd1 vssd1
+ vccd1 vccd1 genblk1\[6\].osc.clkdiv_C.cnt\[17\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11619_ net991 _05507_ _05445_ _05525_ vssd1 vssd1 vccd1 vccd1 _00838_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12599_ clknet_leaf_21_clk genblk1\[3\].osc.clkdiv_C.next_cnt\[2\] net97 vssd1 vssd1
+ vccd1 vccd1 genblk1\[3\].osc.clkdiv_C.cnt\[2\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_106_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold506 genblk2\[10\].wave_shpr.div.quo\[2\] vssd1 vssd1 vccd1 vccd1 net724 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold517 _00514_ vssd1 vssd1 vccd1 vccd1 net735 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11995__S _05802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold528 genblk2\[9\].wave_shpr.div.quo\[0\] vssd1 vssd1 vccd1 vccd1 net746 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold539 genblk2\[1\].wave_shpr.div.i\[2\] vssd1 vssd1 vccd1 vccd1 net757 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07927__C1 genblk1\[8\].osc.clkdiv_C.cnt\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08830_ _03482_ _03530_ _03529_ vssd1 vssd1 vccd1 vccd1 _03537_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_148_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_877 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07942__A2 _01311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_888 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08761_ net10 _02744_ _03467_ vssd1 vssd1 vccd1 vccd1 _03468_ sky130_fd_sc_hd__and3_1
XTAP_899 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07712_ _02418_ vssd1 vssd1 vccd1 vccd1 _02419_ sky130_fd_sc_hd__buf_2
X_08692_ _03187_ _03194_ vssd1 vssd1 vccd1 vccd1 _03399_ sky130_fd_sc_hd__xnor2_1
X_07643_ genblk1\[11\].osc.clkdiv_C.cnt\[16\] genblk1\[11\].osc.clkdiv_C.cnt\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02350_ sky130_fd_sc_hd__nor2_4
XANTENNA_fanout169_A net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07574_ _01336_ _01437_ _01226_ genblk1\[9\].osc.clkdiv_C.cnt\[5\] vssd1 vssd1 vccd1
+ vccd1 _02281_ sky130_fd_sc_hd__o31a_1
X_09313_ _03782_ _03897_ vssd1 vssd1 vccd1 vccd1 _03898_ sky130_fd_sc_hd__xnor2_1
X_06525_ _01450_ vssd1 vssd1 vccd1 vccd1 _01451_ sky130_fd_sc_hd__buf_2
XFILLER_0_8_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_60_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_60_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_118_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09244_ net543 _03845_ _03847_ genblk2\[0\].wave_shpr.div.quo\[14\] _03850_ vssd1
+ vssd1 vccd1 vccd1 _00138_ sky130_fd_sc_hd__a221o_1
XFILLER_0_134_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06456_ genblk1\[1\].osc.clkdiv_C.cnt\[8\] genblk1\[1\].osc.clkdiv_C.cnt\[7\] _01387_
+ vssd1 vssd1 vccd1 vccd1 _01392_ sky130_fd_sc_hd__and3_1
XANTENNA__07949__A _01172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09175_ _03814_ vssd1 vssd1 vccd1 vccd1 _00105_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06681__A2 _01362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06387_ genblk1\[1\].osc.clkdiv_C.cnt\[3\] _01323_ _01329_ _01330_ vssd1 vssd1 vccd1
+ vccd1 _01331_ sky130_fd_sc_hd__a22o_1
X_08126_ genblk1\[4\].osc.clkdiv_C.cnt\[7\] _01340_ _02829_ vssd1 vssd1 vccd1 vccd1
+ _02833_ sky130_fd_sc_hd__a21o_1
XFILLER_0_16_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09080__B1 _03733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08057_ genblk1\[5\].osc.clkdiv_C.cnt\[7\] _01223_ vssd1 vssd1 vccd1 vccd1 _02764_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_98_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07008_ genblk1\[7\].osc.clkdiv_C.cnt\[7\] _01832_ genblk1\[7\].osc.clkdiv_C.cnt\[8\]
+ vssd1 vssd1 vccd1 vccd1 _01836_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11190__A1 _03831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08959_ sig_norm.quo\[4\] _03647_ _02248_ vssd1 vssd1 vccd1 vccd1 _03648_ sky130_fd_sc_hd__mux2_1
X_11970_ genblk2\[10\].wave_shpr.div.fin_quo\[2\] net220 _00003_ vssd1 vssd1 vccd1
+ vccd1 _05790_ sky130_fd_sc_hd__mux2_1
X_10921_ _05045_ vssd1 vssd1 vccd1 vccd1 _00620_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13640_ clknet_leaf_94_clk net683 net160 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.quo\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10852_ genblk2\[6\].wave_shpr.div.b1\[7\] genblk2\[6\].wave_shpr.div.acc\[7\] vssd1
+ vssd1 vccd1 vccd1 _04996_ sky130_fd_sc_hd__and2b_1
XFILLER_0_66_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10783_ _04938_ _04939_ vssd1 vssd1 vccd1 vccd1 _04940_ sky130_fd_sc_hd__nand2_1
XPHY_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13571_ clknet_leaf_56_clk _00886_ net182 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.quo\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_51_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_51_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_26_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08110__A2 _01313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12522_ clknet_leaf_103_clk PWM.next_counter\[6\] net156 vssd1 vssd1 vccd1 vccd1
+ PWM.counter\[6\] sky130_fd_sc_hd__dfrtp_1
XPHY_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12453_ clknet_leaf_42_clk net5 net123 vssd1 vssd1 vccd1 vccd1 modein.delay_octave_up_in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07578__B _01234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11404_ genblk2\[8\].wave_shpr.div.b1\[3\] genblk2\[8\].wave_shpr.div.acc\[3\] vssd1
+ vssd1 vccd1 vccd1 _05380_ sky130_fd_sc_hd__and2b_1
XFILLER_0_105_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_256 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12384_ _05959_ _05933_ vssd1 vssd1 vccd1 vccd1 _06060_ sky130_fd_sc_hd__or2b_1
XFILLER_0_62_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09071__B1 _01302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11335_ _05325_ _05212_ vssd1 vssd1 vccd1 vccd1 _05326_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_120_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11266_ _05219_ _05220_ vssd1 vssd1 vccd1 vccd1 _05273_ sky130_fd_sc_hd__nor2_2
XFILLER_0_120_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09374__A1 _03942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10217_ genblk2\[3\].wave_shpr.div.acc\[19\] _04538_ vssd1 vssd1 vccd1 vccd1 _04541_
+ sky130_fd_sc_hd__or2_1
X_13005_ clknet_leaf_138_clk _00334_ net40 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.acc\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11197_ _01859_ vssd1 vssd1 vccd1 vccd1 _05239_ sky130_fd_sc_hd__inv_2
XANTENNA__11181__A1 _03819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10148_ net976 _04488_ _04420_ vssd1 vssd1 vccd1 vccd1 _04489_ sky130_fd_sc_hd__mux2_1
XANTENNA__11844__A _03693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10079_ _03833_ net1227 vssd1 vssd1 vccd1 vccd1 _04450_ sky130_fd_sc_hd__and2_1
XFILLER_0_89_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13769_ clknet_leaf_71_clk _01080_ net217 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.acc\[21\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_42_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_42_clk sky130_fd_sc_hd__clkbuf_16
X_06310_ genblk1\[0\].osc.clkdiv_C.cnt\[1\] genblk1\[0\].osc.clkdiv_C.cnt\[0\] vssd1
+ vssd1 vccd1 vccd1 _01271_ sky130_fd_sc_hd__or2_1
X_07290_ _02027_ _02056_ _02057_ vssd1 vssd1 vccd1 vccd1 genblk1\[10\].osc.clkdiv_C.next_cnt\[14\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_57_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06241_ _01201_ genblk1\[0\].osc.clkdiv_C.cnt\[7\] genblk1\[0\].osc.clkdiv_C.cnt\[8\]
+ vssd1 vssd1 vccd1 vccd1 _01203_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_127_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_41_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06172_ _01141_ _01143_ _01119_ _01126_ vssd1 vssd1 vccd1 vccd1 _01144_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_53_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08404__A3 _01362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold303 genblk2\[10\].wave_shpr.div.quo\[13\] vssd1 vssd1 vccd1 vccd1 net521 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold314 _00476_ vssd1 vssd1 vccd1 vccd1 net532 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold325 genblk2\[0\].wave_shpr.div.quo\[15\] vssd1 vssd1 vccd1 vccd1 net543 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold336 _00303_ vssd1 vssd1 vccd1 vccd1 net554 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold347 genblk2\[9\].wave_shpr.div.quo\[23\] vssd1 vssd1 vccd1 vccd1 net565 sky130_fd_sc_hd__dlygate4sd3_1
Xhold358 genblk2\[11\].wave_shpr.div.acc\[18\] vssd1 vssd1 vccd1 vccd1 net576 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09931_ _04210_ net22 vssd1 vssd1 vccd1 vccd1 _04339_ sky130_fd_sc_hd__nor2_1
Xhold369 _00870_ vssd1 vssd1 vccd1 vccd1 net587 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09862_ _04179_ _04170_ vssd1 vssd1 vccd1 vccd1 _04286_ sky130_fd_sc_hd__or2b_1
XANTENNA__06690__A2_N _01209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08813_ _03511_ _03515_ _03513_ _03514_ vssd1 vssd1 vccd1 vccd1 _03520_ sky130_fd_sc_hd__o211ai_2
Xhold1003 _01059_ vssd1 vssd1 vccd1 vccd1 net1221 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09969__B_N genblk2\[3\].wave_shpr.div.b1\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1014 genblk2\[4\].wave_shpr.div.b1\[10\] vssd1 vssd1 vccd1 vccd1 net1232 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09793_ _02164_ vssd1 vssd1 vccd1 vccd1 _04247_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1025 genblk2\[0\].wave_shpr.div.b1\[1\] vssd1 vssd1 vccd1 vccd1 net1243 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1036 genblk2\[10\].wave_shpr.div.b1\[7\] vssd1 vssd1 vccd1 vccd1 net1254 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1047 genblk2\[11\].wave_shpr.div.b1\[3\] vssd1 vssd1 vccd1 vccd1 net1265 sky130_fd_sc_hd__dlygate4sd3_1
X_08744_ _03422_ _03427_ _03449_ _03450_ vssd1 vssd1 vccd1 vccd1 _03451_ sky130_fd_sc_hd__a211oi_2
Xhold1058 genblk2\[0\].wave_shpr.div.b1\[9\] vssd1 vssd1 vccd1 vccd1 net1276 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1069 genblk2\[5\].wave_shpr.div.b1\[4\] vssd1 vssd1 vccd1 vccd1 net1287 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08675_ _03359_ _03380_ _03379_ vssd1 vssd1 vccd1 vccd1 _03382_ sky130_fd_sc_hd__o21a_1
XTAP_1807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07626_ _02081_ _01241_ _02331_ _02332_ vssd1 vssd1 vccd1 vccd1 _02333_ sky130_fd_sc_hd__a211o_1
XTAP_1829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06351__A1 genblk1\[0\].osc.clkdiv_C.cnt\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07557_ genblk2\[9\].wave_shpr.div.fin_quo\[3\] _02263_ vssd1 vssd1 vccd1 vccd1 _02264_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_119_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_33_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_33_clk sky130_fd_sc_hd__clkbuf_16
X_06508_ _01201_ _01410_ _01432_ _01412_ genblk1\[2\].osc.clkdiv_C.cnt\[7\] vssd1
+ vssd1 vccd1 vccd1 _01434_ sky130_fd_sc_hd__a221o_1
XFILLER_0_63_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07679__A _01489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07488_ genblk2\[11\].wave_shpr.div.busy _02211_ vssd1 vssd1 vccd1 vccd1 _02212_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_64_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09840__A2 _04247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06439_ genblk1\[1\].osc.clkdiv_C.cnt\[3\] _01378_ vssd1 vssd1 vccd1 vccd1 _01380_
+ sky130_fd_sc_hd__and2_1
X_09227_ net277 _03836_ _03840_ net379 vssd1 vssd1 vccd1 vccd1 _00131_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09158_ _03805_ vssd1 vssd1 vccd1 vccd1 _00097_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08109_ genblk1\[4\].osc.clkdiv_C.cnt\[9\] _01323_ _02811_ _02815_ vssd1 vssd1 vccd1
+ vccd1 _02816_ sky130_fd_sc_hd__a211o_1
XANTENNA__06406__A2 genblk1\[1\].osc.clkdiv_C.cnt\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09089_ _03737_ modein.delay_octave_down_in\[1\] _01197_ _03738_ vssd1 vssd1 vccd1
+ vccd1 _03740_ sky130_fd_sc_hd__or4_1
X_11120_ genblk2\[7\].wave_shpr.div.acc\[3\] genblk2\[7\].wave_shpr.div.b1\[3\] vssd1
+ vssd1 vccd1 vccd1 _05180_ sky130_fd_sc_hd__or2b_1
Xhold870 sig_norm.b1\[3\] vssd1 vssd1 vccd1 vccd1 net1088 sky130_fd_sc_hd__dlygate4sd3_1
Xhold881 genblk2\[3\].wave_shpr.div.b1\[5\] vssd1 vssd1 vccd1 vccd1 net1099 sky130_fd_sc_hd__dlygate4sd3_1
Xhold892 genblk2\[2\].wave_shpr.div.i\[1\] vssd1 vssd1 vccd1 vccd1 net1110 sky130_fd_sc_hd__dlygate4sd3_1
X_11051_ _05009_ _05127_ vssd1 vssd1 vccd1 vccd1 _05128_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11163__A1 _05222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10002_ _04369_ _04396_ _04397_ vssd1 vssd1 vccd1 vccd1 _04398_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11953_ _05734_ _05773_ _05774_ vssd1 vssd1 vccd1 vccd1 _05775_ sky130_fd_sc_hd__a21o_1
XFILLER_0_86_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10904_ net1200 _01799_ _04848_ vssd1 vssd1 vccd1 vccd1 _05036_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11884_ net892 _03696_ _03694_ _05714_ vssd1 vssd1 vccd1 vccd1 _00914_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13623_ clknet_leaf_85_clk _00936_ net204 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.b1\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11218__A2 _05246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10835_ genblk2\[6\].wave_shpr.div.acc\[4\] genblk2\[6\].wave_shpr.div.b1\[4\] vssd1
+ vssd1 vccd1 vccd1 _04979_ sky130_fd_sc_hd__or2b_1
XFILLER_0_104_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_24_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_24_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_109_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13554_ clknet_leaf_100_clk _00869_ net164 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.quo\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12451__CLK clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10766_ _04807_ _04926_ vssd1 vssd1 vccd1 vccd1 _04927_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12505_ clknet_leaf_104_clk _00067_ net154 vssd1 vssd1 vccd1 vccd1 PWM.final_in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13485_ clknet_leaf_97_clk _00802_ net167 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10697_ _04869_ genblk1\[5\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 _04876_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_89_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_120_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12436_ net619 _06072_ _06073_ _06098_ vssd1 vssd1 vccd1 vccd1 _01082_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12367_ _05951_ _05937_ vssd1 vssd1 vccd1 vccd1 _06047_ sky130_fd_sc_hd__or2b_1
XFILLER_0_22_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11318_ _05204_ _05312_ vssd1 vssd1 vccd1 vccd1 _05313_ sky130_fd_sc_hd__xnor2_1
X_12298_ _03941_ vssd1 vssd1 vccd1 vccd1 _06010_ sky130_fd_sc_hd__buf_4
X_11249_ net400 _05255_ _05256_ net585 _05264_ vssd1 vssd1 vccd1 vccd1 _00729_ sky130_fd_sc_hd__a221o_1
XFILLER_0_129_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09743__S _00009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06790_ genblk1\[5\].osc.clkdiv_C.cnt\[5\] net36 vssd1 vssd1 vccd1 vccd1 _01662_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08460_ _03165_ _03166_ vssd1 vssd1 vccd1 vccd1 _03167_ sky130_fd_sc_hd__nor2_1
XFILLER_0_148_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_77_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07411_ genblk2\[0\].wave_shpr.div.start vssd1 vssd1 vccd1 vccd1 _02155_ sky130_fd_sc_hd__buf_8
XFILLER_0_148_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08391_ _01412_ _01302_ vssd1 vssd1 vccd1 vccd1 _03098_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_15_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_15_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_18_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07499__A net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07342_ genblk1\[11\].osc.clkdiv_C.cnt\[3\] _02097_ vssd1 vssd1 vccd1 vccd1 _02103_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_57_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11090__A0 _05054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07273_ genblk1\[10\].osc.clkdiv_C.cnt\[7\] _02041_ net1183 vssd1 vssd1 vccd1 vccd1
+ _02047_ sky130_fd_sc_hd__a21oi_1
X_09012_ genblk2\[9\].wave_shpr.div.i\[0\] _02202_ vssd1 vssd1 vccd1 vccd1 _03686_
+ sky130_fd_sc_hd__nand2_1
X_06224_ _01179_ vssd1 vssd1 vccd1 vccd1 _01186_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_131_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold100 _00718_ vssd1 vssd1 vccd1 vccd1 net318 sky130_fd_sc_hd__dlygate4sd3_1
X_06155_ _01124_ _01125_ vssd1 vssd1 vccd1 vccd1 _01127_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_226 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold111 genblk2\[8\].wave_shpr.div.quo\[9\] vssd1 vssd1 vccd1 vccd1 net329 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout201_A net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold122 genblk2\[1\].wave_shpr.div.quo\[22\] vssd1 vssd1 vccd1 vccd1 net340 sky130_fd_sc_hd__dlygate4sd3_1
Xhold133 genblk2\[11\].wave_shpr.div.quo\[15\] vssd1 vssd1 vccd1 vccd1 net351 sky130_fd_sc_hd__dlygate4sd3_1
Xhold144 genblk2\[9\].wave_shpr.div.quo\[19\] vssd1 vssd1 vccd1 vccd1 net362 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09219__A _03838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold155 genblk2\[10\].wave_shpr.div.quo\[14\] vssd1 vssd1 vccd1 vccd1 net373 sky130_fd_sc_hd__dlygate4sd3_1
Xhold166 genblk2\[11\].wave_shpr.div.b1\[14\] vssd1 vssd1 vccd1 vccd1 net384 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold177 smpl_rt_clkdiv.clkDiv_inst.cnt\[7\] vssd1 vssd1 vccd1 vccd1 net395 sky130_fd_sc_hd__dlygate4sd3_1
Xhold188 genblk2\[1\].wave_shpr.div.b1\[15\] vssd1 vssd1 vccd1 vccd1 net406 sky130_fd_sc_hd__dlygate4sd3_1
X_09914_ _04203_ _04158_ vssd1 vssd1 vccd1 vccd1 _04326_ sky130_fd_sc_hd__or2b_1
Xhold199 genblk2\[1\].wave_shpr.div.quo\[19\] vssd1 vssd1 vccd1 vccd1 net417 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09845_ _04269_ genblk1\[2\].osc.clkdiv_C.cnt\[16\] vssd1 vssd1 vccd1 vccd1 _04274_
+ sky130_fd_sc_hd__and2_1
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09776_ _04237_ vssd1 vssd1 vccd1 vccd1 _00283_ sky130_fd_sc_hd__clkbuf_1
X_06988_ net1058 _01823_ vssd1 vssd1 vccd1 vccd1 genblk1\[7\].osc.clkdiv_C.next_cnt\[0\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__07311__A2_N _01211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08727_ _03113_ _03117_ genblk2\[2\].wave_shpr.div.fin_quo\[4\] vssd1 vssd1 vccd1
+ vccd1 _03434_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_69_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13546__RESET_B net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08658_ genblk2\[3\].wave_shpr.div.fin_quo\[3\] _02467_ _03364_ _02592_ vssd1 vssd1
+ vccd1 vccd1 _03365_ sky130_fd_sc_hd__a22o_1
XTAP_1615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07609_ _02222_ vssd1 vssd1 vccd1 vccd1 _02316_ sky130_fd_sc_hd__clkbuf_4
XTAP_1648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08589_ _03275_ _03276_ _03295_ vssd1 vssd1 vccd1 vccd1 _03296_ sky130_fd_sc_hd__and3_1
XFILLER_0_92_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10620_ _01730_ vssd1 vssd1 vccd1 vccd1 _04836_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10551_ genblk2\[5\].wave_shpr.div.acc\[3\] genblk2\[5\].wave_shpr.div.b1\[3\] vssd1
+ vssd1 vccd1 vccd1 _04779_ sky130_fd_sc_hd__or2b_1
XFILLER_0_52_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13270_ clknet_leaf_1_clk _00593_ net43 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.acc\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10482_ _04609_ _04726_ vssd1 vssd1 vccd1 vccd1 _04727_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12221_ genblk2\[11\].wave_shpr.div.b1\[9\] genblk2\[11\].wave_shpr.div.acc\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05959_ sky130_fd_sc_hd__and2b_1
XANTENNA__11659__A _03690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12152_ net1135 _05876_ _05883_ _05902_ vssd1 vssd1 vccd1 vccd1 _00994_ sky130_fd_sc_hd__a22o_1
X_11103_ net280 _05162_ _05163_ vssd1 vssd1 vccd1 vccd1 _00684_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_102_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12083_ net969 _05844_ _05817_ _05849_ vssd1 vssd1 vccd1 vccd1 _00978_ sky130_fd_sc_hd__a22o_1
XFILLER_0_102_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11034_ genblk2\[6\].wave_shpr.div.acc\[10\] _05114_ _05105_ vssd1 vssd1 vccd1 vccd1
+ _05115_ sky130_fd_sc_hd__mux2_1
XANTENNA__07591__B _01801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12985_ clknet_leaf_13_clk _00314_ net69 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.quo\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09501__A1 _03831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09799__A _04250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11936_ _03821_ genblk2\[10\].wave_shpr.div.acc\[6\] _05757_ vssd1 vssd1 vccd1 vccd1
+ _05758_ sky130_fd_sc_hd__o21a_1
XANTENNA__08907__S _01157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11867_ genblk2\[9\].wave_shpr.div.acc\[17\] _05702_ _05673_ vssd1 vssd1 vccd1 vccd1
+ _05703_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08068__A1 _01196_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13606_ clknet_leaf_67_clk _00919_ net194 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.i\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10818_ _04855_ _04961_ _04963_ _04858_ net783 vssd1 vssd1 vccd1 vccd1 _00599_ sky130_fd_sc_hd__a32o_1
XANTENNA__09804__A2 _04248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11798_ _05575_ _05649_ vssd1 vssd1 vccd1 vccd1 _05650_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13537_ clknet_leaf_81_clk _00852_ net200 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.i\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10749_ genblk2\[5\].wave_shpr.div.acc\[10\] _04913_ _04907_ vssd1 vssd1 vccd1 vccd1
+ _04914_ sky130_fd_sc_hd__mux2_1
XFILLER_0_54_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13468_ clknet_leaf_75_clk _00785_ net203 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.b1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07766__B _01255_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12419_ genblk2\[11\].wave_shpr.div.acc\[17\] _06086_ _05981_ vssd1 vssd1 vccd1 vccd1
+ _06087_ sky130_fd_sc_hd__mux2_1
X_13399_ clknet_leaf_119_clk net318 net139 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_457 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07043__A2 _01487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09039__A _02147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07960_ genblk1\[7\].osc.clkdiv_C.cnt\[9\] _01514_ _02651_ _02665_ _02666_ vssd1
+ vssd1 vccd1 vccd1 _02667_ sky130_fd_sc_hd__a221o_1
Xclkbuf_leaf_4_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_4_clk sky130_fd_sc_hd__clkbuf_16
X_06911_ genblk1\[6\].osc.clkdiv_C.cnt\[2\] genblk1\[6\].osc.clkdiv_C.cnt\[1\] genblk1\[6\].osc.clkdiv_C.cnt\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01763_ sky130_fd_sc_hd__and3_1
X_07891_ _02509_ _02597_ vssd1 vssd1 vccd1 vccd1 _02598_ sky130_fd_sc_hd__or2_1
X_09630_ genblk2\[1\].wave_shpr.div.acc\[16\] _04124_ _04095_ vssd1 vssd1 vccd1 vccd1
+ _04125_ sky130_fd_sc_hd__mux2_1
X_06842_ genblk1\[5\].osc.clkdiv_C.cnt\[7\] _01705_ _01694_ vssd1 vssd1 vccd1 vccd1
+ _01707_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06398__A _01188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06773_ _01599_ _01646_ _01648_ vssd1 vssd1 vccd1 vccd1 _01649_ sky130_fd_sc_hd__and3_1
X_09561_ genblk2\[1\].wave_shpr.div.b1\[0\] net752 _04011_ vssd1 vssd1 vccd1 vccd1
+ _04072_ sky130_fd_sc_hd__nand3_1
XFILLER_0_78_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08512_ _03204_ _03217_ _03127_ _03218_ vssd1 vssd1 vccd1 vccd1 _03219_ sky130_fd_sc_hd__o211a_1
X_09492_ _01411_ vssd1 vssd1 vccd1 vccd1 _04036_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10102__A2 _04457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08443_ _03145_ _03149_ vssd1 vssd1 vccd1 vccd1 _03150_ sky130_fd_sc_hd__xor2_2
XANTENNA_fanout151_A net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08374_ _02520_ net1354 _03080_ _02600_ vssd1 vssd1 vccd1 vccd1 _03081_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_147_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12939__RESET_B net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07325_ genblk1\[11\].osc.clkdiv_C.cnt\[1\] _01321_ _01925_ genblk1\[11\].osc.clkdiv_C.cnt\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02089_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_129_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09271__A3 _03804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07256_ genblk1\[10\].osc.clkdiv_C.cnt\[3\] _02032_ vssd1 vssd1 vccd1 vccd1 _02035_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06207_ genblk1\[0\].osc.clkdiv_C.cnt\[10\] vssd1 vssd1 vccd1 vccd1 _01169_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10383__A _04058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07187_ genblk1\[9\].osc.clkdiv_C.cnt\[10\] _01974_ _01976_ _01954_ vssd1 vssd1 vccd1
+ vccd1 genblk1\[9\].osc.clkdiv_C.next_cnt\[10\] sky130_fd_sc_hd__o211a_1
XFILLER_0_14_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06138_ _01108_ _01109_ vssd1 vssd1 vccd1 vccd1 _01110_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08534__A2 _02526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09828_ net393 _04257_ _04259_ net573 _04264_ vssd1 vssd1 vccd1 vccd1 _00308_ sky130_fd_sc_hd__a221o_1
X_09759_ _04228_ vssd1 vssd1 vccd1 vccd1 _00275_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_96_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12770_ clknet_leaf_93_clk _00103_ net148 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.fin_quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11721_ _05612_ vssd1 vssd1 vccd1 vccd1 _05613_ sky130_fd_sc_hd__buf_4
XTAP_2179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11652_ _05449_ _05546_ _05547_ _05448_ net1098 vssd1 vssd1 vccd1 vccd1 _00849_ sky130_fd_sc_hd__a32o_1
XANTENNA__08028__A genblk2\[6\].wave_shpr.div.fin_quo\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout50 net85 vssd1 vssd1 vccd1 vccd1 net50 sky130_fd_sc_hd__clkbuf_2
Xfanout61 net62 vssd1 vssd1 vccd1 vccd1 net61 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10603_ _04826_ vssd1 vssd1 vccd1 vccd1 _00521_ sky130_fd_sc_hd__clkbuf_1
Xfanout72 net75 vssd1 vssd1 vccd1 vccd1 net72 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09798__B2 _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout83 net84 vssd1 vssd1 vccd1 vccd1 net83 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_153_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11583_ _05390_ _05367_ vssd1 vssd1 vccd1 vccd1 _05498_ sky130_fd_sc_hd__or2b_1
Xfanout94 net98 vssd1 vssd1 vccd1 vccd1 net94 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13322_ clknet_leaf_26_clk _00643_ net87 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.quo\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10534_ net281 _04761_ _04762_ vssd1 vssd1 vccd1 vccd1 _00516_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_107_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13253_ clknet_leaf_1_clk _00576_ net41 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.acc\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10465_ genblk2\[4\].wave_shpr.div.acc\[10\] _04713_ _04704_ vssd1 vssd1 vccd1 vccd1
+ _04714_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12204_ genblk2\[11\].wave_shpr.div.acc\[0\] genblk2\[11\].wave_shpr.div.b1\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05942_ sky130_fd_sc_hd__and2b_1
XANTENNA__08222__A1 _02789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13184_ clknet_leaf_112_clk _00509_ net129 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.acc\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10396_ genblk2\[4\].wave_shpr.div.quo\[15\] _04661_ _04663_ net596 _04666_ vssd1
+ vssd1 vccd1 vccd1 _00474_ sky130_fd_sc_hd__a221o_1
X_12135_ net944 _05876_ _05883_ _05889_ vssd1 vssd1 vccd1 vccd1 _00990_ sky130_fd_sc_hd__a22o_1
XANTENNA__06784__A1 _01436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09293__S _03804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12306__B1 _06010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12066_ _05835_ genblk1\[10\].osc.clkdiv_C.cnt\[15\] vssd1 vssd1 vccd1 vccd1 _05838_
+ sky130_fd_sc_hd__and2_1
X_11017_ genblk2\[6\].wave_shpr.div.acc\[6\] _05101_ _05023_ vssd1 vssd1 vccd1 vccd1
+ _05102_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12968_ clknet_leaf_111_clk _00297_ net130 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_0_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11919_ genblk2\[10\].wave_shpr.div.acc\[7\] genblk2\[10\].wave_shpr.div.b1\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05741_ sky130_fd_sc_hd__or2b_1
XTAP_2680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12899_ clknet_leaf_30_clk net341 net102 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.quo\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07110_ genblk1\[8\].osc.clkdiv_C.cnt\[14\] _01910_ _01913_ vssd1 vssd1 vccd1 vccd1
+ genblk1\[8\].osc.clkdiv_C.next_cnt\[14\] sky130_fd_sc_hd__o21a_1
XFILLER_0_55_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08090_ net11 _02364_ _02365_ vssd1 vssd1 vccd1 vccd1 _02797_ sky130_fd_sc_hd__and3_1
XANTENNA__07777__A genblk1\[0\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07041_ _01439_ _01576_ vssd1 vssd1 vccd1 vccd1 _01859_ sky130_fd_sc_hd__nand2_2
XFILLER_0_2_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_152_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08992_ _03134_ _03571_ _03009_ vssd1 vssd1 vccd1 vccd1 _03675_ sky130_fd_sc_hd__o21a_1
XANTENNA__10931__A _02171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07943_ genblk1\[7\].osc.clkdiv_C.cnt\[11\] _01925_ _02649_ vssd1 vssd1 vccd1 vccd1
+ _02650_ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout199_A net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07874_ _02517_ _02579_ _02577_ vssd1 vssd1 vccd1 vccd1 _02581_ sky130_fd_sc_hd__and3_1
XANTENNA__07724__B1 _01313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09613_ genblk2\[1\].wave_shpr.div.acc\[12\] _04111_ _04095_ vssd1 vssd1 vccd1 vccd1
+ _04112_ sky130_fd_sc_hd__mux2_1
X_06825_ genblk1\[5\].osc.clkdiv_C.cnt\[1\] genblk1\[5\].osc.clkdiv_C.cnt\[0\] vssd1
+ vssd1 vccd1 vccd1 _01696_ sky130_fd_sc_hd__nand2_1
X_09544_ _04055_ genblk1\[1\].osc.clkdiv_C.cnt\[10\] vssd1 vssd1 vccd1 vccd1 _04063_
+ sky130_fd_sc_hd__and2_1
X_06756_ genblk1\[4\].osc.clkdiv_C.cnt\[10\] _01631_ _01635_ _01600_ vssd1 vssd1 vccd1
+ vccd1 genblk1\[4\].osc.clkdiv_C.next_cnt\[10\] sky130_fd_sc_hd__o211a_1
XFILLER_0_78_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09475_ genblk2\[2\].wave_shpr.div.b1\[5\] _01248_ _04024_ vssd1 vssd1 vccd1 vccd1
+ _04026_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06687_ _01576_ vssd1 vssd1 vccd1 vccd1 _01577_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__06575__B _01327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08426_ _03131_ _03132_ vssd1 vssd1 vccd1 vccd1 _03133_ sky130_fd_sc_hd__and2b_1
XFILLER_0_19_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08357_ genblk2\[4\].wave_shpr.div.fin_quo\[5\] _02521_ _02838_ _03063_ vssd1 vssd1
+ vccd1 vccd1 _03064_ sky130_fd_sc_hd__a211o_1
XFILLER_0_117_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07308_ genblk1\[11\].osc.clkdiv_C.cnt\[4\] _01513_ _02070_ _02071_ vssd1 vssd1 vccd1
+ vccd1 _02072_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08288_ _02972_ _02991_ vssd1 vssd1 vccd1 vccd1 _02995_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07239_ genblk1\[10\].osc.clkdiv_C.cnt\[10\] _01215_ vssd1 vssd1 vccd1 vccd1 _02021_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10250_ _03690_ _04562_ _04563_ vssd1 vssd1 vccd1 vccd1 _00431_ sky130_fd_sc_hd__nor3_1
X_10181_ genblk2\[3\].wave_shpr.div.acc\[10\] _04513_ _04507_ vssd1 vssd1 vccd1 vccd1
+ _04514_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10052__S _04238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12822_ clknet_leaf_62_clk _00155_ net189 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.acc\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09468__B1 _03733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10078__A1 _03714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12753_ clknet_leaf_51_clk genblk1\[11\].osc.clkdiv_C.next_cnt\[12\] net110 vssd1
+ vssd1 vccd1 vccd1 genblk1\[11\].osc.clkdiv_C.cnt\[12\] sky130_fd_sc_hd__dfrtp_4
XTAP_1231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_97_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06485__B _01337_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11704_ genblk2\[9\].wave_shpr.div.b1\[12\] genblk2\[9\].wave_shpr.div.acc\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05596_ sky130_fd_sc_hd__and2b_1
XTAP_1275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12684_ clknet_leaf_120_clk genblk1\[7\].osc.clkdiv_C.next_cnt\[15\] net141 vssd1
+ vssd1 vccd1 vccd1 genblk1\[7\].osc.clkdiv_C.cnt\[15\] sky130_fd_sc_hd__dfrtp_4
XTAP_1286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11635_ genblk2\[8\].wave_shpr.div.acc\[21\] _05534_ vssd1 vssd1 vccd1 vccd1 _05537_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_112_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11566_ _05382_ _05371_ vssd1 vssd1 vccd1 vccd1 _05485_ sky130_fd_sc_hd__or2b_1
X_13305_ clknet_leaf_96_clk _00626_ net161 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.b1\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08994__A2 _01099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10517_ _04750_ _04621_ _04751_ vssd1 vssd1 vccd1 vccd1 _04752_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_122_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11497_ _05444_ vssd1 vssd1 vccd1 vccd1 _05446_ sky130_fd_sc_hd__clkbuf_4
X_13236_ clknet_leaf_15_clk _00559_ net74 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.quo\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10448_ genblk2\[4\].wave_shpr.div.acc\[6\] _04700_ _04623_ vssd1 vssd1 vccd1 vccd1
+ _04701_ sky130_fd_sc_hd__mux2_1
XANTENNA__13649__RESET_B net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13167_ clknet_leaf_123_clk net972 net76 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.acc\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10379_ net251 _04652_ _04656_ net408 vssd1 vssd1 vccd1 vccd1 _00467_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12118_ _05812_ vssd1 vssd1 vccd1 vccd1 _05876_ sky130_fd_sc_hd__clkbuf_4
X_13098_ clknet_leaf_137_clk _00425_ net39 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.acc\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12049_ _05819_ genblk1\[10\].osc.clkdiv_C.cnt\[7\] vssd1 vssd1 vccd1 vccd1 _05829_
+ sky130_fd_sc_hd__and2_1
XANTENNA__09036__B _01432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_66 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06610_ genblk1\[3\].osc.clkdiv_C.cnt\[10\] _01231_ _01515_ _01516_ _01517_ vssd1
+ vssd1 vccd1 vccd1 _01518_ sky130_fd_sc_hd__o2111a_1
X_07590_ genblk1\[9\].osc.clkdiv_C.cnt\[9\] _01991_ _01923_ genblk1\[9\].osc.clkdiv_C.cnt\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02297_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_62_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10069__A1 _04444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06541_ genblk1\[2\].osc.clkdiv_C.cnt\[6\] _01459_ vssd1 vssd1 vccd1 vccd1 _01461_
+ sky130_fd_sc_hd__and2_1
XANTENNA__09052__A _03689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06472_ genblk1\[1\].osc.clkdiv_C.cnt\[13\] _01399_ _01402_ vssd1 vssd1 vccd1 vccd1
+ genblk1\[1\].osc.clkdiv_C.next_cnt\[13\] sky130_fd_sc_hd__o21a_1
X_09260_ genblk2\[0\].wave_shpr.div.quo\[22\] _03835_ _03847_ net265 _03859_ vssd1
+ vssd1 vccd1 vccd1 _00145_ sky130_fd_sc_hd__a221o_1
XFILLER_0_75_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08211_ _02916_ _02917_ vssd1 vssd1 vccd1 vccd1 _02918_ sky130_fd_sc_hd__or2b_1
XFILLER_0_118_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09191_ _03823_ vssd1 vssd1 vccd1 vccd1 _00112_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__06693__B1 _01340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08142_ _02848_ vssd1 vssd1 vccd1 vccd1 _02849_ sky130_fd_sc_hd__inv_2
XFILLER_0_114_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07300__A _01182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08073_ _02761_ _02762_ _02779_ _02764_ vssd1 vssd1 vccd1 vccd1 _02780_ sky130_fd_sc_hd__a31o_1
XFILLER_0_114_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout114_A net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07024_ genblk1\[7\].osc.clkdiv_C.cnt\[14\] genblk1\[7\].osc.clkdiv_C.cnt\[13\] _01842_
+ vssd1 vssd1 vccd1 vccd1 _01846_ sky130_fd_sc_hd__and3_1
XFILLER_0_101_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07954__B _01805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11741__A1 _02248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07945__B1 _01805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08131__A _02221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08975_ sig_norm.quo\[7\] vssd1 vssd1 vccd1 vccd1 _03661_ sky130_fd_sc_hd__inv_2
Xhold15 genblk2\[5\].wave_shpr.div.quo\[19\] vssd1 vssd1 vccd1 vccd1 net233 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 _00878_ vssd1 vssd1 vccd1 vccd1 net244 sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 genblk2\[4\].wave_shpr.div.quo\[18\] vssd1 vssd1 vccd1 vccd1 net255 sky130_fd_sc_hd__dlygate4sd3_1
X_07926_ _02607_ _02608_ vssd1 vssd1 vccd1 vccd1 _02633_ sky130_fd_sc_hd__or2b_1
Xhold48 _00145_ vssd1 vssd1 vccd1 vccd1 net266 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 genblk2\[0\].wave_shpr.div.quo\[8\] vssd1 vssd1 vccd1 vccd1 net277 sky130_fd_sc_hd__dlygate4sd3_1
X_07857_ genblk2\[0\].wave_shpr.div.fin_quo\[0\] genblk2\[0\].wave_shpr.div.fin_quo\[1\]
+ _02510_ _02316_ vssd1 vssd1 vccd1 vccd1 _02564_ sky130_fd_sc_hd__a31oi_1
XANTENNA__11492__A _05441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10600__S _00015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06808_ genblk1\[5\].osc.clkdiv_C.cnt\[15\] _01359_ vssd1 vssd1 vccd1 vccd1 _01680_
+ sky130_fd_sc_hd__or2_1
XANTENNA__06586__A _01342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07788_ _02493_ _02494_ vssd1 vssd1 vccd1 vccd1 _02495_ sky130_fd_sc_hd__or2_1
XANTENNA__11257__B1 _05249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09527_ _04046_ vssd1 vssd1 vccd1 vccd1 _04053_ sky130_fd_sc_hd__buf_2
XFILLER_0_149_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06739_ _01600_ _01621_ _01622_ vssd1 vssd1 vccd1 vccd1 _01623_ sky130_fd_sc_hd__and3_1
XFILLER_0_79_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08122__B1 _01304_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09458_ genblk2\[1\].wave_shpr.div.fin_quo\[5\] net414 _00007_ vssd1 vssd1 vccd1
+ vccd1 _04017_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08409_ genblk2\[2\].wave_shpr.div.fin_quo\[2\] _03115_ vssd1 vssd1 vccd1 vccd1 _03116_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_19_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09389_ net288 _03952_ _03953_ vssd1 vssd1 vccd1 vccd1 _00180_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_108_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11420_ genblk2\[8\].wave_shpr.div.b1\[11\] genblk2\[8\].wave_shpr.div.acc\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05396_ sky130_fd_sc_hd__and2b_1
XFILLER_0_105_811 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11351_ _05336_ _05337_ vssd1 vssd1 vccd1 vccd1 _05338_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11980__A1 genblk2\[10\].wave_shpr.div.quo\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10302_ _04449_ genblk2\[4\].wave_shpr.div.acc\[16\] vssd1 vssd1 vccd1 vccd1 _04614_
+ sky130_fd_sc_hd__and2_1
X_11282_ genblk2\[7\].wave_shpr.div.acc\[3\] _05285_ _05222_ vssd1 vssd1 vccd1 vccd1
+ _05286_ sky130_fd_sc_hd__mux2_1
X_13021_ clknet_leaf_122_clk _00348_ net76 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.i\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10233_ genblk2\[3\].wave_shpr.div.acc\[24\] vssd1 vssd1 vccd1 vccd1 _04552_ sky130_fd_sc_hd__inv_2
XFILLER_0_120_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10164_ genblk2\[3\].wave_shpr.div.acc\[6\] _04500_ _04420_ vssd1 vssd1 vccd1 vccd1
+ _04501_ sky130_fd_sc_hd__mux2_1
XANTENNA__07951__A3 _01564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10095_ genblk2\[3\].wave_shpr.div.quo\[8\] _04452_ _04456_ net401 vssd1 vssd1 vccd1
+ vccd1 _00383_ sky130_fd_sc_hd__a22o_1
XANTENNA__11496__B1 _05417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12805_ clknet_leaf_59_clk net544 net187 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.quo\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_812 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10997_ _05051_ vssd1 vssd1 vccd1 vccd1 _05086_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__08113__B1 _01592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12624__RESET_B net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12736_ clknet_leaf_37_clk genblk1\[10\].osc.clkdiv_C.next_cnt\[13\] net114 vssd1
+ vssd1 vccd1 vccd1 genblk1\[10\].osc.clkdiv_C.cnt\[13\] sky130_fd_sc_hd__dfrtp_4
XTAP_1061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09861__B1 _04252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12667_ clknet_leaf_24_clk genblk1\[6\].osc.clkdiv_C.next_cnt\[16\] net88 vssd1 vssd1
+ vccd1 vccd1 genblk1\[6\].osc.clkdiv_C.cnt\[16\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_25_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11618_ genblk2\[8\].wave_shpr.div.acc\[16\] _05524_ _05416_ vssd1 vssd1 vccd1 vccd1
+ _05525_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12598_ clknet_leaf_21_clk genblk1\[3\].osc.clkdiv_C.next_cnt\[1\] net97 vssd1 vssd1
+ vccd1 vccd1 genblk1\[3\].osc.clkdiv_C.cnt\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_13_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07120__A _01432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11549_ genblk2\[8\].wave_shpr.div.acc\[0\] _00020_ _05471_ net274 _05472_ vssd1
+ vssd1 vccd1 vccd1 _00821_ sky130_fd_sc_hd__o221a_1
XFILLER_0_123_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold507 genblk2\[3\].wave_shpr.div.i\[2\] vssd1 vssd1 vccd1 vccd1 net725 sky130_fd_sc_hd__dlygate4sd3_1
Xhold518 genblk2\[7\].wave_shpr.div.quo\[10\] vssd1 vssd1 vccd1 vccd1 net736 sky130_fd_sc_hd__dlygate4sd3_1
Xhold529 genblk2\[6\].wave_shpr.div.b1\[14\] vssd1 vssd1 vccd1 vccd1 net747 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13219_ clknet_leaf_3_clk _00542_ net47 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.b1\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07774__B _01215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07927__B1 _01362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09047__A _01248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_867 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08760_ genblk2\[4\].wave_shpr.div.fin_quo\[0\] _02521_ _02838_ vssd1 vssd1 vccd1
+ vccd1 _03467_ sky130_fd_sc_hd__a21o_1
XTAP_889 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07711_ net2 net163 _02312_ vssd1 vssd1 vccd1 vccd1 _02418_ sky130_fd_sc_hd__and3_1
X_08691_ _03340_ _03350_ _03349_ vssd1 vssd1 vccd1 vccd1 _03398_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_79_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_79_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07642_ net33 vssd1 vssd1 vccd1 vccd1 _02349_ sky130_fd_sc_hd__clkbuf_4
X_07573_ _02278_ _02279_ vssd1 vssd1 vccd1 vccd1 _02280_ sky130_fd_sc_hd__nand2_1
XANTENNA__08104__B1 _01592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09312_ _03783_ _03753_ vssd1 vssd1 vccd1 vccd1 _03897_ sky130_fd_sc_hd__or2b_1
X_06524_ _01410_ _01231_ _01413_ _01429_ _01449_ vssd1 vssd1 vccd1 vccd1 _01450_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_146_711 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09510__A _04046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06666__B1 _01223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09243_ _03725_ genblk1\[0\].osc.clkdiv_C.cnt\[6\] vssd1 vssd1 vccd1 vccd1 _03850_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_146_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06455_ _01391_ vssd1 vssd1 vccd1 vccd1 genblk1\[1\].osc.clkdiv_C.next_cnt\[7\] sky130_fd_sc_hd__clkbuf_1
XANTENNA__07949__B _02011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10656__A _04856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06386_ genblk1\[1\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 _01330_ sky130_fd_sc_hd__inv_2
X_09174_ genblk2\[10\].wave_shpr.div.b1\[0\] _03813_ _03722_ vssd1 vssd1 vccd1 vccd1
+ _03814_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08125_ _01570_ _01870_ _02829_ _02830_ _02831_ vssd1 vssd1 vccd1 vccd1 _02832_ sky130_fd_sc_hd__o2111ai_1
XFILLER_0_133_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09080__A1 _03732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08056_ _02761_ _02762_ vssd1 vssd1 vccd1 vccd1 _02763_ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07007_ genblk1\[7\].osc.clkdiv_C.cnt\[8\] genblk1\[7\].osc.clkdiv_C.cnt\[7\] _01832_
+ vssd1 vssd1 vccd1 vccd1 _01835_ sky130_fd_sc_hd__and3_1
XFILLER_0_113_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12082__S _05787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10391__A _04058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08958_ _03565_ _03646_ vssd1 vssd1 vccd1 vccd1 _03647_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07501__A_N net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07909_ genblk1\[8\].osc.clkdiv_C.cnt\[11\] _01869_ _02613_ _02614_ _02615_ vssd1
+ vssd1 vccd1 vccd1 _02616_ sky130_fd_sc_hd__o221a_1
X_08889_ sig_norm.acc\[11\] sig_norm.acc\[12\] _03591_ _03594_ vssd1 vssd1 vccd1 vccd1
+ _03595_ sky130_fd_sc_hd__or4_1
X_10920_ genblk2\[7\].wave_shpr.div.b1\[11\] _02433_ _05042_ vssd1 vssd1 vccd1 vccd1
+ _05045_ sky130_fd_sc_hd__mux2_1
X_10851_ _04977_ _04993_ _04994_ vssd1 vssd1 vccd1 vccd1 _04995_ sky130_fd_sc_hd__a21o_1
XFILLER_0_85_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13570_ clknet_leaf_56_clk net363 net182 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.quo\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10782_ _04815_ _04880_ net630 vssd1 vssd1 vccd1 vccd1 _04939_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_39_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12521_ clknet_leaf_103_clk PWM.next_counter\[5\] net156 vssd1 vssd1 vccd1 vccd1
+ PWM.counter\[5\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_40_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12452_ clknet_leaf_116_clk net222 net150 vssd1 vssd1 vccd1 vccd1 modein.delay_in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11403_ _05373_ _05377_ _05378_ vssd1 vssd1 vccd1 vccd1 _05379_ sky130_fd_sc_hd__a21o_1
XFILLER_0_152_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12383_ net762 _06039_ _06040_ _06059_ vssd1 vssd1 vccd1 vccd1 _01068_ sky130_fd_sc_hd__a22o_1
XANTENNA__09071__A1 _03726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09071__B2 _03727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11334_ _05213_ _05165_ vssd1 vssd1 vccd1 vccd1 _05325_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07621__A2 _01430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_55_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11265_ _03819_ net1255 _00018_ genblk2\[7\].wave_shpr.div.acc\[0\] _05272_ vssd1
+ vssd1 vccd1 vccd1 _00737_ sky130_fd_sc_hd__o221a_1
X_13004_ clknet_leaf_138_clk _00333_ net39 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.acc\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10216_ net904 _04518_ _04522_ _04540_ vssd1 vssd1 vccd1 vccd1 _00420_ sky130_fd_sc_hd__a22o_1
X_11196_ _05238_ vssd1 vssd1 vccd1 vccd1 _00702_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11181__A2 _01242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10147_ _04383_ _04487_ vssd1 vssd1 vccd1 vccd1 _04488_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_113_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10078_ _03714_ _04449_ _03736_ vssd1 vssd1 vccd1 vccd1 _00373_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07688__A2 _01215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07115__A genblk1\[8\].osc.clkdiv_C.cnt\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_128_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13768_ clknet_leaf_71_clk _01079_ net217 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.acc\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08637__A1 _02592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12719_ clknet_leaf_86_clk genblk1\[9\].osc.clkdiv_C.next_cnt\[14\] net181 vssd1
+ vssd1 vccd1 vccd1 genblk1\[9\].osc.clkdiv_C.cnt\[14\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_127_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_0_clk clk vssd1 vssd1 vccd1 vccd1 clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__10476__A _04654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13699_ clknet_leaf_94_clk _01010_ net160 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.fin_quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_254 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06240_ _01201_ genblk1\[0\].osc.clkdiv_C.cnt\[7\] genblk1\[0\].osc.clkdiv_C.cnt\[8\]
+ vssd1 vssd1 vccd1 vccd1 _01202_ sky130_fd_sc_hd__a21o_1
XFILLER_0_155_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06171_ _01121_ _01123_ _01142_ vssd1 vssd1 vccd1 vccd1 _01143_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_131_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold304 genblk2\[0\].wave_shpr.div.quo\[16\] vssd1 vssd1 vccd1 vccd1 net522 sky130_fd_sc_hd__dlygate4sd3_1
Xhold315 genblk2\[9\].wave_shpr.div.quo\[20\] vssd1 vssd1 vccd1 vccd1 net533 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold326 _00138_ vssd1 vssd1 vccd1 vccd1 net544 sky130_fd_sc_hd__dlygate4sd3_1
Xhold337 genblk2\[10\].wave_shpr.div.quo\[5\] vssd1 vssd1 vccd1 vccd1 net555 sky130_fd_sc_hd__dlygate4sd3_1
Xhold348 genblk2\[5\].wave_shpr.div.acc\[21\] vssd1 vssd1 vccd1 vccd1 net566 sky130_fd_sc_hd__dlygate4sd3_1
X_09930_ net605 _04315_ _04322_ _04338_ vssd1 vssd1 vccd1 vccd1 _00336_ sky130_fd_sc_hd__a22o_1
Xhold359 genblk2\[0\].wave_shpr.div.b1\[15\] vssd1 vssd1 vccd1 vccd1 net577 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09861_ net918 _04282_ _04252_ _04285_ vssd1 vssd1 vccd1 vccd1 _00320_ sky130_fd_sc_hd__a22o_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08812_ _03517_ _03518_ vssd1 vssd1 vccd1 vccd1 _03519_ sky130_fd_sc_hd__or2b_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09792_ _04246_ vssd1 vssd1 vccd1 vccd1 _00290_ sky130_fd_sc_hd__clkbuf_1
Xhold1004 genblk2\[8\].wave_shpr.div.acc\[18\] vssd1 vssd1 vccd1 vccd1 net1222 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1015 genblk2\[6\].wave_shpr.div.b1\[11\] vssd1 vssd1 vccd1 vccd1 net1233 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1026 genblk2\[10\].wave_shpr.div.b1\[8\] vssd1 vssd1 vccd1 vccd1 net1244 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08743_ _03447_ _03448_ _03445_ _03446_ vssd1 vssd1 vccd1 vccd1 _03450_ sky130_fd_sc_hd__a211oi_4
Xhold1037 genblk1\[7\].osc.clkdiv_C.cnt\[17\] vssd1 vssd1 vccd1 vccd1 net1255 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11754__B genblk1\[9\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09505__A _04042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1048 genblk2\[5\].wave_shpr.div.b1\[11\] vssd1 vssd1 vccd1 vccd1 net1266 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1059 genblk2\[2\].wave_shpr.div.b1\[12\] vssd1 vssd1 vccd1 vccd1 net1277 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout181_A net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08325__B1 _02223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08674_ _03359_ _03379_ _03380_ vssd1 vssd1 vccd1 vccd1 _03381_ sky130_fd_sc_hd__nor3_2
XFILLER_0_95_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07625_ genblk1\[11\].osc.clkdiv_C.cnt\[13\] _01208_ _01576_ genblk1\[11\].osc.clkdiv_C.cnt\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02332_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07556_ genblk2\[9\].wave_shpr.div.fin_quo\[2\] _02262_ vssd1 vssd1 vccd1 vccd1 _02263_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_76_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06507_ _01200_ _01432_ vssd1 vssd1 vccd1 vccd1 _01433_ sky130_fd_sc_hd__nand2_2
XFILLER_0_118_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07487_ genblk2\[11\].wave_shpr.div.i\[1\] _02210_ genblk2\[11\].wave_shpr.div.i\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02211_ sky130_fd_sc_hd__or3b_1
XANTENNA__06583__B _01250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_591 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10986__A2 _05051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09226_ genblk2\[0\].wave_shpr.div.quo\[7\] _03836_ _03840_ net269 vssd1 vssd1 vccd1
+ vccd1 _00130_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06438_ _01373_ _01378_ _01379_ vssd1 vssd1 vccd1 vccd1 genblk1\[1\].osc.clkdiv_C.next_cnt\[2\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_106_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09157_ genblk2\[0\].wave_shpr.div.fin_quo\[0\] _03804_ _00001_ vssd1 vssd1 vccd1
+ vccd1 _03805_ sky130_fd_sc_hd__mux2_1
X_06369_ _01192_ _01208_ vssd1 vssd1 vccd1 vccd1 _01313_ sky130_fd_sc_hd__nand2_4
X_08108_ _02812_ _02809_ _02813_ _02814_ vssd1 vssd1 vccd1 vccd1 _02815_ sky130_fd_sc_hd__or4_1
XFILLER_0_133_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09088_ _03737_ modein.delay_octave_down_in\[1\] _01591_ _03738_ vssd1 vssd1 vccd1
+ vccd1 _03739_ sky130_fd_sc_hd__o211a_1
XFILLER_0_114_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08039_ _02741_ _02743_ _02745_ vssd1 vssd1 vccd1 vccd1 _02746_ sky130_fd_sc_hd__o21a_1
Xhold860 genblk2\[11\].wave_shpr.div.acc\[25\] vssd1 vssd1 vccd1 vccd1 net1078 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout94_A net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold871 genblk1\[0\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 net1089 sky130_fd_sc_hd__dlygate4sd3_1
Xhold882 genblk2\[4\].wave_shpr.div.b1\[1\] vssd1 vssd1 vccd1 vccd1 net1100 sky130_fd_sc_hd__dlygate4sd3_1
Xhold893 PWM.final_sample_in\[0\] vssd1 vssd1 vccd1 vccd1 net1111 sky130_fd_sc_hd__dlygate4sd3_1
X_11050_ _05010_ _04969_ vssd1 vssd1 vccd1 vccd1 _05127_ sky130_fd_sc_hd__or2b_1
XFILLER_0_102_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10001_ genblk2\[3\].wave_shpr.div.b1\[9\] genblk2\[3\].wave_shpr.div.acc\[9\] vssd1
+ vssd1 vccd1 vccd1 _04397_ sky130_fd_sc_hd__and2b_1
XANTENNA__07772__D1 _02336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11952_ genblk2\[10\].wave_shpr.div.b1\[14\] genblk2\[10\].wave_shpr.div.acc\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05774_ sky130_fd_sc_hd__and2b_1
XFILLER_0_98_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10903_ _05035_ vssd1 vssd1 vccd1 vccd1 _00612_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_58_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_86_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11883_ net646 _05609_ _05713_ vssd1 vssd1 vccd1 vccd1 _05714_ sky130_fd_sc_hd__a21o_1
XFILLER_0_39_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13622_ clknet_leaf_75_clk _00935_ net204 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.b1\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10834_ genblk2\[6\].wave_shpr.div.acc\[5\] genblk2\[6\].wave_shpr.div.b1\[5\] vssd1
+ vssd1 vccd1 vccd1 _04978_ sky130_fd_sc_hd__or2b_1
XFILLER_0_13_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13553_ clknet_leaf_100_clk net687 net164 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10765_ _04808_ _04766_ vssd1 vssd1 vccd1 vccd1 _04926_ sky130_fd_sc_hd__or2b_1
XFILLER_0_81_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12504_ clknet_leaf_106_clk _00066_ net154 vssd1 vssd1 vccd1 vccd1 PWM.final_in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13484_ clknet_leaf_99_clk _00801_ net168 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10696_ genblk2\[5\].wave_shpr.div.quo\[22\] _02183_ _04856_ net245 _04875_ vssd1
+ vssd1 vccd1 vccd1 _00565_ sky130_fd_sc_hd__a221o_1
XFILLER_0_152_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12435_ genblk2\[11\].wave_shpr.div.acc\[22\] _06096_ vssd1 vssd1 vccd1 vccd1 _06098_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_140_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12366_ net958 _06039_ _06040_ _06046_ vssd1 vssd1 vccd1 vccd1 _01064_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11317_ _05205_ _05169_ vssd1 vssd1 vccd1 vccd1 _05312_ sky130_fd_sc_hd__or2b_1
XFILLER_0_50_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12297_ _03942_ vssd1 vssd1 vccd1 vccd1 _06009_ sky130_fd_sc_hd__buf_4
XFILLER_0_129_25 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11248_ _05260_ genblk1\[7\].osc.clkdiv_C.cnt\[9\] vssd1 vssd1 vccd1 vccd1 _05264_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_120_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10362__B1 _03736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11179_ _03831_ net864 _03705_ vssd1 vssd1 vccd1 vccd1 _00693_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_89_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07410_ _02154_ vssd1 vssd1 vccd1 vccd1 _00001_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08390_ genblk1\[2\].osc.clkdiv_C.cnt\[8\] _01442_ _02011_ genblk1\[2\].osc.clkdiv_C.cnt\[7\]
+ vssd1 vssd1 vccd1 vccd1 _03097_ sky130_fd_sc_hd__a22o_1
XANTENNA__09807__B1 _04252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07341_ _02101_ vssd1 vssd1 vccd1 vccd1 _02102_ sky130_fd_sc_hd__inv_2
XANTENNA__11090__A1 _05051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07272_ genblk1\[10\].osc.clkdiv_C.cnt\[8\] genblk1\[10\].osc.clkdiv_C.cnt\[7\] _02041_
+ vssd1 vssd1 vccd1 vccd1 _02046_ sky130_fd_sc_hd__and3_1
XFILLER_0_73_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07833__A2 _02539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09011_ _03685_ vssd1 vssd1 vccd1 vccd1 _00070_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06223_ _01184_ vssd1 vssd1 vccd1 vccd1 _01185_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10934__A _05051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06154_ _01124_ _01125_ vssd1 vssd1 vccd1 vccd1 _01126_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold101 genblk2\[8\].wave_shpr.div.i\[4\] vssd1 vssd1 vccd1 vccd1 net319 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_112_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold112 _00805_ vssd1 vssd1 vccd1 vccd1 net330 sky130_fd_sc_hd__dlygate4sd3_1
Xhold123 _00230_ vssd1 vssd1 vccd1 vccd1 net341 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_124_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_238 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold134 _01049_ vssd1 vssd1 vccd1 vccd1 net352 sky130_fd_sc_hd__dlygate4sd3_1
Xhold145 _00885_ vssd1 vssd1 vccd1 vccd1 net363 sky130_fd_sc_hd__dlygate4sd3_1
Xhold156 genblk2\[9\].wave_shpr.div.b1\[14\] vssd1 vssd1 vccd1 vccd1 net374 sky130_fd_sc_hd__dlygate4sd3_1
Xhold167 genblk2\[6\].wave_shpr.div.quo\[23\] vssd1 vssd1 vccd1 vccd1 net385 sky130_fd_sc_hd__dlygate4sd3_1
Xhold178 genblk2\[0\].wave_shpr.div.b1\[16\] vssd1 vssd1 vccd1 vccd1 net396 sky130_fd_sc_hd__dlygate4sd3_1
X_09913_ net1036 _04315_ _04322_ _04325_ vssd1 vssd1 vccd1 vccd1 _00332_ sky130_fd_sc_hd__a22o_1
Xhold189 smpl_rt_clkdiv.clkDiv_inst.cnt\[5\] vssd1 vssd1 vccd1 vccd1 net407 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09844_ net259 _04247_ _04250_ net520 _04273_ vssd1 vssd1 vccd1 vccd1 _00315_ sky130_fd_sc_hd__a221o_1
XANTENNA__07962__B _01361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08010__A2 _01365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09775_ genblk2\[3\].wave_shpr.div.b1\[10\] _02336_ _04039_ vssd1 vssd1 vccd1 vccd1
+ _04237_ sky130_fd_sc_hd__mux2_1
X_06987_ _01822_ vssd1 vssd1 vccd1 vccd1 _01823_ sky130_fd_sc_hd__clkbuf_4
X_08726_ _03397_ _03400_ _03432_ vssd1 vssd1 vccd1 vccd1 _03433_ sky130_fd_sc_hd__a21oi_1
XTAP_2306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08657_ genblk2\[3\].wave_shpr.div.fin_quo\[2\] _03363_ vssd1 vssd1 vccd1 vccd1 _03364_
+ sky130_fd_sc_hd__xnor2_1
XTAP_1605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07608_ _02306_ _02311_ _02314_ vssd1 vssd1 vccd1 vccd1 _02315_ sky130_fd_sc_hd__o21a_1
XTAP_1638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08588_ _03293_ _03294_ vssd1 vssd1 vccd1 vccd1 _03295_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_76_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07539_ PWM.final_sample_in\[1\] net1103 PWM.start vssd1 vssd1 vccd1 vccd1 _02253_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10550_ _04776_ _04777_ vssd1 vssd1 vccd1 vccd1 _04778_ sky130_fd_sc_hd__nand2_1
XFILLER_0_107_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09209_ _03714_ _03832_ _03736_ vssd1 vssd1 vccd1 vccd1 _00121_ sky130_fd_sc_hd__o21ai_1
X_10481_ _04610_ _04568_ vssd1 vssd1 vccd1 vccd1 _04726_ sky130_fd_sc_hd__or2b_1
XFILLER_0_17_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12220_ _05934_ _05956_ _05957_ vssd1 vssd1 vccd1 vccd1 _05958_ sky130_fd_sc_hd__a21o_1
XFILLER_0_121_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12030__B1 _05817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08314__A _02216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12151_ _05900_ _05901_ vssd1 vssd1 vccd1 vccd1 _05902_ sky130_fd_sc_hd__nand2_1
XFILLER_0_20_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10055__S _04238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11102_ net280 _05162_ _03855_ vssd1 vssd1 vccd1 vccd1 _05163_ sky130_fd_sc_hd__o21ai_1
X_12082_ genblk2\[10\].wave_shpr.div.acc\[2\] _05848_ _05787_ vssd1 vssd1 vccd1 vccd1
+ _05849_ sky130_fd_sc_hd__mux2_1
Xhold690 genblk2\[8\].wave_shpr.div.acc\[10\] vssd1 vssd1 vccd1 vccd1 net908 sky130_fd_sc_hd__dlygate4sd3_1
X_11033_ _05001_ _05113_ vssd1 vssd1 vccd1 vccd1 _05114_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08001__A2 _01577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12984_ clknet_leaf_13_clk net262 net69 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.quo\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_11935_ _05742_ _05755_ _05756_ vssd1 vssd1 vccd1 vccd1 _05757_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_115_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11866_ _05605_ _05701_ vssd1 vssd1 vccd1 vccd1 _05702_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12344__B_N _03941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13605_ clknet_leaf_59_clk _00918_ net193 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.i\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_145_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10817_ _04962_ vssd1 vssd1 vccd1 vccd1 _04963_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11797_ genblk2\[9\].wave_shpr.div.b1\[0\] _05573_ _05574_ vssd1 vssd1 vccd1 vccd1
+ _05649_ sky130_fd_sc_hd__and3_1
XFILLER_0_131_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13536_ clknet_leaf_81_clk _00851_ net199 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.i\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10748_ _04799_ _04912_ vssd1 vssd1 vccd1 vccd1 _04913_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13467_ clknet_leaf_75_clk _00784_ net203 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.b1\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10679_ net249 _04861_ _04862_ net294 _04866_ vssd1 vssd1 vccd1 vccd1 _00557_ sky130_fd_sc_hd__a221o_1
XFILLER_0_125_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12021__B1 _05787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12418_ _05974_ _06085_ vssd1 vssd1 vccd1 vccd1 _06086_ sky130_fd_sc_hd__xnor2_1
X_13398_ clknet_leaf_117_clk _00717_ net140 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12349_ genblk2\[11\].wave_shpr.div.acc\[1\] _05981_ vssd1 vssd1 vccd1 vccd1 _06033_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12891__RESET_B net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06910_ _01761_ _01762_ vssd1 vssd1 vccd1 vccd1 genblk1\[6\].osc.clkdiv_C.next_cnt\[1\]
+ sky130_fd_sc_hd__nor2_1
X_07890_ genblk2\[0\].wave_shpr.div.fin_quo\[7\] _02539_ _02596_ _02592_ vssd1 vssd1
+ vccd1 vccd1 _02597_ sky130_fd_sc_hd__a22o_1
X_06841_ _01693_ _01705_ _01706_ vssd1 vssd1 vccd1 vccd1 genblk1\[5\].osc.clkdiv_C.next_cnt\[6\]
+ sky130_fd_sc_hd__nor3_1
X_09560_ _03819_ genblk1\[1\].osc.clkdiv_C.cnt\[17\] _00006_ net752 _04071_ vssd1
+ vssd1 vccd1 vccd1 _00233_ sky130_fd_sc_hd__o221a_1
X_06772_ _01647_ vssd1 vssd1 vccd1 vccd1 _01648_ sky130_fd_sc_hd__inv_2
X_08511_ _03079_ _03126_ _03125_ vssd1 vssd1 vccd1 vccd1 _03218_ sky130_fd_sc_hd__o21ai_1
X_09491_ _04035_ vssd1 vssd1 vccd1 vccd1 _00200_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08442_ _02416_ _03148_ _02419_ vssd1 vssd1 vccd1 vccd1 _03149_ sky130_fd_sc_hd__o21a_1
XFILLER_0_81_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08373_ _02599_ vssd1 vssd1 vccd1 vccd1 _03080_ sky130_fd_sc_hd__inv_2
XANTENNA__08059__A2 _01238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout144_A net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07324_ genblk1\[11\].osc.clkdiv_C.cnt\[3\] _01334_ _02086_ _01197_ _02087_ vssd1
+ vssd1 vccd1 vccd1 _02088_ sky130_fd_sc_hd__o221a_1
XFILLER_0_90_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07255_ genblk1\[10\].osc.clkdiv_C.cnt\[3\] _02032_ vssd1 vssd1 vccd1 vccd1 _02034_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_6_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12355__S _05982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06206_ net399 _01166_ vssd1 vssd1 vccd1 vccd1 PWM.next_counter\[7\] sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07186_ genblk1\[9\].osc.clkdiv_C.cnt\[10\] _01974_ vssd1 vssd1 vccd1 vccd1 _01976_
+ sky130_fd_sc_hd__nand2_1
X_06137_ net1 net7 vssd1 vssd1 vccd1 vccd1 _01109_ sky130_fd_sc_hd__or2_1
XANTENNA__11495__A _05444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07692__B _02011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09827_ _04058_ _01412_ vssd1 vssd1 vccd1 vccd1 _04264_ sky130_fd_sc_hd__nor2_1
XANTENNA__12079__B1 _05817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09758_ genblk2\[3\].wave_shpr.div.b1\[2\] _04227_ _04039_ vssd1 vssd1 vccd1 vccd1
+ _04228_ sky130_fd_sc_hd__mux2_1
XTAP_2103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout57_A net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08709_ _03114_ _03415_ _03122_ vssd1 vssd1 vccd1 vccd1 _03416_ sky130_fd_sc_hd__o21a_1
XTAP_2114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09495__A1 net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09689_ genblk2\[2\].wave_shpr.div.acc\[4\] genblk2\[2\].wave_shpr.div.b1\[4\] vssd1
+ vssd1 vccd1 vccd1 _04169_ sky130_fd_sc_hd__or2b_1
XTAP_2136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11720_ _05610_ _05611_ vssd1 vssd1 vccd1 vccd1 _05612_ sky130_fd_sc_hd__or2_1
XFILLER_0_84_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11651_ genblk2\[8\].wave_shpr.div.i\[1\] genblk2\[8\].wave_shpr.div.i\[0\] vssd1
+ vssd1 vccd1 vccd1 _05547_ sky130_fd_sc_hd__nand2_1
XTAP_1479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_111 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout40 net44 vssd1 vssd1 vccd1 vccd1 net40 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_49_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08028__B genblk2\[6\].wave_shpr.div.fin_quo\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout51 net53 vssd1 vssd1 vccd1 vccd1 net51 sky130_fd_sc_hd__buf_4
XFILLER_0_153_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_138_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout62 net63 vssd1 vssd1 vccd1 vccd1 net62 sky130_fd_sc_hd__clkbuf_4
X_10602_ genblk2\[5\].wave_shpr.div.fin_quo\[4\] net1326 _00015_ vssd1 vssd1 vccd1
+ vccd1 _04826_ sky130_fd_sc_hd__mux2_1
XANTENNA__09798__A2 _04248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout73 net74 vssd1 vssd1 vccd1 vccd1 net73 sky130_fd_sc_hd__clkbuf_4
X_11582_ net978 _05447_ _05484_ _05497_ vssd1 vssd1 vccd1 vccd1 _00829_ sky130_fd_sc_hd__a22o_1
Xfanout84 net85 vssd1 vssd1 vccd1 vccd1 net84 sky130_fd_sc_hd__buf_2
XFILLER_0_92_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout95 net98 vssd1 vssd1 vccd1 vccd1 net95 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_119_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13321_ clknet_leaf_26_clk _00642_ net87 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.quo\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10533_ net281 _04761_ _03855_ vssd1 vssd1 vccd1 vccd1 _04762_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_52_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12265__S _05802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13252_ clknet_leaf_1_clk _00575_ net41 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.acc\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10464_ _04601_ _04712_ vssd1 vssd1 vccd1 vccd1 _04713_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_150_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12203_ genblk2\[11\].wave_shpr.div.acc\[1\] genblk2\[11\].wave_shpr.div.b1\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05941_ sky130_fd_sc_hd__xor2_1
XFILLER_0_33_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13183_ clknet_leaf_112_clk _00508_ net129 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.acc\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10395_ _04477_ genblk1\[4\].osc.clkdiv_C.cnt\[6\] vssd1 vssd1 vccd1 vccd1 _04666_
+ sky130_fd_sc_hd__and2_1
X_12134_ genblk2\[10\].wave_shpr.div.acc\[14\] _05888_ _05865_ vssd1 vssd1 vccd1 vccd1
+ _05889_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06784__A2 _01304_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12306__B2 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12065_ genblk2\[10\].wave_shpr.div.quo\[23\] _05812_ _05815_ net474 _05837_ vssd1
+ vssd1 vccd1 vccd1 _00972_ sky130_fd_sc_hd__a221o_1
XFILLER_0_19_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11016_ _04993_ _05100_ vssd1 vssd1 vccd1 vccd1 _05101_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_126_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12967_ clknet_leaf_111_clk net697 net130 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11918_ genblk2\[10\].wave_shpr.div.acc\[8\] genblk2\[10\].wave_shpr.div.b1\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05740_ sky130_fd_sc_hd__or2b_1
XFILLER_0_59_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12898_ clknet_leaf_31_clk _00229_ net102 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.quo\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07123__A _01432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_146 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11849_ _05598_ _05558_ vssd1 vssd1 vccd1 vccd1 _05689_ sky130_fd_sc_hd__or2b_1
XFILLER_0_28_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09749__S _00009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13519_ clknet_leaf_79_clk _00836_ net206 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.acc\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07040_ _01489_ _01344_ vssd1 vssd1 vccd1 vccd1 _01858_ sky130_fd_sc_hd__nand2_4
XANTENNA__06472__A1 genblk1\[1\].osc.clkdiv_C.cnt\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11114__B_N genblk2\[7\].wave_shpr.div.b1\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_377 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08991_ _03674_ vssd1 vssd1 vccd1 vccd1 _00061_ sky130_fd_sc_hd__clkbuf_1
X_07942_ genblk1\[7\].osc.clkdiv_C.cnt\[10\] _01311_ _01925_ genblk1\[7\].osc.clkdiv_C.cnt\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02649_ sky130_fd_sc_hd__o22a_1
XANTENNA__11264__B_N _05249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07873_ _02517_ _02577_ _02579_ vssd1 vssd1 vccd1 vccd1 _02580_ sky130_fd_sc_hd__a21o_1
X_09612_ _03993_ _04110_ vssd1 vssd1 vccd1 vccd1 _04111_ sky130_fd_sc_hd__xnor2_1
X_06824_ genblk1\[5\].osc.clkdiv_C.cnt\[1\] genblk1\[5\].osc.clkdiv_C.cnt\[0\] vssd1
+ vssd1 vccd1 vccd1 _01695_ sky130_fd_sc_hd__or2_1
XANTENNA__11762__B genblk1\[9\].osc.clkdiv_C.cnt\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09543_ net426 _04052_ _04053_ genblk2\[1\].wave_shpr.div.quo\[17\] _04062_ vssd1
+ vssd1 vccd1 vccd1 _00225_ sky130_fd_sc_hd__a221o_1
X_06755_ genblk1\[4\].osc.clkdiv_C.cnt\[10\] _01631_ vssd1 vssd1 vccd1 vccd1 _01635_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09477__A1 _01437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09474_ _04025_ vssd1 vssd1 vccd1 vccd1 _00193_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06686_ _01575_ vssd1 vssd1 vccd1 vccd1 _01576_ sky130_fd_sc_hd__buf_4
XFILLER_0_148_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08425_ _03011_ _03128_ vssd1 vssd1 vccd1 vccd1 _03132_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08356_ _03061_ _03062_ vssd1 vssd1 vccd1 vccd1 _03063_ sky130_fd_sc_hd__nor2_1
XANTENNA__06872__A _01441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07307_ genblk1\[11\].osc.clkdiv_C.cnt\[0\] _01223_ _01678_ vssd1 vssd1 vccd1 vccd1
+ _02071_ sky130_fd_sc_hd__or3_1
XFILLER_0_144_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08287_ _02964_ _02958_ _02963_ vssd1 vssd1 vccd1 vccd1 _02994_ sky130_fd_sc_hd__a21o_1
XFILLER_0_117_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06463__A1 genblk1\[1\].osc.clkdiv_C.cnt\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07238_ genblk1\[10\].osc.clkdiv_C.cnt\[12\] _02011_ _02012_ _02014_ _02019_ vssd1
+ vssd1 vccd1 vccd1 _02020_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07169_ _01964_ vssd1 vssd1 vccd1 vccd1 genblk1\[9\].osc.clkdiv_C.next_cnt\[4\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10180_ _04398_ _04512_ vssd1 vssd1 vccd1 vccd1 _04513_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07963__A1 _01200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11511__A2 _05448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12821_ clknet_leaf_67_clk net824 net196 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.acc\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09468__A1 _03732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12752_ clknet_leaf_50_clk genblk1\[11\].osc.clkdiv_C.next_cnt\[11\] net111 vssd1
+ vssd1 vccd1 vccd1 genblk1\[11\].osc.clkdiv_C.cnt\[11\] sky130_fd_sc_hd__dfrtp_1
XTAP_1221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11703_ _05560_ _05593_ _05594_ vssd1 vssd1 vccd1 vccd1 _05595_ sky130_fd_sc_hd__a21o_1
XTAP_1254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12683_ clknet_leaf_120_clk genblk1\[7\].osc.clkdiv_C.next_cnt\[14\] net81 vssd1
+ vssd1 vccd1 vccd1 genblk1\[7\].osc.clkdiv_C.cnt\[14\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_84_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11634_ genblk2\[8\].wave_shpr.div.acc\[21\] _05534_ vssd1 vssd1 vccd1 vccd1 _05536_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11565_ _05444_ vssd1 vssd1 vccd1 vccd1 _05484_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_64_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13304_ clknet_leaf_96_clk _00625_ net161 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.b1\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10516_ _04750_ _04748_ vssd1 vssd1 vccd1 vccd1 _04751_ sky130_fd_sc_hd__nand2_1
X_11496_ net743 _05442_ _05417_ _05445_ vssd1 vssd1 vccd1 vccd1 _00795_ sky130_fd_sc_hd__a22o_1
X_13235_ clknet_leaf_15_clk net250 net73 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.quo\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10447_ _04593_ _04699_ vssd1 vssd1 vccd1 vccd1 _04700_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_32_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13166_ clknet_leaf_127_clk _00491_ net79 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.acc\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10378_ net408 _04652_ _04656_ net508 vssd1 vssd1 vccd1 vccd1 _00466_ sky130_fd_sc_hd__a22o_1
X_12117_ net844 _05844_ _05850_ _05875_ vssd1 vssd1 vccd1 vccd1 _00986_ sky130_fd_sc_hd__a22o_1
XANTENNA__11750__A2 _05623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13097_ clknet_leaf_137_clk _00424_ net41 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.acc\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08221__B _02789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12048_ net357 _05823_ _05825_ net373 _05828_ vssd1 vssd1 vccd1 vccd1 _00964_ sky130_fd_sc_hd__a221o_1
XANTENNA__06509__A2 _01365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08903__B1 _01157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06676__B _01565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06540_ _01452_ _01459_ _01460_ vssd1 vssd1 vccd1 vccd1 genblk1\[2\].osc.clkdiv_C.next_cnt\[5\]
+ sky130_fd_sc_hd__nor3_1
XANTENNA__09052__B _01242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_55 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06471_ _01373_ _01401_ vssd1 vssd1 vccd1 vccd1 _01402_ sky130_fd_sc_hd__nor2_1
X_08210_ _02315_ _02421_ vssd1 vssd1 vccd1 vccd1 _02917_ sky130_fd_sc_hd__xor2_1
X_09190_ net1254 _03706_ _03822_ vssd1 vssd1 vccd1 vccd1 _03823_ sky130_fd_sc_hd__mux2_1
XANTENNA_hold82_A genblk2\[2\].wave_shpr.div.quo\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08141_ _02799_ _02847_ vssd1 vssd1 vccd1 vccd1 _02848_ sky130_fd_sc_hd__xor2_2
XFILLER_0_16_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12844__D _00007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08072_ genblk1\[5\].osc.clkdiv_C.cnt\[6\] _01309_ _01180_ _02767_ _02766_ vssd1
+ vssd1 vccd1 vccd1 _02779_ sky130_fd_sc_hd__a311o_1
XANTENNA__07300__B _01226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07023_ genblk1\[7\].osc.clkdiv_C.cnt\[13\] _01842_ genblk1\[7\].osc.clkdiv_C.cnt\[14\]
+ vssd1 vssd1 vccd1 vccd1 _01845_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10529__B1 _04657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout107_A net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10153__S _04420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08974_ _03660_ vssd1 vssd1 vccd1 vccd1 _00058_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08131__B _02837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold16 _00563_ vssd1 vssd1 vccd1 vccd1 net234 sky130_fd_sc_hd__dlygate4sd3_1
Xhold27 genblk2\[5\].wave_shpr.div.quo\[21\] vssd1 vssd1 vccd1 vccd1 net245 sky130_fd_sc_hd__dlygate4sd3_1
X_07925_ _02609_ _02616_ _02629_ _02631_ vssd1 vssd1 vccd1 vccd1 _02632_ sky130_fd_sc_hd__o22a_1
Xhold38 _00478_ vssd1 vssd1 vccd1 vccd1 net256 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 genblk2\[9\].wave_shpr.div.quo\[6\] vssd1 vssd1 vccd1 vccd1 net267 sky130_fd_sc_hd__buf_1
XANTENNA__11773__A _04676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold1124_A genblk2\[5\].wave_shpr.div.quo\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07856_ genblk2\[0\].wave_shpr.div.fin_quo\[0\] net31 genblk2\[0\].wave_shpr.div.fin_quo\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02563_ sky130_fd_sc_hd__a21o_1
X_06807_ genblk1\[5\].osc.clkdiv_C.cnt\[9\] _01678_ vssd1 vssd1 vccd1 vccd1 _01679_
+ sky130_fd_sc_hd__nor2_1
X_07787_ genblk1\[0\].osc.clkdiv_C.cnt\[8\] _01193_ _01184_ genblk1\[0\].osc.clkdiv_C.cnt\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02494_ sky130_fd_sc_hd__a22o_1
XANTENNA__06586__B _01248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09526_ _04042_ vssd1 vssd1 vccd1 vccd1 _04052_ sky130_fd_sc_hd__buf_2
X_06738_ genblk1\[4\].osc.clkdiv_C.cnt\[6\] _01616_ vssd1 vssd1 vccd1 vccd1 _01622_
+ sky130_fd_sc_hd__or2_1
XPHY_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09457_ _04016_ vssd1 vssd1 vccd1 vccd1 _00185_ sky130_fd_sc_hd__clkbuf_1
X_06669_ _01349_ _01180_ vssd1 vssd1 vccd1 vccd1 _01559_ sky130_fd_sc_hd__nand2_2
XFILLER_0_109_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_149_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08408_ genblk2\[2\].wave_shpr.div.fin_quo\[0\] genblk2\[2\].wave_shpr.div.fin_quo\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03115_ sky130_fd_sc_hd__or2_1
XFILLER_0_93_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10480__A2 _04715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09388_ net288 _03952_ _03819_ vssd1 vssd1 vccd1 vccd1 _03953_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_124_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08339_ genblk2\[6\].wave_shpr.div.fin_quo\[5\] _02467_ _02742_ vssd1 vssd1 vccd1
+ vccd1 _03046_ sky130_fd_sc_hd__a21o_1
XANTENNA__10328__S _04440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10232__A2 _04454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11350_ genblk2\[7\].wave_shpr.div.acc\[20\] _05334_ vssd1 vssd1 vccd1 vccd1 _05337_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__07633__B1 _01494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10301_ _04567_ _04611_ _04612_ vssd1 vssd1 vccd1 vccd1 _04613_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_61_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11281_ _05187_ _05284_ vssd1 vssd1 vccd1 vccd1 _05285_ sky130_fd_sc_hd__xnor2_1
X_13020_ clknet_leaf_123_clk _00347_ net77 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.i\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10232_ _04418_ _04454_ _04551_ _04457_ net1064 vssd1 vssd1 vccd1 vccd1 _00425_ sky130_fd_sc_hd__a32o_1
XFILLER_0_30_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10163_ _04390_ _04499_ vssd1 vssd1 vccd1 vccd1 _04500_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10940__B1 _05056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08041__B _01576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10094_ net401 _04452_ _04456_ net820 vssd1 vssd1 vccd1 vccd1 _00382_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11999__B1_N _03705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12804_ clknet_leaf_59_clk net496 net188 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.quo\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12445__B1 _03944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10996_ _05055_ _05083_ _05085_ _05057_ net1165 vssd1 vssd1 vccd1 vccd1 _00655_ sky130_fd_sc_hd__a32o_1
XFILLER_0_85_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12735_ clknet_leaf_38_clk genblk1\[10\].osc.clkdiv_C.next_cnt\[12\] net114 vssd1
+ vssd1 vccd1 vccd1 genblk1\[10\].osc.clkdiv_C.cnt\[12\] sky130_fd_sc_hd__dfrtp_2
XTAP_1062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10471__A2 _04715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12666_ clknet_leaf_25_clk genblk1\[6\].osc.clkdiv_C.next_cnt\[15\] net88 vssd1 vssd1
+ vccd1 vccd1 genblk1\[6\].osc.clkdiv_C.cnt\[15\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_154_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12664__RESET_B net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11617_ _05523_ _05405_ vssd1 vssd1 vccd1 vccd1 _05524_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12597_ clknet_leaf_21_clk genblk1\[3\].osc.clkdiv_C.next_cnt\[0\] net97 vssd1 vssd1
+ vccd1 vccd1 genblk1\[3\].osc.clkdiv_C.cnt\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_154_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07120__B _01221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11548_ _03719_ genblk1\[8\].osc.clkdiv_C.cnt\[17\] vssd1 vssd1 vccd1 vccd1 _05472_
+ sky130_fd_sc_hd__or2_1
XANTENNA__07624__B1 _01172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold508 genblk2\[8\].wave_shpr.div.i\[2\] vssd1 vssd1 vccd1 vccd1 net726 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold519 genblk2\[3\].wave_shpr.div.quo\[2\] vssd1 vssd1 vccd1 vccd1 net737 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11479_ _05436_ vssd1 vssd1 vccd1 vccd1 _00787_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13218_ clknet_leaf_5_clk _00541_ net46 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.b1\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08232__A _02225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07927__A1 _01200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13149_ clknet_leaf_121_clk net597 net80 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.quo\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09047__B _02374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09762__S _04039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_868 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_879 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07710_ genblk2\[10\].wave_shpr.div.fin_quo\[7\] _02362_ _02416_ vssd1 vssd1 vccd1
+ vccd1 _02417_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07790__B _01996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08690_ _02798_ _03370_ _03375_ _03396_ vssd1 vssd1 vccd1 vccd1 _03397_ sky130_fd_sc_hd__a31o_1
XANTENNA__06687__A _01576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07641_ _02330_ _02335_ _02343_ _02347_ vssd1 vssd1 vccd1 vccd1 _02348_ sky130_fd_sc_hd__o31ai_4
XFILLER_0_79_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07572_ genblk1\[9\].osc.clkdiv_C.cnt\[5\] _01186_ _01437_ _01225_ vssd1 vssd1 vccd1
+ vccd1 _02279_ sky130_fd_sc_hd__or4_1
XFILLER_0_87_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09311_ net934 _03870_ _03877_ _03896_ vssd1 vssd1 vccd1 vccd1 _00159_ sky130_fd_sc_hd__a22o_1
X_06523_ genblk1\[2\].osc.clkdiv_C.cnt\[10\] _01431_ _01448_ vssd1 vssd1 vccd1 vccd1
+ _01449_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_146_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10937__A _05054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_723 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09852__B2 _04248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09242_ genblk2\[0\].wave_shpr.div.quo\[14\] _03845_ _03847_ net495 _03849_ vssd1
+ vssd1 vccd1 vccd1 _00137_ sky130_fd_sc_hd__a221o_1
XFILLER_0_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06454_ _01374_ _01389_ _01390_ vssd1 vssd1 vccd1 vccd1 _01391_ sky130_fd_sc_hd__and3_1
XFILLER_0_145_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08407__A _02221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09173_ _01342_ _01441_ vssd1 vssd1 vccd1 vccd1 _03813_ sky130_fd_sc_hd__nor2_2
XANTENNA__10148__S _04420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06385_ _01326_ _01328_ vssd1 vssd1 vccd1 vccd1 _01329_ sky130_fd_sc_hd__and2_2
XFILLER_0_44_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08124_ genblk1\[4\].osc.clkdiv_C.cnt\[7\] _01340_ _01304_ genblk1\[4\].osc.clkdiv_C.cnt\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02831_ sky130_fd_sc_hd__a22oi_1
XANTENNA__10214__A2 _04480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_62 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08055_ _01309_ _01180_ genblk1\[5\].osc.clkdiv_C.cnt\[6\] vssd1 vssd1 vccd1 vccd1
+ _02762_ sky130_fd_sc_hd__a21o_1
XANTENNA__07091__A1 genblk1\[8\].osc.clkdiv_C.cnt\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10672__A _04672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xoutput17 net17 vssd1 vssd1 vccd1 vccd1 mode_out[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_141_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07006_ _01823_ _01834_ vssd1 vssd1 vccd1 vccd1 genblk1\[7\].osc.clkdiv_C.next_cnt\[7\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__09238__A _03838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08957_ _03506_ _03566_ vssd1 vssd1 vccd1 vccd1 _03646_ sky130_fd_sc_hd__nor2_1
X_07908_ genblk1\[8\].osc.clkdiv_C.cnt\[10\] _01870_ _02610_ vssd1 vssd1 vccd1 vccd1
+ _02615_ sky130_fd_sc_hd__or3_1
XANTENNA__11478__A1 _01227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08888_ _03582_ _03581_ _03593_ vssd1 vssd1 vccd1 vccd1 _03594_ sky130_fd_sc_hd__nor3_1
X_07839_ _02541_ _02545_ _02529_ _02518_ vssd1 vssd1 vccd1 vccd1 _02546_ sky130_fd_sc_hd__and4b_1
X_10850_ genblk2\[6\].wave_shpr.div.b1\[6\] genblk2\[6\].wave_shpr.div.acc\[6\] vssd1
+ vssd1 vccd1 vccd1 _04994_ sky130_fd_sc_hd__and2b_1
XFILLER_0_67_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09509_ _04044_ vssd1 vssd1 vccd1 vccd1 _04046_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_149_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10781_ _04816_ _04880_ vssd1 vssd1 vccd1 vccd1 _04938_ sky130_fd_sc_hd__or2_1
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12520_ clknet_leaf_104_clk PWM.next_counter\[4\] net157 vssd1 vssd1 vccd1 vccd1
+ PWM.counter\[4\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_581 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12451_ clknet_4_0_0_clk net6 net38 vssd1 vssd1 vccd1 vccd1 modein.delay_in\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_81_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11402_ genblk2\[8\].wave_shpr.div.b1\[2\] genblk2\[8\].wave_shpr.div.acc\[2\] vssd1
+ vssd1 vccd1 vccd1 _05378_ sky130_fd_sc_hd__and2b_1
XFILLER_0_90_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12382_ genblk2\[11\].wave_shpr.div.acc\[8\] _06058_ _06055_ vssd1 vssd1 vccd1 vccd1
+ _06059_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11333_ net1010 _05311_ _05315_ _05324_ vssd1 vssd1 vccd1 vccd1 _00753_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11264_ net540 _05249_ vssd1 vssd1 vccd1 vccd1 _05272_ sky130_fd_sc_hd__or2b_1
XANTENNA__07909__A1 genblk1\[8\].osc.clkdiv_C.cnt\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13003_ clknet_leaf_133_clk _00332_ net59 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.acc\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10215_ _04538_ _04539_ vssd1 vssd1 vccd1 vccd1 _04540_ sky130_fd_sc_hd__nand2_1
X_11195_ net1246 _05236_ _05237_ vssd1 vssd1 vccd1 vccd1 _05238_ sky130_fd_sc_hd__mux2_1
XANTENNA__11181__A3 _02064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10146_ _04384_ _04378_ vssd1 vssd1 vccd1 vccd1 _04487_ sky130_fd_sc_hd__or2b_1
XFILLER_0_118_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06593__B1 _01500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10077_ net667 vssd1 vssd1 vccd1 vccd1 _04449_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_134_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13767_ clknet_leaf_71_clk _01078_ net214 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.acc\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10979_ _05074_ genblk1\[6\].osc.clkdiv_C.cnt\[13\] vssd1 vssd1 vccd1 vccd1 _05075_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_84_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12718_ clknet_leaf_86_clk genblk1\[9\].osc.clkdiv_C.next_cnt\[13\] net181 vssd1
+ vssd1 vccd1 vccd1 genblk1\[9\].osc.clkdiv_C.cnt\[13\] sky130_fd_sc_hd__dfrtp_4
X_13698_ clknet_leaf_94_clk _01009_ net160 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.fin_quo\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_127_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_5_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12649_ clknet_leaf_10_clk genblk1\[5\].osc.clkdiv_C.next_cnt\[16\] net55 vssd1 vssd1
+ vccd1 vccd1 genblk1\[5\].osc.clkdiv_C.cnt\[16\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_111_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06170_ _01119_ _01126_ vssd1 vssd1 vccd1 vccd1 _01142_ sky130_fd_sc_hd__xor2_1
XFILLER_0_87_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold305 genblk2\[6\].wave_shpr.div.quo\[7\] vssd1 vssd1 vccd1 vccd1 net523 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold316 genblk2\[7\].wave_shpr.div.quo\[24\] vssd1 vssd1 vccd1 vccd1 net534 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_472 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold327 genblk2\[3\].wave_shpr.div.quo\[20\] vssd1 vssd1 vccd1 vccd1 net545 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_7_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold338 genblk2\[9\].wave_shpr.div.acc\[21\] vssd1 vssd1 vccd1 vccd1 net556 sky130_fd_sc_hd__dlygate4sd3_1
Xhold349 genblk2\[6\].wave_shpr.div.quo\[20\] vssd1 vssd1 vccd1 vccd1 net567 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09058__A _02170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13633__RESET_B net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09860_ genblk2\[2\].wave_shpr.div.acc\[2\] _04284_ _04214_ vssd1 vssd1 vccd1 vccd1
+ _04285_ sky130_fd_sc_hd__mux2_1
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08811_ _03512_ _03516_ _03223_ _03509_ vssd1 vssd1 vccd1 vccd1 _03518_ sky130_fd_sc_hd__a211o_1
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09791_ _03833_ net1190 vssd1 vssd1 vccd1 vccd1 _04246_ sky130_fd_sc_hd__and2_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1005 genblk2\[5\].wave_shpr.div.b1\[17\] vssd1 vssd1 vccd1 vccd1 net1223 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1016 genblk2\[7\].wave_shpr.div.b1\[17\] vssd1 vssd1 vccd1 vccd1 net1234 sky130_fd_sc_hd__dlygate4sd3_1
X_08742_ _03445_ _03446_ _03447_ _03448_ vssd1 vssd1 vccd1 vccd1 _03449_ sky130_fd_sc_hd__o211a_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1027 genblk2\[3\].wave_shpr.div.b1\[4\] vssd1 vssd1 vccd1 vccd1 net1245 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1038 genblk1\[2\].osc.clkdiv_C.cnt\[12\] vssd1 vssd1 vccd1 vccd1 net1256 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1049 genblk2\[1\].wave_shpr.div.b1\[4\] vssd1 vssd1 vccd1 vccd1 net1267 sky130_fd_sc_hd__dlygate4sd3_1
X_08673_ _03357_ _03358_ _03334_ _03335_ vssd1 vssd1 vccd1 vccd1 _03380_ sky130_fd_sc_hd__o211a_1
XFILLER_0_108_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06210__A _01171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout174_A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07624_ genblk1\[11\].osc.clkdiv_C.cnt\[14\] _02085_ _01172_ vssd1 vssd1 vccd1 vccd1
+ _02331_ sky130_fd_sc_hd__o21a_1
XTAP_1809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12586__RESET_B net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07555_ genblk2\[9\].wave_shpr.div.fin_quo\[0\] genblk2\[9\].wave_shpr.div.fin_quo\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02262_ sky130_fd_sc_hd__or2_1
X_06506_ _01230_ vssd1 vssd1 vccd1 vccd1 _01432_ sky130_fd_sc_hd__buf_8
XFILLER_0_118_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07836__B1 _02261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07486_ genblk2\[11\].wave_shpr.div.i\[2\] genblk2\[11\].wave_shpr.div.i\[3\] genblk2\[11\].wave_shpr.div.i\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02210_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_76_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09225_ net269 _03836_ _03840_ net652 vssd1 vssd1 vccd1 vccd1 _00129_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07041__A _01439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06437_ genblk1\[1\].osc.clkdiv_C.cnt\[1\] genblk1\[1\].osc.clkdiv_C.cnt\[0\] genblk1\[1\].osc.clkdiv_C.cnt\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01379_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_106_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09156_ _03803_ vssd1 vssd1 vccd1 vccd1 _03804_ sky130_fd_sc_hd__buf_4
X_06368_ _01309_ _01221_ vssd1 vssd1 vccd1 vccd1 _01312_ sky130_fd_sc_hd__and2_2
X_08107_ _01192_ _01208_ _01588_ vssd1 vssd1 vccd1 vccd1 _02814_ sky130_fd_sc_hd__a21oi_1
X_09087_ modein.delay_octave_up_in\[1\] modein.delay_octave_up_in\[0\] vssd1 vssd1
+ vccd1 vccd1 _03738_ sky130_fd_sc_hd__and2b_1
XANTENNA__10606__S _00015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_110_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_110_clk
+ sky130_fd_sc_hd__clkbuf_16
X_06299_ _01176_ _01178_ _01194_ vssd1 vssd1 vccd1 vccd1 _01261_ sky130_fd_sc_hd__mux2_1
XFILLER_0_4_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08038_ net12 _02744_ _02365_ vssd1 vssd1 vccd1 vccd1 _02745_ sky130_fd_sc_hd__and3_2
Xhold850 genblk2\[4\].wave_shpr.div.acc\[3\] vssd1 vssd1 vccd1 vccd1 net1068 sky130_fd_sc_hd__dlygate4sd3_1
Xhold861 genblk2\[3\].wave_shpr.div.i\[1\] vssd1 vssd1 vccd1 vccd1 net1079 sky130_fd_sc_hd__dlygate4sd3_1
Xhold872 genblk2\[10\].wave_shpr.div.i\[1\] vssd1 vssd1 vccd1 vccd1 net1090 sky130_fd_sc_hd__dlygate4sd3_1
Xhold883 genblk1\[3\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 net1101 sky130_fd_sc_hd__dlygate4sd3_1
Xhold894 _02252_ vssd1 vssd1 vccd1 vccd1 net1112 sky130_fd_sc_hd__dlygate4sd3_1
X_10000_ _04370_ _04394_ _04395_ vssd1 vssd1 vccd1 vccd1 _04396_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout87_A net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09989_ _04378_ _04383_ _04384_ vssd1 vssd1 vccd1 vccd1 _04385_ sky130_fd_sc_hd__a21o_1
XANTENNA__09513__B1 _04047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11951_ _05735_ _05771_ _05772_ vssd1 vssd1 vccd1 vccd1 _05773_ sky130_fd_sc_hd__a21o_1
XANTENNA__11320__B1 _05283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10902_ net1250 _01923_ _04848_ vssd1 vssd1 vccd1 vccd1 _05035_ sky130_fd_sc_hd__mux2_1
X_11882_ _05610_ _05611_ vssd1 vssd1 vccd1 vccd1 _05713_ sky130_fd_sc_hd__and2b_1
X_10833_ genblk2\[6\].wave_shpr.div.acc\[6\] genblk2\[6\].wave_shpr.div.b1\[6\] vssd1
+ vssd1 vccd1 vccd1 _04977_ sky130_fd_sc_hd__or2b_1
X_13621_ clknet_leaf_74_clk _00934_ net212 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.b1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10764_ net902 _04918_ _04922_ _04925_ vssd1 vssd1 vccd1 vccd1 _00583_ sky130_fd_sc_hd__a22o_1
X_13552_ clknet_leaf_100_clk net650 net165 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.quo\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12503_ clknet_leaf_106_clk _00065_ net154 vssd1 vssd1 vccd1 vccd1 PWM.final_in\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_13483_ clknet_leaf_99_clk _00800_ net168 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10695_ _04869_ genblk1\[5\].osc.clkdiv_C.cnt\[13\] vssd1 vssd1 vccd1 vccd1 _04875_
+ sky130_fd_sc_hd__and2_1
X_12434_ net955 _06072_ _06073_ _06097_ vssd1 vssd1 vccd1 vccd1 _01081_ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12365_ genblk2\[11\].wave_shpr.div.acc\[4\] _06045_ _05982_ vssd1 vssd1 vccd1 vccd1
+ _06046_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_101_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_101_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_105_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11316_ _05245_ vssd1 vssd1 vccd1 vccd1 _05311_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12296_ _03687_ net409 _03735_ vssd1 vssd1 vccd1 vccd1 _01032_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_10_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11247_ genblk2\[7\].wave_shpr.div.quo\[17\] _05255_ _05256_ net548 _05263_ vssd1
+ vssd1 vccd1 vccd1 _00728_ sky130_fd_sc_hd__a221o_1
XFILLER_0_129_37 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11178_ net1216 vssd1 vssd1 vccd1 vccd1 _00692_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10362__A1 _03726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10129_ net490 _04451_ _04455_ net529 _04475_ vssd1 vssd1 vccd1 vccd1 _00398_ sky130_fd_sc_hd__a221o_1
XANTENNA__12032__A _02155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07678__A2_N _01215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11311__B1 _05283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06965__A _01213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09807__A1 genblk2\[2\].wave_shpr.div.quo\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07340_ genblk1\[11\].osc.clkdiv_C.cnt\[3\] _02097_ vssd1 vssd1 vccd1 vccd1 _02101_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_128_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07271_ _02045_ vssd1 vssd1 vccd1 vccd1 genblk1\[10\].osc.clkdiv_C.next_cnt\[7\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09010_ net1128 sig_norm.quo\[6\] _01154_ vssd1 vssd1 vccd1 vccd1 _03685_ sky130_fd_sc_hd__mux2_1
X_06222_ _01172_ _01180_ _01183_ vssd1 vssd1 vccd1 vccd1 _01184_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_115_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06153_ net3 _01100_ _01101_ vssd1 vssd1 vccd1 vccd1 _01125_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_131_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold102 genblk2\[10\].wave_shpr.div.quo\[7\] vssd1 vssd1 vccd1 vccd1 net320 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold113 genblk2\[7\].wave_shpr.div.quo\[3\] vssd1 vssd1 vccd1 vccd1 net331 sky130_fd_sc_hd__dlygate4sd3_1
Xhold124 genblk2\[11\].wave_shpr.div.quo\[13\] vssd1 vssd1 vccd1 vccd1 net342 sky130_fd_sc_hd__dlygate4sd3_1
Xhold135 genblk2\[10\].wave_shpr.div.quo\[16\] vssd1 vssd1 vccd1 vccd1 net353 sky130_fd_sc_hd__dlygate4sd3_1
Xhold146 smpl_rt_clkdiv.clkDiv_inst.cnt\[1\] vssd1 vssd1 vccd1 vccd1 net364 sky130_fd_sc_hd__dlygate4sd3_1
Xhold157 genblk2\[3\].wave_shpr.div.acc\[26\] vssd1 vssd1 vccd1 vccd1 net375 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold168 _00651_ vssd1 vssd1 vccd1 vccd1 net386 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09912_ genblk2\[2\].wave_shpr.div.acc\[14\] _04324_ _04301_ vssd1 vssd1 vccd1 vccd1
+ _04325_ sky130_fd_sc_hd__mux2_1
Xhold179 genblk2\[11\].wave_shpr.div.quo\[6\] vssd1 vssd1 vccd1 vccd1 net397 sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09843_ _04269_ genblk1\[2\].osc.clkdiv_C.cnt\[15\] vssd1 vssd1 vccd1 vccd1 _04273_
+ sky130_fd_sc_hd__and2_1
XANTENNA__11765__B genblk1\[9\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09774_ _03831_ net614 _03733_ vssd1 vssd1 vccd1 vccd1 _00282_ sky130_fd_sc_hd__a21bo_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06986_ genblk1\[7\].osc.clkdiv_C.cnt\[2\] _01227_ _01793_ _01821_ vssd1 vssd1 vccd1
+ vccd1 _01822_ sky130_fd_sc_hd__o211a_2
X_08725_ _03399_ _03398_ vssd1 vssd1 vccd1 vccd1 _03432_ sky130_fd_sc_hd__and2b_1
XTAP_2307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08656_ _03188_ _03189_ _02885_ vssd1 vssd1 vccd1 vccd1 _03363_ sky130_fd_sc_hd__a21o_1
XTAP_2329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_54_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07607_ _02313_ vssd1 vssd1 vccd1 vccd1 _02314_ sky130_fd_sc_hd__buf_2
XTAP_1628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08587_ _03237_ _03239_ _03243_ vssd1 vssd1 vccd1 vccd1 _03294_ sky130_fd_sc_hd__a21bo_1
XANTENNA__10397__A _04477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07538_ net1112 vssd1 vssd1 vccd1 vccd1 _00030_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_687 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_134 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07469_ _02198_ vssd1 vssd1 vccd1 vccd1 _00020_ sky130_fd_sc_hd__inv_2
XFILLER_0_91_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_69_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09208_ net959 vssd1 vssd1 vccd1 vccd1 _03832_ sky130_fd_sc_hd__inv_2
XFILLER_0_63_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10480_ net850 _04715_ _04722_ _04725_ vssd1 vssd1 vccd1 vccd1 _00499_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_112_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09139_ genblk2\[0\].wave_shpr.div.b1\[12\] genblk2\[0\].wave_shpr.div.acc\[12\]
+ vssd1 vssd1 vccd1 vccd1 _03787_ sky130_fd_sc_hd__and2b_1
XFILLER_0_134_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10336__S _04440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12030__A1 genblk2\[10\].wave_shpr.div.quo\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12150_ _05781_ _05899_ genblk2\[10\].wave_shpr.div.acc\[18\] vssd1 vssd1 vccd1 vccd1
+ _05901_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_60_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11101_ _03690_ _05161_ _05162_ vssd1 vssd1 vccd1 vccd1 _00683_ sky130_fd_sc_hd__nor3_1
XFILLER_0_130_773 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12081_ _05749_ _05847_ vssd1 vssd1 vccd1 vccd1 _05848_ sky130_fd_sc_hd__xnor2_1
XANTENNA_clkbuf_leaf_127_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold680 genblk2\[8\].wave_shpr.div.acc\[5\] vssd1 vssd1 vccd1 vccd1 net898 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_5_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold691 genblk2\[8\].wave_shpr.div.acc\[12\] vssd1 vssd1 vccd1 vccd1 net909 sky130_fd_sc_hd__dlygate4sd3_1
X_11032_ _05002_ _04973_ vssd1 vssd1 vccd1 vccd1 _05113_ sky130_fd_sc_hd__or2b_1
XANTENNA__10071__S _04440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09860__S _04214_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12983_ clknet_leaf_125_clk _00312_ net69 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.quo\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_11934_ genblk2\[10\].wave_shpr.div.b1\[5\] genblk2\[10\].wave_shpr.div.acc\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05756_ sky130_fd_sc_hd__and2b_1
XTAP_2830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11865_ _05606_ _05554_ vssd1 vssd1 vccd1 vccd1 _05701_ sky130_fd_sc_hd__or2b_1
X_13604_ clknet_leaf_97_clk _00003_ net166 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.done
+ sky130_fd_sc_hd__dfrtp_1
X_10816_ genblk2\[5\].wave_shpr.div.i\[1\] genblk2\[5\].wave_shpr.div.i\[0\] genblk2\[5\].wave_shpr.div.i\[2\]
+ genblk2\[5\].wave_shpr.div.i\[3\] vssd1 vssd1 vccd1 vccd1 _04962_ sky130_fd_sc_hd__and4_1
XFILLER_0_95_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11796_ _03694_ _05647_ _05648_ _03696_ net1059 vssd1 vssd1 vccd1 vccd1 _00892_ sky130_fd_sc_hd__a32o_1
XFILLER_0_54_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13535_ clknet_leaf_81_clk _00850_ net199 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.i\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10747_ _04800_ _04770_ vssd1 vssd1 vccd1 vccd1 _04912_ sky130_fd_sc_hd__or2b_1
XFILLER_0_54_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10678_ _04672_ genblk1\[5\].osc.clkdiv_C.cnt\[5\] vssd1 vssd1 vccd1 vccd1 _04866_
+ sky130_fd_sc_hd__and2_1
X_13466_ clknet_leaf_75_clk _00783_ net203 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.b1\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_36_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12021__A1 genblk2\[10\].wave_shpr.div.quo\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12417_ _05975_ _05925_ vssd1 vssd1 vccd1 vccd1 _06085_ sky130_fd_sc_hd__or2b_1
XANTENNA__12021__B2 _05816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13397_ clknet_leaf_117_clk net662 net140 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12348_ _03944_ _06031_ _06032_ _03947_ net1044 vssd1 vssd1 vccd1 vccd1 _01060_ sky130_fd_sc_hd__a32o_1
XFILLER_0_121_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12279_ _01308_ genblk2\[1\].wave_shpr.div.b1\[8\] _03719_ vssd1 vssd1 vccd1 vccd1
+ _06001_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06840_ genblk1\[5\].osc.clkdiv_C.cnt\[6\] _01703_ vssd1 vssd1 vccd1 vccd1 _01706_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__09770__S _04039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06771_ genblk1\[4\].osc.clkdiv_C.cnt\[14\] genblk1\[4\].osc.clkdiv_C.cnt\[13\] _01641_
+ vssd1 vssd1 vccd1 vccd1 _01647_ sky130_fd_sc_hd__and3_1
X_08510_ _03204_ _03205_ _03216_ vssd1 vssd1 vccd1 vccd1 _03217_ sky130_fd_sc_hd__nor3b_2
XANTENNA__11805__S _05613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09490_ genblk2\[2\].wave_shpr.div.b1\[11\] _04034_ _04024_ vssd1 vssd1 vccd1 vccd1
+ _04035_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08441_ _02525_ _03146_ _03147_ _02361_ genblk2\[10\].wave_shpr.div.fin_quo\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03148_ sky130_fd_sc_hd__a32o_1
XFILLER_0_93_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08372_ _03055_ _03077_ _03001_ _03078_ vssd1 vssd1 vccd1 vccd1 _03079_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_46_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07323_ genblk1\[11\].osc.clkdiv_C.cnt\[3\] _01334_ _01321_ genblk1\[11\].osc.clkdiv_C.cnt\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02087_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_73_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_85_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout137_A net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07254_ _02027_ _02032_ _02033_ vssd1 vssd1 vccd1 vccd1 genblk1\[10\].osc.clkdiv_C.next_cnt\[2\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_155_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08415__A net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06205_ _01168_ vssd1 vssd1 vccd1 vccd1 PWM.next_counter\[6\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10156__S _04420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07185_ _01953_ _01974_ _01975_ vssd1 vssd1 vccd1 vccd1 genblk1\[9\].osc.clkdiv_C.next_cnt\[9\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_143_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06136_ net1 net7 vssd1 vssd1 vccd1 vccd1 _01108_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10680__A _04676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09192__A1 _02002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09826_ genblk2\[2\].wave_shpr.div.quo\[16\] _04257_ _04259_ net315 _04263_ vssd1
+ vssd1 vccd1 vccd1 _00307_ sky130_fd_sc_hd__a221o_1
X_09757_ _01496_ vssd1 vssd1 vccd1 vccd1 _04227_ sky130_fd_sc_hd__inv_2
X_06969_ _01179_ _01233_ vssd1 vssd1 vccd1 vccd1 _01805_ sky130_fd_sc_hd__or2_2
XTAP_2104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08708_ _03413_ _03414_ genblk2\[2\].wave_shpr.div.fin_quo\[4\] _02468_ vssd1 vssd1
+ vccd1 vccd1 _03415_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_69_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12400__A _03942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09688_ genblk2\[2\].wave_shpr.div.acc\[5\] genblk2\[2\].wave_shpr.div.b1\[5\] vssd1
+ vssd1 vccd1 vccd1 _04168_ sky130_fd_sc_hd__or2b_1
XTAP_2137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08639_ _02685_ _02681_ _02686_ _02526_ vssd1 vssd1 vccd1 vccd1 _03346_ sky130_fd_sc_hd__o31a_1
XTAP_1425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08309__B _02361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11650_ genblk2\[8\].wave_shpr.div.i\[1\] genblk2\[8\].wave_shpr.div.i\[0\] vssd1
+ vssd1 vccd1 vccd1 _05546_ sky130_fd_sc_hd__or2_1
XTAP_1469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout41 net43 vssd1 vssd1 vccd1 vccd1 net41 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10601_ _04825_ vssd1 vssd1 vccd1 vccd1 _00520_ sky130_fd_sc_hd__clkbuf_1
Xfanout52 net53 vssd1 vssd1 vccd1 vccd1 net52 sky130_fd_sc_hd__clkbuf_4
Xfanout63 net85 vssd1 vssd1 vccd1 vccd1 net63 sky130_fd_sc_hd__buf_2
X_11581_ genblk2\[8\].wave_shpr.div.acc\[7\] _05496_ _05493_ vssd1 vssd1 vccd1 vccd1
+ _05497_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_454 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout74 net75 vssd1 vssd1 vccd1 vccd1 net74 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_80_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_135_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout85 net16 vssd1 vssd1 vccd1 vccd1 net85 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10532_ _03690_ _04760_ _04761_ vssd1 vssd1 vccd1 vccd1 _00515_ sky130_fd_sc_hd__nor3_1
XFILLER_0_52_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13320_ clknet_leaf_26_clk net499 net87 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.quo\[14\]
+ sky130_fd_sc_hd__dfrtp_1
Xfanout96 net98 vssd1 vssd1 vccd1 vccd1 net96 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_135_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13251_ clknet_leaf_2_clk _00574_ net41 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.acc\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10463_ _04602_ _04572_ vssd1 vssd1 vccd1 vccd1 _04712_ sky130_fd_sc_hd__or2b_1
XANTENNA__10066__S _04440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09955__B1 _04253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12202_ genblk2\[11\].wave_shpr.div.b1\[2\] vssd1 vssd1 vccd1 vccd1 _05940_ sky130_fd_sc_hd__inv_2
X_13182_ clknet_leaf_130_clk net473 net129 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.acc\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_682 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10394_ net596 _04661_ _04663_ net637 _04665_ vssd1 vssd1 vccd1 vccd1 _00473_ sky130_fd_sc_hd__a221o_1
X_12133_ _05773_ _05887_ vssd1 vssd1 vccd1 vccd1 _05888_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08979__B _01157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12306__A2 _06009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12064_ _03833_ _01995_ vssd1 vssd1 vccd1 vccd1 _05837_ sky130_fd_sc_hd__nor2_1
X_11015_ _04994_ _04977_ vssd1 vssd1 vccd1 vccd1 _05100_ sky130_fd_sc_hd__or2b_1
XFILLER_0_126_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12966_ clknet_leaf_111_clk net337 net130 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.quo\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_11917_ genblk2\[10\].wave_shpr.div.acc\[9\] genblk2\[10\].wave_shpr.div.b1\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05739_ sky130_fd_sc_hd__or2b_1
XTAP_2660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12897_ clknet_leaf_31_clk net258 net99 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.quo\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07123__B _01344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11848_ net967 _05684_ _05685_ _05688_ vssd1 vssd1 vccd1 vccd1 _00904_ sky130_fd_sc_hd__a22o_1
XTAP_1970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11779_ _05631_ genblk1\[9\].osc.clkdiv_C.cnt\[11\] vssd1 vssd1 vccd1 vccd1 _05639_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_144_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06962__B _01797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13518_ clknet_leaf_78_clk _00835_ net206 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.acc\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_126 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13449_ clknet_leaf_91_clk _00766_ net144 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.i\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_340 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08749__A1 genblk2\[8\].wave_shpr.div.fin_quo\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__09946__B1 _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11753__B1 _05624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08990_ net1261 _03673_ _01158_ vssd1 vssd1 vccd1 vccd1 _03674_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07941_ _02646_ _02647_ vssd1 vssd1 vccd1 vccd1 _02648_ sky130_fd_sc_hd__nor2_2
XFILLER_0_76_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09174__A1 _03813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07872_ _02469_ _02578_ _02529_ vssd1 vssd1 vccd1 vccd1 _02579_ sky130_fd_sc_hd__o21a_1
XANTENNA__07724__A2 _01323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09611_ _03994_ _03959_ vssd1 vssd1 vccd1 vccd1 _04110_ sky130_fd_sc_hd__or2b_1
X_06823_ net1355 vssd1 vssd1 vccd1 vccd1 _01694_ sky130_fd_sc_hd__inv_2
X_06754_ _01634_ vssd1 vssd1 vccd1 vccd1 genblk1\[4\].osc.clkdiv_C.next_cnt\[9\] sky130_fd_sc_hd__clkbuf_1
X_09542_ _04055_ genblk1\[1\].osc.clkdiv_C.cnt\[9\] vssd1 vssd1 vccd1 vccd1 _04062_
+ sky130_fd_sc_hd__and2_1
X_09473_ genblk2\[2\].wave_shpr.div.b1\[4\] _04023_ _04024_ vssd1 vssd1 vccd1 vccd1
+ _04025_ sky130_fd_sc_hd__mux2_1
X_06685_ _01194_ _01175_ _01191_ vssd1 vssd1 vccd1 vccd1 _01575_ sky130_fd_sc_hd__or3_1
Xclkbuf_leaf_90_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_90_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_93_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08424_ _03083_ _03124_ _03130_ vssd1 vssd1 vccd1 vccd1 _03131_ sky130_fd_sc_hd__o21a_1
XFILLER_0_148_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08355_ genblk2\[4\].wave_shpr.div.fin_quo\[4\] _02932_ _02841_ _02222_ vssd1 vssd1
+ vccd1 vccd1 _03062_ sky130_fd_sc_hd__a31o_1
XFILLER_0_129_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08437__B1 _02361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07306_ _01223_ _01678_ genblk1\[11\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1
+ _02070_ sky130_fd_sc_hd__o21ai_1
X_08286_ _02964_ _02958_ _02963_ vssd1 vssd1 vccd1 vccd1 _02993_ sky130_fd_sc_hd__nand3_1
XFILLER_0_61_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07237_ _01242_ _02015_ _02017_ _01197_ _02018_ vssd1 vssd1 vccd1 vccd1 _02019_ sky130_fd_sc_hd__o221a_1
XFILLER_0_143_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07168_ _01954_ _01962_ _01963_ vssd1 vssd1 vccd1 vccd1 _01964_ sky130_fd_sc_hd__and3_1
XFILLER_0_131_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06119_ net365 _01088_ vssd1 vssd1 vccd1 vccd1 smpl_rt_clkdiv.clkDiv_inst.next_cnt\[6\]
+ sky130_fd_sc_hd__xor2_1
X_07099_ genblk1\[8\].osc.clkdiv_C.cnt\[11\] _01904_ vssd1 vssd1 vccd1 vccd1 _01906_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_100_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09809_ _04069_ genblk1\[2\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 _04254_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_97_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12820_ clknet_leaf_66_clk _00153_ net196 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.acc\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12751_ clknet_leaf_50_clk genblk1\[11\].osc.clkdiv_C.next_cnt\[10\] net111 vssd1
+ vssd1 vccd1 vccd1 genblk1\[11\].osc.clkdiv_C.cnt\[10\] sky130_fd_sc_hd__dfrtp_2
XTAP_1222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_81_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_81_clk sky130_fd_sc_hd__clkbuf_16
XTAP_1244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11702_ genblk2\[9\].wave_shpr.div.b1\[11\] genblk2\[9\].wave_shpr.div.acc\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05594_ sky130_fd_sc_hd__and2b_1
XTAP_1255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12682_ clknet_leaf_120_clk genblk1\[7\].osc.clkdiv_C.next_cnt\[13\] net81 vssd1
+ vssd1 vccd1 vccd1 genblk1\[7\].osc.clkdiv_C.cnt\[13\] sky130_fd_sc_hd__dfrtp_4
XTAP_1277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11633_ net1018 _05507_ _05445_ _05535_ vssd1 vssd1 vccd1 vccd1 _00842_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11564_ net980 _05447_ _05446_ _05483_ vssd1 vssd1 vccd1 vccd1 _00825_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11983__B1 _05796_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13303_ clknet_leaf_87_clk _00624_ net201 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.b1\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10515_ genblk2\[4\].wave_shpr.div.acc\[24\] vssd1 vssd1 vccd1 vccd1 _04750_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11495_ _05444_ vssd1 vssd1 vccd1 vccd1 _05445_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_150_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10446_ _04594_ _04576_ vssd1 vssd1 vccd1 vccd1 _04699_ sky130_fd_sc_hd__or2b_1
X_13234_ clknet_leaf_16_clk net295 net73 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.quo\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13165_ clknet_leaf_127_clk _00490_ net68 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.acc\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10377_ net508 _04652_ _04656_ net781 vssd1 vssd1 vccd1 vccd1 _00465_ sky130_fd_sc_hd__a22o_1
XANTENNA__11204__A1_N _03727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12116_ genblk2\[10\].wave_shpr.div.acc\[10\] _05874_ _05865_ vssd1 vssd1 vccd1 vccd1
+ _05875_ sky130_fd_sc_hd__mux2_1
X_13096_ clknet_leaf_137_clk _00423_ net41 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.acc\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12452__RESET_B net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12047_ _05819_ genblk1\[10\].osc.clkdiv_C.cnt\[6\] vssd1 vssd1 vccd1 vccd1 _05828_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_1_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12949_ clknet_leaf_121_clk _00278_ net77 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.b1\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_72_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_72_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_141_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06470_ genblk1\[1\].osc.clkdiv_C.cnt\[13\] genblk1\[1\].osc.clkdiv_C.cnt\[12\] _01398_
+ vssd1 vssd1 vccd1 vccd1 _01401_ sky130_fd_sc_hd__and3_1
XFILLER_0_146_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_62_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07890__B2 _02592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08140_ _02838_ _02845_ _02846_ vssd1 vssd1 vccd1 vccd1 _02847_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_43_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08071_ _02772_ _02774_ _02776_ _02777_ vssd1 vssd1 vccd1 vccd1 _02778_ sky130_fd_sc_hd__o31a_1
XFILLER_0_125_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07022_ genblk1\[7\].osc.clkdiv_C.cnt\[13\] _01842_ _01844_ vssd1 vssd1 vccd1 vccd1
+ genblk1\[7\].osc.clkdiv_C.next_cnt\[13\] sky130_fd_sc_hd__o21a_1
XFILLER_0_102_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06609__A2_N _01514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10529__A1 _04655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08973_ net1300 _03659_ _01158_ vssd1 vssd1 vccd1 vccd1 _03660_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold17 genblk2\[5\].wave_shpr.div.quo\[17\] vssd1 vssd1 vccd1 vccd1 net235 sky130_fd_sc_hd__dlygate4sd3_1
Xhold28 _00565_ vssd1 vssd1 vccd1 vccd1 net246 sky130_fd_sc_hd__dlygate4sd3_1
X_07924_ _02609_ _02613_ _02630_ _02614_ vssd1 vssd1 vccd1 vccd1 _02631_ sky130_fd_sc_hd__or4b_1
Xhold39 genblk2\[1\].wave_shpr.div.quo\[20\] vssd1 vssd1 vccd1 vccd1 net257 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09524__A _03853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07855_ _02509_ _02551_ _02554_ _02560_ _02518_ vssd1 vssd1 vccd1 vccd1 _02562_ sky130_fd_sc_hd__o311a_1
X_06806_ _01336_ _01564_ vssd1 vssd1 vccd1 vccd1 _01678_ sky130_fd_sc_hd__nor2_4
X_07786_ genblk1\[0\].osc.clkdiv_C.cnt\[8\] _01193_ _01184_ genblk1\[0\].osc.clkdiv_C.cnt\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02493_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_79_866 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09525_ net645 _04048_ _04045_ net610 _04051_ vssd1 vssd1 vccd1 vccd1 _00218_ sky130_fd_sc_hd__a221o_1
XFILLER_0_149_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11257__A2 _05245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06737_ _01620_ vssd1 vssd1 vccd1 vccd1 _01621_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_63_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_63_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__08122__A2 _01340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07979__A genblk2\[7\].wave_shpr.div.fin_quo\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_78_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09456_ genblk2\[1\].wave_shpr.div.fin_quo\[4\] net1316 _00007_ vssd1 vssd1 vccd1
+ vccd1 _04016_ sky130_fd_sc_hd__mux2_1
X_06668_ genblk1\[4\].osc.clkdiv_C.cnt\[6\] _01557_ vssd1 vssd1 vccd1 vccd1 _01558_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_148_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08407_ _02221_ _03113_ vssd1 vssd1 vccd1 vccd1 _03114_ sky130_fd_sc_hd__nor2_2
X_06599_ _01441_ _01249_ vssd1 vssd1 vccd1 vccd1 _01507_ sky130_fd_sc_hd__nor2_2
X_09387_ _03726_ _03951_ _03952_ vssd1 vssd1 vccd1 vccd1 _00179_ sky130_fd_sc_hd__nor3_1
XFILLER_0_47_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_136_459 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08338_ _03043_ _03044_ vssd1 vssd1 vccd1 vccd1 _03045_ sky130_fd_sc_hd__nor2_1
XFILLER_0_117_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_871 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08269_ _02973_ _02974_ _02975_ _02360_ vssd1 vssd1 vccd1 vccd1 _02976_ sky130_fd_sc_hd__o211a_1
X_10300_ genblk2\[4\].wave_shpr.div.b1\[15\] genblk2\[4\].wave_shpr.div.acc\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04612_ sky130_fd_sc_hd__and2b_1
XFILLER_0_62_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_868 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11280_ _05188_ _05180_ vssd1 vssd1 vccd1 vccd1 _05284_ sky130_fd_sc_hd__or2b_1
X_10231_ _04549_ _04550_ vssd1 vssd1 vccd1 vccd1 _04551_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10162_ _04391_ _04372_ vssd1 vssd1 vccd1 vccd1 _04499_ sky130_fd_sc_hd__or2b_1
XANTENNA__10940__B2 net792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10093_ genblk2\[3\].wave_shpr.div.quo\[6\] _04452_ _04456_ net814 vssd1 vssd1 vccd1
+ vccd1 _00381_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06496__C _01327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12803_ clknet_leaf_59_clk _00136_ net188 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.quo\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10995_ _05023_ _05084_ vssd1 vssd1 vccd1 vccd1 _05085_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_54_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_54_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__08113__A2 _01323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12734_ clknet_leaf_38_clk genblk1\[10\].osc.clkdiv_C.next_cnt\[11\] net113 vssd1
+ vssd1 vccd1 vccd1 genblk1\[10\].osc.clkdiv_C.cnt\[11\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_32_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_123_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12665_ clknet_leaf_25_clk genblk1\[6\].osc.clkdiv_C.next_cnt\[14\] net86 vssd1 vssd1
+ vccd1 vccd1 genblk1\[6\].osc.clkdiv_C.cnt\[14\] sky130_fd_sc_hd__dfrtp_4
XTAP_1096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11616_ _05406_ _05359_ vssd1 vssd1 vccd1 vccd1 _05523_ sky130_fd_sc_hd__or2b_1
XFILLER_0_65_593 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12596_ clknet_leaf_15_clk genblk1\[2\].osc.clkdiv_C.next_cnt\[17\] net73 vssd1 vssd1
+ vccd1 vccd1 genblk1\[2\].osc.clkdiv_C.cnt\[17\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_80_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11547_ _05444_ vssd1 vssd1 vccd1 vccd1 _05471_ sky130_fd_sc_hd__inv_2
Xhold509 genblk2\[0\].wave_shpr.div.b1\[5\] vssd1 vssd1 vccd1 vccd1 net727 sky130_fd_sc_hd__dlygate4sd3_1
X_11478_ net1231 _01227_ _05433_ vssd1 vssd1 vccd1 vccd1 _05436_ sky130_fd_sc_hd__mux2_1
XFILLER_0_111_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12633__RESET_B net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13217_ clknet_leaf_6_clk _00540_ net48 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.b1\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10429_ net937 _04683_ _04656_ _04686_ vssd1 vssd1 vccd1 vccd1 _00487_ sky130_fd_sc_hd__a22o_1
XFILLER_0_110_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08232__B _02885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07927__A2 genblk1\[8\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13148_ clknet_leaf_121_clk _00473_ net81 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.quo\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13079_ clknet_leaf_125_clk _00406_ net61 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.acc\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_869 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07790__C _01801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08352__A2 _02521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07640_ _02335_ _02344_ _02345_ _02346_ vssd1 vssd1 vccd1 vccd1 _02347_ sky130_fd_sc_hd__o211a_1
XFILLER_0_88_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07560__B1 _01328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07571_ genblk1\[9\].osc.clkdiv_C.cnt\[4\] _01186_ _01355_ vssd1 vssd1 vccd1 vccd1
+ _02278_ sky130_fd_sc_hd__or3_1
XANTENNA__08104__A2 _01323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_45_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_45_clk sky130_fd_sc_hd__clkbuf_16
X_09310_ genblk2\[0\].wave_shpr.div.acc\[9\] _03895_ _03889_ vssd1 vssd1 vccd1 vccd1
+ _03896_ sky130_fd_sc_hd__mux2_1
X_06522_ genblk1\[2\].osc.clkdiv_C.cnt\[10\] _01431_ _01447_ vssd1 vssd1 vccd1 vccd1
+ _01448_ sky130_fd_sc_hd__o21bai_1
XANTENNA__07312__B1 _01578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06453_ genblk1\[1\].osc.clkdiv_C.cnt\[7\] _01387_ vssd1 vssd1 vccd1 vccd1 _01390_
+ sky130_fd_sc_hd__or2_1
X_09241_ _03725_ genblk1\[0\].osc.clkdiv_C.cnt\[5\] vssd1 vssd1 vccd1 vccd1 _03849_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_146_735 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06666__A2 _01221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09172_ net1219 vssd1 vssd1 vccd1 vccd1 _00104_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06384_ _01186_ _01327_ vssd1 vssd1 vccd1 vccd1 _01328_ sky130_fd_sc_hd__nor2_4
XFILLER_0_7_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08123_ genblk1\[4\].osc.clkdiv_C.cnt\[5\] _01224_ _01249_ _01565_ genblk1\[4\].osc.clkdiv_C.cnt\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02830_ sky130_fd_sc_hd__o32a_1
XFILLER_0_32_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout217_A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08054_ genblk1\[5\].osc.clkdiv_C.cnt\[7\] _01223_ vssd1 vssd1 vccd1 vccd1 _02761_
+ sky130_fd_sc_hd__or2_1
XANTENNA__09519__A _04042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07005_ genblk1\[7\].osc.clkdiv_C.cnt\[7\] _01832_ vssd1 vssd1 vccd1 vccd1 _01834_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_113_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xoutput18 net18 vssd1 vssd1 vccd1 vccd1 mode_out[1] sky130_fd_sc_hd__clkbuf_4
XANTENNA__10164__S _04420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07039__A genblk1\[8\].osc.clkdiv_C.cnt\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire32_A _02302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10922__A1 _01811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08956_ _03645_ vssd1 vssd1 vccd1 vccd1 _00055_ sky130_fd_sc_hd__clkbuf_1
X_07907_ genblk1\[8\].osc.clkdiv_C.cnt\[8\] _01865_ _01859_ genblk1\[8\].osc.clkdiv_C.cnt\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02614_ sky130_fd_sc_hd__o22a_1
X_08887_ sig_norm.b1\[0\] _03578_ _03592_ vssd1 vssd1 vccd1 vccd1 _03593_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06597__B _01197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07838_ genblk2\[0\].wave_shpr.div.fin_quo\[5\] _02539_ _02509_ _02544_ vssd1 vssd1
+ vccd1 vccd1 _02545_ sky130_fd_sc_hd__a211o_1
X_07769_ genblk1\[0\].osc.clkdiv_C.cnt\[13\] _01256_ _01240_ genblk1\[0\].osc.clkdiv_C.cnt\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02476_ sky130_fd_sc_hd__o22a_1
Xclkbuf_leaf_36_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_36_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_78_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09508_ genblk2\[1\].wave_shpr.div.quo\[0\] _04043_ _04011_ _04045_ vssd1 vssd1 vccd1
+ vccd1 _00207_ sky130_fd_sc_hd__a22o_1
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10780_ net630 _04918_ _04922_ _04937_ vssd1 vssd1 vccd1 vccd1 _00587_ sky130_fd_sc_hd__a22o_1
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07303__B1 _01595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07502__A _02222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09439_ _03955_ _04001_ _04002_ vssd1 vssd1 vccd1 vccd1 _04003_ sky130_fd_sc_hd__o21bai_1
XPHY_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12450_ clknet_leaf_107_clk _00029_ net153 vssd1 vssd1 vccd1 vccd1 sig_norm.i\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_47_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11401_ _05374_ _05375_ _05376_ vssd1 vssd1 vccd1 vccd1 _05377_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_152_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12381_ _05956_ _06057_ vssd1 vssd1 vccd1 vccd1 _06058_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11332_ genblk2\[7\].wave_shpr.div.acc\[15\] _05323_ _05300_ vssd1 vssd1 vccd1 vccd1
+ _05324_ sky130_fd_sc_hd__mux2_1
X_11263_ net540 _05245_ _05249_ net534 _05271_ vssd1 vssd1 vccd1 vccd1 _00736_ sky130_fd_sc_hd__a221o_1
XFILLER_0_104_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13002_ clknet_leaf_133_clk _00331_ net59 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.acc\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07909__A2 _01869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10214_ _04414_ _04480_ genblk2\[3\].wave_shpr.div.acc\[18\] vssd1 vssd1 vccd1 vccd1
+ _04539_ sky130_fd_sc_hd__o21ai_1
X_11194_ _03707_ vssd1 vssd1 vccd1 vccd1 _05237_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__10913__A1 _01819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10145_ _04451_ vssd1 vssd1 vccd1 vccd1 _04486_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__06788__A _01179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10076_ _04448_ vssd1 vssd1 vccd1 vccd1 _00372_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10103__A _04451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_27_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_27_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_134_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13766_ clknet_leaf_69_clk _01077_ net213 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.acc\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10978_ _04268_ vssd1 vssd1 vccd1 vccd1 _05074_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_58_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12717_ clknet_leaf_86_clk genblk1\[9\].osc.clkdiv_C.next_cnt\[12\] net181 vssd1
+ vssd1 vccd1 vccd1 genblk1\[9\].osc.clkdiv_C.cnt\[12\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_155_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_57_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13697_ clknet_leaf_96_clk _01008_ net160 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.fin_quo\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_72_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07131__B _01250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12648_ clknet_leaf_9_clk genblk1\[5\].osc.clkdiv_C.next_cnt\[15\] net54 vssd1 vssd1
+ vccd1 vccd1 genblk1\[5\].osc.clkdiv_C.cnt\[15\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_26_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_749 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12579_ clknet_leaf_14_clk genblk1\[2\].osc.clkdiv_C.next_cnt\[0\] net70 vssd1 vssd1
+ vccd1 vccd1 genblk1\[2\].osc.clkdiv_C.cnt\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_80_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold306 genblk2\[3\].wave_shpr.div.acc\[21\] vssd1 vssd1 vccd1 vccd1 net524 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08243__A _02225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold317 _00735_ vssd1 vssd1 vccd1 vccd1 net535 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold328 _00396_ vssd1 vssd1 vccd1 vccd1 net546 sky130_fd_sc_hd__dlygate4sd3_1
Xhold339 genblk2\[9\].wave_shpr.div.quo\[10\] vssd1 vssd1 vccd1 vccd1 net557 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_99 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10904__A1 _01799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08810_ _03223_ _03509_ _03512_ _03516_ vssd1 vssd1 vccd1 vccd1 _03517_ sky130_fd_sc_hd__o211a_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09770__A1 _02077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09790_ _03714_ _04245_ _03736_ vssd1 vssd1 vccd1 vccd1 _00289_ sky130_fd_sc_hd__o21ai_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1006 genblk2\[10\].wave_shpr.div.b1\[10\] vssd1 vssd1 vccd1 vccd1 net1224 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06584__B2 _01490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1017 genblk2\[1\].wave_shpr.div.b1\[3\] vssd1 vssd1 vccd1 vccd1 net1235 sky130_fd_sc_hd__dlygate4sd3_1
X_08741_ _03410_ _03417_ vssd1 vssd1 vccd1 vccd1 _03448_ sky130_fd_sc_hd__or2_2
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1028 genblk2\[8\].wave_shpr.div.b1\[9\] vssd1 vssd1 vccd1 vccd1 net1246 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1039 genblk2\[10\].wave_shpr.div.acc\[22\] vssd1 vssd1 vccd1 vccd1 net1257 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08672_ _03361_ _03378_ vssd1 vssd1 vccd1 vccd1 _03379_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07623_ _02317_ _02328_ _02329_ vssd1 vssd1 vccd1 vccd1 _02330_ sky130_fd_sc_hd__a21oi_2
XANTENNA__06887__A2 _01738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10948__A _05051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_18_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_18_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_48_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout167_A net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07554_ _02223_ vssd1 vssd1 vccd1 vccd1 _02261_ sky130_fd_sc_hd__buf_4
XANTENNA__08089__B2 _02527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06505_ _01362_ _01430_ _01196_ vssd1 vssd1 vccd1 vccd1 _01431_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_146_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07485_ _02209_ vssd1 vssd1 vccd1 vccd1 _00003_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_75_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09224_ genblk2\[0\].wave_shpr.div.quo\[5\] _03836_ _03840_ net600 vssd1 vssd1 vccd1
+ vccd1 _00128_ sky130_fd_sc_hd__a22o_1
XANTENNA__07041__B _01576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06487__A2_N _01411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06436_ genblk1\[1\].osc.clkdiv_C.cnt\[2\] genblk1\[1\].osc.clkdiv_C.cnt\[1\] genblk1\[1\].osc.clkdiv_C.cnt\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01378_ sky130_fd_sc_hd__and3_1
XFILLER_0_134_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_733 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_498 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09155_ genblk2\[0\].wave_shpr.div.acc\[25\] genblk2\[0\].wave_shpr.div.acc\[24\]
+ genblk2\[0\].wave_shpr.div.acc\[26\] _03802_ vssd1 vssd1 vccd1 vccd1 _03803_ sky130_fd_sc_hd__or4_2
X_06367_ _01310_ vssd1 vssd1 vccd1 vccd1 _01311_ sky130_fd_sc_hd__buf_4
XFILLER_0_17_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08106_ genblk1\[4\].osc.clkdiv_C.cnt\[11\] _01574_ vssd1 vssd1 vccd1 vccd1 _02813_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09249__A _03707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09086_ modein.delay_octave_down_in\[0\] vssd1 vssd1 vccd1 vccd1 _03737_ sky130_fd_sc_hd__inv_2
X_06298_ genblk1\[0\].osc.clkdiv_C.cnt\[14\] _01256_ _01240_ genblk1\[0\].osc.clkdiv_C.cnt\[13\]
+ _01259_ vssd1 vssd1 vccd1 vccd1 _01260_ sky130_fd_sc_hd__o221ai_1
XFILLER_0_31_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08037_ _02364_ vssd1 vssd1 vccd1 vccd1 _02744_ sky130_fd_sc_hd__buf_2
XFILLER_0_4_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold840 genblk1\[7\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 net1058 sky130_fd_sc_hd__dlygate4sd3_1
Xhold851 sig_norm.acc\[2\] vssd1 vssd1 vccd1 vccd1 net1069 sky130_fd_sc_hd__dlygate4sd3_1
Xhold862 genblk1\[10\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 net1080 sky130_fd_sc_hd__dlygate4sd3_1
Xhold873 genblk2\[1\].wave_shpr.div.i\[1\] vssd1 vssd1 vccd1 vccd1 net1091 sky130_fd_sc_hd__dlygate4sd3_1
Xhold884 PWM.final_in\[2\] vssd1 vssd1 vccd1 vccd1 net1102 sky130_fd_sc_hd__dlygate4sd3_1
Xhold895 genblk2\[7\].wave_shpr.div.i\[1\] vssd1 vssd1 vccd1 vccd1 net1113 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06425__A2_N _01368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09988_ genblk2\[3\].wave_shpr.div.b1\[2\] genblk2\[3\].wave_shpr.div.acc\[2\] vssd1
+ vssd1 vccd1 vccd1 _04384_ sky130_fd_sc_hd__and2b_1
XANTENNA__07772__B1 net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08939_ sig_norm.quo\[1\] _03631_ _00024_ vssd1 vssd1 vccd1 vccd1 _03632_ sky130_fd_sc_hd__mux2_1
XFILLER_0_99_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10659__B1 _04857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11950_ genblk2\[10\].wave_shpr.div.b1\[13\] genblk2\[10\].wave_shpr.div.acc\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05772_ sky130_fd_sc_hd__and2b_1
XANTENNA__07216__B _01442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold546_A genblk2\[1\].wave_shpr.div.quo\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10901_ _05034_ vssd1 vssd1 vccd1 vccd1 _00611_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11881_ net646 _05684_ _05685_ _05712_ vssd1 vssd1 vccd1 vccd1 _00913_ sky130_fd_sc_hd__a22o_1
XFILLER_0_98_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13620_ clknet_leaf_75_clk _00933_ net204 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.b1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10832_ genblk2\[6\].wave_shpr.div.acc\[7\] genblk2\[6\].wave_shpr.div.b1\[7\] vssd1
+ vssd1 vccd1 vccd1 _04976_ sky130_fd_sc_hd__or2b_1
X_13551_ clknet_leaf_100_clk _00866_ net165 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.quo\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10069__S _04440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10763_ genblk2\[5\].wave_shpr.div.acc\[13\] _04924_ _04907_ vssd1 vssd1 vccd1 vccd1
+ _04925_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12502_ clknet_leaf_106_clk _00064_ net154 vssd1 vssd1 vccd1 vccd1 PWM.final_in\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09029__B1 _03696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13482_ clknet_leaf_99_clk net347 net168 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.quo\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10694_ net245 _02183_ _04856_ net503 _04874_ vssd1 vssd1 vccd1 vccd1 _00564_ sky130_fd_sc_hd__a221o_1
XFILLER_0_81_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12433_ genblk2\[11\].wave_shpr.div.acc\[21\] _06095_ _06096_ vssd1 vssd1 vccd1 vccd1
+ _06097_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_63_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06790__B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12364_ _06044_ _05948_ vssd1 vssd1 vccd1 vccd1 _06045_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11315_ net852 _05279_ _05283_ _05310_ vssd1 vssd1 vccd1 vccd1 _00749_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12295_ _03687_ net425 _03716_ vssd1 vssd1 vccd1 vccd1 _01031_ sky130_fd_sc_hd__a21bo_1
X_11246_ _05260_ genblk1\[7\].osc.clkdiv_C.cnt\[8\] vssd1 vssd1 vccd1 vccd1 _05263_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_120_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09752__A1 _04223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11177_ net1215 genblk2\[7\].wave_shpr.div.quo\[6\] _00019_ vssd1 vssd1 vccd1 vccd1
+ _05230_ sky130_fd_sc_hd__mux2_1
X_10128_ _04465_ genblk1\[3\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 _04475_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_145_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10059_ net1206 _01263_ _04238_ vssd1 vssd1 vccd1 vccd1 _04439_ sky130_fd_sc_hd__mux2_1
XANTENNA__06965__B _01344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09807__A2 _04248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_70_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07142__A genblk1\[9\].osc.clkdiv_C.cnt\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13749_ clknet_leaf_75_clk _01060_ net211 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.acc\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07270_ _02028_ _02043_ _02044_ vssd1 vssd1 vccd1 vccd1 _02045_ sky130_fd_sc_hd__and3_1
XANTENNA__09768__S _04039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06221_ _01181_ _01182_ vssd1 vssd1 vccd1 vccd1 _01183_ sky130_fd_sc_hd__nor2_8
XFILLER_0_155_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06152_ _01121_ _01123_ vssd1 vssd1 vccd1 vccd1 _01124_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09069__A _03701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold103 _00957_ vssd1 vssd1 vccd1 vccd1 net321 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10050__A1 _01248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold114 _00715_ vssd1 vssd1 vccd1 vccd1 net332 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold125 _01047_ vssd1 vssd1 vccd1 vccd1 net343 sky130_fd_sc_hd__dlygate4sd3_1
Xhold136 _00966_ vssd1 vssd1 vccd1 vccd1 net354 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_7_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_7_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_1_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold147 smpl_rt_clkdiv.clkDiv_inst.cnt\[6\] vssd1 vssd1 vccd1 vccd1 net365 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold158 genblk2\[3\].wave_shpr.div.quo\[16\] vssd1 vssd1 vccd1 vccd1 net376 sky130_fd_sc_hd__dlygate4sd3_1
X_09911_ _04200_ _04323_ vssd1 vssd1 vccd1 vccd1 _04324_ sky130_fd_sc_hd__xnor2_1
Xhold169 genblk2\[3\].wave_shpr.div.quo\[12\] vssd1 vssd1 vccd1 vccd1 net387 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09842_ net520 _04247_ _04250_ net639 _04272_ vssd1 vssd1 vccd1 vccd1 _00314_ sky130_fd_sc_hd__a221o_1
XFILLER_0_95_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09773_ _04236_ vssd1 vssd1 vccd1 vccd1 _00281_ sky130_fd_sc_hd__clkbuf_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06221__A _01181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06985_ _01795_ _01796_ _01798_ _01818_ _01820_ vssd1 vssd1 vccd1 vccd1 _01821_ sky130_fd_sc_hd__o2111a_1
X_08724_ _03429_ _03430_ vssd1 vssd1 vccd1 vccd1 _03431_ sky130_fd_sc_hd__xnor2_2
XTAP_2308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08655_ _03263_ _03274_ _03273_ vssd1 vssd1 vccd1 vccd1 _03362_ sky130_fd_sc_hd__a21boi_1
XANTENNA__10678__A _04672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12369__S _05982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07606_ net15 net163 _02312_ vssd1 vssd1 vccd1 vccd1 _02313_ sky130_fd_sc_hd__and3_1
XFILLER_0_49_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08586_ _03280_ _03292_ vssd1 vssd1 vccd1 vccd1 _03293_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_48_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07052__A _01441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07537_ net1111 PWM.final_in\[0\] PWM.start vssd1 vssd1 vccd1 vccd1 _02252_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07809__B2 _02468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07987__A _02225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07468_ _02147_ _02197_ vssd1 vssd1 vccd1 vccd1 _02198_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09207_ _03831_ net674 _03717_ vssd1 vssd1 vccd1 vccd1 _00120_ sky130_fd_sc_hd__a21bo_1
XANTENNA__06493__B1 _01418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06419_ _01362_ vssd1 vssd1 vccd1 vccd1 _01363_ sky130_fd_sc_hd__buf_4
X_07399_ _02146_ vssd1 vssd1 vccd1 vccd1 genblk1\[11\].osc.clkdiv_C.next_cnt\[16\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09138_ _03752_ _03784_ _03785_ vssd1 vssd1 vccd1 vccd1 _03786_ sky130_fd_sc_hd__a21o_1
XANTENNA__08234__A1 _02885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_719 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12030__A2 _05813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09069_ _03701_ _01221_ vssd1 vssd1 vccd1 vccd1 _03727_ sky130_fd_sc_hd__nand2_8
X_11100_ genblk2\[6\].wave_shpr.div.i\[3\] _02187_ _05159_ vssd1 vssd1 vccd1 vccd1
+ _05162_ sky130_fd_sc_hd__and3_1
XANTENNA__07993__B1 _01519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12080_ _05750_ _05745_ vssd1 vssd1 vccd1 vccd1 _05847_ sky130_fd_sc_hd__or2b_1
Xhold670 genblk2\[5\].wave_shpr.div.acc\[4\] vssd1 vssd1 vccd1 vccd1 net888 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold681 genblk2\[6\].wave_shpr.div.acc\[17\] vssd1 vssd1 vccd1 vccd1 net899 sky130_fd_sc_hd__dlygate4sd3_1
Xhold692 genblk2\[5\].wave_shpr.div.acc\[2\] vssd1 vssd1 vccd1 vccd1 net910 sky130_fd_sc_hd__dlygate4sd3_1
X_11031_ net1003 _05086_ _05093_ _05112_ vssd1 vssd1 vccd1 vccd1 _00663_ sky130_fd_sc_hd__a22o_1
XANTENNA__10352__S _04637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07745__B1 _01337_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06131__A net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12982_ clknet_leaf_125_clk net323 net70 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.quo\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_11933_ _05743_ _05753_ _05754_ vssd1 vssd1 vccd1 vccd1 _05755_ sky130_fd_sc_hd__o21ba_1
XTAP_2820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12279__S _03719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11183__S _05042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06785__B _01483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08170__B1 _01507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11864_ net987 _05684_ _05685_ _05700_ vssd1 vssd1 vccd1 vccd1 _00908_ sky130_fd_sc_hd__a22o_1
XFILLER_0_86_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12477__RESET_B net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13603_ clknet_leaf_45_clk _00002_ net121 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.busy
+ sky130_fd_sc_hd__dfrtp_1
X_10815_ genblk2\[5\].wave_shpr.div.i\[1\] genblk2\[5\].wave_shpr.div.i\[0\] genblk2\[5\].wave_shpr.div.i\[2\]
+ genblk2\[5\].wave_shpr.div.i\[3\] vssd1 vssd1 vccd1 vccd1 _04961_ sky130_fd_sc_hd__a31o_1
XFILLER_0_94_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11795_ genblk2\[9\].wave_shpr.div.b1\[0\] _05613_ genblk2\[9\].wave_shpr.div.acc\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05648_ sky130_fd_sc_hd__a21o_1
XANTENNA__10804__B1 _04855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13534_ clknet_leaf_81_clk _00849_ net199 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.i\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10746_ genblk2\[5\].wave_shpr.div.acc\[10\] _04886_ _04890_ _04911_ vssd1 vssd1
+ vccd1 vccd1 _00579_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09670__B1 _04048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_36_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13465_ clknet_leaf_75_clk _00782_ net203 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.b1\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10677_ net294 _04861_ _04862_ net453 _04865_ vssd1 vssd1 vccd1 vccd1 _00556_ sky130_fd_sc_hd__a221o_1
XFILLER_0_153_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11212__A _05245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12416_ net878 _06072_ _06073_ _06084_ vssd1 vssd1 vccd1 vccd1 _01076_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12021__A2 _05813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13396_ clknet_leaf_117_clk net332 net140 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.quo\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12347_ genblk2\[11\].wave_shpr.div.b1\[0\] _05982_ genblk2\[11\].wave_shpr.div.acc\[0\]
+ vssd1 vssd1 vccd1 vccd1 _06032_ sky130_fd_sc_hd__a21o_1
XFILLER_0_121_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12309__B1 _03944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08521__A _02216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12278_ _06000_ vssd1 vssd1 vccd1 vccd1 _01022_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__13265__RESET_B net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11229_ _05074_ genblk1\[7\].osc.clkdiv_C.cnt\[1\] vssd1 vssd1 vccd1 vccd1 _05253_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_4_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12043__A _04676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07137__A genblk1\[9\].osc.clkdiv_C.cnt\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12088__A2 _05844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06770_ genblk1\[4\].osc.clkdiv_C.cnt\[13\] genblk1\[4\].osc.clkdiv_C.cnt\[12\] _01637_
+ genblk1\[4\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 _01646_ sky130_fd_sc_hd__a31o_1
XFILLER_0_77_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06695__B _01323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08440_ _02407_ _02403_ genblk2\[10\].wave_shpr.div.fin_quo\[2\] vssd1 vssd1 vccd1
+ vccd1 _03147_ sky130_fd_sc_hd__or3b_1
XFILLER_0_148_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_93_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08371_ _02998_ _03000_ _02999_ vssd1 vssd1 vccd1 vccd1 _03078_ sky130_fd_sc_hd__o21a_1
XFILLER_0_147_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09498__S _04039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07322_ genblk1\[11\].osc.clkdiv_C.cnt\[16\] _02085_ vssd1 vssd1 vccd1 vccd1 _02086_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__09661__B1 _04045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07600__A net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07253_ genblk1\[10\].osc.clkdiv_C.cnt\[1\] genblk1\[10\].osc.clkdiv_C.cnt\[0\] genblk1\[10\].osc.clkdiv_C.cnt\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02033_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_143_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_639 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06204_ _01166_ _01167_ vssd1 vssd1 vccd1 vccd1 _01168_ sky130_fd_sc_hd__and2_1
X_07184_ genblk1\[9\].osc.clkdiv_C.cnt\[9\] _01972_ vssd1 vssd1 vccd1 vccd1 _01975_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06135_ net11 _01106_ vssd1 vssd1 vccd1 vccd1 _01107_ sky130_fd_sc_hd__xor2_1
XANTENNA__11220__B1 _05250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09527__A _04046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09825_ _04069_ genblk1\[2\].osc.clkdiv_C.cnt\[7\] vssd1 vssd1 vccd1 vccd1 _04263_
+ sky130_fd_sc_hd__and2_1
XANTENNA__07047__A _01336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09756_ _04226_ vssd1 vssd1 vccd1 vccd1 _00274_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10900__S _04848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06968_ genblk1\[7\].osc.clkdiv_C.cnt\[1\] _01801_ _01803_ vssd1 vssd1 vccd1 vccd1
+ _01804_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12079__A2 _05844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08707_ genblk2\[2\].wave_shpr.div.fin_quo\[3\] net25 _03116_ _02224_ vssd1 vssd1
+ vccd1 vccd1 _03414_ sky130_fd_sc_hd__a31o_1
XFILLER_0_69_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12099__S _05787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09687_ genblk2\[2\].wave_shpr.div.acc\[6\] genblk2\[2\].wave_shpr.div.b1\[6\] vssd1
+ vssd1 vccd1 vccd1 _04167_ sky130_fd_sc_hd__or2b_1
XTAP_2116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06899_ genblk1\[6\].osc.clkdiv_C.cnt\[7\] vssd1 vssd1 vccd1 vccd1 _01753_ sky130_fd_sc_hd__inv_2
XANTENNA__08152__B1 _01250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08638_ _02682_ _02686_ _02685_ vssd1 vssd1 vccd1 vccd1 _03345_ sky130_fd_sc_hd__o21ai_1
XTAP_1415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08569_ _03273_ _03274_ _03263_ vssd1 vssd1 vccd1 vccd1 _03276_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10600_ genblk2\[5\].wave_shpr.div.fin_quo\[3\] genblk2\[5\].wave_shpr.div.quo\[2\]
+ _00015_ vssd1 vssd1 vccd1 vccd1 _04825_ sky130_fd_sc_hd__mux2_1
Xfanout42 net43 vssd1 vssd1 vccd1 vccd1 net42 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_647 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout53 net58 vssd1 vssd1 vccd1 vccd1 net53 sky130_fd_sc_hd__buf_2
XFILLER_0_119_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11580_ _05387_ _05495_ vssd1 vssd1 vccd1 vccd1 _05496_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout64 net65 vssd1 vssd1 vccd1 vccd1 net64 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_107_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09201__S _03822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout75 net84 vssd1 vssd1 vccd1 vccd1 net75 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_36_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout86 net88 vssd1 vssd1 vccd1 vccd1 net86 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_107_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10531_ genblk2\[4\].wave_shpr.div.i\[3\] _02176_ _04758_ vssd1 vssd1 vccd1 vccd1
+ _04761_ sky130_fd_sc_hd__and3_1
XFILLER_0_64_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout97 net98 vssd1 vssd1 vccd1 vccd1 net97 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10347__S _04637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13250_ clknet_leaf_2_clk _00573_ net43 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.acc\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10462_ net1024 _04683_ _04690_ _04711_ vssd1 vssd1 vccd1 vccd1 _00495_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06126__A _01097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06218__B1 _01179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12201_ genblk2\[11\].wave_shpr.div.acc\[3\] genblk2\[11\].wave_shpr.div.b1\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05939_ sky130_fd_sc_hd__or2b_1
XANTENNA__09955__A1 _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13181_ clknet_leaf_112_clk _00506_ net68 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.acc\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10393_ _04477_ genblk1\[4\].osc.clkdiv_C.cnt\[5\] vssd1 vssd1 vccd1 vccd1 _04665_
+ sky130_fd_sc_hd__and2_1
XANTENNA__07966__B1 _01675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12132_ _05774_ _05734_ vssd1 vssd1 vccd1 vccd1 _05887_ sky130_fd_sc_hd__or2b_1
XFILLER_0_103_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12063_ genblk2\[10\].wave_shpr.div.quo\[22\] _05812_ _05825_ net334 _05836_ vssd1
+ vssd1 vccd1 vccd1 _00971_ sky130_fd_sc_hd__a221o_1
XANTENNA__08060__B _01238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06499__C net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11014_ net819 _05086_ _05093_ _05099_ vssd1 vssd1 vccd1 vccd1 _00659_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11278__B1 _05250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12965_ clknet_leaf_110_clk _00294_ net130 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_11916_ genblk2\[10\].wave_shpr.div.acc\[10\] genblk2\[10\].wave_shpr.div.b1\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05738_ sky130_fd_sc_hd__or2b_1
XTAP_2650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12896_ clknet_leaf_32_clk _00227_ net99 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.quo\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09900__A _04247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11847_ genblk2\[9\].wave_shpr.div.acc\[12\] _05687_ _05673_ vssd1 vssd1 vccd1 vccd1
+ _05688_ sky130_fd_sc_hd__mux2_1
XTAP_1960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11778_ net362 _05628_ _05629_ net513 _05638_ vssd1 vssd1 vccd1 vccd1 _00884_ sky130_fd_sc_hd__a221o_1
XFILLER_0_16_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13517_ clknet_leaf_77_clk _00834_ net208 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.acc\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06457__B1 genblk1\[1\].osc.clkdiv_C.cnt\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10729_ net863 _04886_ _04890_ _04898_ vssd1 vssd1 vccd1 vccd1 _00575_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_319 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13448_ clknet_leaf_91_clk _00765_ net147 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.i\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08749__A2 _02309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13379_ clknet_leaf_81_clk _00698_ net199 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.b1\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11753__A1 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_9 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_53_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07940_ net13 _02364_ vssd1 vssd1 vccd1 vccd1 _02647_ sky130_fd_sc_hd__nand2_1
X_07871_ genblk2\[1\].wave_shpr.div.fin_quo\[0\] _02524_ _02307_ genblk2\[1\].wave_shpr.div.fin_quo\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02578_ sky130_fd_sc_hd__a22o_1
XANTENNA__08382__B1 _01418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09610_ _04042_ vssd1 vssd1 vccd1 vccd1 _04109_ sky130_fd_sc_hd__buf_2
XANTENNA__11816__S _05613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06822_ net1120 _01693_ vssd1 vssd1 vccd1 vccd1 genblk1\[5\].osc.clkdiv_C.next_cnt\[0\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_leaf_68_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_111_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09541_ net552 _04052_ _04053_ net462 _04061_ vssd1 vssd1 vccd1 vccd1 _00224_ sky130_fd_sc_hd__a221o_1
X_06753_ _01599_ _01632_ _01633_ vssd1 vssd1 vccd1 vccd1 _01634_ sky130_fd_sc_hd__and3_1
X_09472_ _03701_ vssd1 vssd1 vccd1 vccd1 _04024_ sky130_fd_sc_hd__clkbuf_4
X_06684_ _01173_ _01187_ _01188_ vssd1 vssd1 vccd1 vccd1 _01574_ sky130_fd_sc_hd__mux2_4
XFILLER_0_116_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08423_ _03085_ _03123_ vssd1 vssd1 vccd1 vccd1 _03130_ sky130_fd_sc_hd__or2_1
XANTENNA__06696__B1 _01574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10956__A _05051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_126_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08354_ _02932_ _02841_ genblk2\[4\].wave_shpr.div.fin_quo\[4\] vssd1 vssd1 vccd1
+ vccd1 _03061_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08437__A1 _02525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07305_ _02063_ _02066_ _02067_ _02068_ vssd1 vssd1 vccd1 vccd1 _02069_ sky130_fd_sc_hd__or4_1
XFILLER_0_18_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08285_ _02972_ _02991_ vssd1 vssd1 vccd1 vccd1 _02992_ sky130_fd_sc_hd__and2b_1
XFILLER_0_132_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_285 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11992__A1 _01855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07236_ genblk1\[10\].osc.clkdiv_C.cnt\[1\] _02001_ _02002_ _02003_ vssd1 vssd1 vccd1
+ vccd1 _02018_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_33_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_14_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07167_ genblk1\[9\].osc.clkdiv_C.cnt\[4\] _01960_ vssd1 vssd1 vccd1 vccd1 _01963_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_132_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09257__A _03853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06118_ _01088_ _01092_ vssd1 vssd1 vccd1 vccd1 smpl_rt_clkdiv.clkDiv_inst.next_cnt\[5\]
+ sky130_fd_sc_hd__nor2_1
X_07098_ genblk1\[8\].osc.clkdiv_C.cnt\[10\] _01902_ _01905_ vssd1 vssd1 vccd1 vccd1
+ genblk1\[8\].osc.clkdiv_C.next_cnt\[10\] sky130_fd_sc_hd__o21a_1
XFILLER_0_112_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07963__A3 _01361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout210 net218 vssd1 vssd1 vccd1 vccd1 net210 sky130_fd_sc_hd__buf_2
XANTENNA__11726__S _00023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09808_ _04247_ vssd1 vssd1 vccd1 vccd1 _04253_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__10630__S _04834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout62_A net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09739_ genblk2\[2\].wave_shpr.div.fin_quo\[2\] net1343 _00009_ vssd1 vssd1 vccd1
+ vccd1 _04217_ sky130_fd_sc_hd__mux2_1
X_12750_ clknet_leaf_46_clk genblk1\[11\].osc.clkdiv_C.next_cnt\[9\] net119 vssd1
+ vssd1 vccd1 vccd1 genblk1\[11\].osc.clkdiv_C.cnt\[9\] sky130_fd_sc_hd__dfrtp_2
XTAP_1201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11701_ _05561_ _05591_ _05592_ vssd1 vssd1 vccd1 vccd1 _05593_ sky130_fd_sc_hd__a21o_1
XTAP_1245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12681_ clknet_leaf_120_clk genblk1\[7\].osc.clkdiv_C.next_cnt\[12\] net82 vssd1
+ vssd1 vccd1 vccd1 genblk1\[7\].osc.clkdiv_C.cnt\[12\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_139_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11632_ genblk2\[8\].wave_shpr.div.acc\[20\] _05533_ _05534_ vssd1 vssd1 vccd1 vccd1
+ _05535_ sky130_fd_sc_hd__a21o_1
XFILLER_0_108_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11563_ genblk2\[8\].wave_shpr.div.acc\[3\] _05482_ _05417_ vssd1 vssd1 vccd1 vccd1
+ _05483_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13302_ clknet_leaf_87_clk _00623_ net179 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.b1\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11983__A1 _03732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10514_ net1144 _04657_ _04655_ _04749_ vssd1 vssd1 vccd1 vccd1 _00509_ sky130_fd_sc_hd__a22o_1
XFILLER_0_135_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11494_ _05443_ vssd1 vssd1 vccd1 vccd1 _05444_ sky130_fd_sc_hd__buf_2
XFILLER_0_107_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13233_ clknet_leaf_15_clk _00556_ net73 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.quo\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10445_ net998 _04683_ _04690_ _04698_ vssd1 vssd1 vccd1 vccd1 _00491_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13164_ clknet_leaf_127_clk net843 net67 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.acc\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10376_ genblk2\[4\].wave_shpr.div.quo\[5\] _04652_ _04656_ net749 vssd1 vssd1 vccd1
+ vccd1 _00464_ sky130_fd_sc_hd__a22o_1
X_12115_ _05765_ _05873_ vssd1 vssd1 vccd1 vccd1 _05874_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06611__B1 _01171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13095_ clknet_leaf_1_clk _00422_ net41 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.acc\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_12046_ net373 _05823_ _05825_ net521 _05827_ vssd1 vssd1 vccd1 vccd1 _00963_ sky130_fd_sc_hd__a221o_1
XANTENNA__11499__B1 _05446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07415__A _02155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12948_ clknet_leaf_125_clk _00277_ net71 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.b1\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08667__B2 _02362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12879_ clknet_leaf_119_clk _00210_ net139 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07890__A2 _02539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08070_ _02770_ _02771_ _02775_ vssd1 vssd1 vccd1 vccd1 _02777_ sky130_fd_sc_hd__a21o_1
XFILLER_0_114_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07021_ genblk1\[7\].osc.clkdiv_C.cnt\[13\] _01842_ _01822_ vssd1 vssd1 vccd1 vccd1
+ _01844_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_140_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11400__A genblk2\[8\].wave_shpr.div.b1\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08972_ _03657_ _03658_ sig_norm.quo\[6\] _01098_ vssd1 vssd1 vccd1 vccd1 _03659_
+ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__07309__B _01430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07923_ genblk1\[8\].osc.clkdiv_C.cnt\[8\] _01865_ vssd1 vssd1 vccd1 vccd1 _02630_
+ sky130_fd_sc_hd__and2_1
Xhold18 _00561_ vssd1 vssd1 vccd1 vccd1 net236 sky130_fd_sc_hd__dlygate4sd3_1
Xhold29 genblk2\[10\].wave_shpr.div.acc_next\[0\] vssd1 vssd1 vccd1 vccd1 net247 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08355__B1 _02222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout197_A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07854_ _02518_ _02555_ _02560_ vssd1 vssd1 vccd1 vccd1 _02561_ sky130_fd_sc_hd__a21oi_1
X_06805_ genblk1\[5\].osc.clkdiv_C.cnt\[9\] _01362_ _01226_ vssd1 vssd1 vccd1 vccd1
+ _01677_ sky130_fd_sc_hd__and3_1
X_07785_ _02482_ _02488_ _02491_ vssd1 vssd1 vccd1 vccd1 _02492_ sky130_fd_sc_hd__o21ba_1
X_09524_ _03853_ genblk1\[1\].osc.clkdiv_C.cnt\[2\] vssd1 vssd1 vccd1 vccd1 _04051_
+ sky130_fd_sc_hd__and2_1
X_06736_ genblk1\[4\].osc.clkdiv_C.cnt\[6\] _01616_ vssd1 vssd1 vccd1 vccd1 _01620_
+ sky130_fd_sc_hd__and2_1
XANTENNA__08658__B2 _02592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09540__A _04058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09455_ _04015_ vssd1 vssd1 vccd1 vccd1 _00184_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06667_ _01556_ _01344_ vssd1 vssd1 vccd1 vccd1 _01557_ sky130_fd_sc_hd__nand2_1
XFILLER_0_149_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08406_ net25 vssd1 vssd1 vccd1 vccd1 _03113_ sky130_fd_sc_hd__buf_2
XFILLER_0_143_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09386_ genblk2\[11\].wave_shpr.div.i\[3\] _02212_ _03949_ vssd1 vssd1 vccd1 vccd1
+ _03952_ sky130_fd_sc_hd__and3_1
XFILLER_0_81_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06598_ genblk1\[3\].osc.clkdiv_C.cnt\[16\] _01197_ vssd1 vssd1 vccd1 vccd1 _01506_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07060__A genblk1\[8\].osc.clkdiv_C.cnt\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08337_ genblk2\[6\].wave_shpr.div.fin_quo\[4\] _02734_ _02737_ _02261_ vssd1 vssd1
+ vccd1 vccd1 _03044_ sky130_fd_sc_hd__a31o_1
XANTENNA__09428__A_N genblk2\[1\].wave_shpr.div.b1\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08268_ genblk2\[11\].wave_shpr.div.fin_quo\[5\] _02361_ vssd1 vssd1 vccd1 vccd1
+ _02975_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07219_ _01358_ net37 vssd1 vssd1 vccd1 vccd1 _02001_ sky130_fd_sc_hd__nand2_2
X_08199_ _02404_ _02410_ _02405_ vssd1 vssd1 vccd1 vccd1 _02906_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_132_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10230_ genblk2\[3\].wave_shpr.div.acc\[23\] _04417_ vssd1 vssd1 vccd1 vccd1 _04550_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_30_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06404__A genblk1\[1\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10161_ net941 _04486_ _04490_ _04498_ vssd1 vssd1 vccd1 vccd1 _00407_ sky130_fd_sc_hd__a22o_1
XANTENNA__07219__B net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_hold576_A genblk2\[3\].wave_shpr.div.quo\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10940__A2 _05052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10092_ net814 _04452_ _04456_ net849 vssd1 vssd1 vccd1 vccd1 _00380_ sky130_fd_sc_hd__a22o_1
XANTENNA__07149__B2 genblk1\[9\].osc.clkdiv_C.cnt\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12802_ clknet_leaf_59_clk _00135_ net193 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.quo\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09846__B1 _04250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10994_ _04982_ _04983_ vssd1 vssd1 vccd1 vccd1 _05084_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12445__A2 _03947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12733_ clknet_leaf_38_clk genblk1\[10\].osc.clkdiv_C.next_cnt\[10\] net115 vssd1
+ vssd1 vccd1 vccd1 genblk1\[10\].osc.clkdiv_C.cnt\[10\] sky130_fd_sc_hd__dfrtp_4
XTAP_1020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06793__B _01592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11191__S _05042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12664_ clknet_leaf_26_clk genblk1\[6\].osc.clkdiv_C.next_cnt\[13\] net88 vssd1 vssd1
+ vccd1 vccd1 genblk1\[6\].osc.clkdiv_C.cnt\[13\] sky130_fd_sc_hd__dfrtp_4
XTAP_1086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_764 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11615_ net802 _05507_ _05445_ _05522_ vssd1 vssd1 vccd1 vccd1 _00837_ sky130_fd_sc_hd__a22o_1
XFILLER_0_143_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09074__A1 _01592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12595_ clknet_leaf_11_clk genblk1\[2\].osc.clkdiv_C.next_cnt\[16\] net56 vssd1 vssd1
+ vccd1 vccd1 genblk1\[2\].osc.clkdiv_C.cnt\[16\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_93_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09596__S _04095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11546_ net274 _05441_ _05444_ net445 _05470_ vssd1 vssd1 vccd1 vccd1 _00820_ sky130_fd_sc_hd__a221o_1
XFILLER_0_53_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11477_ _03704_ net1042 _04233_ vssd1 vssd1 vccd1 vccd1 _00786_ sky130_fd_sc_hd__a21o_1
XFILLER_0_123_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13216_ clknet_leaf_6_clk _00539_ net46 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.b1\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10428_ genblk2\[4\].wave_shpr.div.acc\[1\] _04685_ _04623_ vssd1 vssd1 vccd1 vccd1
+ _04686_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13147_ clknet_leaf_121_clk net638 net80 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.quo\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10359_ genblk2\[5\].wave_shpr.div.b1\[15\] _01365_ _04637_ vssd1 vssd1 vccd1 vccd1
+ _04648_ sky130_fd_sc_hd__mux2_1
XANTENNA__07129__B _01801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13078_ clknet_leaf_125_clk _00405_ net61 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.acc\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08337__B1 _02261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12029_ net320 _05813_ _05817_ genblk2\[10\].wave_shpr.div.quo\[6\] vssd1 vssd1 vccd1
+ vccd1 _00956_ sky130_fd_sc_hd__a22o_1
XANTENNA__12051__A _03833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10144__B1 _04456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11892__B1 _03694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07560__A1 genblk1\[9\].osc.clkdiv_C.cnt\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07570_ _02267_ _02273_ _02276_ vssd1 vssd1 vccd1 vccd1 _02277_ sky130_fd_sc_hd__a21o_1
X_06521_ _01433_ _01434_ _01435_ _01436_ _01446_ vssd1 vssd1 vccd1 vccd1 _01447_ sky130_fd_sc_hd__a221o_1
XFILLER_0_88_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09240_ net495 _03845_ _03847_ net584 _03848_ vssd1 vssd1 vccd1 vccd1 _00136_ sky130_fd_sc_hd__a221o_1
X_06452_ genblk1\[1\].osc.clkdiv_C.cnt\[7\] _01387_ vssd1 vssd1 vccd1 vccd1 _01389_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_146_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09171_ net1218 genblk2\[0\].wave_shpr.div.quo\[6\] _00001_ vssd1 vssd1 vccd1 vccd1
+ _03812_ sky130_fd_sc_hd__mux2_1
X_06383_ _01254_ vssd1 vssd1 vccd1 vccd1 _01327_ sky130_fd_sc_hd__clkbuf_8
X_08122_ genblk1\[4\].osc.clkdiv_C.cnt\[7\] _01340_ _01304_ genblk1\[4\].osc.clkdiv_C.cnt\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02829_ sky130_fd_sc_hd__o22a_1
XFILLER_0_43_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08053_ _02756_ _02757_ _02758_ _02759_ vssd1 vssd1 vccd1 vccd1 _02760_ sky130_fd_sc_hd__or4_1
XFILLER_0_31_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout112_A net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07004_ _01823_ _01832_ _01833_ vssd1 vssd1 vccd1 vccd1 genblk1\[7\].osc.clkdiv_C.next_cnt\[6\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_102_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput19 net19 vssd1 vssd1 vccd1 vccd1 sigout sky130_fd_sc_hd__buf_2
XANTENNA__06224__A _01179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08576__B1 _02361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07039__B _01487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09535__A _03719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08955_ net1339 _03644_ _00024_ vssd1 vssd1 vccd1 vccd1 _03645_ sky130_fd_sc_hd__mux2_1
X_07906_ genblk1\[8\].osc.clkdiv_C.cnt\[9\] _01859_ _02610_ _02611_ _02612_ vssd1
+ vssd1 vccd1 vccd1 _02613_ sky130_fd_sc_hd__a2111o_1
X_08886_ sig_norm.b1\[3\] sig_norm.acc\[3\] vssd1 vssd1 vccd1 vccd1 _03592_ sky130_fd_sc_hd__xnor2_1
X_07837_ _02542_ _02543_ vssd1 vssd1 vccd1 vccd1 _02544_ sky130_fd_sc_hd__nor2_1
X_07768_ _02472_ _02473_ _02474_ vssd1 vssd1 vccd1 vccd1 _02475_ sky130_fd_sc_hd__or3b_1
XANTENNA__13549__RESET_B net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09507_ _04044_ vssd1 vssd1 vccd1 vccd1 _04045_ sky130_fd_sc_hd__clkbuf_4
X_06719_ genblk1\[4\].osc.clkdiv_C.cnt\[1\] genblk1\[4\].osc.clkdiv_C.cnt\[0\] genblk1\[4\].osc.clkdiv_C.cnt\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01607_ sky130_fd_sc_hd__a21o_1
XFILLER_0_39_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07699_ genblk2\[10\].wave_shpr.div.fin_quo\[3\] vssd1 vssd1 vccd1 vccd1 _02406_
+ sky130_fd_sc_hd__inv_2
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09438_ genblk2\[1\].wave_shpr.div.b1\[16\] genblk2\[1\].wave_shpr.div.acc\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04002_ sky130_fd_sc_hd__and2b_1
XPHY_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09369_ _03937_ _03938_ vssd1 vssd1 vccd1 vccd1 _03939_ sky130_fd_sc_hd__nand2_1
XFILLER_0_136_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09056__A1 _01201_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11400_ genblk2\[8\].wave_shpr.div.b1\[1\] genblk2\[8\].wave_shpr.div.acc\[1\] vssd1
+ vssd1 vccd1 vccd1 _05376_ sky130_fd_sc_hd__or2b_1
XFILLER_0_124_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12380_ _05957_ _05934_ vssd1 vssd1 vccd1 vccd1 _06057_ sky130_fd_sc_hd__or2b_1
XFILLER_0_62_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10610__A1 _01189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11331_ _05210_ _05322_ vssd1 vssd1 vccd1 vccd1 _05323_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10355__S _04637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11040__A _05051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11262_ _04676_ _01813_ vssd1 vssd1 vccd1 vccd1 _05271_ sky130_fd_sc_hd__nor2_1
XFILLER_0_104_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13001_ clknet_leaf_133_clk _00330_ net59 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.acc\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10213_ _04415_ _04480_ vssd1 vssd1 vccd1 vccd1 _04538_ sky130_fd_sc_hd__or2_1
X_11193_ _01865_ vssd1 vssd1 vccd1 vccd1 _05236_ sky130_fd_sc_hd__inv_2
X_10144_ net976 _04452_ _04456_ _04485_ vssd1 vssd1 vccd1 vccd1 _00403_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08319__B1 _02316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06788__B _01262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11186__S _05042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10075_ genblk2\[4\].wave_shpr.div.b1\[15\] _01365_ _04440_ vssd1 vssd1 vccd1 vccd1
+ _04448_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13765_ clknet_leaf_69_clk _01076_ net213 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.acc\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10977_ genblk2\[6\].wave_shpr.div.quo\[21\] _05062_ _05064_ net567 _05073_ vssd1
+ vssd1 vccd1 vccd1 _00648_ sky130_fd_sc_hd__a221o_1
XFILLER_0_97_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12716_ clknet_leaf_56_clk genblk1\[9\].osc.clkdiv_C.next_cnt\[11\] net175 vssd1
+ vssd1 vccd1 vccd1 genblk1\[9\].osc.clkdiv_C.cnt\[11\] sky130_fd_sc_hd__dfrtp_4
X_13696_ clknet_leaf_96_clk _01007_ net161 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.fin_quo\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_127_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12647_ clknet_leaf_9_clk genblk1\[5\].osc.clkdiv_C.next_cnt\[14\] net54 vssd1 vssd1
+ vccd1 vccd1 genblk1\[5\].osc.clkdiv_C.cnt\[14\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_26_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07058__B1 _01246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12578_ clknet_leaf_29_clk genblk1\[1\].osc.clkdiv_C.next_cnt\[17\] net96 vssd1 vssd1
+ vccd1 vccd1 genblk1\[1\].osc.clkdiv_C.cnt\[17\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__08524__A _02216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11529_ net263 _05454_ _05458_ net502 _05461_ vssd1 vssd1 vccd1 vccd1 _00812_ sky130_fd_sc_hd__a221o_1
XFILLER_0_80_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold307 genblk2\[3\].wave_shpr.div.quo\[11\] vssd1 vssd1 vccd1 vccd1 net525 sky130_fd_sc_hd__clkdlybuf4s25_1
XFILLER_0_40_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold318 genblk2\[10\].wave_shpr.div.acc\[24\] vssd1 vssd1 vccd1 vccd1 net536 sky130_fd_sc_hd__dlygate4sd3_1
Xhold329 genblk2\[10\].wave_shpr.div.quo\[17\] vssd1 vssd1 vccd1 vccd1 net547 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_68_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08558__B1 _02223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_67 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06584__A2 _01231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08740_ _03412_ _03416_ vssd1 vssd1 vccd1 vccd1 _03447_ sky130_fd_sc_hd__nand2_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1007 genblk2\[4\].wave_shpr.div.b1\[7\] vssd1 vssd1 vccd1 vccd1 net1225 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1018 genblk2\[9\].wave_shpr.div.b1\[8\] vssd1 vssd1 vccd1 vccd1 net1236 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1029 genblk2\[2\].wave_shpr.div.b1\[1\] vssd1 vssd1 vccd1 vccd1 net1247 sky130_fd_sc_hd__dlygate4sd3_1
X_08671_ _03362_ _03377_ vssd1 vssd1 vccd1 vccd1 _03378_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11824__S _05613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07622_ genblk1\[11\].osc.clkdiv_C.cnt\[7\] _01211_ vssd1 vssd1 vccd1 vccd1 _02329_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07603__A _02221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07553_ _01157_ vssd1 vssd1 vccd1 vccd1 _02260_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__08089__A2 _02309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06504_ _01224_ vssd1 vssd1 vccd1 vccd1 _01430_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_146_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07484_ _02206_ _02153_ genblk2\[10\].wave_shpr.div.busy vssd1 vssd1 vccd1 vccd1
+ _02209_ sky130_fd_sc_hd__and3b_2
XANTENNA__06219__A _01174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_146_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09223_ net600 _03836_ _03840_ net728 vssd1 vssd1 vccd1 vccd1 _00127_ sky130_fd_sc_hd__a22o_1
X_06435_ _01377_ vssd1 vssd1 vccd1 vccd1 genblk1\[1\].osc.clkdiv_C.next_cnt\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_745 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09154_ genblk2\[0\].wave_shpr.div.acc\[23\] _03801_ vssd1 vssd1 vccd1 vccd1 _03802_
+ sky130_fd_sc_hd__or2_2
XFILLER_0_146_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06366_ _01308_ _01309_ vssd1 vssd1 vccd1 vccd1 _01310_ sky130_fd_sc_hd__nand2_1
X_08105_ _01588_ _01192_ _01208_ vssd1 vssd1 vccd1 vccd1 _02812_ sky130_fd_sc_hd__and3_1
X_09085_ _03714_ _03734_ _03736_ vssd1 vssd1 vccd1 vccd1 _00093_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_114_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06297_ genblk1\[0\].osc.clkdiv_C.cnt\[2\] _01190_ _01258_ genblk1\[0\].osc.clkdiv_C.cnt\[5\]
+ vssd1 vssd1 vccd1 vccd1 _01259_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_130_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06272__A1 _01229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08036_ genblk2\[6\].wave_shpr.div.fin_quo\[7\] _02539_ _02742_ vssd1 vssd1 vccd1
+ vccd1 _02743_ sky130_fd_sc_hd__a21o_1
XFILLER_0_114_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold830 genblk2\[7\].wave_shpr.div.acc\[19\] vssd1 vssd1 vccd1 vccd1 net1048 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold841 genblk2\[9\].wave_shpr.div.acc\[1\] vssd1 vssd1 vccd1 vccd1 net1059 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12345__A1 _03819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold852 genblk2\[7\].wave_shpr.div.acc\[1\] vssd1 vssd1 vccd1 vccd1 net1070 sky130_fd_sc_hd__dlygate4sd3_1
Xhold863 genblk2\[10\].wave_shpr.div.acc\[26\] vssd1 vssd1 vccd1 vccd1 net1081 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08013__A2 _01367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold874 genblk1\[8\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 net1092 sky130_fd_sc_hd__dlygate4sd3_1
Xhold885 PWM.final_in\[1\] vssd1 vssd1 vccd1 vccd1 net1103 sky130_fd_sc_hd__dlygate4sd3_1
Xhold896 genblk2\[8\].wave_shpr.div.acc\[19\] vssd1 vssd1 vccd1 vccd1 net1114 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09265__A _03853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09987_ _04379_ genblk2\[3\].wave_shpr.div.acc\[1\] _04382_ vssd1 vssd1 vccd1 vccd1
+ _04383_ sky130_fd_sc_hd__a21o_1
X_08938_ sig_norm.quo\[0\] _01098_ _03629_ _03630_ vssd1 vssd1 vccd1 vccd1 _03631_
+ sky130_fd_sc_hd__a22o_1
XANTENNA__07323__A2_N _01334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09513__A2 _04043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08869_ sig_norm.b1\[3\] vssd1 vssd1 vccd1 vccd1 _03575_ sky130_fd_sc_hd__inv_2
XFILLER_0_98_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11734__S _00023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10900_ net1288 _01991_ _04848_ vssd1 vssd1 vccd1 vccd1 _05034_ sky130_fd_sc_hd__mux2_1
X_11880_ _05609_ _05646_ _05709_ genblk2\[9\].wave_shpr.div.acc\[21\] vssd1 vssd1
+ vccd1 vccd1 _05712_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_86_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10831_ genblk2\[6\].wave_shpr.div.acc\[8\] genblk2\[6\].wave_shpr.div.b1\[8\] vssd1
+ vssd1 vccd1 vccd1 _04975_ sky130_fd_sc_hd__or2b_1
XFILLER_0_39_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13550_ clknet_leaf_100_clk _00865_ net170 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.quo\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10762_ _04805_ _04923_ vssd1 vssd1 vccd1 vccd1 _04924_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06129__A net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07827__A2 _02309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06594__A2_N _01500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12501_ clknet_leaf_106_clk _00063_ net153 vssd1 vssd1 vccd1 vccd1 PWM.final_in\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_13481_ clknet_leaf_100_clk _00798_ net168 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09029__A1 _03694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10693_ _04869_ genblk1\[5\].osc.clkdiv_C.cnt\[12\] vssd1 vssd1 vccd1 vccd1 _04874_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12432_ genblk2\[11\].wave_shpr.div.acc\[21\] genblk2\[11\].wave_shpr.div.acc\[20\]
+ _05978_ net20 vssd1 vssd1 vccd1 vccd1 _06096_ sky130_fd_sc_hd__or4_1
XFILLER_0_81_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12363_ _05949_ _05938_ vssd1 vssd1 vccd1 vccd1 _06044_ sky130_fd_sc_hd__or2b_1
XANTENNA__08063__B _01238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11314_ genblk2\[7\].wave_shpr.div.acc\[11\] _05309_ _05300_ vssd1 vssd1 vccd1 vccd1
+ _05310_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12294_ _03732_ net406 _03733_ vssd1 vssd1 vccd1 vccd1 _01030_ sky130_fd_sc_hd__o21a_1
XFILLER_0_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11245_ net548 _05255_ _05256_ net550 _05262_ vssd1 vssd1 vccd1 vccd1 _00727_ sky130_fd_sc_hd__a221o_1
XANTENNA__09201__A1 _01183_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08004__A2 _01519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07212__B1 _01214_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11176_ _05229_ vssd1 vssd1 vccd1 vccd1 _00691_ sky130_fd_sc_hd__clkbuf_1
X_10127_ net529 _04451_ _04455_ net607 _04474_ vssd1 vssd1 vccd1 vccd1 _00397_ sky130_fd_sc_hd__a221o_1
XFILLER_0_145_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10058_ _04438_ vssd1 vssd1 vccd1 vccd1 _00364_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11311__A2 _05279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08519__A _02216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07142__B _01514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13748_ clknet_leaf_85_clk net1221 net184 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.acc\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_57_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13679_ clknet_leaf_43_clk net860 net190 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.acc\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06220_ _01177_ vssd1 vssd1 vccd1 vccd1 _01182_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_26_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12024__B1 _05817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06151_ _01107_ _01110_ _01122_ vssd1 vssd1 vccd1 vccd1 _01123_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_81_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09069__B _01221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold104 genblk2\[2\].wave_shpr.div.quo\[19\] vssd1 vssd1 vccd1 vccd1 net322 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold115 genblk2\[3\].wave_shpr.div.i\[4\] vssd1 vssd1 vccd1 vccd1 net333 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold126 genblk2\[6\].wave_shpr.div.quo\[10\] vssd1 vssd1 vccd1 vccd1 net344 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold137 genblk2\[11\].wave_shpr.div.quo\[8\] vssd1 vssd1 vccd1 vccd1 net355 sky130_fd_sc_hd__clkbuf_2
Xhold148 genblk2\[1\].wave_shpr.div.acc\[11\] vssd1 vssd1 vccd1 vccd1 net366 sky130_fd_sc_hd__dlygate4sd3_1
X_09910_ _04201_ _04159_ vssd1 vssd1 vccd1 vccd1 _04323_ sky130_fd_sc_hd__or2b_1
XFILLER_0_1_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold159 _00392_ vssd1 vssd1 vccd1 vccd1 net377 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09841_ _04269_ genblk1\[2\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 _04272_
+ sky130_fd_sc_hd__and2_1
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11550__A2 _05417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09772_ net1298 _01256_ _04039_ vssd1 vssd1 vccd1 vccd1 _04236_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06984_ genblk1\[7\].osc.clkdiv_C.cnt\[8\] _01819_ vssd1 vssd1 vccd1 vccd1 _01820_
+ sky130_fd_sc_hd__xnor2_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06221__B _01182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08723_ _02536_ _02586_ vssd1 vssd1 vccd1 vccd1 _03430_ sky130_fd_sc_hd__and2b_1
XANTENNA__09813__A _04058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10959__A _05054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08654_ _03320_ _03325_ _03360_ vssd1 vssd1 vccd1 vccd1 _03361_ sky130_fd_sc_hd__o21bai_2
XTAP_2309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07605_ net17 net18 vssd1 vssd1 vccd1 vccd1 _02312_ sky130_fd_sc_hd__or2_2
XTAP_1608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08585_ _03284_ _03291_ vssd1 vssd1 vccd1 vccd1 _03292_ sky130_fd_sc_hd__xnor2_2
XTAP_1619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07536_ net279 _02249_ _02251_ vssd1 vssd1 vccd1 vccd1 _00029_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07052__B _01226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07467_ genblk2\[8\].wave_shpr.div.busy _02196_ vssd1 vssd1 vccd1 vccd1 _02197_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_146_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_64_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_147_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09206_ _02171_ vssd1 vssd1 vccd1 vccd1 _03831_ sky130_fd_sc_hd__buf_8
XFILLER_0_151_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06493__A1 _01197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06418_ _01361_ vssd1 vssd1 vccd1 vccd1 _01362_ sky130_fd_sc_hd__buf_4
XANTENNA__08164__A _01181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07398_ _02091_ _02144_ _02145_ vssd1 vssd1 vccd1 vccd1 _02146_ sky130_fd_sc_hd__and3_1
X_09137_ genblk2\[0\].wave_shpr.div.b1\[11\] genblk2\[0\].wave_shpr.div.acc\[11\]
+ vssd1 vssd1 vccd1 vccd1 _03785_ sky130_fd_sc_hd__and2b_1
XFILLER_0_45_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06349_ genblk1\[0\].osc.clkdiv_C.cnt\[15\] _01295_ vssd1 vssd1 vccd1 vccd1 _01296_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_44_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09068_ _03725_ vssd1 vssd1 vccd1 vccd1 _03726_ sky130_fd_sc_hd__buf_8
X_08019_ genblk1\[6\].osc.clkdiv_C.cnt\[8\] _01732_ _02725_ _01753_ vssd1 vssd1 vccd1
+ vccd1 _02726_ sky130_fd_sc_hd__o2bb2a_1
Xhold660 genblk2\[11\].wave_shpr.div.acc\[17\] vssd1 vssd1 vccd1 vccd1 net878 sky130_fd_sc_hd__dlygate4sd3_1
Xhold671 genblk2\[0\].wave_shpr.div.acc\[12\] vssd1 vssd1 vccd1 vccd1 net889 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08611__B _02223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold682 genblk2\[6\].wave_shpr.div.acc\[11\] vssd1 vssd1 vccd1 vccd1 net900 sky130_fd_sc_hd__dlygate4sd3_1
X_11030_ genblk2\[6\].wave_shpr.div.acc\[9\] _05111_ _05105_ vssd1 vssd1 vccd1 vccd1
+ _05112_ sky130_fd_sc_hd__mux2_1
Xhold693 _00571_ vssd1 vssd1 vccd1 vccd1 net911 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06412__A _01226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07745__A1 genblk1\[1\].osc.clkdiv_C.cnt\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07745__B2 genblk1\[1\].osc.clkdiv_C.cnt\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12981_ clknet_leaf_124_clk _00310_ net75 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.quo\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09498__A1 _01327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11932_ genblk2\[10\].wave_shpr.div.b1\[4\] genblk2\[10\].wave_shpr.div.acc\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05754_ sky130_fd_sc_hd__and2b_1
XFILLER_0_87_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11863_ genblk2\[9\].wave_shpr.div.acc\[16\] _05699_ _05673_ vssd1 vssd1 vccd1 vccd1
+ _05700_ sky130_fd_sc_hd__mux2_1
XANTENNA__09869__S _04214_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10814_ _04855_ _04959_ _04960_ _04858_ net1154 vssd1 vssd1 vccd1 vccd1 _00598_ sky130_fd_sc_hd__a32o_1
X_13602_ clknet_leaf_77_clk _00917_ net209 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.acc\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11794_ _05646_ _05573_ genblk2\[9\].wave_shpr.div.b1\[0\] vssd1 vssd1 vccd1 vccd1
+ _05647_ sky130_fd_sc_hd__or3b_1
XFILLER_0_27_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10745_ net772 _04910_ _04907_ vssd1 vssd1 vccd1 vccd1 _04911_ sky130_fd_sc_hd__mux2_1
X_13533_ clknet_leaf_81_clk _00848_ net199 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.i\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__09670__A1 _04045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_40_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13464_ clknet_leaf_83_clk _00781_ net203 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.b1\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10676_ _04672_ genblk1\[5\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 _04865_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_125_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12415_ genblk2\[11\].wave_shpr.div.acc\[16\] _06083_ _06055_ vssd1 vssd1 vccd1 vccd1
+ _06084_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_523 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13395_ clknet_leaf_116_clk _00714_ net140 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10109__A _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12346_ genblk2\[11\].wave_shpr.div.b1\[0\] genblk2\[11\].wave_shpr.div.acc\[0\]
+ _05982_ vssd1 vssd1 vccd1 vccd1 _06031_ sky130_fd_sc_hd__nand3_1
XFILLER_0_23_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12309__B2 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12277_ net1274 _02001_ _05994_ vssd1 vssd1 vccd1 vccd1 _06000_ sky130_fd_sc_hd__mux2_1
XANTENNA__12324__A _03689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07418__A _02160_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11228_ net302 _05251_ _05248_ net492 _05252_ vssd1 vssd1 vccd1 vccd1 _00720_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11159_ genblk2\[7\].wave_shpr.div.acc\[22\] _05218_ vssd1 vssd1 vccd1 vccd1 _05219_
+ sky130_fd_sc_hd__or2_2
XFILLER_0_65_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06976__B _01811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_147_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08370_ _03054_ _03075_ _03076_ vssd1 vssd1 vccd1 vccd1 _03077_ sky130_fd_sc_hd__or3_2
XFILLER_0_58_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07321_ genblk1\[11\].osc.clkdiv_C.cnt\[15\] _01359_ vssd1 vssd1 vccd1 vccd1 _02085_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06475__A1 genblk1\[1\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07600__B net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07252_ genblk1\[10\].osc.clkdiv_C.cnt\[2\] genblk1\[10\].osc.clkdiv_C.cnt\[1\] genblk1\[10\].osc.clkdiv_C.cnt\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02032_ sky130_fd_sc_hd__and3_1
XFILLER_0_45_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06203_ PWM.counter\[6\] _01164_ vssd1 vssd1 vccd1 vccd1 _01167_ sky130_fd_sc_hd__or2_1
XANTENNA__08415__C _02365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07183_ genblk1\[9\].osc.clkdiv_C.cnt\[9\] _01972_ vssd1 vssd1 vccd1 vccd1 _01974_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_60_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06227__A1 _01174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06134_ _01104_ _01105_ vssd1 vssd1 vccd1 vccd1 _01106_ sky130_fd_sc_hd__nand2_1
XANTENNA__09808__A _04247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10453__S _04704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09824_ net315 _04257_ _04259_ net480 _04262_ vssd1 vssd1 vccd1 vccd1 _00306_ sky130_fd_sc_hd__a221o_1
XANTENNA__07047__B _01223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09755_ genblk2\[3\].wave_shpr.div.b1\[1\] _04225_ _04039_ vssd1 vssd1 vccd1 vccd1
+ _04226_ sky130_fd_sc_hd__mux2_1
X_06967_ genblk1\[7\].osc.clkdiv_C.cnt\[7\] _01574_ _01802_ genblk1\[7\].osc.clkdiv_C.cnt\[6\]
+ vssd1 vssd1 vccd1 vccd1 _01803_ sky130_fd_sc_hd__a22o_1
X_08706_ _03113_ _03116_ genblk2\[2\].wave_shpr.div.fin_quo\[3\] vssd1 vssd1 vccd1
+ vccd1 _03413_ sky130_fd_sc_hd__a21oi_1
X_09686_ genblk2\[2\].wave_shpr.div.acc\[7\] genblk2\[2\].wave_shpr.div.b1\[7\] vssd1
+ vssd1 vccd1 vccd1 _04166_ sky130_fd_sc_hd__or2b_1
XTAP_2106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08159__A _01489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06898_ genblk1\[6\].osc.clkdiv_C.cnt\[6\] _01367_ _01750_ genblk1\[6\].osc.clkdiv_C.cnt\[7\]
+ _01751_ vssd1 vssd1 vccd1 vccd1 _01752_ sky130_fd_sc_hd__a221o_1
XTAP_2117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08637_ _02592_ _03342_ _03343_ _02636_ vssd1 vssd1 vccd1 vccd1 _03344_ sky130_fd_sc_hd__a211o_1
XTAP_2139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08568_ _03263_ _03273_ _03274_ vssd1 vssd1 vccd1 vccd1 _03275_ sky130_fd_sc_hd__nand3_1
XFILLER_0_49_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07519_ _01163_ PWM.final_sample_in\[4\] _02233_ _02238_ vssd1 vssd1 vccd1 vccd1
+ _02239_ sky130_fd_sc_hd__a22o_1
Xfanout43 net44 vssd1 vssd1 vccd1 vccd1 net43 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_732 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08499_ _02547_ _02586_ _02588_ vssd1 vssd1 vccd1 vccd1 _03206_ sky130_fd_sc_hd__a21o_1
XFILLER_0_76_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout54 net58 vssd1 vssd1 vccd1 vccd1 net54 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10628__S _04834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout65 net68 vssd1 vssd1 vccd1 vccd1 net65 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout76 net84 vssd1 vssd1 vccd1 vccd1 net76 sky130_fd_sc_hd__clkbuf_4
X_10530_ _00012_ _04758_ net1160 vssd1 vssd1 vccd1 vccd1 _04760_ sky130_fd_sc_hd__a21oi_1
Xfanout87 net88 vssd1 vssd1 vccd1 vccd1 net87 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07663__B1 _01241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout98 net127 vssd1 vssd1 vccd1 vccd1 net98 sky130_fd_sc_hd__buf_2
XFILLER_0_134_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10461_ genblk2\[4\].wave_shpr.div.acc\[9\] _04710_ _04704_ vssd1 vssd1 vccd1 vccd1
+ _04711_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06218__A1 _01174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12200_ genblk2\[11\].wave_shpr.div.acc\[4\] genblk2\[11\].wave_shpr.div.b1\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05938_ sky130_fd_sc_hd__or2b_1
XFILLER_0_33_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13180_ clknet_leaf_130_clk _00505_ net68 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.acc\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_115_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10392_ net637 _04661_ _04663_ genblk2\[4\].wave_shpr.div.quo\[12\] _04664_ vssd1
+ vssd1 vccd1 vccd1 _00472_ sky130_fd_sc_hd__a221o_1
X_12131_ net945 _05876_ _05883_ _05886_ vssd1 vssd1 vccd1 vccd1 _00989_ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12062_ _05835_ genblk1\[10\].osc.clkdiv_C.cnt\[13\] vssd1 vssd1 vccd1 vccd1 _05836_
+ sky130_fd_sc_hd__and2_1
Xhold490 genblk2\[5\].wave_shpr.div.b1\[6\] vssd1 vssd1 vccd1 vccd1 net708 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06142__A net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11013_ genblk2\[6\].wave_shpr.div.acc\[5\] _05098_ _05023_ vssd1 vssd1 vccd1 vccd1
+ _05099_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12964_ clknet_leaf_111_clk _00293_ net130 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.quo\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_11915_ genblk2\[10\].wave_shpr.div.acc\[11\] genblk2\[10\].wave_shpr.div.b1\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05737_ sky130_fd_sc_hd__or2b_1
XTAP_2640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12895_ clknet_leaf_32_clk _00226_ net99 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.quo\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_51_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11846_ _05595_ _05686_ vssd1 vssd1 vccd1 vccd1 _05687_ sky130_fd_sc_hd__xnor2_1
XTAP_2695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11777_ _04676_ _02268_ vssd1 vssd1 vccd1 vccd1 _05638_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06457__A1 genblk1\[1\].osc.clkdiv_C.cnt\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10728_ genblk2\[5\].wave_shpr.div.acc\[5\] _04897_ _04821_ vssd1 vssd1 vccd1 vccd1
+ _04898_ sky130_fd_sc_hd__mux2_1
X_13516_ clknet_leaf_78_clk _00833_ net208 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.acc\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10659_ net745 _04853_ _04857_ net882 vssd1 vssd1 vccd1 vccd1 _00546_ sky130_fd_sc_hd__a22o_1
X_13447_ clknet_leaf_90_clk _00764_ net144 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.i\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_3_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09946__A2 _04253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13378_ clknet_leaf_81_clk _00697_ net205 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.b1\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10781__B _04880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11753__A2 _05623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12329_ net509 _06014_ _06015_ net510 _06022_ vssd1 vssd1 vccd1 vccd1 _01051_ sky130_fd_sc_hd__a221o_1
XANTENNA__07148__A genblk1\[9\].osc.clkdiv_C.cnt\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07870_ _02221_ _02510_ _02576_ vssd1 vssd1 vccd1 vccd1 _02577_ sky130_fd_sc_hd__o21bai_1
X_06821_ net27 vssd1 vssd1 vccd1 vccd1 _01693_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__11269__A1 _05248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09540_ _04058_ _02444_ vssd1 vssd1 vccd1 vccd1 _04061_ sky130_fd_sc_hd__nor2_1
X_06752_ genblk1\[4\].osc.clkdiv_C.cnt\[9\] _01627_ vssd1 vssd1 vccd1 vccd1 _01633_
+ sky130_fd_sc_hd__or2_1
X_09471_ _01418_ vssd1 vssd1 vccd1 vccd1 _04023_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06683_ _01566_ _01567_ _01569_ _01572_ vssd1 vssd1 vccd1 vccd1 _01573_ sky130_fd_sc_hd__or4b_1
XFILLER_0_92_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08422_ _03011_ _03128_ vssd1 vssd1 vccd1 vccd1 _03129_ sky130_fd_sc_hd__and2b_1
XFILLER_0_25_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10492__A2 _04715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_762 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_447 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08353_ _03058_ _03059_ _02798_ vssd1 vssd1 vccd1 vccd1 _03060_ sky130_fd_sc_hd__o21a_1
XFILLER_0_19_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout142_A net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07304_ genblk1\[11\].osc.clkdiv_C.cnt\[5\] _02064_ _01925_ genblk1\[11\].osc.clkdiv_C.cnt\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02068_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_117_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08284_ _02984_ _02989_ _02990_ vssd1 vssd1 vccd1 vccd1 _02991_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_116_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07235_ genblk1\[10\].osc.clkdiv_C.cnt\[16\] _02016_ vssd1 vssd1 vccd1 vccd1 _02017_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_26_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11787__B genblk1\[9\].osc.clkdiv_C.cnt\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07166_ genblk1\[9\].osc.clkdiv_C.cnt\[4\] _01960_ vssd1 vssd1 vccd1 vccd1 _01962_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06117_ net380 _01087_ net407 vssd1 vssd1 vccd1 vccd1 _01092_ sky130_fd_sc_hd__a21oi_1
X_07097_ _01887_ _01904_ vssd1 vssd1 vccd1 vccd1 _01905_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08161__B _01498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout200 net210 vssd1 vssd1 vccd1 vccd1 net200 sky130_fd_sc_hd__buf_2
Xfanout211 net212 vssd1 vssd1 vccd1 vccd1 net211 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10911__S _04848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09807_ genblk2\[2\].wave_shpr.div.quo\[8\] _04248_ _04252_ net275 vssd1 vssd1 vccd1
+ vccd1 _00299_ sky130_fd_sc_hd__a22o_1
X_07999_ _01200_ genblk1\[6\].osc.clkdiv_C.cnt\[15\] _01361_ _02704_ _02705_ vssd1
+ vssd1 vccd1 vccd1 _02706_ sky130_fd_sc_hd__o311a_1
XANTENNA__07581__C1 genblk1\[9\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09738_ _04216_ vssd1 vssd1 vccd1 vccd1 _00266_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_fanout55_A net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09669_ _04151_ vssd1 vssd1 vccd1 vccd1 _04152_ sky130_fd_sc_hd__inv_2
XFILLER_0_69_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11700_ genblk2\[9\].wave_shpr.div.b1\[10\] genblk2\[9\].wave_shpr.div.acc\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05592_ sky130_fd_sc_hd__and2b_1
XTAP_1235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12680_ clknet_leaf_120_clk genblk1\[7\].osc.clkdiv_C.next_cnt\[11\] net82 vssd1
+ vssd1 vccd1 vccd1 genblk1\[7\].osc.clkdiv_C.cnt\[11\] sky130_fd_sc_hd__dfrtp_4
XTAP_1246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11631_ _05410_ _05416_ vssd1 vssd1 vccd1 vccd1 _05534_ sky130_fd_sc_hd__and2b_1
XTAP_1279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_108_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11562_ _05379_ _05481_ vssd1 vssd1 vccd1 vccd1 _05482_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_92_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06137__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10513_ genblk2\[4\].wave_shpr.div.acc\[23\] _04620_ _04748_ vssd1 vssd1 vccd1 vccd1
+ _04749_ sky130_fd_sc_hd__a21o_1
X_13301_ clknet_leaf_84_clk _00622_ net202 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.b1\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11493_ _02152_ genblk2\[8\].wave_shpr.div.busy _02196_ vssd1 vssd1 vccd1 vccd1 _05443_
+ sky130_fd_sc_hd__and3_1
X_13232_ clknet_leaf_15_clk net501 net73 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.quo\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10444_ genblk2\[4\].wave_shpr.div.acc\[5\] _04697_ _04623_ vssd1 vssd1 vccd1 vccd1
+ _04698_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13163_ clknet_leaf_114_clk _00488_ net67 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.acc\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10375_ genblk2\[4\].wave_shpr.div.quo\[4\] _04652_ _04656_ net732 vssd1 vssd1 vccd1
+ vccd1 _00463_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10943__B1 _05056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12114_ _05766_ _05738_ vssd1 vssd1 vccd1 vccd1 _05873_ sky130_fd_sc_hd__or2b_1
XFILLER_0_20_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13094_ clknet_leaf_1_clk _00421_ net38 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.acc\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_12045_ _05819_ genblk1\[10\].osc.clkdiv_C.cnt\[5\] vssd1 vssd1 vccd1 vccd1 _05827_
+ sky130_fd_sc_hd__and2_1
XANTENNA__12160__A2 _05818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06600__A _01241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10122__A _04058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12947_ clknet_leaf_125_clk _00276_ net69 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.b1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12878_ clknet_leaf_119_clk net685 net143 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.quo\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07431__A _02152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11829_ genblk2\[9\].wave_shpr.div.acc\[8\] _05672_ _05673_ vssd1 vssd1 vccd1 vccd1
+ _05674_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07627__B1 _01256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_3_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07020_ net1189 _01841_ _01843_ vssd1 vssd1 vccd1 vccd1 genblk1\[7\].osc.clkdiv_C.next_cnt\[12\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_141_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08971_ _03656_ _03523_ _01098_ vssd1 vssd1 vccd1 vccd1 _03658_ sky130_fd_sc_hd__a21o_1
X_07922_ _02624_ _02626_ _02627_ _02628_ vssd1 vssd1 vccd1 vccd1 _02629_ sky130_fd_sc_hd__o211a_1
Xhold19 genblk2\[8\].wave_shpr.div.quo\[14\] vssd1 vssd1 vccd1 vccd1 net237 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07606__A net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07853_ _02558_ _02559_ _02424_ vssd1 vssd1 vccd1 vccd1 _02560_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06510__A _01349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06804_ genblk1\[5\].osc.clkdiv_C.cnt\[15\] _01362_ genblk1\[5\].osc.clkdiv_C.cnt\[17\]
+ vssd1 vssd1 vccd1 vccd1 _01676_ sky130_fd_sc_hd__a21o_1
X_07784_ genblk1\[0\].osc.clkdiv_C.cnt\[5\] _02486_ _02489_ _02490_ vssd1 vssd1 vccd1
+ vccd1 _02491_ sky130_fd_sc_hd__o31ai_1
XANTENNA__12439__B1 _03944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08107__A1 _01192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09821__A _04069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06735_ _01619_ vssd1 vssd1 vccd1 vccd1 genblk1\[4\].osc.clkdiv_C.next_cnt\[5\] sky130_fd_sc_hd__clkbuf_1
X_09523_ net610 _04048_ _04045_ net517 _04050_ vssd1 vssd1 vccd1 vccd1 _00217_ sky130_fd_sc_hd__a221o_1
XANTENNA__08658__A2 _02467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09454_ genblk2\[1\].wave_shpr.div.fin_quo\[3\] genblk2\[1\].wave_shpr.div.quo\[2\]
+ _00007_ vssd1 vssd1 vccd1 vccd1 _04015_ sky130_fd_sc_hd__mux2_1
X_06666_ _01230_ _01221_ _01223_ vssd1 vssd1 vccd1 vccd1 _01556_ sky130_fd_sc_hd__a21o_4
XPHY_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08405_ genblk1\[2\].osc.clkdiv_C.cnt\[16\] _01578_ _03111_ genblk1\[2\].osc.clkdiv_C.cnt\[17\]
+ vssd1 vssd1 vccd1 vccd1 _03112_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_93_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09385_ _00004_ _03949_ net1163 vssd1 vssd1 vccd1 vccd1 _03951_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_143_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_220 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06597_ genblk1\[3\].osc.clkdiv_C.cnt\[16\] _01197_ vssd1 vssd1 vccd1 vccd1 _01505_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_19_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08336_ _02734_ _02737_ genblk2\[6\].wave_shpr.div.fin_quo\[4\] vssd1 vssd1 vccd1
+ vccd1 _03043_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_426 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08267_ genblk2\[11\].wave_shpr.div.fin_quo\[4\] net33 _02350_ _02354_ _02222_ vssd1
+ vssd1 vccd1 vccd1 _02974_ sky130_fd_sc_hd__a41o_1
XFILLER_0_61_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07218_ genblk1\[10\].osc.clkdiv_C.cnt\[14\] _01246_ _01442_ genblk1\[10\].osc.clkdiv_C.cnt\[13\]
+ _01999_ vssd1 vssd1 vccd1 vccd1 _02000_ sky130_fd_sc_hd__a221o_1
XANTENNA__09268__A _02171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08198_ _02902_ _02903_ _02904_ _02360_ vssd1 vssd1 vccd1 vccd1 _02905_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_61_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07149_ genblk1\[9\].osc.clkdiv_C.cnt\[12\] _01799_ _01947_ genblk1\[9\].osc.clkdiv_C.cnt\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01949_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_132_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06404__B _01327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10160_ genblk2\[3\].wave_shpr.div.acc\[5\] _04497_ _04420_ vssd1 vssd1 vccd1 vccd1
+ _04498_ sky130_fd_sc_hd__mux2_1
XFILLER_0_100_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10091_ genblk2\[3\].wave_shpr.div.quo\[4\] _04452_ _04456_ net779 vssd1 vssd1 vccd1
+ vccd1 _00379_ sky130_fd_sc_hd__a22o_1
XFILLER_0_16_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12801_ clknet_leaf_59_clk net570 net193 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.quo\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10993_ genblk2\[6\].wave_shpr.div.acc\[1\] _05022_ vssd1 vssd1 vccd1 vccd1 _05083_
+ sky130_fd_sc_hd__or2_1
XANTENNA__11102__B1 _03855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12732_ clknet_leaf_38_clk genblk1\[10\].osc.clkdiv_C.next_cnt\[9\] net115 vssd1
+ vssd1 vccd1 vccd1 genblk1\[10\].osc.clkdiv_C.cnt\[9\] sky130_fd_sc_hd__dfrtp_4
XTAP_1021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07857__B1 _02316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold903_A genblk2\[1\].wave_shpr.div.b1\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_52_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12663_ clknet_leaf_26_clk genblk1\[6\].osc.clkdiv_C.next_cnt\[12\] net88 vssd1 vssd1
+ vccd1 vccd1 genblk1\[6\].osc.clkdiv_C.cnt\[12\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_84_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09877__S _04214_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11614_ genblk2\[8\].wave_shpr.div.acc\[15\] _05521_ _05493_ vssd1 vssd1 vccd1 vccd1
+ _05522_ sky130_fd_sc_hd__mux2_1
X_12594_ clknet_leaf_12_clk genblk1\[2\].osc.clkdiv_C.next_cnt\[15\] net52 vssd1 vssd1
+ vccd1 vccd1 genblk1\[2\].osc.clkdiv_C.cnt\[15\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_53_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11545_ _05464_ genblk1\[8\].osc.clkdiv_C.cnt\[16\] vssd1 vssd1 vccd1 vccd1 _05470_
+ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_131_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_131_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_clkbuf_leaf_67_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13760__RESET_B net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11476_ _05435_ vssd1 vssd1 vccd1 vccd1 _00785_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_123_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_110_clk_A clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_40_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10427_ _04585_ _04684_ vssd1 vssd1 vccd1 vccd1 _04685_ sky130_fd_sc_hd__nor2_1
X_13215_ clknet_leaf_6_clk _00538_ net48 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.b1\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_892 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10358_ _03704_ net800 _04647_ vssd1 vssd1 vccd1 vccd1 _00455_ sky130_fd_sc_hd__a21o_1
X_13146_ clknet_leaf_121_clk _00471_ net81 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.quo\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13077_ clknet_leaf_125_clk _00404_ net62 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.acc\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10289_ _04573_ _04599_ _04600_ vssd1 vssd1 vccd1 vccd1 _04601_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_125_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12332__A _03833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12028_ genblk2\[10\].wave_shpr.div.quo\[6\] _05813_ _05817_ net555 vssd1 vssd1 vccd1
+ vccd1 _00955_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06984__B _01819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06520_ _01438_ _01443_ _01444_ _01445_ vssd1 vssd1 vccd1 vccd1 _01446_ sky130_fd_sc_hd__or4_1
XFILLER_0_87_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07312__A2 _01210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06451_ _01373_ _01387_ _01388_ vssd1 vssd1 vccd1 vccd1 genblk1\[1\].osc.clkdiv_C.next_cnt\[6\]
+ sky130_fd_sc_hd__nor3_1
XANTENNA__09787__S _04238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09170_ _03811_ vssd1 vssd1 vccd1 vccd1 _00103_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06382_ _01229_ _01325_ vssd1 vssd1 vccd1 vccd1 _01326_ sky130_fd_sc_hd__nand2_4
X_08121_ genblk1\[4\].osc.clkdiv_C.cnt\[3\] _01439_ _02827_ vssd1 vssd1 vccd1 vccd1
+ _02828_ sky130_fd_sc_hd__a21o_1
XFILLER_0_7_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_122_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_122_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_114_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08052_ _01489_ genblk1\[5\].osc.clkdiv_C.cnt\[9\] net37 _01667_ genblk1\[5\].osc.clkdiv_C.cnt\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02759_ sky130_fd_sc_hd__a32o_1
XFILLER_0_113_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07003_ genblk1\[7\].osc.clkdiv_C.cnt\[6\] _01830_ vssd1 vssd1 vccd1 vccd1 _01833_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__08576__A1 _02525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09816__A _04058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10461__S _04704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08954_ sig_norm.quo\[3\] _03643_ _02248_ vssd1 vssd1 vccd1 vccd1 _03644_ sky130_fd_sc_hd__mux2_1
XANTENNA__09525__B1 _04045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07905_ genblk1\[8\].osc.clkdiv_C.cnt\[10\] _01870_ vssd1 vssd1 vccd1 vccd1 _02612_
+ sky130_fd_sc_hd__xnor2_1
X_08885_ sig_norm.acc\[10\] _03590_ vssd1 vssd1 vccd1 vccd1 _03591_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_80 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_99_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07055__B _01430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07836_ genblk2\[0\].wave_shpr.div.fin_quo\[4\] _02510_ _02512_ _02261_ vssd1 vssd1
+ vccd1 vccd1 _02543_ sky130_fd_sc_hd__a31o_1
X_07767_ genblk1\[0\].osc.clkdiv_C.cnt\[15\] _01309_ _01208_ genblk1\[0\].osc.clkdiv_C.cnt\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02474_ sky130_fd_sc_hd__o22a_1
X_09506_ _02170_ genblk2\[1\].wave_shpr.div.busy _02157_ vssd1 vssd1 vccd1 vccd1 _04044_
+ sky130_fd_sc_hd__and3_1
X_06718_ _01605_ vssd1 vssd1 vccd1 vccd1 _01606_ sky130_fd_sc_hd__inv_2
X_07698_ genblk2\[10\].wave_shpr.div.fin_quo\[5\] vssd1 vssd1 vccd1 vccd1 _02405_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_63_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09437_ _03956_ _03999_ _04000_ vssd1 vssd1 vccd1 vccd1 _04001_ sky130_fd_sc_hd__a21oi_1
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06649_ genblk1\[3\].osc.clkdiv_C.cnt\[12\] _01543_ vssd1 vssd1 vccd1 vccd1 _01545_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_137_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09368_ genblk2\[0\].wave_shpr.div.acc\[25\] _03802_ genblk2\[0\].wave_shpr.div.acc\[24\]
+ genblk2\[0\].wave_shpr.div.acc\[26\] vssd1 vssd1 vccd1 vccd1 _03938_ sky130_fd_sc_hd__or4b_1
XFILLER_0_93_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08319_ genblk2\[9\].wave_shpr.div.fin_quo\[3\] _02303_ _02263_ _02316_ vssd1 vssd1
+ vccd1 vccd1 _03026_ sky130_fd_sc_hd__a31o_1
XFILLER_0_151_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_113_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_113_clk
+ sky130_fd_sc_hd__clkbuf_16
X_09299_ _03777_ _03756_ vssd1 vssd1 vccd1 vccd1 _03887_ sky130_fd_sc_hd__or2b_1
XFILLER_0_90_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_117_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11321__A _05249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11330_ _05211_ _05166_ vssd1 vssd1 vccd1 vccd1 _05322_ sky130_fd_sc_hd__or2b_1
XFILLER_0_22_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11261_ net534 _05245_ _05249_ genblk2\[7\].wave_shpr.div.quo\[23\] _05270_ vssd1
+ vssd1 vccd1 vccd1 _00735_ sky130_fd_sc_hd__a221o_1
XANTENNA__08016__B1 _01739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10212_ net657 _04518_ _04522_ _04537_ vssd1 vssd1 vccd1 vccd1 _00419_ sky130_fd_sc_hd__a22o_1
X_13000_ clknet_leaf_132_clk _00329_ net63 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.acc\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07568__A2_N _01349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11192_ _05235_ vssd1 vssd1 vccd1 vccd1 _00701_ sky130_fd_sc_hd__clkbuf_1
X_10143_ genblk2\[3\].wave_shpr.div.acc\[1\] _04484_ _04420_ vssd1 vssd1 vccd1 vccd1
+ _04485_ sky130_fd_sc_hd__mux2_1
XANTENNA__09516__B1 _04047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10074_ _04447_ vssd1 vssd1 vccd1 vccd1 _00371_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13764_ clknet_leaf_69_clk _01075_ net214 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.acc\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10976_ _05059_ genblk1\[6\].osc.clkdiv_C.cnt\[12\] vssd1 vssd1 vccd1 vccd1 _05073_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_57_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12715_ clknet_leaf_54_clk genblk1\[9\].osc.clkdiv_C.next_cnt\[10\] net175 vssd1
+ vssd1 vccd1 vccd1 genblk1\[9\].osc.clkdiv_C.cnt\[10\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_85_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13695_ clknet_leaf_45_clk _01006_ net188 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.i\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12646_ clknet_leaf_24_clk genblk1\[5\].osc.clkdiv_C.next_cnt\[13\] net92 vssd1 vssd1
+ vccd1 vccd1 genblk1\[5\].osc.clkdiv_C.cnt\[13\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_81_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07058__A1 genblk1\[8\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_104_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_104_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_5_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07058__B2 genblk1\[8\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12577_ clknet_leaf_21_clk genblk1\[1\].osc.clkdiv_C.next_cnt\[16\] net95 vssd1 vssd1
+ vccd1 vccd1 genblk1\[1\].osc.clkdiv_C.cnt\[16\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_108_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11231__A _05074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_418 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11528_ _05450_ genblk1\[8\].osc.clkdiv_C.cnt\[8\] vssd1 vssd1 vccd1 vccd1 _05461_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_40_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold308 genblk2\[9\].wave_shpr.div.quo\[8\] vssd1 vssd1 vccd1 vccd1 net526 sky130_fd_sc_hd__buf_1
XANTENNA__08007__B1 _01735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold319 genblk2\[1\].wave_shpr.div.quo\[12\] vssd1 vssd1 vccd1 vccd1 net537 sky130_fd_sc_hd__dlygate4sd3_1
X_11459_ _05426_ vssd1 vssd1 vccd1 vccd1 _00777_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08558__A1 genblk2\[8\].wave_shpr.div.fin_quo\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13129_ clknet_leaf_3_clk _00454_ net46 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.b1\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07156__A genblk1\[9\].osc.clkdiv_C.cnt\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1008 genblk2\[10\].wave_shpr.div.acc\[25\] vssd1 vssd1 vccd1 vccd1 net1226 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_84_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1019 genblk1\[3\].osc.clkdiv_C.cnt\[15\] vssd1 vssd1 vccd1 vccd1 net1237 sky130_fd_sc_hd__dlygate4sd3_1
X_08670_ _03366_ _03376_ vssd1 vssd1 vccd1 vccd1 _03377_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09371__A _02170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07621_ genblk1\[11\].osc.clkdiv_C.cnt\[6\] _01430_ _02326_ _02327_ vssd1 vssd1 vccd1
+ vccd1 _02328_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_49_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07552_ _02259_ vssd1 vssd1 vccd1 vccd1 _00037_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07603__B net32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06503_ genblk1\[2\].osc.clkdiv_C.cnt\[12\] _01411_ _01415_ _01419_ _01428_ vssd1
+ vssd1 vccd1 vccd1 _01429_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_76_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12290__A1 _01249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07483_ _02208_ vssd1 vssd1 vccd1 vccd1 _00002_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_29_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09222_ genblk2\[0\].wave_shpr.div.quo\[3\] _03836_ _03840_ net558 vssd1 vssd1 vccd1
+ vccd1 _00126_ sky130_fd_sc_hd__a22o_1
X_06434_ _01374_ _01375_ _01376_ vssd1 vssd1 vccd1 vccd1 _01377_ sky130_fd_sc_hd__and3_1
XFILLER_0_146_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09153_ genblk2\[0\].wave_shpr.div.acc\[22\] genblk2\[0\].wave_shpr.div.acc\[21\]
+ genblk2\[0\].wave_shpr.div.acc\[20\] _03800_ vssd1 vssd1 vccd1 vccd1 _03801_ sky130_fd_sc_hd__or4_1
XANTENNA__07049__A1 genblk1\[8\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06365_ _01171_ vssd1 vssd1 vccd1 vccd1 _01309_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_99_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08104_ genblk1\[4\].osc.clkdiv_C.cnt\[9\] _01323_ _01592_ genblk1\[4\].osc.clkdiv_C.cnt\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02811_ sky130_fd_sc_hd__o22a_1
XFILLER_0_72_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09084_ _03735_ vssd1 vssd1 vccd1 vccd1 _03736_ sky130_fd_sc_hd__buf_8
XFILLER_0_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06235__A _01196_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06296_ _01238_ _01257_ vssd1 vssd1 vccd1 vccd1 _01258_ sky130_fd_sc_hd__or2_2
XFILLER_0_31_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_31_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08035_ _02221_ _02733_ vssd1 vssd1 vccd1 vccd1 _02742_ sky130_fd_sc_hd__nor2_2
XFILLER_0_130_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold820 genblk2\[5\].wave_shpr.div.acc\[24\] vssd1 vssd1 vccd1 vccd1 net1038 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold831 genblk2\[0\].wave_shpr.div.acc\[8\] vssd1 vssd1 vccd1 vccd1 net1049 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12345__A2 net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold842 genblk2\[9\].wave_shpr.div.acc\[16\] vssd1 vssd1 vccd1 vccd1 net1060 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold853 genblk2\[4\].wave_shpr.div.b1\[0\] vssd1 vssd1 vccd1 vccd1 net1071 sky130_fd_sc_hd__dlygate4sd3_1
Xhold864 genblk2\[0\].wave_shpr.div.acc\[25\] vssd1 vssd1 vccd1 vccd1 net1082 sky130_fd_sc_hd__dlygate4sd3_1
Xhold875 genblk2\[6\].wave_shpr.div.acc\[16\] vssd1 vssd1 vccd1 vccd1 net1093 sky130_fd_sc_hd__dlygate4sd3_1
Xhold886 genblk1\[6\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 net1104 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold897 genblk1\[5\].osc.clkdiv_C.cnt\[15\] vssd1 vssd1 vccd1 vccd1 net1115 sky130_fd_sc_hd__dlygate4sd3_1
X_09986_ genblk2\[3\].wave_shpr.div.b1\[0\] _04380_ _04381_ vssd1 vssd1 vccd1 vccd1
+ _04382_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07772__A2 _01190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08937_ _01098_ _03550_ vssd1 vssd1 vccd1 vccd1 _03630_ sky130_fd_sc_hd__nor2_1
XANTENNA__06980__B1 _01574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10659__A2 _04853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08868_ _01156_ vssd1 vssd1 vccd1 vccd1 _03574_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07819_ _02525_ vssd1 vssd1 vccd1 vccd1 _02526_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08799_ _03500_ _03504_ _03427_ _03505_ vssd1 vssd1 vccd1 vccd1 _03506_ sky130_fd_sc_hd__o211a_1
XANTENNA__11316__A _05245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10830_ genblk2\[6\].wave_shpr.div.acc\[9\] genblk2\[6\].wave_shpr.div.b1\[9\] vssd1
+ vssd1 vccd1 vccd1 _04974_ sky130_fd_sc_hd__or2b_1
XFILLER_0_39_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10761_ _04806_ _04767_ vssd1 vssd1 vccd1 vccd1 _04923_ sky130_fd_sc_hd__or2b_1
XFILLER_0_109_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12281__A1 _02013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06129__B net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12500_ clknet_leaf_102_clk net429 net156 vssd1 vssd1 vccd1 vccd1 sig_norm.acc_next\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13480_ clknet_leaf_99_clk _00797_ net168 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.quo\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10692_ genblk2\[5\].wave_shpr.div.quo\[20\] _04861_ _04862_ net233 _04873_ vssd1
+ vssd1 vccd1 vccd1 _00563_ sky130_fd_sc_hd__a221o_1
XFILLER_0_48_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12431_ genblk2\[11\].wave_shpr.div.acc\[20\] _05978_ net20 vssd1 vssd1 vccd1 vccd1
+ _06095_ sky130_fd_sc_hd__or3_1
XFILLER_0_63_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_23_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12362_ net985 _06039_ _06040_ _06043_ vssd1 vssd1 vccd1 vccd1 _01063_ sky130_fd_sc_hd__a22o_1
XANTENNA__06145__A _01114_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06799__B1 _01304_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08063__C net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11313_ _05202_ _05308_ vssd1 vssd1 vccd1 vccd1 _05309_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_105_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12293_ _06008_ vssd1 vssd1 vccd1 vccd1 _01029_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11244_ _05260_ genblk1\[7\].osc.clkdiv_C.cnt\[7\] vssd1 vssd1 vccd1 vccd1 _05262_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_31_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08360__A _02885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10347__A1 _01658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07212__A1 _01308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11175_ genblk2\[7\].wave_shpr.div.fin_quo\[6\] net754 _00019_ vssd1 vssd1 vccd1
+ vccd1 _05229_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07763__A2 _02468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10126_ _04465_ genblk1\[3\].osc.clkdiv_C.cnt\[13\] vssd1 vssd1 vccd1 vccd1 _04474_
+ sky130_fd_sc_hd__and2_1
XANTENNA__06971__B1 _01805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10057_ net1225 _01329_ _04238_ vssd1 vssd1 vccd1 vccd1 _04438_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07920__C1 _01441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11226__A _05245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13747_ clknet_leaf_51_clk net413 net111 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.acc_next\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10959_ _05054_ vssd1 vssd1 vccd1 vccd1 _05064_ sky130_fd_sc_hd__buf_2
XFILLER_0_70_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13678_ clknet_leaf_42_clk _00991_ net125 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.acc\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12629_ clknet_leaf_120_clk genblk1\[4\].osc.clkdiv_C.next_cnt\[14\] net82 vssd1
+ vssd1 vccd1 vccd1 genblk1\[4\].osc.clkdiv_C.cnt\[14\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_5_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06150_ _01103_ _01111_ vssd1 vssd1 vccd1 vccd1 _01122_ sky130_fd_sc_hd__and2b_1
XFILLER_0_108_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold105 _00311_ vssd1 vssd1 vccd1 vccd1 net323 sky130_fd_sc_hd__dlygate4sd3_1
Xhold116 genblk2\[10\].wave_shpr.div.quo\[21\] vssd1 vssd1 vccd1 vccd1 net334 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold127 _00638_ vssd1 vssd1 vccd1 vccd1 net345 sky130_fd_sc_hd__dlygate4sd3_1
Xhold138 _01042_ vssd1 vssd1 vccd1 vccd1 net356 sky130_fd_sc_hd__dlygate4sd3_1
Xhold149 _00245_ vssd1 vssd1 vccd1 vccd1 net367 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10338__A1 _03831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09840_ genblk2\[2\].wave_shpr.div.quo\[22\] _04247_ _04259_ net261 _04271_ vssd1
+ vssd1 vccd1 vccd1 _00313_ sky130_fd_sc_hd__a221o_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08400__B1 _01591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09771_ _04235_ vssd1 vssd1 vccd1 vccd1 _00280_ sky130_fd_sc_hd__clkbuf_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06983_ _01436_ _01334_ vssd1 vssd1 vccd1 vccd1 _01819_ sky130_fd_sc_hd__nand2_2
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08722_ _02588_ _02546_ vssd1 vssd1 vccd1 vccd1 _03429_ sky130_fd_sc_hd__nor2_1
XANTENNA__07506__A2 _02221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08653_ _03313_ _03326_ vssd1 vssd1 vccd1 vccd1 _03360_ sky130_fd_sc_hd__and2b_1
XFILLER_0_14_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07604_ genblk2\[9\].wave_shpr.div.fin_quo\[7\] _02309_ _02310_ vssd1 vssd1 vccd1
+ vccd1 _02311_ sky130_fd_sc_hd__a21o_1
XTAP_1609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08584_ _03289_ _03290_ _02419_ vssd1 vssd1 vccd1 vccd1 _03291_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_95_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07535_ net279 _02249_ _01099_ vssd1 vssd1 vccd1 vccd1 _02251_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12263__A1 _01263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07466_ _02195_ genblk2\[8\].wave_shpr.div.i\[1\] genblk2\[8\].wave_shpr.div.i\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02196_ sky130_fd_sc_hd__or3b_1
XFILLER_0_147_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09205_ _03704_ net759 _03728_ vssd1 vssd1 vccd1 vccd1 _00119_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_45_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06417_ _01360_ vssd1 vssd1 vccd1 vccd1 _01361_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_91_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07397_ genblk1\[11\].osc.clkdiv_C.cnt\[16\] _02143_ vssd1 vssd1 vccd1 vccd1 _02145_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_151_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09136_ _03753_ _03782_ _03783_ vssd1 vssd1 vccd1 vccd1 _03784_ sky130_fd_sc_hd__a21o_1
XFILLER_0_44_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06348_ _01269_ _01294_ _01295_ vssd1 vssd1 vccd1 vccd1 genblk1\[0\].osc.clkdiv_C.next_cnt\[14\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_60_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09067_ _02155_ vssd1 vssd1 vccd1 vccd1 _03725_ sky130_fd_sc_hd__buf_2
X_06279_ _01237_ vssd1 vssd1 vccd1 vccd1 _01241_ sky130_fd_sc_hd__buf_4
XANTENNA__06607__A2_N _01513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07993__A2 _01484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08018_ _01739_ vssd1 vssd1 vccd1 vccd1 _02725_ sky130_fd_sc_hd__inv_2
XFILLER_0_130_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold650 genblk2\[10\].wave_shpr.div.acc\[4\] vssd1 vssd1 vccd1 vccd1 net868 sky130_fd_sc_hd__dlygate4sd3_1
Xhold661 genblk2\[5\].wave_shpr.div.quo\[1\] vssd1 vssd1 vccd1 vccd1 net879 sky130_fd_sc_hd__dlygate4sd3_1
Xhold672 genblk2\[3\].wave_shpr.div.acc\[7\] vssd1 vssd1 vccd1 vccd1 net890 sky130_fd_sc_hd__dlygate4sd3_1
Xhold683 genblk2\[4\].wave_shpr.div.acc\[13\] vssd1 vssd1 vccd1 vccd1 net901 sky130_fd_sc_hd__dlygate4sd3_1
Xhold694 genblk2\[9\].wave_shpr.div.acc\[15\] vssd1 vssd1 vccd1 vccd1 net912 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06412__B _01355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout85_A net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07745__A2 _01344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09969_ genblk2\[3\].wave_shpr.div.acc\[13\] genblk2\[3\].wave_shpr.div.b1\[13\]
+ vssd1 vssd1 vccd1 vccd1 _04365_ sky130_fd_sc_hd__or2b_1
X_12980_ clknet_leaf_14_clk _00309_ net72 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.quo\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_11931_ _05744_ _05751_ _05752_ vssd1 vssd1 vccd1 vccd1 _05753_ sky130_fd_sc_hd__a21oi_1
XTAP_2800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08170__A2 _01508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_24_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11862_ _05698_ _05603_ vssd1 vssd1 vccd1 vccd1 _05699_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13601_ clknet_leaf_77_clk _00916_ net209 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.acc\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10813_ genblk2\[5\].wave_shpr.div.i\[1\] genblk2\[5\].wave_shpr.div.i\[0\] genblk2\[5\].wave_shpr.div.i\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04960_ sky130_fd_sc_hd__nand3_1
X_11793_ _05610_ _05611_ vssd1 vssd1 vccd1 vccd1 _05646_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13532_ clknet_leaf_97_clk _00023_ net166 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.done
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10804__A2 _04858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10744_ _04797_ _04909_ vssd1 vssd1 vccd1 vccd1 _04910_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_82_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12006__A1 _01494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13463_ clknet_leaf_83_clk _00780_ net203 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.b1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10675_ net453 _04861_ _04862_ net500 _04864_ vssd1 vssd1 vccd1 vccd1 _00555_ sky130_fd_sc_hd__a221o_1
X_12414_ _05926_ _05972_ vssd1 vssd1 vccd1 vccd1 _06083_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13394_ clknet_leaf_116_clk net564 net145 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.quo\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12345_ _03819_ net1220 _00004_ genblk2\[11\].wave_shpr.div.acc\[0\] _06030_ vssd1
+ vssd1 vccd1 vccd1 _01059_ sky130_fd_sc_hd__o221a_1
XANTENNA__08630__B1 _02261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12309__A2 _03947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08090__A net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12276_ _05999_ vssd1 vssd1 vccd1 vccd1 _01021_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_120_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09186__A1 _03704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11227_ _05074_ genblk1\[7\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 _05252_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_120_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_120_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06322__B genblk1\[0\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11158_ genblk2\[7\].wave_shpr.div.acc\[21\] genblk2\[7\].wave_shpr.div.acc\[20\]
+ genblk2\[7\].wave_shpr.div.acc\[19\] _05217_ vssd1 vssd1 vccd1 vccd1 _05218_ sky130_fd_sc_hd__or4_1
X_10109_ _04268_ vssd1 vssd1 vccd1 vccd1 _04465_ sky130_fd_sc_hd__clkbuf_2
X_11089_ net1043 _05057_ _05055_ _05154_ vssd1 vssd1 vccd1 vccd1 _00679_ sky130_fd_sc_hd__a22o_1
XANTENNA__12340__A _03833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07434__A _02171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08449__B1 _02316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12245__A1 _05982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07320_ genblk1\[11\].osc.clkdiv_C.cnt\[4\] _01513_ _02076_ _02079_ _02083_ vssd1
+ vssd1 vccd1 vccd1 _02084_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_45_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09661__A2 _04048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07121__B1 _01855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07251_ _02031_ vssd1 vssd1 vccd1 vccd1 genblk1\[10\].osc.clkdiv_C.next_cnt\[1\]
+ sky130_fd_sc_hd__clkbuf_1
X_06202_ PWM.counter\[6\] _01164_ vssd1 vssd1 vccd1 vccd1 _01166_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07182_ _01953_ _01972_ _01973_ vssd1 vssd1 vccd1 vccd1 genblk1\[9\].osc.clkdiv_C.next_cnt\[8\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_42_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06133_ net8 net9 vssd1 vssd1 vccd1 vccd1 _01105_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11220__A2 _05246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07609__A _02222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06513__A _01213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12181__B1 _05818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07727__A2 _02433_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09823_ _04069_ genblk1\[2\].osc.clkdiv_C.cnt\[6\] vssd1 vssd1 vccd1 vccd1 _04262_
+ sky130_fd_sc_hd__and2_1
XANTENNA__06593__A2_N _01498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09754_ _01436_ _01925_ vssd1 vssd1 vccd1 vccd1 _04225_ sky130_fd_sc_hd__nand2_2
X_06966_ _01192_ _01245_ vssd1 vssd1 vccd1 vccd1 _01802_ sky130_fd_sc_hd__nand2_1
X_08705_ _03361_ _03378_ _03411_ vssd1 vssd1 vccd1 vccd1 _03412_ sky130_fd_sc_hd__a21o_1
X_09685_ genblk2\[2\].wave_shpr.div.acc\[8\] genblk2\[2\].wave_shpr.div.b1\[8\] vssd1
+ vssd1 vccd1 vccd1 _04165_ sky130_fd_sc_hd__or2b_1
XFILLER_0_96_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06897_ genblk1\[6\].osc.clkdiv_C.cnt\[6\] _01367_ _01750_ genblk1\[6\].osc.clkdiv_C.cnt\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01751_ sky130_fd_sc_hd__o22ai_1
XTAP_2107 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_93_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_93_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__08152__A2 _01500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2118 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2129 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08636_ _02216_ _02552_ genblk2\[8\].wave_shpr.div.fin_quo\[3\] vssd1 vssd1 vccd1
+ vccd1 _03343_ sky130_fd_sc_hd__and3_1
XTAP_1406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08567_ _02946_ _03272_ _03268_ vssd1 vssd1 vccd1 vccd1 _03274_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07998__B _01361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10909__S _04848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10247__B1 _04457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07518_ _02232_ PWM.final_sample_in\[3\] PWM.final_sample_in\[2\] _02234_ _02237_
+ vssd1 vssd1 vccd1 vccd1 _02238_ sky130_fd_sc_hd__a221o_1
XFILLER_0_64_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout44 net85 vssd1 vssd1 vccd1 vccd1 net44 sky130_fd_sc_hd__clkbuf_2
X_08498_ _03077_ _03203_ _03175_ _03202_ vssd1 vssd1 vccd1 vccd1 _03205_ sky130_fd_sc_hd__a211oi_1
XANTENNA__09652__A2 _04048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout55 net58 vssd1 vssd1 vccd1 vccd1 net55 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_147_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout66 net68 vssd1 vssd1 vccd1 vccd1 net66 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_91_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout77 net84 vssd1 vssd1 vccd1 vccd1 net77 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07663__A1 _01360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07449_ _02180_ _02153_ genblk2\[5\].wave_shpr.div.busy vssd1 vssd1 vccd1 vccd1 _02184_
+ sky130_fd_sc_hd__and3b_1
Xfanout88 net91 vssd1 vssd1 vccd1 vccd1 net88 sky130_fd_sc_hd__clkbuf_4
Xfanout99 net101 vssd1 vssd1 vccd1 vccd1 net99 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_107_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10460_ _04599_ _04709_ vssd1 vssd1 vccd1 vccd1 _04710_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_150_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_91_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11747__B1 _05624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09119_ _03761_ genblk2\[0\].wave_shpr.div.acc\[2\] _03766_ vssd1 vssd1 vccd1 vccd1
+ _03767_ sky130_fd_sc_hd__o21a_1
XFILLER_0_122_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10391_ _04058_ _01570_ vssd1 vssd1 vccd1 vccd1 _04664_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_60_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12130_ genblk2\[10\].wave_shpr.div.acc\[13\] _05885_ _05865_ vssd1 vssd1 vccd1 vccd1
+ _05886_ sky130_fd_sc_hd__mux2_1
XANTENNA__07966__A2 _01214_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_102_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11739__A1_N _01099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12061_ _02155_ vssd1 vssd1 vccd1 vccd1 _05835_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold480 genblk2\[4\].wave_shpr.div.quo\[23\] vssd1 vssd1 vccd1 vccd1 net698 sky130_fd_sc_hd__dlygate4sd3_1
Xhold491 genblk2\[8\].wave_shpr.div.quo\[2\] vssd1 vssd1 vccd1 vccd1 net709 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12172__B1 _05816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11012_ _05097_ _04991_ vssd1 vssd1 vccd1 vccd1 _05098_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12963_ clknet_leaf_111_clk _00292_ net130 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.quo\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11278__A2 _05279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_84_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_84_clk sky130_fd_sc_hd__clkbuf_16
X_11914_ genblk2\[10\].wave_shpr.div.acc\[12\] genblk2\[10\].wave_shpr.div.b1\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05736_ sky130_fd_sc_hd__or2b_1
XFILLER_0_59_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12894_ clknet_leaf_32_clk net427 net99 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.quo\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11845_ _05596_ _05559_ vssd1 vssd1 vccd1 vccd1 _05686_ sky130_fd_sc_hd__or2b_1
XTAP_2685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_142_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10238__B1 _04454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11776_ net513 _05628_ _05629_ net530 _05637_ vssd1 vssd1 vccd1 vccd1 _00883_ sky130_fd_sc_hd__a221o_1
XTAP_1995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_144_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13515_ clknet_leaf_78_clk _00832_ net206 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.acc\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10727_ _04896_ _04789_ vssd1 vssd1 vccd1 vccd1 _04897_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09909__A _04250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13446_ clknet_leaf_99_clk _00021_ net166 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.done
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12667__RESET_B net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10658_ genblk2\[5\].wave_shpr.div.quo\[2\] _04853_ _04857_ net879 vssd1 vssd1 vccd1
+ vccd1 _00545_ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_51_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13377_ clknet_leaf_81_clk _00696_ net199 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.b1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10589_ genblk2\[5\].wave_shpr.div.acc\[21\] genblk2\[5\].wave_shpr.div.acc\[20\]
+ genblk2\[5\].wave_shpr.div.acc\[19\] _04816_ vssd1 vssd1 vccd1 vccd1 _04817_ sky130_fd_sc_hd__or4_1
XANTENNA__07429__A _02155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12328_ _03689_ genblk1\[11\].osc.clkdiv_C.cnt\[9\] vssd1 vssd1 vccd1 vccd1 _06022_
+ sky130_fd_sc_hd__and2_1
XANTENNA__09159__A1 genblk2\[0\].wave_shpr.div.quo\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12259_ genblk2\[11\].wave_shpr.div.fin_quo\[7\] net1341 _00005_ vssd1 vssd1 vccd1
+ vccd1 _05990_ sky130_fd_sc_hd__mux2_1
XANTENNA__08959__S _02248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08382__A2 _02336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06820_ _01656_ _01657_ _01664_ _01691_ vssd1 vssd1 vccd1 vccd1 _01692_ sky130_fd_sc_hd__nor4_1
XANTENNA__12070__A _05815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07590__B1 _01923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07164__A genblk1\[9\].osc.clkdiv_C.cnt\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06751_ _01631_ vssd1 vssd1 vccd1 vccd1 _01632_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_75_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_75_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_78_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09470_ _04022_ vssd1 vssd1 vccd1 vccd1 _00192_ sky130_fd_sc_hd__clkbuf_1
X_06682_ genblk1\[4\].osc.clkdiv_C.cnt\[4\] _01439_ _01340_ genblk1\[4\].osc.clkdiv_C.cnt\[8\]
+ _01571_ vssd1 vssd1 vccd1 vccd1 _01572_ sky130_fd_sc_hd__o221a_1
X_08421_ _03079_ _03127_ vssd1 vssd1 vccd1 vccd1 _03128_ sky130_fd_sc_hd__or2b_1
XANTENNA__06696__A2 _01326_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08352_ genblk2\[5\].wave_shpr.div.fin_quo\[5\] _02521_ _02791_ vssd1 vssd1 vccd1
+ vccd1 _03059_ sky130_fd_sc_hd__a21o_1
XANTENNA__09095__A0 _01211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07303_ genblk1\[11\].osc.clkdiv_C.cnt\[13\] _01256_ _01595_ genblk1\[11\].osc.clkdiv_C.cnt\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02067_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_116_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08283_ _02366_ _02976_ _02983_ vssd1 vssd1 vccd1 vccd1 _02990_ sky130_fd_sc_hd__or3_1
XFILLER_0_6_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout135_A net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09819__A _04069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07234_ genblk1\[10\].osc.clkdiv_C.cnt\[15\] _01359_ vssd1 vssd1 vccd1 vccd1 _02016_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_693 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_104_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07165_ _01953_ _01960_ _01961_ vssd1 vssd1 vccd1 vccd1 genblk1\[9\].osc.clkdiv_C.next_cnt\[3\]
+ sky130_fd_sc_hd__nor3_1
XANTENNA__09538__B genblk1\[1\].osc.clkdiv_C.cnt\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06116_ net380 _01087_ vssd1 vssd1 vccd1 vccd1 smpl_rt_clkdiv.clkDiv_inst.next_cnt\[4\]
+ sky130_fd_sc_hd__xor2_1
X_07096_ genblk1\[8\].osc.clkdiv_C.cnt\[10\] genblk1\[8\].osc.clkdiv_C.cnt\[9\] _01900_
+ vssd1 vssd1 vccd1 vccd1 _01904_ sky130_fd_sc_hd__and3_1
XFILLER_0_112_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_292 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout201 net210 vssd1 vssd1 vccd1 vccd1 net201 sky130_fd_sc_hd__clkbuf_4
Xfanout212 net213 vssd1 vssd1 vccd1 vccd1 net212 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10704__A1 _03819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09806_ net275 _04248_ _04252_ net449 vssd1 vssd1 vccd1 vccd1 _00298_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07998_ genblk1\[6\].osc.clkdiv_C.cnt\[14\] _01361_ vssd1 vssd1 vccd1 vccd1 _02705_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__07581__B1 _01171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09737_ genblk2\[2\].wave_shpr.div.fin_quo\[1\] net1348 _00009_ vssd1 vssd1 vccd1
+ vccd1 _04216_ sky130_fd_sc_hd__mux2_1
X_06949_ net1356 _01787_ vssd1 vssd1 vccd1 vccd1 _01788_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_66_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_66_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__08125__A2 _01870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09668_ genblk2\[1\].wave_shpr.div.i\[1\] genblk2\[1\].wave_shpr.div.i\[0\] genblk2\[1\].wave_shpr.div.i\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04151_ sky130_fd_sc_hd__and3_1
XANTENNA__09207__B1_N _03717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08530__C1 net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout48_A net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07802__A _02221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08619_ _03320_ _03325_ vssd1 vssd1 vccd1 vccd1 _03326_ sky130_fd_sc_hd__xor2_1
XTAP_1225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10639__S _04834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09599_ _03987_ _04100_ vssd1 vssd1 vccd1 vccd1 _04101_ sky130_fd_sc_hd__xnor2_1
XTAP_1236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11630_ genblk2\[8\].wave_shpr.div.acc\[18\] genblk2\[8\].wave_shpr.div.acc\[19\]
+ _05529_ vssd1 vssd1 vccd1 vccd1 _05533_ sky130_fd_sc_hd__or3_1
XFILLER_0_65_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06418__A _01361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11561_ _05380_ _05372_ vssd1 vssd1 vccd1 vccd1 _05481_ sky130_fd_sc_hd__or2b_1
XANTENNA__06137__B net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_120 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13300_ clknet_leaf_83_clk _00621_ net199 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.b1\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_92_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10512_ genblk2\[4\].wave_shpr.div.acc\[25\] genblk2\[4\].wave_shpr.div.acc\[24\]
+ genblk2\[4\].wave_shpr.div.acc\[26\] _04621_ vssd1 vssd1 vccd1 vccd1 _04748_ sky130_fd_sc_hd__o31a_1
XFILLER_0_80_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11492_ _05441_ vssd1 vssd1 vccd1 vccd1 _05442_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_107_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13231_ clknet_leaf_11_clk _00554_ net73 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.quo\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_134_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10443_ _04696_ _04591_ vssd1 vssd1 vccd1 vccd1 _04697_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13162_ clknet_leaf_115_clk _00487_ net67 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.acc\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10374_ net732 _04652_ _04656_ net793 vssd1 vssd1 vccd1 vccd1 _00462_ sky130_fd_sc_hd__a22o_1
XANTENNA__10009__A_N genblk2\[3\].wave_shpr.div.b1\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_871 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12113_ net951 _05844_ _05850_ _05872_ vssd1 vssd1 vccd1 vccd1 _00985_ sky130_fd_sc_hd__a22o_1
XANTENNA__11994__A _03707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13093_ clknet_leaf_139_clk _00420_ net39 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.acc\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_12044_ net521 _05823_ _05825_ net583 _05826_ vssd1 vssd1 vccd1 vccd1 _00962_ sky130_fd_sc_hd__a221o_1
XANTENNA__10403__A _04058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06600__B _01432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_57_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_57_clk sky130_fd_sc_hd__clkbuf_16
X_12946_ clknet_leaf_125_clk _00275_ net69 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.b1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12877_ clknet_leaf_119_clk _00208_ net141 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.quo\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11234__A _05249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11828_ _05612_ vssd1 vssd1 vccd1 vccd1 _05673_ sky130_fd_sc_hd__buf_4
XTAP_1770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11759_ net481 _03696_ _03694_ net557 _05627_ vssd1 vssd1 vccd1 vccd1 _00876_ sky130_fd_sc_hd__a221o_1
XFILLER_0_55_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13429_ clknet_leaf_83_clk _00748_ net201 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.acc\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08052__A1 _01489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06602__A2 _01484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08970_ _03656_ _03523_ vssd1 vssd1 vccd1 vccd1 _03657_ sky130_fd_sc_hd__nor2_1
XANTENNA__08412__C_N net25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07921_ genblk1\[8\].osc.clkdiv_C.cnt\[7\] _01430_ vssd1 vssd1 vccd1 vccd1 _02628_
+ sky130_fd_sc_hd__or2_1
XANTENNA__10698__B1 _04856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12004__S _05802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07606__B net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07852_ genblk2\[1\].wave_shpr.div.fin_quo\[3\] _02309_ _02469_ vssd1 vssd1 vccd1
+ vccd1 _02559_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07563__B1 _01801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06803_ _01674_ vssd1 vssd1 vccd1 vccd1 _01675_ sky130_fd_sc_hd__buf_4
XFILLER_0_127_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput1 pb[0] vssd1 vssd1 vccd1 vccd1 net1 sky130_fd_sc_hd__buf_2
X_07783_ _01200_ genblk1\[0\].osc.clkdiv_C.cnt\[6\] genblk1\[0\].osc.clkdiv_C.cnt\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02490_ sky130_fd_sc_hd__a21o_1
Xclkbuf_leaf_48_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_48_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_79_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08107__A2 _01208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09522_ _03853_ genblk1\[1\].osc.clkdiv_C.cnt\[1\] vssd1 vssd1 vccd1 vccd1 _04050_
+ sky130_fd_sc_hd__and2_1
X_06734_ _01600_ _01617_ _01618_ vssd1 vssd1 vccd1 vccd1 _01619_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07315__B1 _02077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09453_ _04014_ vssd1 vssd1 vccd1 vccd1 _00183_ sky130_fd_sc_hd__clkbuf_1
X_06665_ net436 _01554_ vssd1 vssd1 vccd1 vccd1 genblk1\[3\].osc.clkdiv_C.next_cnt\[17\]
+ sky130_fd_sc_hd__xnor2_1
XPHY_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_94_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08404_ _01201_ genblk1\[2\].osc.clkdiv_C.cnt\[16\] _01362_ _03109_ _03110_ vssd1
+ vssd1 vccd1 vccd1 _03111_ sky130_fd_sc_hd__o311a_1
XFILLER_0_19_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09384_ _03944_ _03948_ _03950_ _03947_ net741 vssd1 vssd1 vccd1 vccd1 _00178_ sky130_fd_sc_hd__a32o_1
XFILLER_0_52_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06596_ genblk1\[3\].osc.clkdiv_C.cnt\[17\] _01493_ _01495_ _01503_ vssd1 vssd1 vccd1
+ vccd1 _01504_ sky130_fd_sc_hd__or4b_1
XANTENNA__06238__A _01181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08335_ _02604_ _03034_ _03040_ _02648_ vssd1 vssd1 vccd1 vccd1 _03042_ sky130_fd_sc_hd__a22o_1
XANTENNA__10983__A _05074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08266_ _02349_ _02351_ _02354_ genblk2\[11\].wave_shpr.div.fin_quo\[4\] vssd1 vssd1
+ vccd1 vccd1 _02973_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_6_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07217_ _01995_ _01996_ _01997_ _01342_ _01998_ vssd1 vssd1 vccd1 vccd1 _01999_ sky130_fd_sc_hd__a221o_1
XFILLER_0_61_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09268__B genblk1\[0\].osc.clkdiv_C.cnt\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08197_ genblk2\[11\].wave_shpr.div.fin_quo\[6\] _02361_ vssd1 vssd1 vccd1 vccd1
+ _02904_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07148_ genblk1\[9\].osc.clkdiv_C.cnt\[1\] _01947_ vssd1 vssd1 vccd1 vccd1 _01948_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10922__S _05042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07079_ _01887_ _01892_ _01893_ vssd1 vssd1 vccd1 vccd1 genblk1\[8\].osc.clkdiv_C.next_cnt\[3\]
+ sky130_fd_sc_hd__nor3_1
X_10090_ genblk2\[3\].wave_shpr.div.quo\[3\] _04452_ _04456_ net737 vssd1 vssd1 vccd1
+ vccd1 _00378_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_39_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_39_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_97_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12800_ clknet_leaf_59_clk _00133_ net192 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.quo\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10992_ _05081_ _05082_ net1122 _05052_ vssd1 vssd1 vccd1 vccd1 _00654_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_96_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09846__A2 _04247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12731_ clknet_leaf_38_clk genblk1\[10\].osc.clkdiv_C.next_cnt\[8\] net115 vssd1
+ vssd1 vccd1 vccd1 genblk1\[10\].osc.clkdiv_C.cnt\[8\] sky130_fd_sc_hd__dfrtp_1
XTAP_1000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09059__A0 _01229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12941__RESET_B net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12662_ clknet_leaf_25_clk genblk1\[6\].osc.clkdiv_C.next_cnt\[11\] net87 vssd1 vssd1
+ vccd1 vccd1 genblk1\[6\].osc.clkdiv_C.cnt\[11\] sky130_fd_sc_hd__dfrtp_4
XTAP_1066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11613_ _05403_ _05520_ vssd1 vssd1 vccd1 vccd1 _05521_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12593_ clknet_leaf_13_clk genblk1\[2\].osc.clkdiv_C.next_cnt\[14\] net70 vssd1 vssd1
+ vccd1 vccd1 genblk1\[2\].osc.clkdiv_C.cnt\[14\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_93_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11544_ net445 _05441_ _05458_ net505 _05469_ vssd1 vssd1 vccd1 vccd1 _00819_ sky130_fd_sc_hd__a221o_1
XFILLER_0_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11475_ net1236 net34 _05433_ vssd1 vssd1 vccd1 vccd1 _05435_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_111_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_61_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13214_ clknet_leaf_6_clk _00537_ net48 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.b1\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10426_ genblk2\[4\].wave_shpr.div.b1\[0\] _04583_ _04584_ vssd1 vssd1 vccd1 vccd1
+ _04684_ sky130_fd_sc_hd__and3_1
XFILLER_0_111_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10916__A1 _01797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13145_ clknet_leaf_121_clk net603 net81 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.quo\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10357_ _03708_ _01441_ _01367_ vssd1 vssd1 vccd1 vccd1 _04647_ sky130_fd_sc_hd__and3_4
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07707__A _02316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13076_ clknet_leaf_136_clk _00403_ net62 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.acc\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10288_ genblk2\[4\].wave_shpr.div.b1\[9\] genblk2\[4\].wave_shpr.div.acc\[9\] vssd1
+ vssd1 vccd1 vccd1 _04600_ sky130_fd_sc_hd__and2b_1
X_12027_ net555 _05813_ _05817_ net723 vssd1 vssd1 vccd1 vccd1 _00954_ sky130_fd_sc_hd__a22o_1
XANTENNA__11229__A _05074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10133__A _04477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10144__A2 _04452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11892__A2 _03696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12929_ clknet_leaf_123_clk _00008_ net76 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.busy
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11644__A2 _05448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06450_ genblk1\[1\].osc.clkdiv_C.cnt\[6\] _01385_ vssd1 vssd1 vccd1 vccd1 _01388_
+ sky130_fd_sc_hd__nor2_1
XTAP_2290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_118_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06381_ _01324_ vssd1 vssd1 vccd1 vccd1 _01325_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08120_ _01224_ _01249_ genblk1\[4\].osc.clkdiv_C.cnt\[5\] vssd1 vssd1 vccd1 vccd1
+ _02827_ sky130_fd_sc_hd__o21a_1
XFILLER_0_154_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08051_ genblk1\[5\].osc.clkdiv_C.cnt\[10\] _01667_ vssd1 vssd1 vccd1 vccd1 _02758_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_24_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07002_ genblk1\[7\].osc.clkdiv_C.cnt\[6\] _01830_ vssd1 vssd1 vccd1 vccd1 _01832_
+ sky130_fd_sc_hd__and2_1
XANTENNA__09222__B1 _03840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08953_ _03559_ _03642_ vssd1 vssd1 vccd1 vccd1 _03643_ sky130_fd_sc_hd__xnor2_1
X_07904_ genblk1\[8\].osc.clkdiv_C.cnt\[11\] _01869_ vssd1 vssd1 vccd1 vccd1 _02611_
+ sky130_fd_sc_hd__nor2_1
X_08884_ sig_norm.acc\[9\] _03589_ vssd1 vssd1 vccd1 vccd1 _03590_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07835_ _02510_ _02512_ genblk2\[0\].wave_shpr.div.fin_quo\[4\] vssd1 vssd1 vccd1
+ vccd1 _02542_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10978__A _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07766_ genblk1\[0\].osc.clkdiv_C.cnt\[13\] _01255_ vssd1 vssd1 vccd1 vccd1 _02473_
+ sky130_fd_sc_hd__and2_1
XANTENNA__09043__S _03708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09505_ _04042_ vssd1 vssd1 vccd1 vccd1 _04043_ sky130_fd_sc_hd__buf_4
XFILLER_0_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06717_ genblk1\[4\].osc.clkdiv_C.cnt\[2\] genblk1\[4\].osc.clkdiv_C.cnt\[1\] genblk1\[4\].osc.clkdiv_C.cnt\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01605_ sky130_fd_sc_hd__and3_1
X_07697_ _02403_ vssd1 vssd1 vccd1 vccd1 _02404_ sky130_fd_sc_hd__buf_2
XFILLER_0_63_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08167__B _01231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09436_ genblk2\[1\].wave_shpr.div.b1\[15\] genblk2\[1\].wave_shpr.div.acc\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04000_ sky130_fd_sc_hd__and2b_1
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07071__B genblk1\[8\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06648_ _01486_ _01542_ _01544_ vssd1 vssd1 vccd1 vccd1 genblk1\[3\].osc.clkdiv_C.next_cnt\[11\]
+ sky130_fd_sc_hd__a21oi_1
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09367_ genblk2\[0\].wave_shpr.div.acc\[24\] _03802_ genblk2\[0\].wave_shpr.div.acc\[25\]
+ vssd1 vssd1 vccd1 vccd1 _03937_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_81_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06579_ _01172_ _01182_ vssd1 vssd1 vccd1 vccd1 _01487_ sky130_fd_sc_hd__nand2_4
XANTENNA__12225__A_N genblk2\[11\].wave_shpr.div.b1\[11\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_90_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08318_ _02303_ _02263_ genblk2\[9\].wave_shpr.div.fin_quo\[3\] vssd1 vssd1 vccd1
+ vccd1 _03025_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_151_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09298_ net964 _03870_ _03877_ _03886_ vssd1 vssd1 vccd1 vccd1 _00156_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_758 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10071__A1 _01595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08249_ genblk2\[8\].wave_shpr.div.fin_quo\[6\] _02309_ _02636_ vssd1 vssd1 vccd1
+ vccd1 _02956_ sky130_fd_sc_hd__a21o_1
XANTENNA__06814__A2 _01242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12348__B1 _03947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11260_ _05260_ genblk1\[7\].osc.clkdiv_C.cnt\[15\] vssd1 vssd1 vccd1 vccd1 _05270_
+ sky130_fd_sc_hd__and2_1
XANTENNA__13558__RESET_B net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10211_ genblk2\[3\].wave_shpr.div.acc\[17\] _04536_ _04507_ vssd1 vssd1 vccd1 vccd1
+ _04537_ sky130_fd_sc_hd__mux2_1
XANTENNA__09764__A1 _01794_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11191_ net1280 _01556_ _05042_ vssd1 vssd1 vccd1 vccd1 _05235_ sky130_fd_sc_hd__mux2_1
XFILLER_0_101_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10142_ _04382_ _04483_ vssd1 vssd1 vccd1 vccd1 _04484_ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11049__A _05054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09516__A1 net292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10073_ net1262 _04242_ _04440_ vssd1 vssd1 vccd1 vccd1 _04447_ sky130_fd_sc_hd__mux2_1
X_13763_ clknet_leaf_69_clk _01074_ net214 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.acc\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10975_ genblk2\[6\].wave_shpr.div.quo\[20\] _05062_ _05064_ net313 _05072_ vssd1
+ vssd1 vccd1 vccd1 _00647_ sky130_fd_sc_hd__a221o_1
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12714_ clknet_leaf_54_clk genblk1\[9\].osc.clkdiv_C.next_cnt\[9\] net175 vssd1 vssd1
+ vccd1 vccd1 genblk1\[9\].osc.clkdiv_C.cnt\[9\] sky130_fd_sc_hd__dfrtp_2
X_13694_ clknet_leaf_45_clk _01005_ net122 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.i\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12645_ clknet_leaf_24_clk genblk1\[5\].osc.clkdiv_C.next_cnt\[12\] net92 vssd1 vssd1
+ vccd1 vccd1 genblk1\[5\].osc.clkdiv_C.cnt\[12\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_155_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09189__A _03701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07058__A2 _01211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08255__B2 _02539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12576_ clknet_leaf_29_clk genblk1\[1\].osc.clkdiv_C.next_cnt\[15\] net95 vssd1 vssd1
+ vccd1 vccd1 genblk1\[1\].osc.clkdiv_C.cnt\[15\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__06606__A _01234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10062__A1 _01240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11527_ net502 _05454_ _05458_ net611 _05460_ vssd1 vssd1 vccd1 vccd1 _00811_ sky130_fd_sc_hd__a221o_1
XFILLER_0_135_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12339__B1 _03941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold309 genblk2\[7\].wave_shpr.div.quo\[20\] vssd1 vssd1 vccd1 vccd1 net527 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11458_ genblk2\[9\].wave_shpr.div.b1\[0\] _02064_ _05237_ vssd1 vssd1 vccd1 vccd1
+ _05426_ sky130_fd_sc_hd__mux2_1
XANTENNA__09755__A1 _04225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08558__A2 genblk2\[8\].wave_shpr.div.fin_quo\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10409_ genblk2\[4\].wave_shpr.div.quo\[21\] _04661_ _04663_ net626 _04673_ vssd1
+ vssd1 vccd1 vccd1 _00480_ sky130_fd_sc_hd__a221o_1
XFILLER_0_21_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11389_ genblk2\[8\].wave_shpr.div.acc\[10\] genblk2\[8\].wave_shpr.div.b1\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05365_ sky130_fd_sc_hd__or2b_1
XFILLER_0_0_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13128_ clknet_leaf_3_clk _00453_ net46 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.b1\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13059_ clknet_leaf_24_clk _00386_ net92 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.quo\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07156__B genblk1\[9\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1009 genblk2\[4\].wave_shpr.div.b1\[17\] vssd1 vssd1 vccd1 vccd1 net1227 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_17_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07620_ genblk1\[11\].osc.clkdiv_C.cnt\[6\] _01430_ _01595_ genblk1\[11\].osc.clkdiv_C.cnt\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02327_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07551_ net1142 net1128 PWM.start vssd1 vssd1 vccd1 vccd1 _02259_ sky130_fd_sc_hd__mux2_1
XFILLER_0_49_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06502_ genblk1\[2\].osc.clkdiv_C.cnt\[11\] _01420_ _01421_ _01422_ _01427_ vssd1
+ vssd1 vccd1 vccd1 _01428_ sky130_fd_sc_hd__o221a_1
XFILLER_0_124_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07482_ _02147_ _02207_ vssd1 vssd1 vccd1 vccd1 _02208_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09221_ net558 _03836_ _03840_ net655 vssd1 vssd1 vccd1 vccd1 _00125_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06433_ genblk1\[1\].osc.clkdiv_C.cnt\[1\] genblk1\[1\].osc.clkdiv_C.cnt\[0\] vssd1
+ vssd1 vccd1 vccd1 _01376_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09152_ genblk2\[0\].wave_shpr.div.acc\[19\] _03799_ vssd1 vssd1 vccd1 vccd1 _03800_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_146_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06364_ _01178_ vssd1 vssd1 vccd1 vccd1 _01308_ sky130_fd_sc_hd__inv_4
XANTENNA__06254__A2_N _01215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06516__A _01200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08103_ genblk1\[4\].osc.clkdiv_C.cnt\[11\] _01574_ vssd1 vssd1 vccd1 vccd1 _02810_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_32_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06295_ _01188_ _01187_ _01173_ vssd1 vssd1 vccd1 vccd1 _01257_ sky130_fd_sc_hd__o21ba_1
X_09083_ _02170_ _01201_ _01363_ vssd1 vssd1 vccd1 vccd1 _03735_ sky130_fd_sc_hd__or3_4
XANTENNA_fanout215_A net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08034_ _02739_ _02740_ vssd1 vssd1 vccd1 vccd1 _02741_ sky130_fd_sc_hd__and2b_1
XFILLER_0_141_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09827__A _04058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold810 _00043_ vssd1 vssd1 vccd1 vccd1 net1028 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold821 genblk2\[9\].wave_shpr.div.i\[1\] vssd1 vssd1 vccd1 vccd1 net1039 sky130_fd_sc_hd__dlygate4sd3_1
Xhold832 genblk2\[0\].wave_shpr.div.acc\[16\] vssd1 vssd1 vccd1 vccd1 net1050 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11568__S _05417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold843 genblk2\[5\].wave_shpr.div.acc\[11\] vssd1 vssd1 vccd1 vccd1 net1061 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09546__B genblk1\[1\].osc.clkdiv_C.cnt\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold854 genblk1\[5\].osc.clkdiv_C.cnt\[7\] vssd1 vssd1 vccd1 vccd1 net1072 sky130_fd_sc_hd__dlygate4sd3_1
Xhold865 sig_norm.quo\[0\] vssd1 vssd1 vccd1 vccd1 net1083 sky130_fd_sc_hd__dlygate4sd3_1
Xhold876 genblk2\[2\].wave_shpr.div.acc\[25\] vssd1 vssd1 vccd1 vccd1 net1094 sky130_fd_sc_hd__dlygate4sd3_1
Xhold887 genblk1\[5\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 net1105 sky130_fd_sc_hd__dlygate4sd3_1
Xhold898 genblk2\[8\].wave_shpr.div.acc\[1\] vssd1 vssd1 vccd1 vccd1 net1116 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_51_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09985_ genblk2\[3\].wave_shpr.div.b1\[1\] genblk2\[3\].wave_shpr.div.acc\[1\] vssd1
+ vssd1 vccd1 vccd1 _04381_ sky130_fd_sc_hd__xor2_1
XANTENNA__06251__A _01174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08936_ _03529_ _03547_ _03549_ vssd1 vssd1 vccd1 vccd1 _03629_ sky130_fd_sc_hd__a21o_1
X_08867_ net1131 _02260_ _03573_ vssd1 vssd1 vccd1 vccd1 _00038_ sky130_fd_sc_hd__a21o_1
XANTENNA__08182__B1 _02224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_66_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07818_ _02524_ vssd1 vssd1 vccd1 vccd1 _02525_ sky130_fd_sc_hd__clkbuf_4
X_08798_ _03425_ _03426_ _03423_ _03424_ vssd1 vssd1 vccd1 vccd1 _03505_ sky130_fd_sc_hd__o211ai_2
XFILLER_0_79_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07082__A genblk1\[8\].osc.clkdiv_C.cnt\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07749_ _02426_ _02454_ _02428_ _02451_ _02455_ vssd1 vssd1 vccd1 vccd1 _02456_ sky130_fd_sc_hd__a221o_1
X_10760_ _04856_ vssd1 vssd1 vccd1 vccd1 _04922_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_149_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07810__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09419_ _03965_ genblk2\[1\].wave_shpr.div.acc\[6\] _03982_ vssd1 vssd1 vccd1 vccd1
+ _03983_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10691_ _04869_ genblk1\[5\].osc.clkdiv_C.cnt\[11\] vssd1 vssd1 vccd1 vccd1 _04873_
+ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_124_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12430_ net931 _06072_ _06073_ _06094_ vssd1 vssd1 vccd1 vccd1 _01080_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12361_ genblk2\[11\].wave_shpr.div.acc\[3\] _06042_ _05982_ vssd1 vssd1 vccd1 vccd1
+ _06043_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11792__A1 _03819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11312_ _05203_ _05170_ vssd1 vssd1 vccd1 vccd1 _05308_ sky130_fd_sc_hd__or2b_1
XFILLER_0_132_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12292_ net1270 _01327_ _05994_ vssd1 vssd1 vccd1 vccd1 _06008_ sky130_fd_sc_hd__mux2_1
XFILLER_0_120_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_139_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11243_ net550 _05255_ _05256_ net613 _05261_ vssd1 vssd1 vccd1 vccd1 _00726_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_19_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11174_ _05228_ vssd1 vssd1 vccd1 vccd1 _00690_ sky130_fd_sc_hd__clkbuf_1
X_10125_ genblk2\[3\].wave_shpr.div.quo\[21\] _04461_ _04462_ net545 _04473_ vssd1
+ vssd1 vccd1 vccd1 _00396_ sky130_fd_sc_hd__a221o_1
XANTENNA__09472__A _03701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10056_ _04437_ vssd1 vssd1 vccd1 vccd1 _00363_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11507__A _05441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07920__B1 genblk1\[8\].osc.clkdiv_C.cnt\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10807__A0 _04856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13746_ clknet_leaf_51_clk net435 net110 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.quo\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10958_ genblk2\[6\].wave_shpr.div.quo\[12\] _05062_ _05055_ net623 _05063_ vssd1
+ vssd1 vccd1 vccd1 _00639_ sky130_fd_sc_hd__a221o_1
XFILLER_0_85_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13677_ clknet_leaf_42_clk _00990_ net125 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.acc\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10889_ _05028_ vssd1 vssd1 vccd1 vccd1 _00605_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12338__A _03833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12628_ clknet_leaf_18_clk genblk1\[4\].osc.clkdiv_C.next_cnt\[13\] net81 vssd1 vssd1
+ vccd1 vccd1 genblk1\[4\].osc.clkdiv_C.cnt\[13\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__08228__B2 _02362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12024__A2 _05813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11232__B1 _05248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12559_ clknet_leaf_56_clk genblk1\[0\].osc.clkdiv_C.next_cnt\[16\] net181 vssd1
+ vssd1 vccd1 vccd1 genblk1\[0\].osc.clkdiv_C.cnt\[16\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_102_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold106 genblk2\[5\].wave_shpr.div.quo\[24\] vssd1 vssd1 vccd1 vccd1 net324 sky130_fd_sc_hd__dlygate4sd3_1
Xhold117 _00971_ vssd1 vssd1 vccd1 vccd1 net335 sky130_fd_sc_hd__dlygate4sd3_1
Xhold128 genblk2\[8\].wave_shpr.div.quo\[3\] vssd1 vssd1 vccd1 vccd1 net346 sky130_fd_sc_hd__dlygate4sd3_1
Xhold139 genblk2\[10\].wave_shpr.div.quo\[15\] vssd1 vssd1 vccd1 vccd1 net357 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07167__A genblk1\[9\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09770_ genblk2\[3\].wave_shpr.div.b1\[7\] _02077_ _04039_ vssd1 vssd1 vccd1 vccd1
+ _04235_ sky130_fd_sc_hd__mux2_1
X_06982_ _01800_ _01804_ _01807_ _01817_ vssd1 vssd1 vccd1 vccd1 _01818_ sky130_fd_sc_hd__and4_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08721_ _03408_ vssd1 vssd1 vccd1 vccd1 _03428_ sky130_fd_sc_hd__inv_2
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07506__A3 _02224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08652_ _03334_ _03335_ _03357_ _03358_ vssd1 vssd1 vccd1 vccd1 _03359_ sky130_fd_sc_hd__a211oi_4
X_07603_ _02221_ net32 vssd1 vssd1 vccd1 vccd1 _02310_ sky130_fd_sc_hd__nor2_2
XFILLER_0_135_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08583_ genblk2\[10\].wave_shpr.div.fin_quo\[2\] _02308_ _02416_ vssd1 vssd1 vccd1
+ vccd1 _03290_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout165_A net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07534_ _01151_ _02245_ _02250_ vssd1 vssd1 vccd1 vccd1 _00028_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_76_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_37_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07465_ genblk2\[8\].wave_shpr.div.i\[2\] genblk2\[8\].wave_shpr.div.i\[3\] genblk2\[8\].wave_shpr.div.i\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02195_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_9_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09204_ _03830_ vssd1 vssd1 vccd1 vccd1 _00118_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_147_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06416_ _01359_ vssd1 vssd1 vccd1 vccd1 _01360_ sky130_fd_sc_hd__buf_4
XFILLER_0_91_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07396_ genblk1\[11\].osc.clkdiv_C.cnt\[16\] _02143_ vssd1 vssd1 vccd1 vccd1 _02144_
+ sky130_fd_sc_hd__or2_1
XANTENNA__07690__A2 _01991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08164__C _01182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09135_ genblk2\[0\].wave_shpr.div.b1\[10\] genblk2\[0\].wave_shpr.div.acc\[10\]
+ vssd1 vssd1 vccd1 vccd1 _03783_ sky130_fd_sc_hd__and2b_1
XANTENNA__11223__B1 _05250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06347_ genblk1\[0\].osc.clkdiv_C.cnt\[14\] genblk1\[0\].osc.clkdiv_C.cnt\[13\] _01291_
+ vssd1 vssd1 vccd1 vccd1 _01295_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09557__A _04069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09066_ _03724_ vssd1 vssd1 vccd1 vccd1 _00086_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_460 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06278_ _01238_ _01239_ vssd1 vssd1 vccd1 vccd1 _01240_ sky130_fd_sc_hd__nor2_8
X_08017_ _02720_ _02722_ _02723_ vssd1 vssd1 vccd1 vccd1 _02724_ sky130_fd_sc_hd__o21ai_1
Xhold640 genblk2\[10\].wave_shpr.div.acc\[13\] vssd1 vssd1 vccd1 vccd1 net858 sky130_fd_sc_hd__dlygate4sd3_1
Xhold651 _00979_ vssd1 vssd1 vccd1 vccd1 net869 sky130_fd_sc_hd__dlygate4sd3_1
Xhold662 _00545_ vssd1 vssd1 vccd1 vccd1 net880 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07077__A genblk1\[8\].osc.clkdiv_C.cnt\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold673 genblk2\[4\].wave_shpr.div.acc\[8\] vssd1 vssd1 vccd1 vccd1 net891 sky130_fd_sc_hd__dlygate4sd3_1
Xhold684 genblk2\[5\].wave_shpr.div.acc\[14\] vssd1 vssd1 vccd1 vccd1 net902 sky130_fd_sc_hd__dlygate4sd3_1
Xhold695 genblk2\[0\].wave_shpr.div.acc\[14\] vssd1 vssd1 vccd1 vccd1 net913 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06402__B1 _01197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09968_ genblk2\[3\].wave_shpr.div.acc\[14\] genblk2\[3\].wave_shpr.div.b1\[14\]
+ vssd1 vssd1 vccd1 vccd1 _04364_ sky130_fd_sc_hd__or2b_1
X_08919_ sig_norm.acc\[6\] _03614_ net612 vssd1 vssd1 vccd1 vccd1 _03618_ sky130_fd_sc_hd__o21ai_1
X_09899_ net857 _04282_ _04289_ _04314_ vssd1 vssd1 vccd1 vccd1 _00329_ sky130_fd_sc_hd__a22o_1
XANTENNA__08155__B1 _01494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11930_ genblk2\[10\].wave_shpr.div.b1\[3\] genblk2\[10\].wave_shpr.div.acc\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05752_ sky130_fd_sc_hd__and2b_1
XTAP_2801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11861_ _05604_ _05555_ vssd1 vssd1 vccd1 vccd1 _05698_ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13600_ clknet_leaf_76_clk _00915_ net208 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.acc\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10812_ genblk2\[5\].wave_shpr.div.i\[1\] genblk2\[5\].wave_shpr.div.i\[0\] genblk2\[5\].wave_shpr.div.i\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04959_ sky130_fd_sc_hd__a21o_1
XANTENNA__09655__B1 _04048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11792_ _03819_ genblk1\[9\].osc.clkdiv_C.cnt\[17\] _00022_ net1209 _05645_ vssd1
+ vssd1 vccd1 vccd1 _00891_ sky130_fd_sc_hd__o221a_1
XANTENNA__08636__A _02216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13531_ clknet_leaf_84_clk _00022_ net202 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.busy
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_149_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10743_ _04798_ _04771_ vssd1 vssd1 vccd1 vccd1 _04909_ sky130_fd_sc_hd__or2b_1
XFILLER_0_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_116 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13462_ clknet_leaf_83_clk _00779_ net203 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.b1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10674_ _04672_ genblk1\[5\].osc.clkdiv_C.cnt\[3\] vssd1 vssd1 vccd1 vccd1 _04864_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_137_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_152_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12413_ net1125 _06072_ _06073_ _06082_ vssd1 vssd1 vccd1 vccd1 _01075_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13393_ clknet_leaf_118_clk _00712_ net139 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.quo\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12344_ genblk2\[11\].wave_shpr.div.acc_next\[0\] _03941_ vssd1 vssd1 vccd1 vccd1
+ _06030_ sky130_fd_sc_hd__or2b_1
XFILLER_0_51_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12275_ genblk2\[1\].wave_shpr.div.b1\[6\] _01311_ _05994_ vssd1 vssd1 vccd1 vccd1
+ _05999_ sky130_fd_sc_hd__mux2_1
XANTENNA__08090__B _02364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11226_ _05245_ vssd1 vssd1 vccd1 vccd1 _05251_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11157_ genblk2\[7\].wave_shpr.div.acc\[18\] _05216_ vssd1 vssd1 vccd1 vccd1 _05217_
+ sky130_fd_sc_hd__or2_1
X_10108_ genblk2\[3\].wave_shpr.div.quo\[13\] _04461_ _04462_ net387 _04464_ vssd1
+ vssd1 vccd1 vccd1 _00388_ sky130_fd_sc_hd__a221o_1
XFILLER_0_65_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11088_ _05152_ _05153_ vssd1 vssd1 vccd1 vccd1 _05154_ sky130_fd_sc_hd__nand2_1
XANTENNA__11237__A _05074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10039_ genblk2\[3\].wave_shpr.div.fin_quo\[6\] net1346 _04422_ vssd1 vssd1 vccd1
+ vccd1 _04429_ sky130_fd_sc_hd__mux2_1
XANTENNA__08449__A1 genblk2\[8\].wave_shpr.div.fin_quo\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_14_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07450__A _02184_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13729_ clknet_leaf_74_clk _01040_ net212 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11185__A2_N _01432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07121__A1 genblk1\[9\].osc.clkdiv_C.cnt\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07121__B2 genblk1\[9\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07250_ _02028_ _02029_ _02030_ vssd1 vssd1 vccd1 vccd1 _02031_ sky130_fd_sc_hd__and3_1
XFILLER_0_144_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06201_ _01164_ net811 vssd1 vssd1 vccd1 vccd1 PWM.next_counter\[5\] sky130_fd_sc_hd__nor2_1
XFILLER_0_155_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07181_ genblk1\[9\].osc.clkdiv_C.cnt\[7\] _01967_ genblk1\[9\].osc.clkdiv_C.cnt\[8\]
+ vssd1 vssd1 vccd1 vccd1 _01973_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_53_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06132_ net8 net9 vssd1 vssd1 vccd1 vccd1 _01104_ sky130_fd_sc_hd__nand2_1
XFILLER_0_111_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_111_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_485 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08385__B1 _01418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12181__A1 _05816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09822_ genblk2\[2\].wave_shpr.div.quo\[14\] _04257_ _04259_ net457 _04261_ vssd1
+ vssd1 vccd1 vccd1 _00305_ sky130_fd_sc_hd__a221o_1
X_09753_ _04224_ vssd1 vssd1 vccd1 vccd1 _00273_ sky130_fd_sc_hd__clkbuf_1
X_06965_ _01213_ _01344_ vssd1 vssd1 vccd1 vccd1 _01801_ sky130_fd_sc_hd__nand2_2
X_08704_ _03362_ _03377_ vssd1 vssd1 vccd1 vccd1 _03411_ sky130_fd_sc_hd__and2b_1
X_09684_ genblk2\[2\].wave_shpr.div.acc\[9\] genblk2\[2\].wave_shpr.div.b1\[9\] vssd1
+ vssd1 vccd1 vccd1 _04164_ sky130_fd_sc_hd__or2b_1
XFILLER_0_146_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06896_ _01342_ _01439_ vssd1 vssd1 vccd1 vccd1 _01750_ sky130_fd_sc_hd__nand2_2
XTAP_2108 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08635_ genblk2\[8\].wave_shpr.div.fin_quo\[2\] _03341_ vssd1 vssd1 vccd1 vccd1 _03342_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2119 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08566_ _02946_ _03268_ _03272_ vssd1 vssd1 vccd1 vccd1 _03273_ sky130_fd_sc_hd__or3_1
XTAP_1429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10247__A1 _04454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11444__A0 genblk2\[8\].wave_shpr.div.fin_quo\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07517_ _02234_ PWM.final_sample_in\[2\] PWM.final_sample_in\[1\] _02235_ _02236_
+ vssd1 vssd1 vccd1 vccd1 _02237_ sky130_fd_sc_hd__o221a_1
XFILLER_0_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08497_ _03175_ _03202_ _03077_ _03203_ vssd1 vssd1 vccd1 vccd1 _03204_ sky130_fd_sc_hd__o211a_1
XFILLER_0_147_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout45 net47 vssd1 vssd1 vccd1 vccd1 net45 sky130_fd_sc_hd__clkbuf_4
Xfanout56 net58 vssd1 vssd1 vccd1 vccd1 net56 sky130_fd_sc_hd__clkbuf_4
XANTENNA__11995__A1 _02805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout67 net68 vssd1 vssd1 vccd1 vccd1 net67 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_107_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07448_ _02183_ vssd1 vssd1 vccd1 vccd1 _00014_ sky130_fd_sc_hd__inv_2
Xfanout78 net79 vssd1 vssd1 vccd1 vccd1 net78 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07663__A2 _01224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout89 net90 vssd1 vssd1 vccd1 vccd1 net89 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07379_ genblk1\[11\].osc.clkdiv_C.cnt\[12\] _02130_ vssd1 vssd1 vccd1 vccd1 _02131_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_72_480 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09118_ _03764_ _03765_ _03762_ vssd1 vssd1 vccd1 vccd1 _03766_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_44_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10390_ _04654_ vssd1 vssd1 vccd1 vccd1 _04663_ sky130_fd_sc_hd__buf_2
XFILLER_0_115_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09049_ _03713_ vssd1 vssd1 vccd1 vccd1 _00080_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12060_ net334 _05823_ _05825_ net383 _05834_ vssd1 vssd1 vccd1 vccd1 _00970_ sky130_fd_sc_hd__a221o_1
Xhold470 genblk2\[0\].wave_shpr.div.acc\[19\] vssd1 vssd1 vccd1 vccd1 net688 sky130_fd_sc_hd__dlygate4sd3_1
Xhold481 genblk2\[8\].wave_shpr.div.acc\[2\] vssd1 vssd1 vccd1 vccd1 net699 sky130_fd_sc_hd__dlygate4sd3_1
Xhold492 genblk2\[3\].wave_shpr.div.acc\[22\] vssd1 vssd1 vccd1 vccd1 net710 sky130_fd_sc_hd__dlygate4sd3_1
X_11011_ _04992_ _04978_ vssd1 vssd1 vccd1 vccd1 _05097_ sky130_fd_sc_hd__or2b_1
X_12962_ clknet_leaf_130_clk _00291_ net65 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.quo\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_11913_ genblk2\[10\].wave_shpr.div.acc\[13\] genblk2\[10\].wave_shpr.div.b1\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05735_ sky130_fd_sc_hd__or2b_1
XTAP_2620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12893_ clknet_leaf_28_clk _00224_ net91 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.quo\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11844_ _03693_ vssd1 vssd1 vccd1 vccd1 _05685_ sky130_fd_sc_hd__clkbuf_4
XTAP_2664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11775_ _04676_ _01930_ vssd1 vssd1 vccd1 vccd1 _05637_ sky130_fd_sc_hd__nor2_1
XTAP_1974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_82_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11986__A1 _01811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10726_ _04790_ _04775_ vssd1 vssd1 vccd1 vccd1 _04896_ sky130_fd_sc_hd__or2b_1
XFILLER_0_55_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13514_ clknet_leaf_78_clk _00831_ net207 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.acc\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_71_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_302 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13445_ clknet_leaf_81_clk _00020_ net199 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.busy
+ sky130_fd_sc_hd__dfrtp_1
X_10657_ net879 _04853_ _04857_ net1056 vssd1 vssd1 vccd1 vccd1 _00544_ sky130_fd_sc_hd__a22o_1
XFILLER_0_152_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13376_ clknet_leaf_96_clk _00695_ net167 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.b1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10588_ genblk2\[5\].wave_shpr.div.acc\[18\] _04815_ vssd1 vssd1 vccd1 vccd1 _04816_
+ sky130_fd_sc_hd__or2_1
XANTENNA__09800__B1 _04252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06614__B1 _01484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12327_ net510 _06014_ _06015_ net571 _06021_ vssd1 vssd1 vccd1 vccd1 _01050_ sky130_fd_sc_hd__a221o_1
XFILLER_0_133_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12258_ _05989_ vssd1 vssd1 vccd1 vccd1 _01013_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12636__RESET_B net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11209_ _02171_ net1191 vssd1 vssd1 vccd1 vccd1 _05244_ sky130_fd_sc_hd__and2_1
X_12189_ genblk2\[11\].wave_shpr.div.acc\[15\] genblk2\[11\].wave_shpr.div.b1\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05927_ sky130_fd_sc_hd__or2b_1
XANTENNA__12351__A _05982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06750_ genblk1\[4\].osc.clkdiv_C.cnt\[9\] _01627_ vssd1 vssd1 vccd1 vccd1 _01631_
+ sky130_fd_sc_hd__and2_1
X_06681_ genblk1\[4\].osc.clkdiv_C.cnt\[15\] _01362_ _01248_ _01570_ vssd1 vssd1 vccd1
+ vccd1 _01571_ sky130_fd_sc_hd__o22a_1
XFILLER_0_116_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08420_ _03079_ _03125_ _03126_ vssd1 vssd1 vccd1 vccd1 _03127_ sky130_fd_sc_hd__or3_1
XFILLER_0_59_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08351_ genblk2\[5\].wave_shpr.div.fin_quo\[4\] _03056_ _03057_ vssd1 vssd1 vccd1
+ vccd1 _03058_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09095__A1 _01556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_803 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07302_ genblk1\[11\].osc.clkdiv_C.cnt\[13\] _01256_ _02064_ genblk1\[11\].osc.clkdiv_C.cnt\[5\]
+ _02065_ vssd1 vssd1 vccd1 vccd1 _02066_ sky130_fd_sc_hd__a221o_1
XFILLER_0_132_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08282_ _02987_ _02988_ _02314_ vssd1 vssd1 vccd1 vccd1 _02989_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_41_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_116_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07233_ genblk1\[10\].osc.clkdiv_C.cnt\[16\] _01363_ genblk1\[10\].osc.clkdiv_C.cnt\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02015_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_6_555 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_131_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07164_ genblk1\[9\].osc.clkdiv_C.cnt\[3\] _01958_ vssd1 vssd1 vccd1 vccd1 _01961_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06115_ _01087_ _01091_ vssd1 vssd1 vccd1 vccd1 smpl_rt_clkdiv.clkDiv_inst.next_cnt\[3\]
+ sky130_fd_sc_hd__nor2_1
X_07095_ _01887_ _01902_ _01903_ vssd1 vssd1 vccd1 vccd1 genblk1\[8\].osc.clkdiv_C.next_cnt\[9\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_140_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09835__A _02147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout202 net204 vssd1 vssd1 vccd1 vccd1 net202 sky130_fd_sc_hd__clkbuf_4
Xfanout213 net217 vssd1 vssd1 vccd1 vccd1 net213 sky130_fd_sc_hd__clkbuf_4
X_09805_ net449 _04248_ _04252_ net716 vssd1 vssd1 vccd1 vccd1 _00297_ sky130_fd_sc_hd__a22o_1
X_07997_ genblk1\[6\].osc.clkdiv_C.cnt\[14\] _01360_ vssd1 vssd1 vccd1 vccd1 _02704_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_66_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09736_ _04215_ vssd1 vssd1 vccd1 vccd1 _00265_ sky130_fd_sc_hd__clkbuf_1
X_06948_ genblk1\[6\].osc.clkdiv_C.cnt\[15\] genblk1\[6\].osc.clkdiv_C.cnt\[14\] _01783_
+ vssd1 vssd1 vccd1 vccd1 _01787_ sky130_fd_sc_hd__and3_1
XFILLER_0_97_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09667_ genblk2\[1\].wave_shpr.div.i\[1\] genblk2\[1\].wave_shpr.div.i\[0\] genblk2\[1\].wave_shpr.div.i\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04150_ sky130_fd_sc_hd__a21o_1
X_06879_ genblk1\[6\].osc.clkdiv_C.cnt\[4\] _01730_ _01732_ genblk1\[6\].osc.clkdiv_C.cnt\[9\]
+ vssd1 vssd1 vccd1 vccd1 _01733_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__08530__B1 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08618_ _03323_ _03324_ _02846_ vssd1 vssd1 vccd1 vccd1 _03325_ sky130_fd_sc_hd__o21ai_2
XTAP_1204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07802__B net31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09598_ _03988_ _03962_ vssd1 vssd1 vccd1 vccd1 _04100_ sky130_fd_sc_hd__or2b_1
XANTENNA__08186__A net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13165__RESET_B net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08549_ _03253_ _03255_ vssd1 vssd1 vccd1 vccd1 _03256_ sky130_fd_sc_hd__xnor2_1
XTAP_1259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11968__A1 genblk2\[10\].wave_shpr.div.quo\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11560_ net872 _05447_ _05446_ _05480_ vssd1 vssd1 vccd1 vccd1 _00824_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10511_ net787 _04657_ _04722_ _04747_ vssd1 vssd1 vccd1 vccd1 _00508_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11491_ _02198_ vssd1 vssd1 vccd1 vccd1 _05441_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13230_ clknet_leaf_11_clk net311 net73 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.quo\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10442_ _04592_ _04577_ vssd1 vssd1 vccd1 vccd1 _04696_ sky130_fd_sc_hd__or2b_1
XFILLER_0_32_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13161_ clknet_leaf_122_clk _00486_ net79 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.acc\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10373_ genblk2\[4\].wave_shpr.div.quo\[2\] _04652_ _04656_ net464 vssd1 vssd1 vccd1
+ vccd1 _00461_ sky130_fd_sc_hd__a22o_1
XANTENNA__08061__A2 net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12112_ genblk2\[10\].wave_shpr.div.acc\[9\] _05871_ _05865_ vssd1 vssd1 vccd1 vccd1
+ _05872_ sky130_fd_sc_hd__mux2_1
XANTENNA__10943__A2 _05052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_883 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13092_ clknet_leaf_137_clk _00419_ net39 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.acc\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_12043_ _04676_ _01993_ vssd1 vssd1 vccd1 vccd1 _05826_ sky130_fd_sc_hd__nor2_1
XFILLER_0_88_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11656__B1 _05448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12945_ clknet_leaf_13_clk _00274_ net69 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.b1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07324__B2 _01197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08096__A _01174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12876_ clknet_leaf_49_clk _00207_ net113 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.quo\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_2461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10224__A2_N _04480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11827_ _05587_ _05671_ vssd1 vssd1 vccd1 vccd1 _05672_ sky130_fd_sc_hd__xnor2_1
XTAP_1760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11758_ _05464_ genblk1\[9\].osc.clkdiv_C.cnt\[2\] vssd1 vssd1 vccd1 vccd1 _05627_
+ sky130_fd_sc_hd__and2_1
XANTENNA__07627__A2 _01209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10709_ genblk2\[5\].wave_shpr.div.b1\[0\] _04781_ _04782_ vssd1 vssd1 vccd1 vccd1
+ _04883_ sky130_fd_sc_hd__and3_1
X_11689_ _05569_ _05580_ _05567_ vssd1 vssd1 vccd1 vccd1 _05581_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_126_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13428_ clknet_leaf_82_clk net798 net201 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.acc\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13359_ clknet_leaf_91_clk _00018_ net143 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.busy
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07920_ genblk1\[8\].osc.clkdiv_C.cnt\[7\] _01430_ genblk1\[8\].osc.clkdiv_C.cnt\[6\]
+ _01441_ vssd1 vssd1 vccd1 vccd1 _02627_ sky130_fd_sc_hd__a211o_1
X_07851_ _02556_ _02557_ vssd1 vssd1 vccd1 vccd1 _02558_ sky130_fd_sc_hd__or2_1
XANTENNA__11895__A0 _03838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06802_ _01238_ net36 vssd1 vssd1 vccd1 vccd1 _01674_ sky130_fd_sc_hd__nor2_1
X_07782_ genblk1\[0\].osc.clkdiv_C.cnt\[4\] _01241_ _02483_ vssd1 vssd1 vccd1 vccd1
+ _02489_ sky130_fd_sc_hd__o21a_1
Xinput2 pb[10] vssd1 vssd1 vccd1 vccd1 net2 sky130_fd_sc_hd__clkbuf_4
XANTENNA__12439__A2 _03947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09521_ net517 _04048_ _04045_ net460 _04049_ vssd1 vssd1 vccd1 vccd1 _00216_ sky130_fd_sc_hd__a221o_1
X_06733_ genblk1\[4\].osc.clkdiv_C.cnt\[4\] genblk1\[4\].osc.clkdiv_C.cnt\[3\] _01605_
+ genblk1\[4\].osc.clkdiv_C.cnt\[5\] vssd1 vssd1 vccd1 vccd1 _01618_ sky130_fd_sc_hd__a31o_1
XANTENNA__07903__A genblk1\[8\].osc.clkdiv_C.cnt\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09452_ genblk2\[1\].wave_shpr.div.fin_quo\[2\] net1312 _00007_ vssd1 vssd1 vccd1
+ vccd1 _04014_ sky130_fd_sc_hd__mux2_1
X_06664_ _01555_ vssd1 vssd1 vccd1 vccd1 genblk1\[3\].osc.clkdiv_C.next_cnt\[16\]
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07622__B _01211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08403_ _03103_ _03105_ _03106_ _03107_ vssd1 vssd1 vccd1 vccd1 _03110_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_143_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_137_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09383_ _03949_ vssd1 vssd1 vccd1 vccd1 _03950_ sky130_fd_sc_hd__inv_2
XFILLER_0_87_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06595_ genblk1\[3\].osc.clkdiv_C.cnt\[15\] _01363_ _01499_ _01501_ _01502_ vssd1
+ vssd1 vccd1 vccd1 _01503_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_74_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08334_ _02604_ _02648_ _03034_ _03040_ vssd1 vssd1 vccd1 vccd1 _03041_ sky130_fd_sc_hd__nand4_2
XFILLER_0_129_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08265_ _02971_ _02914_ vssd1 vssd1 vccd1 vccd1 _02972_ sky130_fd_sc_hd__xor2_1
XFILLER_0_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07216_ genblk1\[10\].osc.clkdiv_C.cnt\[13\] _01442_ vssd1 vssd1 vccd1 vccd1 _01998_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08196_ genblk2\[11\].wave_shpr.div.fin_quo\[5\] net33 _02350_ _02355_ _02222_ vssd1
+ vssd1 vccd1 vccd1 _02903_ sky130_fd_sc_hd__a41o_1
XFILLER_0_14_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07147_ _01241_ _01946_ vssd1 vssd1 vccd1 vccd1 _01947_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10386__B1 _04655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07078_ genblk1\[8\].osc.clkdiv_C.cnt\[3\] _01890_ vssd1 vssd1 vccd1 vccd1 _01893_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_100_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07085__A genblk1\[8\].osc.clkdiv_C.cnt\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout60_A net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_303 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09719_ genblk2\[2\].wave_shpr.div.b1\[13\] genblk2\[2\].wave_shpr.div.acc\[13\]
+ vssd1 vssd1 vccd1 vccd1 _04199_ sky130_fd_sc_hd__and2b_1
X_10991_ genblk2\[6\].wave_shpr.div.b1\[0\] genblk2\[6\].wave_shpr.div.acc\[0\] _05023_
+ _05079_ vssd1 vssd1 vccd1 vccd1 _05082_ sky130_fd_sc_hd__a31o_1
XANTENNA__07306__A1 _01223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12730_ clknet_leaf_39_clk genblk1\[10\].osc.clkdiv_C.next_cnt\[7\] net115 vssd1
+ vssd1 vccd1 vccd1 genblk1\[10\].osc.clkdiv_C.cnt\[7\] sky130_fd_sc_hd__dfrtp_4
XTAP_1001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12661_ clknet_leaf_26_clk genblk1\[6\].osc.clkdiv_C.next_cnt\[10\] net88 vssd1 vssd1
+ vccd1 vccd1 genblk1\[6\].osc.clkdiv_C.cnt\[10\] sky130_fd_sc_hd__dfrtp_4
XTAP_1056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11612_ _05404_ _05360_ vssd1 vssd1 vccd1 vccd1 _05520_ sky130_fd_sc_hd__or2b_1
XFILLER_0_26_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12592_ clknet_leaf_13_clk genblk1\[2\].osc.clkdiv_C.next_cnt\[13\] net70 vssd1 vssd1
+ vccd1 vccd1 genblk1\[2\].osc.clkdiv_C.cnt\[13\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_108_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11543_ _05464_ genblk1\[8\].osc.clkdiv_C.cnt\[15\] vssd1 vssd1 vccd1 vccd1 _05469_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_107_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12981__RESET_B net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_123_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11474_ _05434_ vssd1 vssd1 vccd1 vccd1 _00784_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13213_ clknet_leaf_7_clk _00536_ net49 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.b1\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10425_ _04651_ vssd1 vssd1 vccd1 vccd1 _04683_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_21_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13144_ clknet_leaf_121_clk net673 net81 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.quo\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07242__B1 _01183_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10356_ _04646_ vssd1 vssd1 vccd1 vccd1 _00454_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_103_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13075_ clknet_leaf_2_clk _00402_ net42 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.acc\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10287_ _04574_ _04597_ _04598_ vssd1 vssd1 vccd1 vccd1 _04599_ sky130_fd_sc_hd__a21o_1
XANTENNA__10129__B1 _04455_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10414__A _03719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12026_ genblk2\[10\].wave_shpr.div.quo\[4\] _05813_ _05817_ net682 vssd1 vssd1 vccd1
+ vccd1 _00953_ sky130_fd_sc_hd__a22o_1
XANTENNA__08019__A2_N _01732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12928_ clknet_leaf_35_clk _00259_ net118 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.acc\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12859_ clknet_leaf_132_clk _00190_ net64 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.b1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06380_ _01178_ _01176_ vssd1 vssd1 vccd1 vccd1 _01324_ sky130_fd_sc_hd__and2_1
XTAP_1590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08050_ genblk1\[5\].osc.clkdiv_C.cnt\[11\] _01355_ vssd1 vssd1 vccd1 vccd1 _02757_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_71_578 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07001_ _01823_ _01830_ _01831_ vssd1 vssd1 vccd1 vccd1 genblk1\[7\].osc.clkdiv_C.next_cnt\[5\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06802__A _01238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08952_ _03564_ _03563_ vssd1 vssd1 vccd1 vccd1 _03642_ sky130_fd_sc_hd__or2b_1
XANTENNA__07228__A2_N _01235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07903_ genblk1\[8\].osc.clkdiv_C.cnt\[11\] _01360_ _02011_ vssd1 vssd1 vccd1 vccd1
+ _02610_ sky130_fd_sc_hd__and3_1
XANTENNA__09525__A2 _04048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08883_ sig_norm.acc\[8\] _03588_ vssd1 vssd1 vccd1 vccd1 _03589_ sky130_fd_sc_hd__or2_1
XANTENNA_fanout195_A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07834_ _02537_ _02538_ _02540_ vssd1 vssd1 vccd1 vccd1 _02541_ sky130_fd_sc_hd__o21a_1
X_07765_ genblk1\[0\].osc.clkdiv_C.cnt\[15\] _01309_ _01208_ genblk1\[0\].osc.clkdiv_C.cnt\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02472_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06716_ _01604_ vssd1 vssd1 vccd1 vccd1 genblk1\[4\].osc.clkdiv_C.next_cnt\[1\] sky130_fd_sc_hd__clkbuf_1
X_09504_ _02159_ vssd1 vssd1 vccd1 vccd1 _04042_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_154_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07696_ _02398_ _02402_ genblk1\[10\].osc.clkdiv_C.cnt\[16\] genblk1\[10\].osc.clkdiv_C.cnt\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02403_ sky130_fd_sc_hd__a211o_4
XANTENNA__06249__A _01182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09435_ _03957_ _03997_ _03998_ vssd1 vssd1 vccd1 vccd1 _03999_ sky130_fd_sc_hd__a21o_1
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06647_ _01522_ _01543_ vssd1 vssd1 vccd1 vccd1 _01544_ sky130_fd_sc_hd__or2_1
XFILLER_0_94_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09366_ net1082 _03841_ _03839_ _03936_ vssd1 vssd1 vccd1 vccd1 _00174_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06578_ genblk1\[3\].osc.clkdiv_C.cnt\[11\] vssd1 vssd1 vccd1 vccd1 _01486_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08317_ _03018_ _03023_ vssd1 vssd1 vccd1 vccd1 _03024_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_35_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09297_ genblk2\[0\].wave_shpr.div.acc\[6\] _03885_ _03804_ vssd1 vssd1 vccd1 vccd1
+ _03886_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_832 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08248_ _02953_ _02954_ vssd1 vssd1 vccd1 vccd1 _02955_ sky130_fd_sc_hd__nor2_1
XFILLER_0_105_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_887 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12348__A1 _03944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08179_ genblk2\[3\].wave_shpr.div.fin_quo\[0\] genblk2\[3\].wave_shpr.div.fin_quo\[1\]
+ genblk2\[3\].wave_shpr.div.fin_quo\[2\] genblk2\[3\].wave_shpr.div.fin_quo\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02886_ sky130_fd_sc_hd__or4_1
XFILLER_0_104_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10210_ _04412_ _04535_ vssd1 vssd1 vccd1 vccd1 _04536_ sky130_fd_sc_hd__xnor2_1
X_11190_ _03831_ net768 _04241_ vssd1 vssd1 vccd1 vccd1 _00700_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_101_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10141_ genblk2\[3\].wave_shpr.div.b1\[0\] _04380_ _04381_ vssd1 vssd1 vccd1 vccd1
+ _04483_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13598__RESET_B net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold574_A genblk2\[6\].wave_shpr.div.quo\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_101_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09516__A2 _04043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10072_ _04446_ vssd1 vssd1 vccd1 vccd1 _00370_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13180__RESET_B net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13762_ clknet_leaf_69_clk net994 net214 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.acc\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10974_ _05059_ genblk1\[6\].osc.clkdiv_C.cnt\[11\] vssd1 vssd1 vccd1 vccd1 _05072_
+ sky130_fd_sc_hd__and2_1
XANTENNA__06159__A _01114_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_97_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12713_ clknet_leaf_55_clk genblk1\[9\].osc.clkdiv_C.next_cnt\[8\] net175 vssd1 vssd1
+ vccd1 vccd1 genblk1\[9\].osc.clkdiv_C.cnt\[8\] sky130_fd_sc_hd__dfrtp_1
X_13693_ clknet_leaf_45_clk _01004_ net122 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.i\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12036__B1 _05816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12644_ clknet_leaf_10_clk genblk1\[5\].osc.clkdiv_C.next_cnt\[11\] net57 vssd1 vssd1
+ vccd1 vccd1 genblk1\[5\].osc.clkdiv_C.cnt\[11\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_155_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12575_ clknet_leaf_29_clk genblk1\[1\].osc.clkdiv_C.next_cnt\[14\] net95 vssd1 vssd1
+ vccd1 vccd1 genblk1\[1\].osc.clkdiv_C.cnt\[14\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_25_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08093__B _01360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11004__S _05023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11526_ _05450_ genblk1\[8\].osc.clkdiv_C.cnt\[7\] vssd1 vssd1 vccd1 vccd1 _05460_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_41_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11457_ _05425_ vssd1 vssd1 vccd1 vccd1 _00776_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10408_ _04672_ genblk1\[4\].osc.clkdiv_C.cnt\[12\] vssd1 vssd1 vccd1 vccd1 _04673_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_123_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07718__A _01360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11388_ genblk2\[8\].wave_shpr.div.acc\[11\] genblk2\[8\].wave_shpr.div.b1\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05364_ sky130_fd_sc_hd__or2b_1
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_103_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10339_ _03732_ net708 _03717_ vssd1 vssd1 vccd1 vccd1 _00447_ sky130_fd_sc_hd__o21a_1
X_13127_ clknet_leaf_3_clk _00452_ net46 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.b1\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__13268__RESET_B net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13058_ clknet_leaf_24_clk _00385_ net92 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.quo\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_12009_ _05809_ vssd1 vssd1 vccd1 vccd1 _00944_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08268__B _02361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07550_ _02258_ vssd1 vssd1 vccd1 vccd1 _00036_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06501_ genblk1\[2\].osc.clkdiv_C.cnt\[15\] _01424_ _01425_ _01426_ vssd1 vssd1 vccd1
+ vccd1 _01427_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_88_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07481_ genblk2\[10\].wave_shpr.div.busy _02206_ vssd1 vssd1 vccd1 vccd1 _02207_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_124_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09220_ net655 _03836_ _03840_ net804 vssd1 vssd1 vccd1 vccd1 _00124_ sky130_fd_sc_hd__a22o_1
X_06432_ genblk1\[1\].osc.clkdiv_C.cnt\[1\] genblk1\[1\].osc.clkdiv_C.cnt\[0\] vssd1
+ vssd1 vccd1 vccd1 _01375_ sky130_fd_sc_hd__or2_1
XANTENNA__12027__B1 _05817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09151_ genblk2\[0\].wave_shpr.div.acc\[18\] _03798_ vssd1 vssd1 vccd1 vccd1 _03799_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_134_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_832 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06363_ genblk1\[1\].osc.clkdiv_C.cnt\[6\] vssd1 vssd1 vccd1 vccd1 _01307_ sky130_fd_sc_hd__inv_2
XFILLER_0_127_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_8_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_854 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08102_ genblk1\[4\].osc.clkdiv_C.cnt\[11\] _01574_ vssd1 vssd1 vccd1 vccd1 _02809_
+ sky130_fd_sc_hd__and2_1
XANTENNA__06516__B _01441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09082_ net702 vssd1 vssd1 vccd1 vccd1 _03734_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06294_ _01255_ vssd1 vssd1 vccd1 vccd1 _01256_ sky130_fd_sc_hd__buf_4
XFILLER_0_13_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08033_ _02699_ _02734_ _02738_ genblk2\[6\].wave_shpr.div.fin_quo\[6\] vssd1 vssd1
+ vccd1 vccd1 _02740_ sky130_fd_sc_hd__a31o_1
Xhold800 genblk2\[8\].wave_shpr.div.acc\[21\] vssd1 vssd1 vccd1 vccd1 net1018 sky130_fd_sc_hd__dlygate4sd3_1
Xhold811 genblk2\[7\].wave_shpr.div.acc\[24\] vssd1 vssd1 vccd1 vccd1 net1029 sky130_fd_sc_hd__dlygate4sd3_1
Xhold822 _00072_ vssd1 vssd1 vccd1 vccd1 net1040 sky130_fd_sc_hd__dlygate4sd3_1
Xhold833 genblk1\[2\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 net1051 sky130_fd_sc_hd__dlygate4sd3_1
Xhold844 genblk2\[5\].wave_shpr.div.acc\[1\] vssd1 vssd1 vccd1 vccd1 net1062 sky130_fd_sc_hd__dlygate4sd3_1
Xhold855 sig_norm.b1\[2\] vssd1 vssd1 vccd1 vccd1 net1073 sky130_fd_sc_hd__dlygate4sd3_1
Xhold866 genblk2\[0\].wave_shpr.div.b1\[11\] vssd1 vssd1 vccd1 vccd1 net1084 sky130_fd_sc_hd__dlygate4sd3_1
Xhold877 genblk1\[3\].osc.clkdiv_C.cnt\[7\] vssd1 vssd1 vccd1 vccd1 net1095 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold888 genblk2\[0\].wave_shpr.div.i\[1\] vssd1 vssd1 vccd1 vccd1 net1106 sky130_fd_sc_hd__dlygate4sd3_1
X_09984_ genblk2\[3\].wave_shpr.div.acc\[0\] vssd1 vssd1 vccd1 vccd1 _04380_ sky130_fd_sc_hd__inv_2
Xhold899 genblk2\[5\].wave_shpr.div.i\[1\] vssd1 vssd1 vccd1 vccd1 net1117 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09843__A _04269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08935_ net1083 _02260_ _03596_ _03574_ vssd1 vssd1 vccd1 vccd1 _00051_ sky130_fd_sc_hd__a22o_1
XANTENNA__06980__A2 _01578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08866_ net428 _02248_ _00024_ _03572_ vssd1 vssd1 vccd1 vccd1 _03573_ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07817_ net17 net18 vssd1 vssd1 vccd1 vccd1 _02524_ sky130_fd_sc_hd__and2b_2
X_08797_ _03501_ _03502_ _03500_ _03503_ vssd1 vssd1 vccd1 vccd1 _03504_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_98_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07082__B genblk1\[8\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07748_ genblk1\[1\].osc.clkdiv_C.cnt\[16\] _01576_ vssd1 vssd1 vccd1 vccd1 _02455_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_67_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07679_ _01489_ genblk1\[10\].osc.clkdiv_C.cnt\[13\] vssd1 vssd1 vccd1 vccd1 _02386_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07810__B net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09418_ _03965_ genblk2\[1\].wave_shpr.div.acc\[6\] _03981_ vssd1 vssd1 vccd1 vccd1
+ _03982_ sky130_fd_sc_hd__o21a_1
X_10690_ net233 _04861_ _04862_ net507 _04872_ vssd1 vssd1 vccd1 vccd1 _00562_ sky130_fd_sc_hd__a221o_1
XANTENNA__08194__A net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09349_ _03924_ _03925_ vssd1 vssd1 vccd1 vccd1 _03926_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12360_ _05946_ _06041_ vssd1 vssd1 vccd1 vccd1 _06042_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_63_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06799__A2 _01210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11311_ net894 _05279_ _05283_ _05307_ vssd1 vssd1 vccd1 vccd1 _00748_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11792__A2 genblk1\[9\].osc.clkdiv_C.cnt\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12291_ _06007_ vssd1 vssd1 vccd1 vccd1 _01028_ sky130_fd_sc_hd__clkbuf_1
X_11242_ _05260_ genblk1\[7\].osc.clkdiv_C.cnt\[6\] vssd1 vssd1 vccd1 vccd1 _05261_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_132_296 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11544__A2 _05441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11173_ genblk2\[7\].wave_shpr.div.fin_quo\[5\] genblk2\[7\].wave_shpr.div.quo\[4\]
+ _00019_ vssd1 vssd1 vccd1 vccd1 _05228_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10124_ _04465_ genblk1\[3\].osc.clkdiv_C.cnt\[12\] vssd1 vssd1 vccd1 vccd1 _04473_
+ sky130_fd_sc_hd__and2_1
X_10055_ net1178 _04436_ _04238_ vssd1 vssd1 vccd1 vccd1 _04437_ sky130_fd_sc_hd__mux2_1
XANTENNA__09370__B1 _03839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07920__A1 genblk1\[8\].osc.clkdiv_C.cnt\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10807__A1 _02183_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13745_ clknet_leaf_51_clk net439 net110 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.quo\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10957_ _05059_ genblk1\[6\].osc.clkdiv_C.cnt\[3\] vssd1 vssd1 vccd1 vccd1 _05063_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_70_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11523__A _05444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07684__A0 _01179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06487__B2 _01183_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11480__A1 _01732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13676_ clknet_leaf_42_clk _00989_ net124 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.acc\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10888_ genblk2\[6\].wave_shpr.div.fin_quo\[4\] net1319 _00017_ vssd1 vssd1 vccd1
+ vccd1 _05028_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12627_ clknet_leaf_120_clk genblk1\[4\].osc.clkdiv_C.next_cnt\[12\] net81 vssd1
+ vssd1 vccd1 vccd1 genblk1\[4\].osc.clkdiv_C.cnt\[12\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_109_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_81_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12558_ clknet_leaf_55_clk genblk1\[0\].osc.clkdiv_C.next_cnt\[15\] net176 vssd1
+ vssd1 vccd1 vccd1 genblk1\[0\].osc.clkdiv_C.cnt\[15\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_112_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11509_ _04268_ vssd1 vssd1 vccd1 vccd1 _05450_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_151_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12489_ clknet_leaf_107_clk _00051_ net151 vssd1 vssd1 vccd1 vccd1 sig_norm.quo\[0\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold107 _00568_ vssd1 vssd1 vccd1 vccd1 net325 sky130_fd_sc_hd__dlygate4sd3_1
Xhold118 genblk2\[2\].wave_shpr.div.quo\[3\] vssd1 vssd1 vccd1 vccd1 net336 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold129 _00799_ vssd1 vssd1 vccd1 vccd1 net347 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07448__A _02183_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07739__A1 genblk1\[1\].osc.clkdiv_C.cnt\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07739__B2 genblk1\[1\].osc.clkdiv_C.cnt\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08978__S _02248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08400__A2 _02425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06981_ _01809_ _01810_ _01812_ _01816_ vssd1 vssd1 vccd1 vccd1 _01817_ sky130_fd_sc_hd__and4b_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08720_ _03423_ _03424_ _03425_ _03426_ vssd1 vssd1 vccd1 vccd1 _03427_ sky130_fd_sc_hd__a211o_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08651_ _03351_ _03352_ _03356_ vssd1 vssd1 vccd1 vccd1 _03358_ sky130_fd_sc_hd__a21oi_2
X_07602_ _02308_ vssd1 vssd1 vccd1 vccd1 _02309_ sky130_fd_sc_hd__buf_4
X_08582_ genblk2\[10\].wave_shpr.div.fin_quo\[1\] _03286_ _03288_ vssd1 vssd1 vccd1
+ vccd1 _03289_ sky130_fd_sc_hd__o21a_1
XFILLER_0_49_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07533_ _02248_ _02249_ vssd1 vssd1 vccd1 vccd1 _02250_ sky130_fd_sc_hd__or2_1
XFILLER_0_49_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_659 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout158_A net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07464_ _02194_ vssd1 vssd1 vccd1 vccd1 _00019_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__07630__B _02336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09203_ net1251 _01302_ _03822_ vssd1 vssd1 vccd1 vccd1 _03830_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06415_ _01358_ vssd1 vssd1 vccd1 vccd1 _01359_ sky130_fd_sc_hd__buf_4
XFILLER_0_147_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07395_ _02080_ _02140_ vssd1 vssd1 vccd1 vccd1 _02143_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09134_ _03754_ _03780_ _03781_ vssd1 vssd1 vccd1 vccd1 _03782_ sky130_fd_sc_hd__a21o_1
X_06346_ genblk1\[0\].osc.clkdiv_C.cnt\[13\] _01291_ genblk1\[0\].osc.clkdiv_C.cnt\[14\]
+ vssd1 vssd1 vccd1 vccd1 _01294_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_127_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09065_ net1184 _01185_ _03722_ vssd1 vssd1 vccd1 vccd1 _03724_ sky130_fd_sc_hd__mux2_1
XANTENNA__10483__S _04704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06277_ _01173_ _01188_ _01191_ vssd1 vssd1 vccd1 vccd1 _01239_ sky130_fd_sc_hd__nor3b_2
XFILLER_0_130_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10982__B1 _05054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08016_ genblk1\[6\].osc.clkdiv_C.cnt\[6\] _01750_ _01739_ genblk1\[6\].osc.clkdiv_C.cnt\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02723_ sky130_fd_sc_hd__o22a_1
XFILLER_0_114_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold630 genblk1\[7\].osc.clkdiv_C.cnt\[17\] vssd1 vssd1 vccd1 vccd1 net848 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold641 genblk2\[10\].wave_shpr.div.acc\[17\] vssd1 vssd1 vccd1 vccd1 net859 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold652 genblk2\[10\].wave_shpr.div.acc\[16\] vssd1 vssd1 vccd1 vccd1 net870 sky130_fd_sc_hd__dlygate4sd3_1
Xhold663 genblk2\[4\].wave_shpr.div.acc\[16\] vssd1 vssd1 vccd1 vccd1 net881 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold674 genblk2\[9\].wave_shpr.div.acc\[23\] vssd1 vssd1 vccd1 vccd1 net892 sky130_fd_sc_hd__dlygate4sd3_1
Xhold685 genblk2\[2\].wave_shpr.div.acc\[8\] vssd1 vssd1 vccd1 vccd1 net903 sky130_fd_sc_hd__dlygate4sd3_1
Xhold696 genblk2\[2\].wave_shpr.div.acc_next\[0\] vssd1 vssd1 vccd1 vccd1 net914 sky130_fd_sc_hd__dlygate4sd3_1
X_09967_ genblk2\[3\].wave_shpr.div.acc\[15\] genblk2\[3\].wave_shpr.div.b1\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04363_ sky130_fd_sc_hd__or2b_1
X_08918_ net612 _02260_ _03617_ _03574_ vssd1 vssd1 vccd1 vccd1 _00045_ sky130_fd_sc_hd__a22o_1
X_09898_ genblk2\[2\].wave_shpr.div.acc\[11\] _04313_ _04301_ vssd1 vssd1 vccd1 vccd1
+ _04314_ sky130_fd_sc_hd__mux2_1
XTAP_990 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08849_ _03498_ _03553_ _03554_ vssd1 vssd1 vccd1 vccd1 _03556_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08384__A_N _01437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07902__A1 genblk1\[8\].osc.clkdiv_C.cnt\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11860_ net1060 _05684_ _05685_ _05697_ vssd1 vssd1 vccd1 vccd1 _00907_ sky130_fd_sc_hd__a22o_1
XTAP_2835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10811_ _04855_ _04957_ _04958_ _04858_ net1117 vssd1 vssd1 vccd1 vccd1 _00597_ sky130_fd_sc_hd__a32o_1
X_11791_ genblk2\[9\].wave_shpr.div.acc_next\[0\] _03693_ vssd1 vssd1 vccd1 vccd1
+ _05645_ sky130_fd_sc_hd__or2b_1
XANTENNA__09037__B1_N _03705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09655__A1 _04045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06469__A1 genblk1\[1\].osc.clkdiv_C.cnt\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13530_ clknet_leaf_98_clk _00847_ net169 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.acc\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11462__A1 _01797_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10742_ net772 _04886_ _04890_ _04908_ vssd1 vssd1 vccd1 vccd1 _00578_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10673_ net500 _04861_ _04862_ net572 _04863_ vssd1 vssd1 vccd1 vccd1 _00554_ sky130_fd_sc_hd__a221o_1
X_13461_ clknet_leaf_84_clk _00778_ net203 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.b1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12412_ genblk2\[11\].wave_shpr.div.acc\[15\] _06081_ _06055_ vssd1 vssd1 vccd1 vccd1
+ _06082_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13392_ clknet_leaf_91_clk _00711_ net143 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.quo\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12343_ genblk2\[11\].wave_shpr.div.acc_next\[0\] _03942_ _03941_ net412 _06029_
+ vssd1 vssd1 vccd1 vccd1 _01058_ sky130_fd_sc_hd__a221o_1
XFILLER_0_133_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08630__A2 _02733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12274_ _05998_ vssd1 vssd1 vccd1 vccd1 _01020_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08090__C _02365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11225_ genblk2\[7\].wave_shpr.div.quo\[8\] _05246_ _05250_ net421 vssd1 vssd1 vccd1
+ vccd1 _00719_ sky130_fd_sc_hd__a22o_1
X_11156_ _05164_ _05214_ _05215_ vssd1 vssd1 vccd1 vccd1 _05216_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10107_ _04269_ genblk1\[3\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 _04464_
+ sky130_fd_sc_hd__and2_1
X_11087_ genblk2\[6\].wave_shpr.div.acc\[25\] _05021_ genblk2\[6\].wave_shpr.div.acc\[24\]
+ genblk2\[6\].wave_shpr.div.acc\[26\] vssd1 vssd1 vccd1 vccd1 _05153_ sky130_fd_sc_hd__or4b_1
X_10038_ _04428_ vssd1 vssd1 vccd1 vccd1 _00354_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08449__A2 net30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11989_ _05799_ vssd1 vssd1 vccd1 vccd1 _00934_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_105_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13728_ clknet_leaf_97_clk _01039_ net167 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06347__A genblk1\[0\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_88 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_50_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13659_ clknet_leaf_47_clk net475 net120 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.quo\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_144_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06200_ PWM.counter\[4\] _01161_ net810 vssd1 vssd1 vccd1 vccd1 _01165_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11205__A1 _03831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07180_ genblk1\[9\].osc.clkdiv_C.cnt\[8\] genblk1\[9\].osc.clkdiv_C.cnt\[7\] _01967_
+ vssd1 vssd1 vccd1 vccd1 _01972_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06131_ net3 _01102_ vssd1 vssd1 vccd1 vccd1 _01103_ sky130_fd_sc_hd__xor2_1
XANTENNA_clkbuf_leaf_65_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12084__A _05815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09821_ _04069_ genblk1\[2\].osc.clkdiv_C.cnt\[5\] vssd1 vssd1 vccd1 vccd1 _04261_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_10_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09752_ genblk2\[3\].wave_shpr.div.b1\[0\] _04223_ _04039_ vssd1 vssd1 vccd1 vccd1
+ _04224_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_123_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10332__A _03717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06964_ genblk1\[7\].osc.clkdiv_C.cnt\[4\] _01799_ vssd1 vssd1 vccd1 vccd1 _01800_
+ sky130_fd_sc_hd__xnor2_1
X_08703_ _02586_ _03409_ vssd1 vssd1 vccd1 vccd1 _03410_ sky130_fd_sc_hd__nand2_1
X_09683_ genblk2\[2\].wave_shpr.div.acc\[10\] genblk2\[2\].wave_shpr.div.b1\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04163_ sky130_fd_sc_hd__or2b_1
X_06895_ genblk1\[6\].osc.clkdiv_C.cnt\[15\] _01362_ vssd1 vssd1 vccd1 vccd1 _01749_
+ sky130_fd_sc_hd__nor2_1
XTAP_2109 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08634_ genblk2\[8\].wave_shpr.div.fin_quo\[0\] genblk2\[8\].wave_shpr.div.fin_quo\[1\]
+ _02638_ vssd1 vssd1 vccd1 vccd1 _03341_ sky130_fd_sc_hd__o21ai_1
XANTENNA_clkbuf_leaf_138_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08565_ _02261_ _03270_ _03271_ _02950_ vssd1 vssd1 vccd1 vccd1 _03272_ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_65_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07516_ PWM.final_sample_in\[1\] _02235_ PWM.counter\[1\] vssd1 vssd1 vccd1 vccd1
+ _02236_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_76_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08496_ _03054_ _03076_ _03075_ vssd1 vssd1 vccd1 vccd1 _03203_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_49_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_18_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout46 net47 vssd1 vssd1 vccd1 vccd1 net46 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_147_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07447_ _02182_ vssd1 vssd1 vccd1 vccd1 _02183_ sky130_fd_sc_hd__clkbuf_4
Xfanout57 net58 vssd1 vssd1 vccd1 vccd1 net57 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_91_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout68 net85 vssd1 vssd1 vccd1 vccd1 net68 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout79 net84 vssd1 vssd1 vccd1 vccd1 net79 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_147_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07378_ _02128_ _02127_ vssd1 vssd1 vccd1 vccd1 _02130_ sky130_fd_sc_hd__nor2_1
XFILLER_0_17_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11747__A2 _05623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11135__A_N genblk2\[7\].wave_shpr.div.b1\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06329_ net592 _01281_ _01283_ vssd1 vssd1 vccd1 vccd1 genblk1\[0\].osc.clkdiv_C.next_cnt\[7\]
+ sky130_fd_sc_hd__a21oi_1
X_09117_ genblk2\[0\].wave_shpr.div.acc\[0\] genblk2\[0\].wave_shpr.div.b1\[0\] vssd1
+ vssd1 vccd1 vccd1 _03765_ sky130_fd_sc_hd__and2b_1
XFILLER_0_115_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08612__A2 _02521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10955__B1 _05055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06704__B _01592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09048_ genblk2\[0\].wave_shpr.div.b1\[4\] _03712_ _03708_ vssd1 vssd1 vccd1 vccd1
+ _03713_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold460 sig_norm.acc\[8\] vssd1 vssd1 vccd1 vccd1 net678 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold471 _00168_ vssd1 vssd1 vccd1 vccd1 net689 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout90_A net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold482 genblk2\[9\].wave_shpr.div.quo\[3\] vssd1 vssd1 vccd1 vccd1 net700 sky130_fd_sc_hd__dlygate4sd3_1
X_11010_ net907 _05086_ _05093_ _05096_ vssd1 vssd1 vccd1 vccd1 _00658_ sky130_fd_sc_hd__a22o_1
XFILLER_0_130_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12172__A2 _05818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold493 genblk2\[2\].wave_shpr.div.i\[2\] vssd1 vssd1 vccd1 vccd1 net711 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06387__B1 _01329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11380__B1 _03855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12961_ clknet_leaf_139_clk _00290_ net39 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.b1\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_11912_ genblk2\[10\].wave_shpr.div.acc\[14\] genblk2\[10\].wave_shpr.div.b1\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05734_ sky130_fd_sc_hd__or2b_1
XTAP_2610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12892_ clknet_leaf_28_clk net463 net91 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.quo\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11843_ _02203_ vssd1 vssd1 vccd1 vccd1 _05684_ sky130_fd_sc_hd__clkbuf_4
XTAP_2665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10238__A2 _04457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11774_ genblk2\[9\].wave_shpr.div.quo\[17\] _05628_ _05629_ net349 _05636_ vssd1
+ vssd1 vccd1 vccd1 _00882_ sky130_fd_sc_hd__a221o_1
XTAP_1975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13513_ clknet_leaf_78_clk _00830_ net205 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.acc\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10725_ net885 _04886_ _04890_ _04895_ vssd1 vssd1 vccd1 vccd1 _00574_ sky130_fd_sc_hd__a22o_1
XTAP_1997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11801__A _02203_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13444_ clknet_leaf_95_clk net382 net149 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.acc\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_10656_ _04856_ vssd1 vssd1 vccd1 vccd1 _04857_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_70_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12108__S _05865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10587_ _04763_ _04813_ _04814_ vssd1 vssd1 vccd1 vccd1 _04815_ sky130_fd_sc_hd__a21o_1
XANTENNA__08603__A2 _02885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13375_ clknet_leaf_86_clk _00694_ net179 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.b1\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_134_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10946__B1 _05056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10417__A _04672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12326_ _03689_ genblk1\[11\].osc.clkdiv_C.cnt\[8\] vssd1 vssd1 vccd1 vccd1 _06021_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_23_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12257_ genblk2\[11\].wave_shpr.div.fin_quo\[6\] net1332 _00005_ vssd1 vssd1 vccd1
+ vccd1 _05989_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12163__A2 _05818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11208_ _03726_ _05243_ _03736_ vssd1 vssd1 vccd1 vccd1 _00709_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07726__A _01342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12188_ genblk2\[11\].wave_shpr.div.b1\[16\] genblk2\[11\].wave_shpr.div.acc\[16\]
+ vssd1 vssd1 vccd1 vccd1 _05926_ sky130_fd_sc_hd__xor2_1
X_11139_ genblk2\[7\].wave_shpr.div.b1\[9\] genblk2\[7\].wave_shpr.div.acc\[9\] vssd1
+ vssd1 vccd1 vccd1 _05199_ sky130_fd_sc_hd__and2b_1
XANTENNA__07590__A2 _01991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06680_ genblk1\[4\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 _01570_ sky130_fd_sc_hd__inv_2
XANTENNA__07461__A _02155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08350_ genblk2\[5\].wave_shpr.div.fin_quo\[4\] _03056_ _02527_ vssd1 vssd1 vccd1
+ vccd1 _03057_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07301_ genblk1\[11\].osc.clkdiv_C.cnt\[6\] _01595_ vssd1 vssd1 vccd1 vccd1 _02065_
+ sky130_fd_sc_hd__nor2_1
X_08281_ genblk2\[9\].wave_shpr.div.fin_quo\[5\] _02521_ _02310_ vssd1 vssd1 vccd1
+ vccd1 _02988_ sky130_fd_sc_hd__a21o_1
XFILLER_0_117_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_62_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07232_ genblk1\[10\].osc.clkdiv_C.cnt\[0\] _01321_ _02013_ genblk1\[10\].osc.clkdiv_C.cnt\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02014_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_143_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07163_ genblk1\[9\].osc.clkdiv_C.cnt\[3\] _01958_ vssd1 vssd1 vccd1 vccd1 _01960_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06114_ net368 _01086_ vssd1 vssd1 vccd1 vccd1 _01091_ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07094_ genblk1\[8\].osc.clkdiv_C.cnt\[9\] _01900_ vssd1 vssd1 vccd1 vccd1 _01903_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10046__B _01996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout203 net204 vssd1 vssd1 vccd1 vccd1 net203 sky130_fd_sc_hd__clkbuf_4
XANTENNA__09555__B1 _04046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout214 net217 vssd1 vssd1 vccd1 vccd1 net214 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_5_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09804_ genblk2\[2\].wave_shpr.div.quo\[5\] _04248_ _04252_ net696 vssd1 vssd1 vccd1
+ vccd1 _00296_ sky130_fd_sc_hd__a22o_1
X_07996_ _02701_ _02702_ vssd1 vssd1 vccd1 vccd1 _02703_ sky130_fd_sc_hd__or2b_1
XANTENNA__07581__A2 _01437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09735_ genblk2\[2\].wave_shpr.div.fin_quo\[0\] _04214_ _00009_ vssd1 vssd1 vccd1
+ vccd1 _04215_ sky130_fd_sc_hd__mux2_1
X_06947_ net1104 _01783_ _01786_ vssd1 vssd1 vccd1 vccd1 genblk1\[6\].osc.clkdiv_C.next_cnt\[14\]
+ sky130_fd_sc_hd__o21a_1
XANTENNA__10997__A _05051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09666_ _04045_ _04148_ _04149_ _04048_ net1091 vssd1 vssd1 vccd1 vccd1 _00261_ sky130_fd_sc_hd__a32o_1
X_06878_ _01731_ vssd1 vssd1 vccd1 vccd1 _01732_ sky130_fd_sc_hd__buf_4
XFILLER_0_96_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08617_ genblk2\[4\].wave_shpr.div.fin_quo\[2\] _02362_ _02838_ vssd1 vssd1 vccd1
+ vccd1 _03324_ sky130_fd_sc_hd__a21o_1
XTAP_1205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09597_ net847 _04076_ _04080_ _04099_ vssd1 vssd1 vccd1 vccd1 _00242_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07090__B genblk1\[8\].osc.clkdiv_C.cnt\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08548_ _02742_ _03254_ _02745_ vssd1 vssd1 vccd1 vccd1 _03255_ sky130_fd_sc_hd__o21a_1
X_08479_ _02838_ _03185_ _02846_ vssd1 vssd1 vccd1 vccd1 _03186_ sky130_fd_sc_hd__o21a_1
X_10510_ _04745_ _04619_ genblk2\[4\].wave_shpr.div.acc\[22\] vssd1 vssd1 vccd1 vccd1
+ _04747_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11490_ _05440_ vssd1 vssd1 vccd1 vccd1 _00794_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10441_ net970 _04683_ _04690_ _04695_ vssd1 vssd1 vccd1 vccd1 _00490_ sky130_fd_sc_hd__a22o_1
XANTENNA__08046__B1 _01666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10372_ genblk2\[4\].wave_shpr.div.quo\[1\] _04652_ _04656_ net418 vssd1 vssd1 vccd1
+ vccd1 _00460_ sky130_fd_sc_hd__a22o_1
X_13160_ clknet_leaf_122_clk _00485_ net78 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.acc\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_60_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12111_ _05763_ _05870_ vssd1 vssd1 vccd1 vccd1 _05871_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_20_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13091_ clknet_leaf_137_clk _00418_ net39 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.acc\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12042_ _05815_ vssd1 vssd1 vccd1 vccd1 _05825_ sky130_fd_sc_hd__clkbuf_4
Xhold290 genblk2\[4\].wave_shpr.div.quo\[6\] vssd1 vssd1 vccd1 vccd1 net508 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_46_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09761__A _01436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12944_ clknet_leaf_2_clk _00273_ net42 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.b1\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11656__A1 _05449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07324__A2 _01334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12875_ clknet_leaf_138_clk _00206_ net39 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.b1\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11826_ _05588_ _05563_ vssd1 vssd1 vccd1 vccd1 _05671_ sky130_fd_sc_hd__or2b_1
XTAP_2495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07088__A1 genblk1\[8\].osc.clkdiv_C.cnt\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_134_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_134_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11757_ genblk2\[9\].wave_shpr.div.quo\[10\] _03696_ _03694_ net290 _05626_ vssd1
+ vssd1 vccd1 vccd1 _00875_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10092__B1 _04456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10708_ _04855_ _04881_ _04882_ _04858_ net1062 vssd1 vssd1 vccd1 vccd1 _00570_ sky130_fd_sc_hd__a32o_1
X_11688_ _05570_ _05578_ _05579_ vssd1 vssd1 vccd1 vccd1 _05580_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_141_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13427_ clknet_leaf_87_clk _00746_ net201 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.acc\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10639_ net1248 _04225_ _04834_ vssd1 vssd1 vccd1 vccd1 _04847_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13358_ clknet_leaf_4_clk _00679_ net46 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.acc\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08052__A3 net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12309_ genblk2\[11\].wave_shpr.div.quo\[9\] _03947_ _03944_ net355 _06011_ vssd1
+ vssd1 vccd1 vccd1 _01042_ sky130_fd_sc_hd__a221o_1
X_13289_ clknet_leaf_92_clk _00610_ net147 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.b1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_07850_ genblk2\[1\].wave_shpr.div.fin_quo\[2\] _02461_ _02462_ _02316_ vssd1 vssd1
+ vccd1 vccd1 _02557_ sky130_fd_sc_hd__a31o_1
XANTENNA__10698__A2 _02183_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07563__A2 _01556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06801_ _01669_ _01559_ _01671_ _01436_ _01672_ vssd1 vssd1 vccd1 vccd1 _01673_ sky130_fd_sc_hd__a221o_1
X_07781_ genblk1\[0\].osc.clkdiv_C.cnt\[5\] _02483_ _02484_ _02486_ _02487_ vssd1
+ vssd1 vccd1 vccd1 _02488_ sky130_fd_sc_hd__a2111o_1
Xinput3 pb[11] vssd1 vssd1 vccd1 vccd1 net3 sky130_fd_sc_hd__clkbuf_4
X_09520_ _03855_ _01330_ vssd1 vssd1 vccd1 vccd1 _04049_ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06732_ _01616_ vssd1 vssd1 vccd1 vccd1 _01617_ sky130_fd_sc_hd__inv_2
XANTENNA__07903__B _01360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07315__A2 _01211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09451_ _04013_ vssd1 vssd1 vccd1 vccd1 _00182_ sky130_fd_sc_hd__clkbuf_1
X_06663_ _01524_ _01553_ _01554_ vssd1 vssd1 vccd1 vccd1 _01555_ sky130_fd_sc_hd__and3_1
XFILLER_0_94_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_819 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08402_ genblk1\[2\].osc.clkdiv_C.cnt\[11\] _01411_ _03102_ _03106_ _03108_ vssd1
+ vssd1 vccd1 vccd1 _03109_ sky130_fd_sc_hd__a2111o_1
X_06594_ genblk1\[3\].osc.clkdiv_C.cnt\[6\] _01500_ _01496_ genblk1\[3\].osc.clkdiv_C.cnt\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01502_ sky130_fd_sc_hd__o2bb2a_1
X_09382_ genblk2\[11\].wave_shpr.div.i\[1\] genblk2\[11\].wave_shpr.div.i\[0\] genblk2\[11\].wave_shpr.div.i\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03949_ sky130_fd_sc_hd__and3_1
XFILLER_0_148_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08333_ _03037_ _03038_ _03039_ _02694_ vssd1 vssd1 vccd1 vccd1 _03040_ sky130_fd_sc_hd__a211o_1
XFILLER_0_52_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_125_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_125_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_19_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout140_A net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08264_ _02915_ _02910_ vssd1 vssd1 vccd1 vccd1 _02971_ sky130_fd_sc_hd__or2b_1
XFILLER_0_74_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_342 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07215_ _01490_ _01993_ genblk1\[10\].osc.clkdiv_C.cnt\[2\] vssd1 vssd1 vccd1 vccd1
+ _01997_ sky130_fd_sc_hd__o21ai_1
X_08195_ _02349_ _02351_ _02355_ genblk2\[11\].wave_shpr.div.fin_quo\[5\] vssd1 vssd1
+ vccd1 vccd1 _02902_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_61_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07146_ _01336_ _01496_ vssd1 vssd1 vccd1 vccd1 _01946_ sky130_fd_sc_hd__nor2_4
XFILLER_0_30_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10491__S _04704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07077_ genblk1\[8\].osc.clkdiv_C.cnt\[3\] _01890_ vssd1 vssd1 vccd1 vccd1 _01892_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_113_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07979_ genblk2\[7\].wave_shpr.div.fin_quo\[0\] genblk2\[7\].wave_shpr.div.fin_quo\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02686_ sky130_fd_sc_hd__nor2_1
X_09718_ _04161_ _04196_ _04197_ vssd1 vssd1 vccd1 vccd1 _04198_ sky130_fd_sc_hd__a21o_1
X_10990_ genblk2\[6\].wave_shpr.div.b1\[0\] _05023_ genblk2\[6\].wave_shpr.div.acc\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05081_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_69_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout53_A net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07306__A2 _01678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09649_ genblk2\[1\].wave_shpr.div.acc\[22\] _04109_ _04113_ _04138_ vssd1 vssd1
+ vccd1 vccd1 _00255_ sky130_fd_sc_hd__a22o_1
XTAP_1002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12660_ clknet_leaf_26_clk genblk1\[6\].osc.clkdiv_C.next_cnt\[9\] net87 vssd1 vssd1
+ vccd1 vccd1 genblk1\[6\].osc.clkdiv_C.cnt\[9\] sky130_fd_sc_hd__dfrtp_4
XTAP_1046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11611_ net947 _05507_ _05445_ _05519_ vssd1 vssd1 vccd1 vccd1 _00836_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08267__B1 _02222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_148_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_116_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_116_clk
+ sky130_fd_sc_hd__clkbuf_16
X_12591_ clknet_leaf_13_clk genblk1\[2\].osc.clkdiv_C.next_cnt\[12\] net70 vssd1 vssd1
+ vccd1 vccd1 genblk1\[2\].osc.clkdiv_C.cnt\[12\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_26_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11542_ genblk2\[8\].wave_shpr.div.quo\[23\] _05441_ _05458_ net229 _05468_ vssd1
+ vssd1 vccd1 vccd1 _00818_ sky130_fd_sc_hd__a221o_1
XFILLER_0_107_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11473_ genblk2\[9\].wave_shpr.div.b1\[7\] _04230_ _05433_ vssd1 vssd1 vccd1 vccd1
+ _05434_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09767__B1 _04233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13212_ clknet_leaf_25_clk _00535_ net86 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.b1\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10424_ _04681_ _04682_ net1129 _04652_ vssd1 vssd1 vccd1 vccd1 _00486_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_104_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08660__A _02789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13143_ clknet_leaf_121_clk net252 net81 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.quo\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10355_ genblk2\[5\].wave_shpr.div.b1\[13\] _04645_ _04637_ vssd1 vssd1 vccd1 vccd1
+ _04646_ sky130_fd_sc_hd__mux2_1
XFILLER_0_131_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10286_ genblk2\[4\].wave_shpr.div.b1\[8\] genblk2\[4\].wave_shpr.div.acc\[8\] vssd1
+ vssd1 vccd1 vccd1 _04598_ sky130_fd_sc_hd__and2b_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13074_ clknet_leaf_11_clk net437 net56 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.acc\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_12025_ net682 _05813_ _05817_ net724 vssd1 vssd1 vccd1 vccd1 _00952_ sky130_fd_sc_hd__a22o_1
XANTENNA__12121__S _05865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12927_ clknet_leaf_35_clk _00258_ net106 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.acc\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06505__B1 _01196_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12858_ clknet_leaf_134_clk _00189_ net60 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.b1\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08835__A net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_206 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__13056__RESET_B net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11809_ genblk2\[9\].wave_shpr.div.acc\[3\] _05658_ _05613_ vssd1 vssd1 vccd1 vccd1
+ _05659_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_107_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_107_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12789_ clknet_leaf_43_clk _00122_ net124 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.b1\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12357__A _03942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_407 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06355__A genblk1\[0\].osc.clkdiv_C.cnt\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_790 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07000_ genblk1\[7\].osc.clkdiv_C.cnt\[4\] _01827_ genblk1\[7\].osc.clkdiv_C.cnt\[5\]
+ vssd1 vssd1 vccd1 vccd1 _01831_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_126_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09222__A2 _03836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06802__B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12109__A2 _05844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08951_ _03641_ vssd1 vssd1 vccd1 vccd1 _00054_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_138_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07902_ genblk1\[8\].osc.clkdiv_C.cnt\[12\] _01328_ _02607_ _02608_ vssd1 vssd1 vccd1
+ vccd1 _02609_ sky130_fd_sc_hd__a211o_1
X_08882_ sig_norm.acc\[7\] sig_norm.acc\[6\] sig_norm.acc\[5\] _03587_ vssd1 vssd1
+ vccd1 vccd1 _03588_ sky130_fd_sc_hd__or4_1
XANTENNA_clkbuf_4_4_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07833_ genblk2\[1\].wave_shpr.div.fin_quo\[5\] _02539_ _02469_ vssd1 vssd1 vccd1
+ vccd1 _02540_ sky130_fd_sc_hd__a21oi_1
XANTENNA_fanout188_A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07764_ _02465_ _02466_ _02470_ vssd1 vssd1 vccd1 vccd1 _02471_ sky130_fd_sc_hd__o21a_1
XFILLER_0_2_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09503_ _03714_ _04041_ _03736_ vssd1 vssd1 vccd1 vccd1 _00206_ sky130_fd_sc_hd__o21ai_1
X_06715_ _01600_ _01602_ _01603_ vssd1 vssd1 vccd1 vccd1 _01604_ sky130_fd_sc_hd__and3_1
XFILLER_0_2_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07695_ _02016_ _02390_ _02393_ _02400_ _02401_ vssd1 vssd1 vccd1 vccd1 _02402_ sky130_fd_sc_hd__a221oi_2
X_09434_ genblk2\[1\].wave_shpr.div.b1\[14\] genblk2\[1\].wave_shpr.div.acc\[14\]
+ vssd1 vssd1 vccd1 vccd1 _03998_ sky130_fd_sc_hd__and2b_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06646_ _01486_ _01542_ vssd1 vssd1 vccd1 vccd1 _01543_ sky130_fd_sc_hd__nor2_1
XFILLER_0_137_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09365_ _03934_ _03802_ genblk2\[0\].wave_shpr.div.acc\[24\] vssd1 vssd1 vccd1 vccd1
+ _03936_ sky130_fd_sc_hd__mux2_1
X_06577_ genblk1\[3\].osc.clkdiv_C.cnt\[8\] vssd1 vssd1 vccd1 vccd1 _01485_ sky130_fd_sc_hd__inv_2
XANTENNA__12267__A _03707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08316_ _02419_ _03022_ vssd1 vssd1 vccd1 vccd1 _03023_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06265__A _01224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09296_ _03774_ _03884_ vssd1 vssd1 vccd1 vccd1 _03885_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08247_ genblk2\[8\].wave_shpr.div.fin_quo\[5\] _02638_ _02952_ _02223_ vssd1 vssd1
+ vccd1 vccd1 _02954_ sky130_fd_sc_hd__a31o_1
XFILLER_0_62_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10359__A1 _01365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08178_ _02853_ _02878_ _02884_ genblk1\[3\].osc.clkdiv_C.cnt\[17\] genblk1\[3\].osc.clkdiv_C.cnt\[16\]
+ vssd1 vssd1 vccd1 vccd1 _02885_ sky130_fd_sc_hd__a311o_4
XANTENNA__11556__B1 _05448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07129_ genblk1\[9\].osc.clkdiv_C.cnt\[9\] _01801_ vssd1 vssd1 vccd1 vccd1 _01929_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10140_ _04454_ _04481_ _04482_ _04457_ net1067 vssd1 vssd1 vccd1 vccd1 _00402_ sky130_fd_sc_hd__a32o_1
XANTENNA__07775__A2 _01227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10234__B _04480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10071_ net1281 _01595_ _04440_ vssd1 vssd1 vccd1 vccd1 _04446_ sky130_fd_sc_hd__mux2_1
XANTENNA__10250__A _03690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap21 net1350 vssd1 vssd1 vccd1 vccd1 net21 sky130_fd_sc_hd__buf_1
XFILLER_0_97_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13761_ clknet_leaf_70_clk _01072_ net214 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.acc\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10973_ net313 _05062_ _05064_ net486 _05071_ vssd1 vssd1 vccd1 vccd1 _00646_ sky130_fd_sc_hd__a221o_1
XFILLER_0_97_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12712_ clknet_leaf_55_clk genblk1\[9\].osc.clkdiv_C.next_cnt\[7\] net175 vssd1 vssd1
+ vccd1 vccd1 genblk1\[9\].osc.clkdiv_C.cnt\[7\] sky130_fd_sc_hd__dfrtp_4
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13692_ clknet_leaf_44_clk _01003_ net122 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.i\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_12643_ clknet_leaf_10_clk genblk1\[5\].osc.clkdiv_C.next_cnt\[10\] net56 vssd1 vssd1
+ vccd1 vccd1 genblk1\[5\].osc.clkdiv_C.cnt\[10\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_38_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12574_ clknet_leaf_29_clk genblk1\[1\].osc.clkdiv_C.next_cnt\[13\] net89 vssd1 vssd1
+ vccd1 vccd1 genblk1\[1\].osc.clkdiv_C.cnt\[13\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_26_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11525_ genblk2\[8\].wave_shpr.div.quo\[15\] _05454_ _05458_ net237 _05459_ vssd1
+ vssd1 vccd1 vccd1 _00810_ sky130_fd_sc_hd__a221o_1
XFILLER_0_92_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12339__A2 _03942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11456_ genblk2\[8\].wave_shpr.div.fin_quo\[7\] net1335 _00021_ vssd1 vssd1 vccd1
+ vccd1 _05425_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07215__A1 _01490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10407_ _04268_ vssd1 vssd1 vccd1 vccd1 _04672_ sky130_fd_sc_hd__buf_2
XANTENNA__12116__S _05865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07718__B _01302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10425__A _04651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11387_ genblk2\[8\].wave_shpr.div.acc\[12\] genblk2\[8\].wave_shpr.div.b1\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05363_ sky130_fd_sc_hd__or2b_1
XFILLER_0_0_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13126_ clknet_leaf_3_clk _00451_ net51 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.b1\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10338_ _03831_ net625 _03733_ vssd1 vssd1 vccd1 vccd1 _00446_ sky130_fd_sc_hd__a21bo_1
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13057_ clknet_leaf_24_clk net539 net92 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.quo\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10269_ genblk2\[4\].wave_shpr.div.acc\[3\] genblk2\[4\].wave_shpr.div.b1\[3\] vssd1
+ vssd1 vccd1 vccd1 _04581_ sky130_fd_sc_hd__or2b_1
XFILLER_0_84_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_84_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12008_ genblk2\[11\].wave_shpr.div.b1\[13\] _01483_ _05802_ vssd1 vssd1 vccd1 vccd1
+ _05809_ sky130_fd_sc_hd__mux2_1
XANTENNA__12275__A1 _01311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06500_ genblk1\[2\].osc.clkdiv_C.cnt\[13\] genblk1\[2\].osc.clkdiv_C.cnt\[0\] net35
+ vssd1 vssd1 vccd1 vccd1 _01426_ sky130_fd_sc_hd__and3_1
X_07480_ genblk2\[10\].wave_shpr.div.i\[1\] _02205_ genblk2\[10\].wave_shpr.div.i\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02206_ sky130_fd_sc_hd__or3b_1
XFILLER_0_124_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06431_ net29 vssd1 vssd1 vccd1 vccd1 _01374_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09150_ _03746_ _03796_ _03797_ vssd1 vssd1 vccd1 vccd1 _03798_ sky130_fd_sc_hd__a21o_1
XFILLER_0_17_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06362_ genblk1\[1\].osc.clkdiv_C.cnt\[5\] _01305_ vssd1 vssd1 vccd1 vccd1 _01306_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_16_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_56_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11786__B1 _03693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08101_ _02804_ _02807_ vssd1 vssd1 vccd1 vccd1 _02808_ sky130_fd_sc_hd__or2_1
X_09081_ _03704_ net396 _03717_ vssd1 vssd1 vccd1 vccd1 _00092_ sky130_fd_sc_hd__a21bo_1
X_06293_ _01196_ _01254_ vssd1 vssd1 vccd1 vccd1 _01255_ sky130_fd_sc_hd__nor2_1
XFILLER_0_154_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_25_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08032_ _02699_ genblk2\[6\].wave_shpr.div.fin_quo\[6\] _02734_ _02738_ _02261_ vssd1
+ vssd1 vccd1 vccd1 _02739_ sky130_fd_sc_hd__a41o_1
XFILLER_0_114_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06813__A genblk1\[5\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold801 genblk2\[1\].wave_shpr.div.acc\[14\] vssd1 vssd1 vccd1 vccd1 net1019 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold812 genblk2\[7\].wave_shpr.div.acc\[5\] vssd1 vssd1 vccd1 vccd1 net1030 sky130_fd_sc_hd__dlygate4sd3_1
Xhold823 genblk2\[5\].wave_shpr.div.acc\[25\] vssd1 vssd1 vccd1 vccd1 net1041 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_114_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold834 genblk2\[8\].wave_shpr.div.acc\[25\] vssd1 vssd1 vccd1 vccd1 net1052 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11387__B_N genblk2\[8\].wave_shpr.div.b1\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold845 genblk1\[6\].osc.clkdiv_C.cnt\[17\] vssd1 vssd1 vccd1 vccd1 net1063 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold856 genblk2\[4\].wave_shpr.div.acc\[18\] vssd1 vssd1 vccd1 vccd1 net1074 sky130_fd_sc_hd__dlygate4sd3_1
Xhold867 genblk2\[9\].wave_shpr.div.quo\[7\] vssd1 vssd1 vccd1 vccd1 net1085 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_149_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold878 genblk2\[6\].wave_shpr.div.b1\[16\] vssd1 vssd1 vccd1 vccd1 net1096 sky130_fd_sc_hd__dlygate4sd3_1
Xhold889 genblk2\[1\].wave_shpr.div.acc\[26\] vssd1 vssd1 vccd1 vccd1 net1107 sky130_fd_sc_hd__dlygate4sd3_1
X_09983_ genblk2\[3\].wave_shpr.div.b1\[1\] vssd1 vssd1 vccd1 vccd1 _04379_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08934_ _01099_ _00024_ _03627_ _03628_ vssd1 vssd1 vccd1 vccd1 _00050_ sky130_fd_sc_hd__a31o_1
XANTENNA__07644__A _02350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08865_ _03009_ _03134_ _03571_ _02248_ vssd1 vssd1 vccd1 vccd1 _03572_ sky130_fd_sc_hd__o31ai_2
X_07816_ genblk2\[1\].wave_shpr.div.fin_quo\[3\] _02522_ vssd1 vssd1 vccd1 vccd1 _02523_
+ sky130_fd_sc_hd__xor2_1
X_08796_ _03395_ _03499_ _03484_ _03498_ vssd1 vssd1 vccd1 vccd1 _03503_ sky130_fd_sc_hd__a211oi_2
X_07747_ genblk1\[1\].osc.clkdiv_C.cnt\[15\] _01172_ vssd1 vssd1 vccd1 vccd1 _02454_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_95_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07678_ genblk1\[10\].osc.clkdiv_C.cnt\[9\] _01215_ _01991_ _02003_ vssd1 vssd1 vccd1
+ vccd1 _02385_ sky130_fd_sc_hd__a2bb2o_1
X_09417_ _03966_ _03979_ _03980_ vssd1 vssd1 vccd1 vccd1 _03981_ sky130_fd_sc_hd__o21bai_1
X_06629_ net1077 _01530_ _01532_ vssd1 vssd1 vccd1 vccd1 genblk1\[3\].osc.clkdiv_C.next_cnt\[4\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_48_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08194__B net163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09348_ _03798_ net23 genblk2\[0\].wave_shpr.div.acc\[18\] vssd1 vssd1 vccd1 vccd1
+ _03925_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_63_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_81_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09279_ _03766_ _03871_ vssd1 vssd1 vccd1 vccd1 _03872_ sky130_fd_sc_hd__xnor2_1
X_11310_ genblk2\[7\].wave_shpr.div.acc\[10\] _05306_ _05300_ vssd1 vssd1 vccd1 vccd1
+ _05307_ sky130_fd_sc_hd__mux2_1
XANTENNA__07819__A _02525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12290_ net1299 _01249_ _05994_ vssd1 vssd1 vccd1 vccd1 _06007_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11241_ _04268_ vssd1 vssd1 vccd1 vccd1 _05260_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_120_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11172_ _05227_ vssd1 vssd1 vccd1 vccd1 _00689_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10792__A2_N _04880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06956__B1 _01732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10123_ genblk2\[3\].wave_shpr.div.quo\[20\] _04461_ _04462_ net296 _04472_ vssd1
+ vssd1 vccd1 vccd1 _00395_ sky130_fd_sc_hd__a221o_1
XANTENNA__06420__A2 _01363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07554__A _02223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10054_ _01557_ vssd1 vssd1 vccd1 vccd1 _04436_ sky130_fd_sc_hd__inv_2
XANTENNA__07920__A2 _01430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13330__RESET_B net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13744_ clknet_leaf_51_clk _01055_ net110 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.quo\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10956_ _05051_ vssd1 vssd1 vccd1 vccd1 _05062_ sky130_fd_sc_hd__buf_2
XANTENNA__09205__B1_N _03728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13675_ clknet_leaf_42_clk _00988_ net125 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.acc\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10887_ _05027_ vssd1 vssd1 vccd1 vccd1 _00604_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12626_ clknet_leaf_16_clk genblk1\[4\].osc.clkdiv_C.next_cnt\[11\] net74 vssd1 vssd1
+ vccd1 vccd1 genblk1\[4\].osc.clkdiv_C.cnt\[11\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_26_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_81_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_54_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12557_ clknet_leaf_55_clk genblk1\[0\].osc.clkdiv_C.next_cnt\[14\] net175 vssd1
+ vssd1 vccd1 vccd1 genblk1\[0\].osc.clkdiv_C.cnt\[14\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_41_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_540 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11508_ _05444_ vssd1 vssd1 vccd1 vccd1 _05449_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_80_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12488_ clknet_leaf_107_clk _00050_ net151 vssd1 vssd1 vccd1 vccd1 sig_norm.acc\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold108 genblk2\[3\].wave_shpr.div.quo\[1\] vssd1 vssd1 vccd1 vccd1 net326 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold119 _00295_ vssd1 vssd1 vccd1 vccd1 net337 sky130_fd_sc_hd__dlygate4sd3_1
X_11439_ genblk2\[8\].wave_shpr.div.acc\[25\] genblk2\[8\].wave_shpr.div.acc\[26\]
+ _05414_ vssd1 vssd1 vccd1 vccd1 _05415_ sky130_fd_sc_hd__or3_1
XFILLER_0_21_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06352__B genblk1\[0\].osc.clkdiv_C.cnt\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07739__A2 _01334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13109_ clknet_leaf_114_clk _00434_ net133 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.fin_quo\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06980_ genblk1\[7\].osc.clkdiv_C.cnt\[16\] _01578_ _01574_ genblk1\[7\].osc.clkdiv_C.cnt\[7\]
+ _01815_ vssd1 vssd1 vccd1 vccd1 _01816_ sky130_fd_sc_hd__o221a_1
XFILLER_0_28_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08650_ _03351_ _03352_ _03356_ vssd1 vssd1 vccd1 vccd1 _03357_ sky130_fd_sc_hd__and3_2
X_07601_ _02307_ vssd1 vssd1 vccd1 vccd1 _02308_ sky130_fd_sc_hd__buf_4
XANTENNA__07911__A2 _01308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08581_ _03285_ _03287_ _02404_ _02525_ vssd1 vssd1 vccd1 vccd1 _03288_ sky130_fd_sc_hd__o31a_1
XFILLER_0_88_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07532_ _01151_ _02245_ vssd1 vssd1 vccd1 vccd1 _02249_ sky130_fd_sc_hd__nor2_1
XANTENNA__13000__RESET_B net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07463_ _02191_ _02153_ genblk2\[7\].wave_shpr.div.busy vssd1 vssd1 vccd1 vccd1 _02194_
+ sky130_fd_sc_hd__and3b_1
XANTENNA__07630__C net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09202_ _03829_ vssd1 vssd1 vccd1 vccd1 _00117_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06414_ _01178_ freq_div.state\[2\] vssd1 vssd1 vccd1 vccd1 _01358_ sky130_fd_sc_hd__or2_1
XFILLER_0_119_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07394_ _02080_ _02140_ _02142_ _02092_ vssd1 vssd1 vccd1 vccd1 genblk1\[11\].osc.clkdiv_C.next_cnt\[15\]
+ sky130_fd_sc_hd__o211a_1
XANTENNA__11759__B1 _03694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_72_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09133_ genblk2\[0\].wave_shpr.div.b1\[9\] genblk2\[0\].wave_shpr.div.acc\[9\] vssd1
+ vssd1 vccd1 vccd1 _03781_ sky130_fd_sc_hd__and2b_1
XANTENNA__11223__A2 _05246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06345_ genblk1\[0\].osc.clkdiv_C.cnt\[13\] _01291_ _01293_ vssd1 vssd1 vccd1 vccd1
+ genblk1\[0\].osc.clkdiv_C.next_cnt\[13\] sky130_fd_sc_hd__o21a_1
XFILLER_0_60_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06276_ _01237_ vssd1 vssd1 vccd1 vccd1 _01238_ sky130_fd_sc_hd__clkbuf_8
X_09064_ _03723_ vssd1 vssd1 vccd1 vccd1 _00085_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08015_ _02721_ _02719_ genblk1\[6\].osc.clkdiv_C.cnt\[6\] _01750_ vssd1 vssd1 vccd1
+ vccd1 _02722_ sky130_fd_sc_hd__a2bb2o_1
Xhold620 genblk2\[6\].wave_shpr.div.acc\[12\] vssd1 vssd1 vccd1 vccd1 net838 sky130_fd_sc_hd__dlygate4sd3_1
Xhold631 genblk2\[3\].wave_shpr.div.quo\[4\] vssd1 vssd1 vccd1 vccd1 net849 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold642 _00992_ vssd1 vssd1 vccd1 vccd1 net860 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold653 genblk2\[8\].wave_shpr.div.quo\[1\] vssd1 vssd1 vccd1 vccd1 net871 sky130_fd_sc_hd__dlygate4sd3_1
Xhold664 genblk2\[5\].wave_shpr.div.quo\[2\] vssd1 vssd1 vccd1 vccd1 net882 sky130_fd_sc_hd__dlygate4sd3_1
Xhold675 genblk2\[7\].wave_shpr.div.acc\[7\] vssd1 vssd1 vccd1 vccd1 net893 sky130_fd_sc_hd__dlygate4sd3_1
Xhold686 genblk2\[3\].wave_shpr.div.acc\[19\] vssd1 vssd1 vccd1 vccd1 net904 sky130_fd_sc_hd__dlygate4sd3_1
Xhold697 _00317_ vssd1 vssd1 vccd1 vccd1 net915 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06402__A2 _01340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09966_ _04245_ genblk2\[3\].wave_shpr.div.acc\[16\] vssd1 vssd1 vccd1 vccd1 _04362_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__09065__S _03722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08917_ sig_norm.acc\[6\] _03614_ vssd1 vssd1 vccd1 vccd1 _03617_ sky130_fd_sc_hd__xnor2_1
X_09897_ _04194_ _04312_ vssd1 vssd1 vccd1 vccd1 _04313_ sky130_fd_sc_hd__xnor2_1
XTAP_980 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_991 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_96_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_96_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_85_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08155__A2 _01483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08848_ _03498_ _03553_ _03554_ vssd1 vssd1 vccd1 vccd1 _03555_ sky130_fd_sc_hd__or3_1
XANTENNA__07902__A2 _01328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08779_ _02518_ _02566_ _02570_ vssd1 vssd1 vccd1 vccd1 _03486_ sky130_fd_sc_hd__a21oi_1
XTAP_2836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10810_ genblk2\[5\].wave_shpr.div.i\[1\] genblk2\[5\].wave_shpr.div.i\[0\] vssd1
+ vssd1 vccd1 vccd1 _04958_ sky130_fd_sc_hd__nand2_1
X_11790_ genblk2\[9\].wave_shpr.div.acc_next\[0\] _02203_ _03693_ net306 _05644_ vssd1
+ vssd1 vccd1 vccd1 _00890_ sky130_fd_sc_hd__a221o_1
XFILLER_0_138_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08636__C genblk2\[8\].wave_shpr.div.fin_quo\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_149_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10741_ genblk2\[5\].wave_shpr.div.acc\[8\] _04906_ _04907_ vssd1 vssd1 vccd1 vccd1
+ _04908_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07666__B2 _01190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13460_ clknet_leaf_84_clk _00777_ net203 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.b1\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_10672_ _04672_ genblk1\[5\].osc.clkdiv_C.cnt\[2\] vssd1 vssd1 vccd1 vccd1 _04863_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_94_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12411_ _05970_ _06080_ vssd1 vssd1 vccd1 vccd1 _06081_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08615__B1 _02223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13391_ clknet_leaf_79_clk _00710_ net206 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.b1\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_20_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_20_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_105_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12342_ _03689_ genblk1\[11\].osc.clkdiv_C.cnt\[16\] vssd1 vssd1 vccd1 vccd1 _06029_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_51_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06453__A genblk1\[1\].osc.clkdiv_C.cnt\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12273_ net1272 _05997_ _05994_ vssd1 vssd1 vccd1 vccd1 _05998_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_4_12_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11224_ genblk2\[7\].wave_shpr.div.quo\[7\] _05246_ _05250_ net317 vssd1 vssd1 vccd1
+ vccd1 _00718_ sky130_fd_sc_hd__a22o_1
X_11155_ genblk2\[7\].wave_shpr.div.b1\[17\] genblk2\[7\].wave_shpr.div.acc\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05215_ sky130_fd_sc_hd__and2b_1
X_10106_ net387 _04461_ _04462_ net525 _04463_ vssd1 vssd1 vccd1 vccd1 _00387_ sky130_fd_sc_hd__a221o_1
X_11086_ genblk2\[6\].wave_shpr.div.acc\[24\] _05021_ genblk2\[6\].wave_shpr.div.acc\[25\]
+ vssd1 vssd1 vccd1 vccd1 _05152_ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_87_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_87_clk sky130_fd_sc_hd__clkbuf_16
X_10037_ genblk2\[3\].wave_shpr.div.fin_quo\[5\] genblk2\[3\].wave_shpr.div.quo\[4\]
+ _04422_ vssd1 vssd1 vccd1 vccd1 _04428_ sky130_fd_sc_hd__mux2_1
XANTENNA__11534__A _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09774__B1_N _03733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11988_ net1265 _01946_ _05433_ vssd1 vssd1 vccd1 vccd1 _05799_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13727_ clknet_leaf_97_clk _01038_ net167 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10939_ _05054_ vssd1 vssd1 vccd1 vccd1 _05056_ sky130_fd_sc_hd__buf_4
XFILLER_0_128_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10661__B1 _04857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13658_ clknet_leaf_44_clk net335 net120 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.quo\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_27_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_38_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_73_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12609_ clknet_leaf_22_clk genblk1\[3\].osc.clkdiv_C.next_cnt\[12\] net94 vssd1 vssd1
+ vccd1 vccd1 genblk1\[3\].osc.clkdiv_C.cnt\[12\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_144_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06880__A2 _01684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13589_ clknet_leaf_72_clk _00904_ net215 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.acc\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_11_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_11_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_81_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06130_ _01100_ _01101_ vssd1 vssd1 vccd1 vccd1 _01102_ sky130_fd_sc_hd__nand2_1
XFILLER_0_54_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10413__B1 _04654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08989__S _01155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12166__B1 _05818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09820_ net457 _04257_ _04259_ net553 _04260_ vssd1 vssd1 vccd1 vccd1 _00304_ sky130_fd_sc_hd__a221o_1
XANTENNA__08385__A2 _01439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06810__B _01326_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07194__A genblk1\[9\].osc.clkdiv_C.cnt\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09751_ _01211_ _01302_ vssd1 vssd1 vccd1 vccd1 _04223_ sky130_fd_sc_hd__nor2_2
X_06963_ _01229_ _01230_ _01238_ vssd1 vssd1 vccd1 vccd1 _01799_ sky130_fd_sc_hd__a21oi_4
Xclkbuf_leaf_78_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_78_clk sky130_fd_sc_hd__clkbuf_16
X_08702_ _02561_ _02585_ _02548_ vssd1 vssd1 vccd1 vccd1 _03409_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_146_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09682_ genblk2\[2\].wave_shpr.div.acc\[11\] genblk2\[2\].wave_shpr.div.b1\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04162_ sky130_fd_sc_hd__or2b_1
X_06894_ genblk1\[6\].osc.clkdiv_C.cnt\[5\] _01747_ vssd1 vssd1 vccd1 vccd1 _01748_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_146_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09613__S _04095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08633_ _02742_ _03338_ _03339_ _02745_ vssd1 vssd1 vccd1 vccd1 _03340_ sky130_fd_sc_hd__o31a_1
XANTENNA_fanout170_A net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08564_ genblk2\[7\].wave_shpr.div.fin_quo\[2\] _02521_ vssd1 vssd1 vccd1 vccd1 _03271_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_147_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07515_ PWM.next_counter\[0\] PWM.final_sample_in\[0\] vssd1 vssd1 vccd1 vccd1 _02235_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_65_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08495_ _03175_ _03200_ _03201_ vssd1 vssd1 vccd1 vccd1 _03202_ sky130_fd_sc_hd__nor3_2
XFILLER_0_9_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_49_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout47 net50 vssd1 vssd1 vccd1 vccd1 net47 sky130_fd_sc_hd__buf_2
XFILLER_0_9_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07446_ _02147_ _02181_ vssd1 vssd1 vccd1 vccd1 _02182_ sky130_fd_sc_hd__nor2_1
Xfanout58 net85 vssd1 vssd1 vccd1 vccd1 net58 sky130_fd_sc_hd__clkbuf_2
XANTENNA__06320__A1 genblk1\[0\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout69 net75 vssd1 vssd1 vccd1 vccd1 net69 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_91_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_909 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07377_ _02128_ _02127_ _02129_ _02092_ vssd1 vssd1 vccd1 vccd1 genblk1\[11\].osc.clkdiv_C.next_cnt\[11\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_128_890 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09116_ _03762_ _03763_ vssd1 vssd1 vccd1 vccd1 _03764_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06328_ genblk1\[0\].osc.clkdiv_C.cnt\[7\] _01281_ _01270_ vssd1 vssd1 vccd1 vccd1
+ _01283_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06273__A _01231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09047_ _01248_ _02374_ vssd1 vssd1 vccd1 vccd1 _03712_ sky130_fd_sc_hd__nor2_2
XFILLER_0_142_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06259_ _01194_ _01175_ vssd1 vssd1 vccd1 vccd1 _01221_ sky130_fd_sc_hd__nand2b_4
XFILLER_0_130_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold450 genblk2\[6\].wave_shpr.div.quo\[24\] vssd1 vssd1 vccd1 vccd1 net668 sky130_fd_sc_hd__dlygate4sd3_1
Xhold461 genblk2\[7\].wave_shpr.div.acc\[21\] vssd1 vssd1 vccd1 vccd1 net679 sky130_fd_sc_hd__dlygate4sd3_1
Xhold472 genblk2\[8\].wave_shpr.div.acc\[20\] vssd1 vssd1 vccd1 vccd1 net690 sky130_fd_sc_hd__dlygate4sd3_1
Xhold483 genblk2\[1\].wave_shpr.div.quo\[3\] vssd1 vssd1 vccd1 vccd1 net701 sky130_fd_sc_hd__dlygate4sd3_1
Xhold494 genblk2\[9\].wave_shpr.div.quo\[5\] vssd1 vssd1 vccd1 vccd1 net712 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout83_A net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09949_ _04349_ _04350_ vssd1 vssd1 vccd1 vccd1 _04351_ sky130_fd_sc_hd__nand2_1
Xclkbuf_leaf_69_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_69_clk sky130_fd_sc_hd__clkbuf_16
X_12960_ clknet_leaf_137_clk _00289_ net39 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.b1\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_11911_ genblk2\[10\].wave_shpr.div.acc\[15\] genblk2\[10\].wave_shpr.div.b1\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05733_ sky130_fd_sc_hd__or2b_1
XANTENNA__07832__A _02309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12891_ clknet_leaf_28_clk net512 net91 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.quo\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11842_ net1046 _05652_ _05653_ _05683_ vssd1 vssd1 vccd1 vccd1 _00903_ sky130_fd_sc_hd__a22o_1
XFILLER_0_67_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_129_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_906 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11773_ _04676_ _01928_ vssd1 vssd1 vccd1 vccd1 _05636_ sky130_fd_sc_hd__nor2_1
XFILLER_0_138_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13512_ clknet_leaf_78_clk _00829_ net205 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.acc\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10724_ genblk2\[5\].wave_shpr.div.acc\[4\] _04894_ _04821_ vssd1 vssd1 vccd1 vccd1
+ _04895_ sky130_fd_sc_hd__mux2_1
XTAP_1987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13443_ clknet_leaf_92_clk _00762_ net149 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.acc\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10655_ _04854_ vssd1 vssd1 vccd1 vccd1 _04856_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_125_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13374_ clknet_leaf_96_clk _00693_ net167 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.b1\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10586_ genblk2\[5\].wave_shpr.div.b1\[17\] genblk2\[5\].wave_shpr.div.acc\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04814_ sky130_fd_sc_hd__and2b_1
XFILLER_0_23_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09800__A2 _04248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12325_ genblk2\[11\].wave_shpr.div.quo\[16\] _06014_ _06015_ net351 _06020_ vssd1
+ vssd1 vccd1 vccd1 _01049_ sky130_fd_sc_hd__a221o_1
XANTENNA__06614__A2 _01483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12256_ _05988_ vssd1 vssd1 vccd1 vccd1 _01012_ sky130_fd_sc_hd__clkbuf_1
X_11207_ net703 vssd1 vssd1 vccd1 vccd1 _05243_ sky130_fd_sc_hd__inv_2
XANTENNA__07726__B _01241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12187_ genblk2\[11\].wave_shpr.div.acc\[17\] genblk2\[11\].wave_shpr.div.b1\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05925_ sky130_fd_sc_hd__or2b_1
X_11138_ _05173_ _05196_ _05197_ vssd1 vssd1 vccd1 vccd1 _05198_ sky130_fd_sc_hd__a21o_1
X_11069_ net622 _05119_ _05126_ _05141_ vssd1 vssd1 vccd1 vccd1 _00672_ sky130_fd_sc_hd__a22o_1
XFILLER_0_92_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_0_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_92_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10882__A0 genblk2\[6\].wave_shpr.div.fin_quo\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_59_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08827__B1 _02468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07300_ _01182_ _01226_ vssd1 vssd1 vccd1 vccd1 _02064_ sky130_fd_sc_hd__nor2_4
XFILLER_0_128_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08280_ _02985_ _02986_ vssd1 vssd1 vccd1 vccd1 _02987_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_490 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07231_ _01225_ _01354_ vssd1 vssd1 vccd1 vccd1 _02013_ sky130_fd_sc_hd__nor2_2
XFILLER_0_128_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_73_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06805__B _01362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08055__A1 _01309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07162_ _01953_ _01958_ _01959_ vssd1 vssd1 vccd1 vccd1 genblk1\[9\].osc.clkdiv_C.next_cnt\[2\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_143_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06113_ _01086_ net360 vssd1 vssd1 vccd1 vccd1 smpl_rt_clkdiv.clkDiv_inst.next_cnt\[2\]
+ sky130_fd_sc_hd__nor2_1
X_07093_ genblk1\[8\].osc.clkdiv_C.cnt\[9\] _01900_ vssd1 vssd1 vccd1 vccd1 _01902_
+ sky130_fd_sc_hd__and2_1
XANTENNA__09608__S _04095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout204 net210 vssd1 vssd1 vccd1 vccd1 net204 sky130_fd_sc_hd__buf_2
Xfanout215 net217 vssd1 vssd1 vccd1 vccd1 net215 sky130_fd_sc_hd__clkbuf_4
X_09803_ genblk2\[2\].wave_shpr.div.quo\[4\] _04248_ _04252_ net336 vssd1 vssd1 vccd1
+ vccd1 _00295_ sky130_fd_sc_hd__a22o_1
X_07995_ genblk1\[6\].osc.clkdiv_C.cnt\[10\] _01484_ _01742_ genblk1\[6\].osc.clkdiv_C.cnt\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02702_ sky130_fd_sc_hd__a22oi_1
X_09734_ _04213_ vssd1 vssd1 vccd1 vccd1 _04214_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__07581__A3 _01226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06946_ net1356 _01785_ vssd1 vssd1 vccd1 vccd1 _01786_ sky130_fd_sc_hd__nor2_1
XANTENNA__08748__A net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12311__B1 _03944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07652__A _02316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09665_ genblk2\[1\].wave_shpr.div.i\[1\] genblk2\[1\].wave_shpr.div.i\[0\] vssd1
+ vssd1 vccd1 vccd1 _04149_ sky130_fd_sc_hd__nand2_1
X_06877_ _01177_ _01249_ vssd1 vssd1 vccd1 vccd1 _01731_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08616_ _03321_ _03322_ vssd1 vssd1 vccd1 vccd1 _03323_ sky130_fd_sc_hd__nor2_1
XTAP_1206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09596_ genblk2\[1\].wave_shpr.div.acc\[8\] _04098_ _04095_ vssd1 vssd1 vccd1 vccd1
+ _04099_ sky130_fd_sc_hd__mux2_1
XTAP_1217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08186__C _02365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08547_ genblk2\[6\].wave_shpr.div.fin_quo\[0\] _02527_ _02309_ genblk2\[6\].wave_shpr.div.fin_quo\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03254_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08478_ _03183_ _03184_ genblk2\[4\].wave_shpr.div.fin_quo\[4\] _02308_ vssd1 vssd1
+ vccd1 vccd1 _03185_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_53_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07429_ _02155_ _02168_ vssd1 vssd1 vccd1 vccd1 _02169_ sky130_fd_sc_hd__nor2_1
XFILLER_0_92_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07099__A genblk1\[8\].osc.clkdiv_C.cnt\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_808 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10440_ genblk2\[4\].wave_shpr.div.acc\[4\] _04694_ _04623_ vssd1 vssd1 vccd1 vccd1
+ _04695_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06882__A2_N _01732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10371_ _04654_ vssd1 vssd1 vccd1 vccd1 _04656_ sky130_fd_sc_hd__buf_2
XFILLER_0_32_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_21_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_131_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12110_ _05764_ _05739_ vssd1 vssd1 vccd1 vccd1 _05870_ sky130_fd_sc_hd__or2b_1
XFILLER_0_103_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13090_ clknet_leaf_137_clk _00417_ net39 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.acc\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_12041_ genblk2\[10\].wave_shpr.div.quo\[12\] _05823_ _05816_ net223 _05824_ vssd1
+ vssd1 vccd1 vccd1 _00961_ sky130_fd_sc_hd__a221o_1
Xhold280 genblk2\[6\].wave_shpr.div.quo\[14\] vssd1 vssd1 vccd1 vccd1 net498 sky130_fd_sc_hd__dlygate4sd3_1
Xhold291 genblk2\[11\].wave_shpr.div.quo\[18\] vssd1 vssd1 vccd1 vccd1 net509 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09761__B _04229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12302__B1 _06010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12943_ clknet_leaf_111_clk _00272_ net130 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.fin_quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_64_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12874_ clknet_leaf_136_clk _00205_ net42 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.b1\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_62_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08096__C _01359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11825_ net839 _05652_ _05653_ _05670_ vssd1 vssd1 vccd1 vccd1 _00899_ sky130_fd_sc_hd__a22o_1
XTAP_2474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11756_ _05464_ genblk1\[9\].osc.clkdiv_C.cnt\[1\] vssd1 vssd1 vccd1 vccd1 _05626_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_138_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_79_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10707_ genblk2\[5\].wave_shpr.div.b1\[0\] _04821_ genblk2\[5\].wave_shpr.div.acc\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04882_ sky130_fd_sc_hd__a21o_1
XFILLER_0_55_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11687_ genblk2\[9\].wave_shpr.div.b1\[3\] genblk2\[9\].wave_shpr.div.acc\[3\] vssd1
+ vssd1 vccd1 vccd1 _05579_ sky130_fd_sc_hd__and2b_1
XFILLER_0_153_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_122_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12346__C _05982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13426_ clknet_leaf_82_clk _00745_ net201 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.acc\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10638_ _04846_ vssd1 vssd1 vccd1 vccd1 _00536_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09234__B1 _03839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09785__A1 _04242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13357_ clknet_leaf_4_clk _00678_ net45 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.acc\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_688 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10569_ _04772_ _04795_ _04796_ vssd1 vssd1 vccd1 vccd1 _04797_ sky130_fd_sc_hd__a21o_1
XFILLER_0_23_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07737__A genblk1\[1\].osc.clkdiv_C.cnt\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12308_ _05835_ genblk1\[11\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 _06011_
+ sky130_fd_sc_hd__and2_1
X_13288_ clknet_leaf_90_clk _00609_ net147 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.b1\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_137_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12239_ genblk2\[11\].wave_shpr.div.acc\[18\] _05976_ vssd1 vssd1 vccd1 vccd1 _05977_
+ sky130_fd_sc_hd__or2_1
XANTENNA__07456__B _02153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_17_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06800_ genblk1\[5\].osc.clkdiv_C.cnt\[11\] _01667_ _01666_ genblk1\[5\].osc.clkdiv_C.cnt\[13\]
+ vssd1 vssd1 vccd1 vccd1 _01672_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__08760__A2 _02521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07563__A3 _01564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07780_ genblk1\[0\].osc.clkdiv_C.cnt\[5\] _02483_ _01215_ genblk1\[0\].osc.clkdiv_C.cnt\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02487_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_36_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput4 pb[12] vssd1 vssd1 vccd1 vccd1 net4 sky130_fd_sc_hd__clkbuf_1
X_06731_ genblk1\[4\].osc.clkdiv_C.cnt\[5\] genblk1\[4\].osc.clkdiv_C.cnt\[4\] _01609_
+ vssd1 vssd1 vccd1 vccd1 _01616_ sky130_fd_sc_hd__and3_1
XANTENNA__11647__A2 _05448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07903__C _02011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09450_ genblk2\[1\].wave_shpr.div.fin_quo\[1\] genblk2\[1\].wave_shpr.div.quo\[0\]
+ _00007_ vssd1 vssd1 vccd1 vccd1 _04013_ sky130_fd_sc_hd__mux2_1
X_06662_ genblk1\[3\].osc.clkdiv_C.cnt\[16\] _01551_ vssd1 vssd1 vccd1 vccd1 _01554_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_149_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07720__B1 _01208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08401_ genblk1\[2\].osc.clkdiv_C.cnt\[12\] _01591_ _03107_ vssd1 vssd1 vccd1 vccd1
+ _03108_ sky130_fd_sc_hd__a21bo_1
X_09381_ genblk2\[11\].wave_shpr.div.i\[1\] genblk2\[11\].wave_shpr.div.i\[0\] genblk2\[11\].wave_shpr.div.i\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03948_ sky130_fd_sc_hd__a21o_1
X_06593_ genblk1\[3\].osc.clkdiv_C.cnt\[14\] _01498_ _01500_ genblk1\[3\].osc.clkdiv_C.cnt\[6\]
+ vssd1 vssd1 vccd1 vccd1 _01501_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_59_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08332_ _02217_ _02553_ genblk2\[7\].wave_shpr.div.fin_quo\[5\] vssd1 vssd1 vccd1
+ vccd1 _03039_ sky130_fd_sc_hd__and3_1
XFILLER_0_129_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08263_ _02899_ _02923_ vssd1 vssd1 vccd1 vccd1 _02970_ sky130_fd_sc_hd__xnor2_1
XANTENNA_clkbuf_4_0_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07214_ _01181_ _01187_ vssd1 vssd1 vccd1 vccd1 _01996_ sky130_fd_sc_hd__nor2_4
XFILLER_0_27_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08194_ net3 net163 _02312_ vssd1 vssd1 vccd1 vccd1 _02901_ sky130_fd_sc_hd__and3_1
XANTENNA__09225__B1 _03840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07145_ genblk1\[9\].osc.clkdiv_C.cnt\[8\] _01514_ _01513_ genblk1\[9\].osc.clkdiv_C.cnt\[7\]
+ vssd1 vssd1 vccd1 vccd1 _01945_ sky130_fd_sc_hd__o22a_1
XFILLER_0_15_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_30_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10386__A2 _04657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07076_ _01887_ _01890_ _01891_ vssd1 vssd1 vccd1 vccd1 genblk1\[8\].osc.clkdiv_C.next_cnt\[2\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_10_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07978_ genblk2\[7\].wave_shpr.div.fin_quo\[2\] vssd1 vssd1 vccd1 vccd1 _02685_ sky130_fd_sc_hd__inv_2
X_09717_ genblk2\[2\].wave_shpr.div.b1\[12\] genblk2\[2\].wave_shpr.div.acc\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04197_ sky130_fd_sc_hd__and2b_1
X_06929_ _01761_ _01773_ _01774_ vssd1 vssd1 vccd1 vccd1 genblk1\[6\].osc.clkdiv_C.next_cnt\[8\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_97_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08197__B _02361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09648_ genblk2\[1\].wave_shpr.div.acc\[21\] _04136_ vssd1 vssd1 vccd1 vccd1 _04138_
+ sky130_fd_sc_hd__xor2_1
XTAP_1003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_78_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09579_ genblk2\[1\].wave_shpr.div.acc\[4\] _04085_ _04011_ vssd1 vssd1 vccd1 vccd1
+ _04086_ sky130_fd_sc_hd__mux2_1
XTAP_1047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_93_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11610_ net846 _05518_ _05493_ vssd1 vssd1 vccd1 vccd1 _05519_ sky130_fd_sc_hd__mux2_1
XTAP_1069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12590_ clknet_leaf_13_clk genblk1\[2\].osc.clkdiv_C.next_cnt\[11\] net70 vssd1 vssd1
+ vccd1 vccd1 genblk1\[2\].osc.clkdiv_C.cnt\[11\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_77_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11541_ _05464_ genblk1\[8\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 _05468_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_93_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11472_ _03707_ vssd1 vssd1 vccd1 vccd1 _05433_ sky130_fd_sc_hd__clkbuf_4
X_13211_ clknet_leaf_25_clk _00534_ net86 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.b1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10423_ genblk2\[4\].wave_shpr.div.b1\[0\] genblk2\[4\].wave_shpr.div.acc\[0\] _04623_
+ _04679_ vssd1 vssd1 vccd1 vccd1 _04682_ sky130_fd_sc_hd__a31o_1
XANTENNA__09767__A1 _03704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_446 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13142_ clknet_leaf_115_clk _00467_ net135 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.quo\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10354_ _01490_ _01242_ vssd1 vssd1 vccd1 vccd1 _04645_ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13073_ clknet_leaf_23_clk net562 net98 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.acc_next\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10285_ _04575_ _04595_ _04596_ vssd1 vssd1 vccd1 vccd1 _04597_ sky130_fd_sc_hd__a21o_1
XANTENNA__10129__A2 _04451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12024_ genblk2\[10\].wave_shpr.div.quo\[2\] _05813_ _05817_ net220 vssd1 vssd1 vccd1
+ vccd1 _00951_ sky130_fd_sc_hd__a22o_1
XANTENNA__11526__B genblk1\[8\].osc.clkdiv_C.cnt\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12926_ clknet_leaf_35_clk _00257_ net106 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.acc\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06505__A1 _01362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12857_ clknet_leaf_91_clk _00188_ net146 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.fin_quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11808_ _05578_ _05657_ vssd1 vssd1 vccd1 vccd1 _05658_ sky130_fd_sc_hd__xnor2_1
X_12788_ clknet_leaf_43_clk _00121_ net124 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.b1\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11739_ _01099_ _01147_ _05622_ net1161 vssd1 vssd1 vccd1 vccd1 _00861_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_83_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_114_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09758__A1 _04227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13409_ clknet_leaf_90_clk net549 net144 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.quo\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_113_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07769__B1 _01240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07233__A2 _01363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08950_ sig_norm.quo\[3\] _03640_ _00024_ vssd1 vssd1 vccd1 vccd1 _03641_ sky130_fd_sc_hd__mux2_1
X_07901_ genblk1\[8\].osc.clkdiv_C.cnt\[13\] _01246_ _01328_ genblk1\[8\].osc.clkdiv_C.cnt\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02608_ sky130_fd_sc_hd__o22ai_1
X_08881_ sig_norm.acc\[4\] _03586_ vssd1 vssd1 vccd1 vccd1 _03587_ sky130_fd_sc_hd__or2_1
XFILLER_0_138_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07832_ _02309_ vssd1 vssd1 vccd1 vccd1 _02539_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_138_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07763_ genblk2\[1\].wave_shpr.div.fin_quo\[6\] _02468_ _02469_ vssd1 vssd1 vccd1
+ vccd1 _02470_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09502_ net761 vssd1 vssd1 vccd1 vccd1 _04041_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06714_ genblk1\[4\].osc.clkdiv_C.cnt\[1\] genblk1\[4\].osc.clkdiv_C.cnt\[0\] vssd1
+ vssd1 vccd1 vccd1 _01603_ sky130_fd_sc_hd__nand2_1
X_07694_ _02386_ _02392_ _02387_ vssd1 vssd1 vccd1 vccd1 _02401_ sky130_fd_sc_hd__and3_1
XFILLER_0_154_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09433_ _03958_ _03995_ _03996_ vssd1 vssd1 vccd1 vccd1 _03997_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06645_ genblk1\[3\].osc.clkdiv_C.cnt\[10\] _01540_ _01542_ _01524_ vssd1 vssd1 vccd1
+ vccd1 genblk1\[3\].osc.clkdiv_C.next_cnt\[10\] sky130_fd_sc_hd__o211a_1
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09364_ net1305 _03841_ _03910_ _03935_ vssd1 vssd1 vccd1 vccd1 _00173_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06576_ _01182_ _01302_ vssd1 vssd1 vccd1 vccd1 _01484_ sky130_fd_sc_hd__or2_2
X_08315_ _03019_ _03020_ _03021_ _02416_ vssd1 vssd1 vccd1 vccd1 _03022_ sky130_fd_sc_hd__a211o_1
XFILLER_0_129_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09295_ _03775_ _03757_ vssd1 vssd1 vccd1 vccd1 _03884_ sky130_fd_sc_hd__or2b_1
XANTENNA__06265__B _01226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09857__A _04247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08246_ _02638_ _02952_ genblk2\[8\].wave_shpr.div.fin_quo\[5\] vssd1 vssd1 vccd1
+ vccd1 _02953_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_90_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08761__A net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11005__B1 _05056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08177_ _02868_ _02879_ _02883_ _02864_ vssd1 vssd1 vccd1 vccd1 _02884_ sky130_fd_sc_hd__a31o_1
XFILLER_0_30_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11556__A1 _05449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07128_ genblk1\[9\].osc.clkdiv_C.cnt\[8\] vssd1 vssd1 vccd1 vccd1 _01928_ sky130_fd_sc_hd__inv_2
X_07059_ genblk1\[8\].osc.clkdiv_C.cnt\[4\] _01866_ _01869_ genblk1\[8\].osc.clkdiv_C.cnt\[12\]
+ vssd1 vssd1 vccd1 vccd1 _01877_ sky130_fd_sc_hd__a22o_1
XFILLER_0_112_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10070_ _04445_ vssd1 vssd1 vccd1 vccd1 _00369_ sky130_fd_sc_hd__clkbuf_1
Xmax_cap22 net1351 vssd1 vssd1 vccd1 vccd1 net22 sky130_fd_sc_hd__buf_1
XFILLER_0_69_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13760_ clknet_leaf_70_clk _01071_ net213 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.acc\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10972_ _05059_ genblk1\[6\].osc.clkdiv_C.cnt\[10\] vssd1 vssd1 vccd1 vccd1 _05071_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_69_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12711_ clknet_leaf_56_clk genblk1\[9\].osc.clkdiv_C.next_cnt\[6\] net175 vssd1 vssd1
+ vccd1 vccd1 genblk1\[9\].osc.clkdiv_C.cnt\[6\] sky130_fd_sc_hd__dfrtp_4
X_13691_ clknet_leaf_44_clk _01002_ net122 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.i\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_69_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12642_ clknet_leaf_10_clk genblk1\[5\].osc.clkdiv_C.next_cnt\[9\] net56 vssd1 vssd1
+ vccd1 vccd1 genblk1\[5\].osc.clkdiv_C.cnt\[9\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_84_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12036__A2 _05818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06456__A genblk1\[1\].osc.clkdiv_C.cnt\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10047__B2 _03687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12573_ clknet_leaf_29_clk genblk1\[1\].osc.clkdiv_C.next_cnt\[12\] net89 vssd1 vssd1
+ vccd1 vccd1 genblk1\[1\].osc.clkdiv_C.cnt\[12\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_108_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_845 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11524_ _05450_ genblk1\[8\].osc.clkdiv_C.cnt\[6\] vssd1 vssd1 vccd1 vccd1 _05459_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_80_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11455_ _05424_ vssd1 vssd1 vccd1 vccd1 _00775_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_40_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_123_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10706__A _04880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06903__B _01327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10406_ net626 _04661_ _04663_ net658 _04671_ vssd1 vssd1 vccd1 vccd1 _00479_ sky130_fd_sc_hd__a221o_1
XFILLER_0_0_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11386_ genblk2\[8\].wave_shpr.div.acc\[13\] genblk2\[8\].wave_shpr.div.b1\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05362_ sky130_fd_sc_hd__or2b_1
X_13125_ clknet_leaf_3_clk _00450_ net51 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.b1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10337_ _04636_ vssd1 vssd1 vccd1 vccd1 _00445_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13056_ clknet_leaf_134_clk _00383_ net63 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.quo\[8\]
+ sky130_fd_sc_hd__dfrtp_2
X_10268_ _04578_ _04579_ vssd1 vssd1 vccd1 vccd1 _04580_ sky130_fd_sc_hd__nand2_1
X_12007_ _05808_ vssd1 vssd1 vccd1 vccd1 _00943_ sky130_fd_sc_hd__clkbuf_1
X_10199_ genblk2\[3\].wave_shpr.div.acc\[14\] _04527_ _04507_ vssd1 vssd1 vccd1 vccd1
+ _04528_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12909_ clknet_leaf_31_clk _00240_ net100 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.acc\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_06430_ net718 _01373_ vssd1 vssd1 vccd1 vccd1 genblk1\[1\].osc.clkdiv_C.next_cnt\[0\]
+ sky130_fd_sc_hd__nor2_1
XTAP_2090 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12027__A2 _05813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06366__A _01308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06361_ _01223_ _01226_ vssd1 vssd1 vccd1 vccd1 _01305_ sky130_fd_sc_hd__or2_2
XANTENNA__13206__RESET_B net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_84_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08100_ genblk1\[4\].osc.clkdiv_C.cnt\[12\] _02805_ _02806_ vssd1 vssd1 vccd1 vccd1
+ _02807_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_127_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09080_ _03732_ net577 _03733_ vssd1 vssd1 vccd1 vccd1 _00091_ sky130_fd_sc_hd__o21a_1
X_06292_ _01176_ _01178_ _01194_ vssd1 vssd1 vccd1 vccd1 _01254_ sky130_fd_sc_hd__and3b_2
XFILLER_0_140_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08031_ genblk2\[6\].wave_shpr.div.fin_quo\[4\] _02737_ vssd1 vssd1 vccd1 vccd1 _02738_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_71_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06813__B _01684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold802 genblk2\[11\].wave_shpr.div.acc\[3\] vssd1 vssd1 vccd1 vccd1 net1020 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07197__A genblk1\[9\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold813 genblk2\[6\].wave_shpr.div.acc\[22\] vssd1 vssd1 vccd1 vccd1 net1031 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_24_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold824 genblk2\[9\].wave_shpr.div.b1\[9\] vssd1 vssd1 vccd1 vccd1 net1042 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold835 genblk2\[7\].wave_shpr.div.acc\[25\] vssd1 vssd1 vccd1 vccd1 net1053 sky130_fd_sc_hd__dlygate4sd3_1
Xhold846 genblk2\[3\].wave_shpr.div.acc\[24\] vssd1 vssd1 vccd1 vccd1 net1064 sky130_fd_sc_hd__dlygate4sd3_1
Xhold857 genblk2\[4\].wave_shpr.div.b1\[2\] vssd1 vssd1 vccd1 vccd1 net1075 sky130_fd_sc_hd__dlygate4sd3_1
X_09982_ genblk2\[3\].wave_shpr.div.acc\[2\] genblk2\[3\].wave_shpr.div.b1\[2\] vssd1
+ vssd1 vccd1 vccd1 _04378_ sky130_fd_sc_hd__or2b_1
Xhold868 genblk2\[11\].wave_shpr.div.b1\[16\] vssd1 vssd1 vccd1 vccd1 net1086 sky130_fd_sc_hd__dlygate4sd3_1
Xhold879 genblk2\[5\].wave_shpr.div.b1\[7\] vssd1 vssd1 vccd1 vccd1 net1097 sky130_fd_sc_hd__dlygate4sd3_1
X_08933_ sig_norm.acc\[12\] _01157_ vssd1 vssd1 vccd1 vccd1 _03628_ sky130_fd_sc_hd__and2_1
XFILLER_0_42_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08864_ _03135_ _03225_ _03570_ vssd1 vssd1 vccd1 vccd1 _03571_ sky130_fd_sc_hd__nor3_1
XANTENNA__10351__A _01355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07815_ genblk2\[1\].wave_shpr.div.fin_quo\[2\] _02462_ _02461_ vssd1 vssd1 vccd1
+ vccd1 _02522_ sky130_fd_sc_hd__o21a_1
X_08795_ _03489_ _03496_ vssd1 vssd1 vccd1 vccd1 _03502_ sky130_fd_sc_hd__or2_1
X_07746_ _02447_ _02446_ _02448_ vssd1 vssd1 vccd1 vccd1 _02453_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_95_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_67_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_79_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07677_ _02377_ _02381_ _02368_ _02382_ _02383_ vssd1 vssd1 vccd1 vccd1 _02384_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_66_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09416_ genblk2\[1\].wave_shpr.div.b1\[5\] genblk2\[1\].wave_shpr.div.acc\[5\] vssd1
+ vssd1 vccd1 vccd1 _03980_ sky130_fd_sc_hd__and2b_1
XFILLER_0_137_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_48_842 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06628_ genblk1\[3\].osc.clkdiv_C.cnt\[4\] _01530_ _01524_ vssd1 vssd1 vccd1 vccd1
+ _01532_ sky130_fd_sc_hd__o21ai_1
XANTENNA__10029__A1 genblk2\[3\].wave_shpr.div.quo\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09347_ _03799_ net23 vssd1 vssd1 vccd1 vccd1 _03924_ sky130_fd_sc_hd__or2_1
X_06559_ _01451_ _01472_ vssd1 vssd1 vccd1 vccd1 _01473_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09278_ genblk2\[0\].wave_shpr.div.b1\[2\] genblk2\[0\].wave_shpr.div.acc\[2\] vssd1
+ vssd1 vccd1 vccd1 _03871_ sky130_fd_sc_hd__xor2_1
XFILLER_0_90_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08229_ _02838_ _02935_ _02846_ vssd1 vssd1 vccd1 vccd1 _02936_ sky130_fd_sc_hd__o21a_1
XFILLER_0_62_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11240_ net613 _05255_ _05256_ net640 _05259_ vssd1 vssd1 vccd1 vccd1 _00725_ sky130_fd_sc_hd__a221o_1
XFILLER_0_105_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11171_ genblk2\[7\].wave_shpr.div.fin_quo\[4\] net1318 _00019_ vssd1 vssd1 vccd1
+ vccd1 _05227_ sky130_fd_sc_hd__mux2_1
XANTENNA__12582__RESET_B net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10122_ _04058_ _01486_ vssd1 vssd1 vccd1 vccd1 _04472_ sky130_fd_sc_hd__nor2_1
XANTENNA__08158__B1 _01858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10053_ _04435_ vssd1 vssd1 vccd1 vccd1 _00362_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09370__A2 _03841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09658__B1 _04045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10955_ genblk2\[6\].wave_shpr.div.quo\[11\] _05057_ _05055_ net344 _05061_ vssd1
+ vssd1 vccd1 vccd1 _00638_ sky130_fd_sc_hd__a221o_1
X_13743_ clknet_leaf_51_clk net240 net110 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.quo\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13674_ clknet_leaf_41_clk _00987_ net125 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.acc\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10886_ genblk2\[6\].wave_shpr.div.fin_quo\[3\] net1320 _00017_ vssd1 vssd1 vccd1
+ vccd1 _05027_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12625_ clknet_leaf_16_clk genblk1\[4\].osc.clkdiv_C.next_cnt\[10\] net74 vssd1 vssd1
+ vccd1 vccd1 genblk1\[4\].osc.clkdiv_C.cnt\[10\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__06892__B1 _01666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09497__A _03701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12556_ clknet_leaf_55_clk genblk1\[0\].osc.clkdiv_C.next_cnt\[13\] net175 vssd1
+ vssd1 vccd1 vccd1 genblk1\[0\].osc.clkdiv_C.cnt\[13\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_109_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11507_ _05441_ vssd1 vssd1 vccd1 vccd1 _05448_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_124_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12487_ clknet_leaf_108_clk _00049_ net151 vssd1 vssd1 vccd1 vccd1 sig_norm.acc\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold109 _00377_ vssd1 vssd1 vccd1 vccd1 net327 sky130_fd_sc_hd__dlygate4sd3_1
X_11438_ genblk2\[8\].wave_shpr.div.acc\[24\] _05413_ vssd1 vssd1 vccd1 vccd1 _05414_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_0_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08397__B1 _02425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11369_ _05349_ vssd1 vssd1 vccd1 vccd1 _00764_ sky130_fd_sc_hd__clkbuf_1
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13108_ clknet_leaf_127_clk _00433_ net133 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.fin_quo\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13039_ clknet_leaf_126_clk _00366_ net61 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.b1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09361__A2 _03841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07600_ net17 net18 vssd1 vssd1 vccd1 vccd1 _02307_ sky130_fd_sc_hd__and2_2
X_08580_ genblk2\[10\].wave_shpr.div.fin_quo\[1\] vssd1 vssd1 vccd1 vccd1 _03287_
+ sky130_fd_sc_hd__inv_2
XANTENNA__07911__A3 _01440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07531_ _01155_ vssd1 vssd1 vccd1 vccd1 _02248_ sky130_fd_sc_hd__buf_4
XFILLER_0_44_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06808__B _01359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07462_ _02193_ vssd1 vssd1 vccd1 vccd1 _00018_ sky130_fd_sc_hd__inv_2
X_09201_ net1199 _01183_ _03822_ vssd1 vssd1 vccd1 vccd1 _03829_ sky130_fd_sc_hd__mux2_1
XFILLER_0_57_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11208__B1 _03736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06413_ genblk1\[1\].osc.clkdiv_C.cnt\[9\] _01356_ vssd1 vssd1 vccd1 vccd1 _01357_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07393_ genblk1\[11\].osc.clkdiv_C.cnt\[15\] _02139_ vssd1 vssd1 vccd1 vccd1 _02142_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_91_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_519 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_268 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09132_ _03755_ _03778_ _03779_ vssd1 vssd1 vccd1 vccd1 _03780_ sky130_fd_sc_hd__a21o_1
X_06344_ genblk1\[0\].osc.clkdiv_C.cnt\[13\] _01291_ _01269_ vssd1 vssd1 vccd1 vccd1
+ _01293_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_115_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_115_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09063_ net1276 _03721_ _03722_ vssd1 vssd1 vccd1 vccd1 _03723_ sky130_fd_sc_hd__mux2_1
X_06275_ _01178_ _01176_ _01194_ vssd1 vssd1 vccd1 vccd1 _01237_ sky130_fd_sc_hd__nor3b_1
XANTENNA_fanout213_A net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10982__A2 _05051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08014_ genblk1\[6\].osc.clkdiv_C.cnt\[5\] _01367_ vssd1 vssd1 vccd1 vccd1 _02721_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold610 genblk2\[5\].wave_shpr.div.acc\[17\] vssd1 vssd1 vccd1 vccd1 net828 sky130_fd_sc_hd__dlygate4sd3_1
Xhold621 genblk2\[9\].wave_shpr.div.acc\[8\] vssd1 vssd1 vccd1 vccd1 net839 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold632 genblk2\[4\].wave_shpr.div.acc\[14\] vssd1 vssd1 vccd1 vccd1 net850 sky130_fd_sc_hd__dlygate4sd3_1
Xhold643 genblk2\[0\].wave_shpr.div.b1\[0\] vssd1 vssd1 vccd1 vccd1 net861 sky130_fd_sc_hd__dlygate4sd3_1
Xhold654 genblk2\[8\].wave_shpr.div.acc\[3\] vssd1 vssd1 vccd1 vccd1 net872 sky130_fd_sc_hd__dlygate4sd3_1
Xhold665 genblk2\[6\].wave_shpr.div.acc\[13\] vssd1 vssd1 vccd1 vccd1 net883 sky130_fd_sc_hd__dlygate4sd3_1
Xhold676 genblk2\[7\].wave_shpr.div.acc\[11\] vssd1 vssd1 vccd1 vccd1 net894 sky130_fd_sc_hd__dlygate4sd3_1
Xhold687 genblk2\[1\].wave_shpr.div.acc\[15\] vssd1 vssd1 vccd1 vccd1 net905 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07655__A _02361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold698 genblk2\[7\].wave_shpr.div.acc\[9\] vssd1 vssd1 vccd1 vccd1 net916 sky130_fd_sc_hd__dlygate4sd3_1
X_09965_ genblk2\[3\].wave_shpr.div.acc\[17\] genblk2\[3\].wave_shpr.div.b1\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04361_ sky130_fd_sc_hd__or2b_1
XANTENNA__11486__B1_N _03717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08916_ net1155 _02260_ _03616_ _03574_ vssd1 vssd1 vccd1 vccd1 _00044_ sky130_fd_sc_hd__a22o_1
X_09896_ _04195_ _04162_ vssd1 vssd1 vccd1 vccd1 _04312_ sky130_fd_sc_hd__or2b_1
XTAP_970 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_992 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08847_ _03536_ _03537_ _03531_ vssd1 vssd1 vccd1 vccd1 _03554_ sky130_fd_sc_hd__a21boi_1
XTAP_2804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08778_ _03333_ _03483_ _03465_ _03482_ vssd1 vssd1 vccd1 vccd1 _03485_ sky130_fd_sc_hd__a211oi_2
XTAP_2815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07729_ _01360_ net37 genblk1\[1\].osc.clkdiv_C.cnt\[6\] vssd1 vssd1 vccd1 vccd1
+ _02436_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10740_ _04820_ vssd1 vssd1 vccd1 vccd1 _04907_ sky130_fd_sc_hd__buf_4
XFILLER_0_138_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10671_ _04854_ vssd1 vssd1 vccd1 vccd1 _04862_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_82_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12410_ _05971_ _05927_ vssd1 vssd1 vccd1 vccd1 _06080_ sky130_fd_sc_hd__or2b_1
XANTENNA__08933__B _01157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13390_ clknet_leaf_79_clk _00709_ net205 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.b1\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09812__B1 _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12341_ net412 _03942_ _03941_ net434 _06028_ vssd1 vssd1 vccd1 vccd1 _01057_ sky130_fd_sc_hd__a221o_1
XFILLER_0_106_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_121_714 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12272_ _01305_ vssd1 vssd1 vccd1 vccd1 _05997_ sky130_fd_sc_hd__inv_2
X_11223_ net317 _05246_ _05250_ net754 vssd1 vssd1 vccd1 vccd1 _00717_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11154_ _05165_ _05212_ _05213_ vssd1 vssd1 vccd1 vccd1 _05214_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_101_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10105_ _04269_ genblk1\[3\].osc.clkdiv_C.cnt\[3\] vssd1 vssd1 vccd1 vccd1 _04463_
+ sky130_fd_sc_hd__and2_1
X_11085_ net1076 _05057_ _05055_ _05151_ vssd1 vssd1 vccd1 vccd1 _00678_ sky130_fd_sc_hd__a22o_1
X_10036_ _04427_ vssd1 vssd1 vccd1 vccd1 _00353_ sky130_fd_sc_hd__clkbuf_1
X_11987_ _05798_ vssd1 vssd1 vccd1 vccd1 _00933_ sky130_fd_sc_hd__clkbuf_1
X_13726_ clknet_leaf_97_clk _01037_ net166 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.quo\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10938_ net792 _05052_ _05023_ _05055_ vssd1 vssd1 vccd1 vccd1 _00627_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_129_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13657_ clknet_leaf_48_clk _00970_ net120 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.quo\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10869_ _04968_ _05011_ _05012_ vssd1 vssd1 vccd1 vccd1 _05013_ sky130_fd_sc_hd__a21o_1
XFILLER_0_85_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12608_ clknet_leaf_23_clk genblk1\[3\].osc.clkdiv_C.next_cnt\[11\] net94 vssd1 vssd1
+ vccd1 vccd1 genblk1\[3\].osc.clkdiv_C.cnt\[11\] sky130_fd_sc_hd__dfrtp_1
XPHY_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09803__B1 _04252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13588_ clknet_leaf_72_clk _00903_ net215 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.acc\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09020__A _02152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12539_ clknet_leaf_62_clk _00091_ net189 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.b1\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12166__A1 _05816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07475__A _02155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09750_ net1198 vssd1 vssd1 vccd1 vccd1 _00272_ sky130_fd_sc_hd__clkbuf_1
X_06962_ genblk1\[7\].osc.clkdiv_C.cnt\[9\] _01797_ vssd1 vssd1 vccd1 vccd1 _01798_
+ sky130_fd_sc_hd__xnor2_1
X_08701_ _03359_ _03381_ _03406_ _03407_ vssd1 vssd1 vccd1 vccd1 _03408_ sky130_fd_sc_hd__o211ai_2
X_09681_ genblk2\[2\].wave_shpr.div.acc\[12\] genblk2\[2\].wave_shpr.div.b1\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04161_ sky130_fd_sc_hd__or2b_1
XFILLER_0_146_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06893_ _01308_ _01577_ vssd1 vssd1 vccd1 vccd1 _01747_ sky130_fd_sc_hd__nand2_2
XANTENNA__08542__B1 _02308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08632_ _02217_ _02553_ genblk2\[6\].wave_shpr.div.fin_quo\[3\] vssd1 vssd1 vccd1
+ vccd1 _03339_ sky130_fd_sc_hd__and3_1
XFILLER_0_146_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08563_ genblk2\[7\].wave_shpr.div.fin_quo\[1\] _03269_ vssd1 vssd1 vccd1 vccd1 _03270_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout163_A net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07514_ PWM.counter\[2\] vssd1 vssd1 vccd1 vccd1 _02234_ sky130_fd_sc_hd__inv_2
X_08494_ _03051_ _03174_ _03154_ _03173_ vssd1 vssd1 vccd1 vccd1 _03201_ sky130_fd_sc_hd__o211a_1
XFILLER_0_76_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07445_ genblk2\[5\].wave_shpr.div.busy _02180_ vssd1 vssd1 vccd1 vccd1 _02181_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout48 net50 vssd1 vssd1 vccd1 vccd1 net48 sky130_fd_sc_hd__clkbuf_4
Xfanout59 net63 vssd1 vssd1 vccd1 vccd1 net59 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_57_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07376_ _02128_ _02127_ vssd1 vssd1 vccd1 vccd1 _02129_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_18_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09115_ genblk2\[0\].wave_shpr.div.acc\[1\] genblk2\[0\].wave_shpr.div.b1\[1\] vssd1
+ vssd1 vccd1 vccd1 _03763_ sky130_fd_sc_hd__or2b_1
X_06327_ _01269_ _01281_ _01282_ vssd1 vssd1 vccd1 vccd1 genblk1\[0\].osc.clkdiv_C.next_cnt\[6\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_17_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06273__B _01234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10955__A2 _05057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09046_ _03711_ vssd1 vssd1 vccd1 vccd1 _00079_ sky130_fd_sc_hd__clkbuf_1
X_06258_ freq_div.state\[1\] _01176_ vssd1 vssd1 vccd1 vccd1 _01220_ sky130_fd_sc_hd__xor2_4
XFILLER_0_103_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold440 genblk2\[4\].wave_shpr.div.quo\[19\] vssd1 vssd1 vccd1 vccd1 net658 sky130_fd_sc_hd__dlygate4sd3_1
X_06189_ net361 vssd1 vssd1 vccd1 vccd1 PWM.next_counter\[0\] sky130_fd_sc_hd__inv_2
XFILLER_0_102_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold451 genblk2\[9\].wave_shpr.div.acc\[18\] vssd1 vssd1 vccd1 vccd1 net669 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09076__S _03722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10707__A2 _04821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold462 genblk2\[4\].wave_shpr.div.quo\[16\] vssd1 vssd1 vccd1 vccd1 net680 sky130_fd_sc_hd__dlygate4sd3_1
Xhold473 genblk1\[8\].osc.clkdiv_C.cnt\[17\] vssd1 vssd1 vccd1 vccd1 net691 sky130_fd_sc_hd__dlygate4sd3_1
Xhold484 genblk2\[0\].wave_shpr.div.b1\[17\] vssd1 vssd1 vccd1 vccd1 net702 sky130_fd_sc_hd__dlygate4sd3_1
Xhold495 genblk2\[9\].wave_shpr.div.b1\[16\] vssd1 vssd1 vccd1 vccd1 net713 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_96_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07584__A1 genblk1\[9\].osc.clkdiv_C.cnt\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06387__A2 _01323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07584__B2 genblk1\[9\].osc.clkdiv_C.cnt\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09948_ genblk2\[2\].wave_shpr.div.acc\[25\] _04212_ genblk2\[2\].wave_shpr.div.acc\[24\]
+ genblk2\[2\].wave_shpr.div.acc\[26\] vssd1 vssd1 vccd1 vccd1 _04350_ sky130_fd_sc_hd__or4b_1
XANTENNA_fanout76_A net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09879_ _04187_ _04166_ vssd1 vssd1 vccd1 vccd1 _04299_ sky130_fd_sc_hd__or2b_1
X_11910_ _03832_ genblk2\[10\].wave_shpr.div.acc\[16\] vssd1 vssd1 vccd1 vccd1 _05732_
+ sky130_fd_sc_hd__nor2_1
XTAP_2601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10340__B1 _04432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12890_ clknet_leaf_28_clk _00221_ net91 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.quo\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11841_ genblk2\[9\].wave_shpr.div.acc\[11\] _05682_ _05673_ vssd1 vssd1 vccd1 vccd1
+ _05683_ sky130_fd_sc_hd__mux2_1
XTAP_2645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11772_ genblk2\[9\].wave_shpr.div.quo\[16\] _05628_ _05629_ net304 _05635_ vssd1
+ vssd1 vccd1 vccd1 _00881_ sky130_fd_sc_hd__a221o_1
XTAP_2689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10723_ _04778_ _04788_ vssd1 vssd1 vccd1 vccd1 _04894_ sky130_fd_sc_hd__xor2_1
XFILLER_0_55_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13511_ clknet_leaf_78_clk _00828_ net205 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.acc\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_95_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10654_ net1342 _04853_ _04821_ _04855_ vssd1 vssd1 vccd1 vccd1 _00543_ sky130_fd_sc_hd__a22o_1
X_13442_ clknet_leaf_92_clk _00761_ net149 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.acc\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13373_ clknet_leaf_117_clk _00692_ net140 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.fin_quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_51_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10585_ _04764_ _04811_ _04812_ vssd1 vssd1 vccd1 vccd1 _04813_ sky130_fd_sc_hd__o21bai_1
XANTENNA__10946__A2 _05052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12324_ _03689_ genblk1\[11\].osc.clkdiv_C.cnt\[7\] vssd1 vssd1 vccd1 vccd1 _06020_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_32_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12255_ genblk2\[11\].wave_shpr.div.fin_quo\[5\] net767 _00005_ vssd1 vssd1 vccd1
+ vccd1 _05988_ sky130_fd_sc_hd__mux2_1
X_11206_ _03831_ net391 _03717_ vssd1 vssd1 vccd1 vccd1 _00708_ sky130_fd_sc_hd__a21bo_1
X_12186_ net289 _05923_ _05924_ vssd1 vssd1 vccd1 vccd1 _01006_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07575__A1 genblk1\[9\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold4_A modein.delay_in\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11137_ genblk2\[7\].wave_shpr.div.b1\[8\] genblk2\[7\].wave_shpr.div.acc\[8\] vssd1
+ vssd1 vccd1 vccd1 _05197_ sky130_fd_sc_hd__and2b_1
X_11068_ _05139_ _05140_ vssd1 vssd1 vccd1 vccd1 _05141_ sky130_fd_sc_hd__nand2_1
XANTENNA__08838__B _03544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10019_ genblk2\[3\].wave_shpr.div.acc\[18\] _04414_ vssd1 vssd1 vccd1 vccd1 _04415_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_149_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10882__A1 genblk2\[6\].wave_shpr.div.quo\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13709_ clknet_leaf_31_clk _01020_ net103 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.b1\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_129_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07230_ genblk1\[10\].osc.clkdiv_C.cnt\[6\] _01432_ vssd1 vssd1 vccd1 vccd1 _02012_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_143_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12614__RESET_B net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06805__C _01226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07161_ genblk1\[9\].osc.clkdiv_C.cnt\[1\] genblk1\[9\].osc.clkdiv_C.cnt\[0\] genblk1\[9\].osc.clkdiv_C.cnt\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01959_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_42_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08055__A2 _01180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_850 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06112_ smpl_rt_clkdiv.clkDiv_inst.cnt\[1\] net338 net359 vssd1 vssd1 vccd1 vccd1
+ _01090_ sky130_fd_sc_hd__a21oi_1
X_07092_ _01887_ _01900_ _01901_ vssd1 vssd1 vccd1 vccd1 genblk1\[8\].osc.clkdiv_C.next_cnt\[8\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_10_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09555__A2 _04042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout205 net209 vssd1 vssd1 vccd1 vccd1 net205 sky130_fd_sc_hd__clkbuf_4
Xfanout216 net217 vssd1 vssd1 vccd1 vccd1 net216 sky130_fd_sc_hd__clkbuf_4
X_09802_ net336 _04248_ _04252_ net719 vssd1 vssd1 vccd1 vccd1 _00294_ sky130_fd_sc_hd__a22o_1
X_07994_ genblk1\[6\].osc.clkdiv_C.cnt\[8\] _01732_ _01742_ genblk1\[6\].osc.clkdiv_C.cnt\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02701_ sky130_fd_sc_hd__o22a_1
XANTENNA__07933__A genblk2\[8\].wave_shpr.div.fin_quo\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_09733_ genblk2\[2\].wave_shpr.div.acc\[25\] genblk2\[2\].wave_shpr.div.acc\[24\]
+ genblk2\[2\].wave_shpr.div.acc\[26\] _04212_ vssd1 vssd1 vccd1 vccd1 _04213_ sky130_fd_sc_hd__or4_2
X_06945_ genblk1\[6\].osc.clkdiv_C.cnt\[14\] _01783_ vssd1 vssd1 vccd1 vccd1 _01785_
+ sky130_fd_sc_hd__and2_1
X_06876_ _01336_ net37 vssd1 vssd1 vccd1 vccd1 _01730_ sky130_fd_sc_hd__or2_1
X_09664_ genblk2\[1\].wave_shpr.div.i\[1\] genblk2\[1\].wave_shpr.div.i\[0\] vssd1
+ vssd1 vccd1 vccd1 _04148_ sky130_fd_sc_hd__or2_1
X_08615_ genblk2\[4\].wave_shpr.div.fin_quo\[0\] genblk2\[4\].wave_shpr.div.fin_quo\[1\]
+ _02932_ _02223_ vssd1 vssd1 vccd1 vccd1 _03322_ sky130_fd_sc_hd__a31o_1
X_09595_ _03985_ _04097_ vssd1 vssd1 vccd1 vccd1 _04098_ sky130_fd_sc_hd__xnor2_1
XTAP_1207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08546_ _03251_ _03252_ vssd1 vssd1 vccd1 vccd1 _03253_ sky130_fd_sc_hd__and2b_1
X_08477_ genblk2\[4\].wave_shpr.div.fin_quo\[3\] _02932_ _02840_ _02222_ vssd1 vssd1
+ vccd1 vccd1 _03184_ sky130_fd_sc_hd__a31o_1
XFILLER_0_77_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07428_ genblk2\[3\].wave_shpr.div.busy _02167_ vssd1 vssd1 vccd1 vccd1 _02168_ sky130_fd_sc_hd__and2_1
XFILLER_0_134_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07359_ genblk1\[11\].osc.clkdiv_C.cnt\[7\] _02112_ vssd1 vssd1 vccd1 vccd1 _02116_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_134_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10389__B1 _04655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10370_ net418 _04652_ _04623_ _04655_ vssd1 vssd1 vccd1 vccd1 _00459_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09029_ _03694_ _03697_ _03699_ _03696_ net789 vssd1 vssd1 vccd1 vccd1 _00074_ sky130_fd_sc_hd__a32o_1
XFILLER_0_131_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12040_ _05819_ genblk1\[10\].osc.clkdiv_C.cnt\[3\] vssd1 vssd1 vccd1 vccd1 _05824_
+ sky130_fd_sc_hd__and2_1
Xhold270 _00734_ vssd1 vssd1 vccd1 vccd1 net488 sky130_fd_sc_hd__dlygate4sd3_1
Xhold281 _00641_ vssd1 vssd1 vccd1 vccd1 net499 sky130_fd_sc_hd__dlygate4sd3_1
Xhold292 genblk2\[11\].wave_shpr.div.quo\[17\] vssd1 vssd1 vccd1 vccd1 net510 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12942_ clknet_leaf_111_clk _00271_ net130 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.fin_quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06459__A genblk1\[1\].osc.clkdiv_C.cnt\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12873_ clknet_leaf_138_clk _00204_ net39 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.b1\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11824_ genblk2\[9\].wave_shpr.div.acc\[7\] _05669_ _05613_ vssd1 vssd1 vccd1 vccd1
+ _05670_ sky130_fd_sc_hd__mux2_1
XTAP_2464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09482__A1 _01183_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11755_ net290 _03696_ _03694_ net526 _05625_ vssd1 vssd1 vccd1 vccd1 _00874_ sky130_fd_sc_hd__a221o_1
XFILLER_0_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10092__A2 _04452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10706_ _04880_ _04781_ genblk2\[5\].wave_shpr.div.b1\[0\] vssd1 vssd1 vccd1 vccd1
+ _04881_ sky130_fd_sc_hd__or3b_1
X_11686_ _05571_ _05576_ _05577_ vssd1 vssd1 vccd1 vccd1 _05578_ sky130_fd_sc_hd__a21o_1
XFILLER_0_125_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13425_ clknet_leaf_87_clk _00744_ net201 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.acc\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10637_ net1233 _04223_ _04834_ vssd1 vssd1 vccd1 vccd1 _04846_ sky130_fd_sc_hd__mux2_1
XFILLER_0_125_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10568_ genblk2\[5\].wave_shpr.div.b1\[8\] genblk2\[5\].wave_shpr.div.acc\[8\] vssd1
+ vssd1 vccd1 vccd1 _04796_ sky130_fd_sc_hd__and2b_1
X_13356_ clknet_leaf_4_clk _00677_ net45 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.acc\[24\]
+ sky130_fd_sc_hd__dfrtp_2
X_12307_ net355 _06009_ _06010_ net358 vssd1 vssd1 vccd1 vccd1 _01041_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10499_ net591 _04715_ _04722_ _04739_ vssd1 vssd1 vccd1 vccd1 _00504_ sky130_fd_sc_hd__a22o_1
X_13287_ clknet_leaf_118_clk _00608_ net138 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.fin_quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_12238_ _05925_ _05974_ _05975_ vssd1 vssd1 vccd1 vccd1 _05976_ sky130_fd_sc_hd__a21o_1
X_12169_ net1226 _05818_ _05816_ _05913_ vssd1 vssd1 vccd1 vccd1 _01000_ sky130_fd_sc_hd__a22o_1
XANTENNA__07753__A _02458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput5 pb[13] vssd1 vssd1 vccd1 vccd1 net5 sky130_fd_sc_hd__clkbuf_1
X_06730_ _01615_ vssd1 vssd1 vccd1 vccd1 genblk1\[4\].osc.clkdiv_C.next_cnt\[4\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_127_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06369__A _01192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06661_ genblk1\[3\].osc.clkdiv_C.cnt\[16\] _01551_ vssd1 vssd1 vccd1 vccd1 _01553_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_148_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08400_ genblk1\[2\].osc.clkdiv_C.cnt\[13\] _02425_ _01591_ genblk1\[2\].osc.clkdiv_C.cnt\[12\]
+ vssd1 vssd1 vccd1 vccd1 _03107_ sky130_fd_sc_hd__o22a_1
XANTENNA__07720__B2 genblk1\[1\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09380_ _03944_ _03945_ _03946_ _03947_ net1124 vssd1 vssd1 vccd1 vccd1 _00177_ sky130_fd_sc_hd__a32o_1
X_06592_ _01233_ _01437_ vssd1 vssd1 vccd1 vccd1 _01500_ sky130_fd_sc_hd__nor2_2
X_08331_ _03036_ _02682_ _03035_ _02526_ vssd1 vssd1 vccd1 vccd1 _03038_ sky130_fd_sc_hd__o31a_1
XANTENNA__09473__A1 _04023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06816__B _01355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08262_ _02945_ _02967_ _02968_ vssd1 vssd1 vccd1 vccd1 _02969_ sky130_fd_sc_hd__a21o_1
XFILLER_0_117_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_27_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07213_ genblk1\[10\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 _01995_ sky130_fd_sc_hd__inv_2
X_08193_ _02423_ _02601_ vssd1 vssd1 vccd1 vccd1 _02900_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09225__A1 net269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout126_A net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07144_ _01933_ _01941_ _01942_ _01943_ vssd1 vssd1 vccd1 vccd1 _01944_ sky130_fd_sc_hd__and4b_1
XANTENNA__07236__B1 _02002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_155 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07075_ _01879_ _01889_ vssd1 vssd1 vccd1 vccd1 _01891_ sky130_fd_sc_hd__and2_1
XFILLER_0_112_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10354__A _01490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08200__A2 _02403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07977_ genblk2\[7\].wave_shpr.div.fin_quo\[3\] vssd1 vssd1 vccd1 vccd1 _02684_ sky130_fd_sc_hd__inv_2
X_09716_ _04162_ _04194_ _04195_ vssd1 vssd1 vccd1 vccd1 _04196_ sky130_fd_sc_hd__a21o_1
X_06928_ genblk1\[6\].osc.clkdiv_C.cnt\[7\] _01770_ genblk1\[6\].osc.clkdiv_C.cnt\[8\]
+ vssd1 vssd1 vccd1 vccd1 _01774_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_93_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09647_ net1109 _04109_ _04113_ _04137_ vssd1 vssd1 vccd1 vccd1 _00254_ sky130_fd_sc_hd__a22o_1
XFILLER_0_96_114 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06859_ _01693_ _01717_ vssd1 vssd1 vccd1 vccd1 _01718_ sky130_fd_sc_hd__nor2_1
XTAP_1004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09578_ _04084_ _03977_ vssd1 vssd1 vccd1 vccd1 _04085_ sky130_fd_sc_hd__xnor2_1
XTAP_1037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_fanout39_A net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08529_ genblk2\[11\].wave_shpr.div.fin_quo\[0\] _02524_ _02307_ genblk2\[11\].wave_shpr.div.fin_quo\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03236_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09464__A1 net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08267__A2 net33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11540_ net229 _05441_ _05458_ net575 _05467_ vssd1 vssd1 vccd1 vccd1 _00817_ sky130_fd_sc_hd__a221o_1
XFILLER_0_107_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11471_ _05432_ vssd1 vssd1 vccd1 vccd1 _00783_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10422_ genblk2\[4\].wave_shpr.div.b1\[0\] _04623_ genblk2\[4\].wave_shpr.div.acc\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04681_ sky130_fd_sc_hd__a21oi_1
X_13210_ clknet_leaf_25_clk _00533_ net86 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.b1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07778__A1 _01181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13141_ clknet_leaf_115_clk _00466_ net135 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10353_ _04644_ vssd1 vssd1 vccd1 vccd1 _00453_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_131_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_hold874_A genblk1\[8\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_103_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13072_ clknet_leaf_23_clk net491 net94 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.quo\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10284_ genblk2\[4\].wave_shpr.div.b1\[7\] genblk2\[4\].wave_shpr.div.acc\[7\] vssd1
+ vssd1 vccd1 vccd1 _04596_ sky130_fd_sc_hd__and2b_1
X_12023_ net220 _05813_ _05817_ net740 vssd1 vssd1 vccd1 vccd1 _00950_ sky130_fd_sc_hd__a22o_1
XANTENNA__07950__A1 _01556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10203__S _04507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12925_ clknet_leaf_35_clk _00256_ net106 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.acc\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06505__A2 _01430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12856_ clknet_leaf_91_clk _00187_ net146 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.fin_quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11807_ _05579_ _05570_ vssd1 vssd1 vccd1 vccd1 _05657_ sky130_fd_sc_hd__or2b_1
XTAP_2294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12787_ clknet_leaf_43_clk _00120_ net124 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.b1\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11738_ _02248_ _01150_ vssd1 vssd1 vccd1 vccd1 _05622_ sky130_fd_sc_hd__nand2_1
XFILLER_0_113_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_83_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09207__A1 _03831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11669_ genblk2\[9\].wave_shpr.div.acc\[10\] genblk2\[9\].wave_shpr.div.b1\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05561_ sky130_fd_sc_hd__or2b_1
XFILLER_0_114_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13408_ clknet_leaf_90_clk _00727_ net142 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.quo\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07218__B1 _01442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_784 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_626 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13339_ clknet_leaf_7_clk _00660_ net49 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.acc\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07900_ genblk1\[8\].osc.clkdiv_C.cnt\[14\] _01172_ _02605_ _02606_ vssd1 vssd1 vccd1
+ vccd1 _02607_ sky130_fd_sc_hd__a211o_1
X_08880_ _03575_ sig_norm.acc\[3\] _03585_ vssd1 vssd1 vccd1 vccd1 _03586_ sky130_fd_sc_hd__a21o_1
XANTENNA__10525__B1 _04657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09174__S _03722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07831_ genblk2\[1\].wave_shpr.div.fin_quo\[4\] _02461_ _02463_ _02224_ vssd1 vssd1
+ vccd1 vccd1 _02538_ sky130_fd_sc_hd__a31o_1
X_07762_ _02458_ _02459_ _02220_ vssd1 vssd1 vccd1 vccd1 _02469_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_79_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09501_ _03831_ net1025 _03717_ vssd1 vssd1 vccd1 vccd1 _00205_ sky130_fd_sc_hd__a21bo_1
X_06713_ genblk1\[4\].osc.clkdiv_C.cnt\[1\] genblk1\[4\].osc.clkdiv_C.cnt\[0\] vssd1
+ vssd1 vccd1 vccd1 _01602_ sky130_fd_sc_hd__or2_1
X_07693_ _02399_ _02394_ _02385_ _02396_ vssd1 vssd1 vccd1 vccd1 _02400_ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09432_ genblk2\[1\].wave_shpr.div.b1\[13\] genblk2\[1\].wave_shpr.div.acc\[13\]
+ vssd1 vssd1 vccd1 vccd1 _03996_ sky130_fd_sc_hd__and2b_1
X_06644_ genblk1\[3\].osc.clkdiv_C.cnt\[10\] _01540_ vssd1 vssd1 vccd1 vccd1 _01542_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_547 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_87_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09363_ genblk2\[0\].wave_shpr.div.acc\[23\] _03801_ _03934_ vssd1 vssd1 vccd1 vccd1
+ _03935_ sky130_fd_sc_hd__a21o_1
X_06575_ _01196_ _01327_ vssd1 vssd1 vccd1 vccd1 _01483_ sky130_fd_sc_hd__or2_4
XFILLER_0_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08249__A2 _02309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08314_ _02216_ _02552_ genblk2\[10\].wave_shpr.div.fin_quo\[4\] vssd1 vssd1 vccd1
+ vccd1 _03021_ sky130_fd_sc_hd__and3_1
X_09294_ net866 _03870_ _03877_ _03883_ vssd1 vssd1 vccd1 vccd1 _00155_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10068__B _01226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08245_ _02641_ vssd1 vssd1 vccd1 vccd1 _02952_ sky130_fd_sc_hd__inv_2
XFILLER_0_6_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08176_ _02880_ _02882_ _02870_ vssd1 vssd1 vccd1 vccd1 _02883_ sky130_fd_sc_hd__a21o_1
X_07127_ genblk1\[9\].osc.clkdiv_C.cnt\[2\] _01920_ _01923_ genblk1\[9\].osc.clkdiv_C.cnt\[11\]
+ _01926_ vssd1 vssd1 vccd1 vccd1 _01927_ sky130_fd_sc_hd__a221oi_1
XANTENNA_clkbuf_leaf_63_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06281__B _01242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07058_ genblk1\[8\].osc.clkdiv_C.cnt\[0\] _01211_ _01246_ genblk1\[8\].osc.clkdiv_C.cnt\[14\]
+ _01875_ vssd1 vssd1 vccd1 vccd1 _01876_ sky130_fd_sc_hd__a221o_1
XFILLER_0_101_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_78_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_121_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap23 net1352 vssd1 vssd1 vccd1 vccd1 net23 sky130_fd_sc_hd__buf_1
X_10971_ net486 _05062_ _05064_ net582 _05070_ vssd1 vssd1 vccd1 vccd1 _00645_ sky130_fd_sc_hd__a221o_1
XFILLER_0_97_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xmax_cap34 _01794_ vssd1 vssd1 vccd1 vccd1 net34 sky130_fd_sc_hd__buf_4
X_12710_ clknet_leaf_56_clk genblk1\[9\].osc.clkdiv_C.next_cnt\[5\] net181 vssd1 vssd1
+ vccd1 vccd1 genblk1\[9\].osc.clkdiv_C.cnt\[5\] sky130_fd_sc_hd__dfrtp_4
X_13690_ clknet_leaf_97_clk _00005_ net166 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.done
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_136_clk_A clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12641_ clknet_leaf_10_clk genblk1\[5\].osc.clkdiv_C.next_cnt\[8\] net56 vssd1 vssd1
+ vccd1 vccd1 genblk1\[5\].osc.clkdiv_C.cnt\[8\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_109_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06456__B genblk1\[1\].osc.clkdiv_C.cnt\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_16_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12572_ clknet_leaf_28_clk genblk1\[1\].osc.clkdiv_C.next_cnt\[11\] net89 vssd1 vssd1
+ vccd1 vccd1 genblk1\[1\].osc.clkdiv_C.cnt\[11\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__12441__B1 _03944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07999__A1 _01200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11795__A2 _05613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11523_ _05444_ vssd1 vssd1 vccd1 vccd1 _05458_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_81_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11454_ genblk2\[8\].wave_shpr.div.fin_quo\[6\] net1325 _00021_ vssd1 vssd1 vccd1
+ vccd1 _05424_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10405_ _04477_ genblk1\[4\].osc.clkdiv_C.cnt\[11\] vssd1 vssd1 vccd1 vccd1 _04671_
+ sky130_fd_sc_hd__and2_1
X_11385_ genblk2\[8\].wave_shpr.div.acc\[14\] genblk2\[8\].wave_shpr.div.b1\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05361_ sky130_fd_sc_hd__or2b_1
XFILLER_0_104_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13124_ clknet_leaf_3_clk _00449_ net51 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.b1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10336_ net1287 _01256_ _04440_ vssd1 vssd1 vccd1 vccd1 _04636_ sky130_fd_sc_hd__mux2_1
XANTENNA__07620__B1 _01595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_9_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_9_0_clk sky130_fd_sc_hd__clkbuf_8
X_10267_ genblk2\[4\].wave_shpr.div.acc\[4\] genblk2\[4\].wave_shpr.div.b1\[4\] vssd1
+ vssd1 vccd1 vccd1 _04579_ sky130_fd_sc_hd__or2b_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13055_ clknet_leaf_113_clk _00382_ net128 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_12006_ genblk2\[11\].wave_shpr.div.b1\[12\] _01494_ _05802_ vssd1 vssd1 vccd1 vccd1
+ _05808_ sky130_fd_sc_hd__mux2_1
XANTENNA__11537__B genblk1\[8\].osc.clkdiv_C.cnt\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10198_ _04406_ _04526_ vssd1 vssd1 vccd1 vccd1 _04527_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12908_ clknet_leaf_36_clk _00239_ net103 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.acc\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_48_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_69_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07151__A2 net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12839_ clknet_leaf_65_clk _00172_ net197 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.acc\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_57_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2080 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2091 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_146_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_29_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06366__B _01309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06360_ _01303_ vssd1 vssd1 vccd1 vccd1 _01304_ sky130_fd_sc_hd__clkbuf_4
XTAP_1390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_90_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11786__A2 _02203_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06291_ genblk1\[0\].osc.clkdiv_C.cnt\[13\] _01240_ _01243_ _01244_ _01252_ vssd1
+ vssd1 vccd1 vccd1 _01253_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08030_ genblk2\[6\].wave_shpr.div.fin_quo\[3\] _02736_ vssd1 vssd1 vccd1 vccd1 _02737_
+ sky130_fd_sc_hd__or2_1
XANTENNA__07478__A _02204_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06382__A _01229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold803 genblk2\[3\].wave_shpr.div.acc\[25\] vssd1 vssd1 vccd1 vccd1 net1021 sky130_fd_sc_hd__dlygate4sd3_1
Xhold814 genblk2\[0\].wave_shpr.div.acc\[21\] vssd1 vssd1 vccd1 vccd1 net1032 sky130_fd_sc_hd__dlygate4sd3_1
Xhold825 genblk2\[6\].wave_shpr.div.acc\[26\] vssd1 vssd1 vccd1 vccd1 net1043 sky130_fd_sc_hd__dlygate4sd3_1
Xhold836 genblk2\[2\].wave_shpr.div.quo\[0\] vssd1 vssd1 vccd1 vccd1 net1054 sky130_fd_sc_hd__buf_1
XFILLER_0_101_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold847 sig_norm.acc\[3\] vssd1 vssd1 vccd1 vccd1 net1065 sky130_fd_sc_hd__dlygate4sd3_1
Xhold858 genblk2\[6\].wave_shpr.div.acc\[25\] vssd1 vssd1 vccd1 vccd1 net1076 sky130_fd_sc_hd__dlygate4sd3_1
Xhold869 genblk2\[10\].wave_shpr.div.acc\[21\] vssd1 vssd1 vccd1 vccd1 net1087 sky130_fd_sc_hd__dlygate4sd3_1
X_09981_ genblk2\[3\].wave_shpr.div.acc\[3\] genblk2\[3\].wave_shpr.div.b1\[3\] vssd1
+ vssd1 vccd1 vccd1 _04377_ sky130_fd_sc_hd__or2b_1
XFILLER_0_40_787 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08932_ _03625_ _03591_ sig_norm.acc\[11\] vssd1 vssd1 vccd1 vccd1 _03627_ sky130_fd_sc_hd__mux2_1
X_08863_ _03525_ _03568_ _03569_ vssd1 vssd1 vccd1 vccd1 _03570_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07914__A1 genblk1\[8\].osc.clkdiv_C.cnt\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07914__B2 _01489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07814_ _02308_ vssd1 vssd1 vccd1 vccd1 _02521_ sky130_fd_sc_hd__buf_4
XFILLER_0_98_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08794_ _03491_ _03495_ vssd1 vssd1 vccd1 vccd1 _03501_ sky130_fd_sc_hd__nand2_1
XFILLER_0_74_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07745_ genblk1\[1\].osc.clkdiv_C.cnt\[12\] _01344_ _01337_ genblk1\[1\].osc.clkdiv_C.cnt\[11\]
+ _02451_ vssd1 vssd1 vccd1 vccd1 _02452_ sky130_fd_sc_hd__a221oi_2
XFILLER_0_79_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07678__B1 _01991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07676_ genblk1\[10\].osc.clkdiv_C.cnt\[7\] _01190_ _01992_ genblk1\[10\].osc.clkdiv_C.cnt\[4\]
+ _02371_ vssd1 vssd1 vccd1 vccd1 _02383_ sky130_fd_sc_hd__a221o_1
X_09415_ _03967_ _03977_ _03978_ vssd1 vssd1 vccd1 vccd1 _03979_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_149_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06627_ _01523_ _01530_ _01531_ vssd1 vssd1 vccd1 vccd1 genblk1\[3\].osc.clkdiv_C.next_cnt\[3\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_137_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10079__A _03833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_71 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09346_ genblk2\[0\].wave_shpr.div.acc\[25\] genblk2\[0\].wave_shpr.div.acc\[24\]
+ genblk2\[0\].wave_shpr.div.acc\[26\] _03802_ vssd1 vssd1 vccd1 vccd1 _03923_ sky130_fd_sc_hd__nor4_1
XFILLER_0_47_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06558_ genblk1\[2\].osc.clkdiv_C.cnt\[12\] genblk1\[2\].osc.clkdiv_C.cnt\[11\] _01468_
+ vssd1 vssd1 vccd1 vccd1 _01472_ sky130_fd_sc_hd__and3_1
XFILLER_0_118_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09277_ _03835_ vssd1 vssd1 vccd1 vccd1 _03870_ sky130_fd_sc_hd__clkbuf_4
X_06489_ genblk1\[2\].osc.clkdiv_C.cnt\[15\] _01414_ _01210_ vssd1 vssd1 vccd1 vccd1
+ _01415_ sky130_fd_sc_hd__mux2_1
XFILLER_0_118_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08228_ _02933_ _02934_ genblk2\[4\].wave_shpr.div.fin_quo\[6\] _02362_ vssd1 vssd1
+ vccd1 vccd1 _02935_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__07850__B1 _02316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08159_ _01489_ genblk1\[3\].osc.clkdiv_C.cnt\[12\] vssd1 vssd1 vccd1 vccd1 _02866_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11170_ _05226_ vssd1 vssd1 vccd1 vccd1 _00688_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__06956__A2 _01311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10121_ net296 _04461_ _04462_ net451 _04471_ vssd1 vssd1 vccd1 vccd1 _00394_ sky130_fd_sc_hd__a221o_1
X_10052_ genblk2\[4\].wave_shpr.div.b1\[5\] _01870_ _04238_ vssd1 vssd1 vccd1 vccd1
+ _04435_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13742_ clknet_leaf_46_clk _01053_ net121 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.quo\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10954_ _04676_ _01729_ vssd1 vssd1 vccd1 vccd1 _05061_ sky130_fd_sc_hd__nor2_1
XFILLER_0_97_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06467__A genblk1\[1\].osc.clkdiv_C.cnt\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07133__A2 _01513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13673_ clknet_leaf_40_clk _00986_ net117 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.acc\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13757__RESET_B net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10885_ _05026_ vssd1 vssd1 vccd1 vccd1 _00603_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_39_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12624_ clknet_leaf_19_clk genblk1\[4\].osc.clkdiv_C.next_cnt\[9\] net109 vssd1 vssd1
+ vccd1 vccd1 genblk1\[4\].osc.clkdiv_C.cnt\[9\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_54_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08094__B1 _01498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12555_ clknet_leaf_55_clk genblk1\[0\].osc.clkdiv_C.next_cnt\[12\] net175 vssd1
+ vssd1 vccd1 vccd1 genblk1\[0\].osc.clkdiv_C.cnt\[12\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_124_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_53_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11506_ genblk2\[8\].wave_shpr.div.quo\[8\] _05447_ _05446_ net404 vssd1 vssd1 vccd1
+ vccd1 _00803_ sky130_fd_sc_hd__a22o_1
X_12486_ clknet_leaf_107_clk _00048_ net151 vssd1 vssd1 vccd1 vccd1 sig_norm.acc\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10991__A3 _05023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11437_ genblk2\[8\].wave_shpr.div.acc\[23\] _05412_ vssd1 vssd1 vccd1 vccd1 _05413_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_1_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11368_ _05249_ _05245_ genblk2\[7\].wave_shpr.div.i\[0\] vssd1 vssd1 vccd1 vccd1
+ _05349_ sky130_fd_sc_hd__mux2_1
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13107_ clknet_leaf_13_clk _00432_ net53 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.i\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11548__A _03719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_95_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10319_ _04627_ vssd1 vssd1 vccd1 vccd1 _00436_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11299_ _05197_ _05173_ vssd1 vssd1 vccd1 vccd1 _05298_ sky130_fd_sc_hd__or2b_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13038_ clknet_leaf_126_clk _00365_ net66 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.b1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07761__A _02467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09452__S _00007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10598__S _00015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_135_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07530_ _02247_ vssd1 vssd1 vccd1 vccd1 _00027_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07461_ _02155_ _02192_ vssd1 vssd1 vccd1 vccd1 _02193_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09200_ _03828_ vssd1 vssd1 vccd1 vccd1 _00116_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06412_ _01226_ _01355_ vssd1 vssd1 vccd1 vccd1 _01356_ sky130_fd_sc_hd__or2_2
XANTENNA__11208__A1 _03726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07392_ _02141_ vssd1 vssd1 vccd1 vccd1 genblk1\[11\].osc.clkdiv_C.next_cnt\[14\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11759__A2 _03696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_134_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06343_ genblk1\[0\].osc.clkdiv_C.cnt\[12\] _01290_ _01292_ vssd1 vssd1 vccd1 vccd1
+ genblk1\[0\].osc.clkdiv_C.next_cnt\[12\] sky130_fd_sc_hd__o21a_1
X_09131_ genblk2\[0\].wave_shpr.div.b1\[8\] genblk2\[0\].wave_shpr.div.acc\[8\] vssd1
+ vssd1 vccd1 vccd1 _03779_ sky130_fd_sc_hd__and2b_1
XFILLER_0_115_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06824__B genblk1\[5\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09062_ _03701_ vssd1 vssd1 vccd1 vccd1 _03722_ sky130_fd_sc_hd__buf_4
X_06274_ genblk1\[0\].osc.clkdiv_C.cnt\[3\] _01227_ _01235_ genblk1\[0\].osc.clkdiv_C.cnt\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01236_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_142_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13080__RESET_B net63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08013_ genblk1\[6\].osc.clkdiv_C.cnt\[5\] _01367_ _02716_ _02718_ _02719_ vssd1
+ vssd1 vccd1 vccd1 _02720_ sky130_fd_sc_hd__o221a_1
XFILLER_0_8_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold600 genblk2\[6\].wave_shpr.div.acc\[15\] vssd1 vssd1 vccd1 vccd1 net818 sky130_fd_sc_hd__dlygate4sd3_1
Xhold611 genblk2\[1\].wave_shpr.div.acc\[4\] vssd1 vssd1 vccd1 vccd1 net829 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold622 genblk2\[0\].wave_shpr.div.acc\[15\] vssd1 vssd1 vccd1 vccd1 net840 sky130_fd_sc_hd__dlygate4sd3_1
Xhold633 genblk1\[4\].osc.clkdiv_C.cnt\[17\] vssd1 vssd1 vccd1 vccd1 net851 sky130_fd_sc_hd__dlygate4sd3_1
Xhold644 genblk2\[3\].wave_shpr.div.acc\[14\] vssd1 vssd1 vccd1 vccd1 net862 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold655 genblk2\[7\].wave_shpr.div.acc\[23\] vssd1 vssd1 vccd1 vccd1 net873 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold666 genblk2\[9\].wave_shpr.div.acc\[10\] vssd1 vssd1 vccd1 vccd1 net884 sky130_fd_sc_hd__dlygate4sd3_1
Xhold677 genblk2\[2\].wave_shpr.div.acc\[9\] vssd1 vssd1 vccd1 vccd1 net895 sky130_fd_sc_hd__dlygate4sd3_1
Xhold688 genblk2\[10\].wave_shpr.div.acc\[23\] vssd1 vssd1 vccd1 vccd1 net906 sky130_fd_sc_hd__dlygate4sd3_1
X_09964_ net282 _04359_ _04360_ vssd1 vssd1 vccd1 vccd1 _00348_ sky130_fd_sc_hd__a21oi_1
Xhold699 genblk2\[8\].wave_shpr.div.acc\[11\] vssd1 vssd1 vccd1 vccd1 net917 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08915_ _03614_ _03615_ vssd1 vssd1 vccd1 vccd1 _03616_ sky130_fd_sc_hd__nand2_1
X_09895_ net830 _04282_ _04289_ _04311_ vssd1 vssd1 vccd1 vccd1 _00328_ sky130_fd_sc_hd__a22o_1
XTAP_960 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_971 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08846_ _03484_ _03485_ _03497_ vssd1 vssd1 vccd1 vccd1 _03553_ sky130_fd_sc_hd__o21ba_1
XTAP_993 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08560__A1 genblk2\[8\].wave_shpr.div.fin_quo\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__07671__A _01308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08777_ _03465_ _03482_ _03333_ _03483_ vssd1 vssd1 vccd1 vccd1 _03484_ sky130_fd_sc_hd__o211a_1
XFILLER_0_79_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07728_ _01342_ genblk1\[1\].osc.clkdiv_C.cnt\[7\] vssd1 vssd1 vccd1 vccd1 _02435_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07659_ net3 _02364_ _02365_ vssd1 vssd1 vccd1 vccd1 _02366_ sky130_fd_sc_hd__nand3_2
XFILLER_0_94_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10670_ _02182_ vssd1 vssd1 vccd1 vccd1 _04861_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_63_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09329_ _03838_ vssd1 vssd1 vccd1 vccd1 _03910_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_146_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10958__B1 _05055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12340_ _03833_ _02080_ vssd1 vssd1 vccd1 vccd1 _06028_ sky130_fd_sc_hd__nor2_1
XFILLER_0_51_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12271_ _05996_ vssd1 vssd1 vccd1 vccd1 _01019_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11222_ genblk2\[7\].wave_shpr.div.quo\[5\] _05246_ _05250_ net661 vssd1 vssd1 vccd1
+ vccd1 _00716_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11153_ _05049_ genblk2\[7\].wave_shpr.div.acc\[16\] vssd1 vssd1 vccd1 vccd1 _05213_
+ sky130_fd_sc_hd__and2_1
X_10104_ _04455_ vssd1 vssd1 vccd1 vccd1 _04462_ sky130_fd_sc_hd__buf_2
X_11084_ _05149_ _05021_ genblk2\[6\].wave_shpr.div.acc\[24\] vssd1 vssd1 vccd1 vccd1
+ _05151_ sky130_fd_sc_hd__mux2_1
X_10035_ genblk2\[3\].wave_shpr.div.fin_quo\[4\] genblk2\[3\].wave_shpr.div.quo\[3\]
+ _04422_ vssd1 vssd1 vccd1 vccd1 _04427_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10211__S _04507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11986_ genblk2\[11\].wave_shpr.div.b1\[2\] _01811_ _05433_ vssd1 vssd1 vccd1 vccd1
+ _05798_ sky130_fd_sc_hd__mux2_1
XANTENNA__09500__B1 _03733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13725_ clknet_leaf_97_clk net403 net166 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10937_ _05054_ vssd1 vssd1 vccd1 vccd1 _05055_ sky130_fd_sc_hd__buf_4
XFILLER_0_86_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_85_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13656_ clknet_leaf_44_clk _00969_ net116 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.quo\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10661__A2 _04853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10868_ genblk2\[6\].wave_shpr.div.b1\[15\] genblk2\[6\].wave_shpr.div.acc\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05012_ sky130_fd_sc_hd__and2b_1
XFILLER_0_128_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_66_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12607_ clknet_leaf_22_clk genblk1\[3\].osc.clkdiv_C.next_cnt\[10\] net94 vssd1 vssd1
+ vccd1 vccd1 genblk1\[3\].osc.clkdiv_C.cnt\[10\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_143_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12138__S _05865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13587_ clknet_leaf_73_clk _00902_ net215 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.acc\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10799_ _04949_ _04950_ vssd1 vssd1 vccd1 vccd1 _04951_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12538_ clknet_leaf_63_clk _00090_ net190 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.b1\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10413__A2 _04651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12469_ clknet_leaf_33_clk smpl_rt_clkdiv.clkDiv_inst.next_cnt\[3\] net101 vssd1
+ vssd1 vccd1 vccd1 smpl_rt_clkdiv.clkDiv_inst.cnt\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06961_ _01432_ _01221_ vssd1 vssd1 vccd1 vccd1 _01797_ sky130_fd_sc_hd__nand2_2
X_08700_ _03405_ _03404_ _03401_ vssd1 vssd1 vccd1 vccd1 _03407_ sky130_fd_sc_hd__a21bo_1
X_09680_ genblk2\[2\].wave_shpr.div.acc\[13\] genblk2\[2\].wave_shpr.div.b1\[13\]
+ vssd1 vssd1 vccd1 vccd1 _04160_ sky130_fd_sc_hd__or2b_1
X_06892_ genblk1\[6\].osc.clkdiv_C.cnt\[14\] _01675_ _01666_ genblk1\[6\].osc.clkdiv_C.cnt\[13\]
+ _01745_ vssd1 vssd1 vccd1 vccd1 _01746_ sky130_fd_sc_hd__o221ai_2
XANTENNA__09182__S _03722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08542__A1 genblk2\[7\].wave_shpr.div.fin_quo\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_146_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08631_ _03336_ _03337_ vssd1 vssd1 vccd1 vccd1 _03338_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08562_ _02676_ _02679_ _02680_ genblk2\[7\].wave_shpr.div.fin_quo\[0\] vssd1 vssd1
+ vccd1 vccd1 _03269_ sky130_fd_sc_hd__o211a_1
XFILLER_0_89_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07513_ _02232_ PWM.final_sample_in\[3\] vssd1 vssd1 vccd1 vccd1 _02233_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08493_ _03196_ _03199_ vssd1 vssd1 vccd1 vccd1 _03200_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_119_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout38 net44 vssd1 vssd1 vccd1 vccd1 net38 sky130_fd_sc_hd__buf_4
X_07444_ genblk2\[5\].wave_shpr.div.i\[1\] _02179_ genblk2\[5\].wave_shpr.div.i\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02180_ sky130_fd_sc_hd__or3b_1
XFILLER_0_18_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13261__RESET_B net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout49 net50 vssd1 vssd1 vccd1 vccd1 net49 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_146_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_64_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09211__A _03833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10357__A _03708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07375_ genblk1\[11\].osc.clkdiv_C.cnt\[11\] vssd1 vssd1 vccd1 vccd1 _02128_ sky130_fd_sc_hd__inv_2
XFILLER_0_146_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09114_ genblk2\[0\].wave_shpr.div.b1\[1\] genblk2\[0\].wave_shpr.div.acc\[1\] vssd1
+ vssd1 vccd1 vccd1 _03762_ sky130_fd_sc_hd__or2b_1
XFILLER_0_60_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06326_ genblk1\[0\].osc.clkdiv_C.cnt\[6\] _01279_ vssd1 vssd1 vccd1 vccd1 _01282_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09270__A2 _03804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06257_ genblk1\[0\].osc.clkdiv_C.cnt\[10\] _01184_ _01206_ _01218_ vssd1 vssd1 vccd1
+ vccd1 _01219_ sky130_fd_sc_hd__o211a_1
XFILLER_0_115_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09045_ net1238 _01991_ _03708_ vssd1 vssd1 vccd1 vccd1 _03711_ sky130_fd_sc_hd__mux2_1
XFILLER_0_143_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09558__B1 _04046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06188_ _01158_ vssd1 vssd1 vccd1 vccd1 _00024_ sky130_fd_sc_hd__clkbuf_4
Xhold430 genblk2\[2\].wave_shpr.div.acc\[20\] vssd1 vssd1 vccd1 vccd1 net648 sky130_fd_sc_hd__dlygate4sd3_1
Xhold441 genblk2\[6\].wave_shpr.div.acc\[23\] vssd1 vssd1 vccd1 vccd1 net659 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11365__B1 _05248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold452 genblk2\[7\].wave_shpr.div.quo\[12\] vssd1 vssd1 vccd1 vccd1 net670 sky130_fd_sc_hd__dlygate4sd3_1
Xhold463 _00475_ vssd1 vssd1 vccd1 vccd1 net681 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold474 genblk2\[5\].wave_shpr.div.b1\[2\] vssd1 vssd1 vccd1 vccd1 net692 sky130_fd_sc_hd__dlygate4sd3_1
Xhold485 genblk2\[8\].wave_shpr.div.b1\[16\] vssd1 vssd1 vccd1 vccd1 net703 sky130_fd_sc_hd__dlygate4sd3_1
Xhold496 genblk2\[4\].wave_shpr.div.quo\[24\] vssd1 vssd1 vccd1 vccd1 net714 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07584__A2 _01234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09947_ genblk2\[2\].wave_shpr.div.acc\[24\] _04212_ genblk2\[2\].wave_shpr.div.acc\[25\]
+ vssd1 vssd1 vccd1 vccd1 _04349_ sky130_fd_sc_hd__o21ai_1
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09878_ net836 _04282_ _04289_ _04298_ vssd1 vssd1 vccd1 vccd1 _00324_ sky130_fd_sc_hd__a22o_1
Xhold1130 genblk2\[2\].wave_shpr.div.quo\[0\] vssd1 vssd1 vccd1 vccd1 net1348 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout69_A net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08829_ _03533_ _03535_ vssd1 vssd1 vccd1 vccd1 _03536_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10340__A1 _03714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10340__B2 _03727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11840_ _05593_ _05681_ vssd1 vssd1 vccd1 vccd1 _05682_ sky130_fd_sc_hd__xnor2_1
XTAP_2635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11771_ _05631_ genblk1\[9\].osc.clkdiv_C.cnt\[7\] vssd1 vssd1 vccd1 vccd1 _05635_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_68_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13510_ clknet_leaf_80_clk _00827_ net205 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.acc\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10722_ net888 _04886_ _04890_ _04893_ vssd1 vssd1 vccd1 vccd1 _00573_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13441_ clknet_leaf_95_clk _00760_ net162 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.acc\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10653_ _04854_ vssd1 vssd1 vccd1 vccd1 _04855_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_82_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13372_ clknet_leaf_115_clk _00691_ net140 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.fin_quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_63_473 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10584_ _04649_ genblk2\[5\].wave_shpr.div.acc\[16\] vssd1 vssd1 vccd1 vccd1 _04812_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_2_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12323_ net351 _06014_ _06015_ net489 _06019_ vssd1 vssd1 vccd1 vccd1 _01048_ sky130_fd_sc_hd__a221o_1
XFILLER_0_50_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12254_ _05987_ vssd1 vssd1 vccd1 vccd1 _01011_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11205_ _03831_ net722 _03728_ vssd1 vssd1 vccd1 vccd1 _00707_ sky130_fd_sc_hd__a21bo_1
X_12185_ net289 _05923_ _03855_ vssd1 vssd1 vccd1 vccd1 _05924_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07575__A2 _01925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09791__A _03833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11136_ _05174_ _05194_ _05195_ vssd1 vssd1 vccd1 vccd1 _05196_ sky130_fd_sc_hd__a21o_1
X_11067_ _05017_ net21 genblk2\[6\].wave_shpr.div.acc\[18\] vssd1 vssd1 vccd1 vccd1
+ _05140_ sky130_fd_sc_hd__o21ai_1
X_10018_ _04361_ _04412_ _04413_ vssd1 vssd1 vccd1 vccd1 _04414_ sky130_fd_sc_hd__a21o_1
XANTENNA__11545__B genblk1\[8\].osc.clkdiv_C.cnt\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10331__A1 _01304_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_137_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_137_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__08827__A2 _02592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11969_ _05789_ vssd1 vssd1 vccd1 vccd1 _00924_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10095__B1 _04456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13708_ clknet_leaf_36_clk _01019_ net104 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.b1\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_144 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09031__A _02155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11485__B1_N _03728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13639_ clknet_leaf_94_clk _00952_ net159 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07160_ genblk1\[9\].osc.clkdiv_C.cnt\[2\] genblk1\[9\].osc.clkdiv_C.cnt\[1\] genblk1\[9\].osc.clkdiv_C.cnt\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01958_ sky130_fd_sc_hd__and3_1
XFILLER_0_109_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_125_862 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06111_ net364 net338 vssd1 vssd1 vccd1 vccd1 smpl_rt_clkdiv.clkDiv_inst.next_cnt\[1\]
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_143_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07091_ genblk1\[8\].osc.clkdiv_C.cnt\[7\] _01897_ genblk1\[8\].osc.clkdiv_C.cnt\[8\]
+ vssd1 vssd1 vccd1 vccd1 _01901_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_124_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_22_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_112_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xfanout206 net209 vssd1 vssd1 vccd1 vccd1 net206 sky130_fd_sc_hd__clkbuf_4
Xfanout217 net218 vssd1 vssd1 vccd1 vccd1 net217 sky130_fd_sc_hd__buf_2
X_09801_ net719 _04248_ _04252_ net812 vssd1 vssd1 vccd1 vccd1 _00293_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07993_ genblk1\[6\].osc.clkdiv_C.cnt\[10\] _01484_ _01519_ genblk1\[6\].osc.clkdiv_C.cnt\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02700_ sky130_fd_sc_hd__o22a_1
X_09732_ genblk2\[2\].wave_shpr.div.acc\[23\] _04211_ vssd1 vssd1 vccd1 vccd1 _04212_
+ sky130_fd_sc_hd__or2_2
X_06944_ net1146 _01781_ _01784_ vssd1 vssd1 vccd1 vccd1 genblk1\[6\].osc.clkdiv_C.next_cnt\[13\]
+ sky130_fd_sc_hd__o21a_1
XANTENNA__12311__A2 _03947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08748__C _02365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09206__A _02171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09663_ _04147_ vssd1 vssd1 vccd1 vccd1 _00260_ sky130_fd_sc_hd__clkbuf_1
X_06875_ genblk1\[6\].osc.clkdiv_C.cnt\[2\] vssd1 vssd1 vccd1 vccd1 _01729_ sky130_fd_sc_hd__inv_2
X_08614_ genblk2\[4\].wave_shpr.div.fin_quo\[0\] _02932_ genblk2\[4\].wave_shpr.div.fin_quo\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03321_ sky130_fd_sc_hd__a21oi_1
X_09594_ _03986_ _03963_ vssd1 vssd1 vccd1 vccd1 _04097_ sky130_fd_sc_hd__or2b_1
XFILLER_0_89_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_49_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08545_ _02604_ _03248_ _03250_ _03247_ vssd1 vssd1 vccd1 vccd1 _03252_ sky130_fd_sc_hd__a22o_1
XANTENNA__08279__B1 _02223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_128_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_128_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__12075__B2 _05813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_420 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08476_ _02932_ _02840_ genblk2\[4\].wave_shpr.div.fin_quo\[3\] vssd1 vssd1 vccd1
+ vccd1 _03183_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_92_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07427_ genblk2\[3\].wave_shpr.div.i\[1\] _02166_ genblk2\[3\].wave_shpr.div.i\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02167_ sky130_fd_sc_hd__or3b_1
XFILLER_0_135_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10087__A _04455_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07358_ _02115_ vssd1 vssd1 vccd1 vccd1 genblk1\[11\].osc.clkdiv_C.next_cnt\[6\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_116_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06309_ _01268_ vssd1 vssd1 vccd1 vccd1 _01270_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07289_ genblk1\[10\].osc.clkdiv_C.cnt\[14\] genblk1\[10\].osc.clkdiv_C.cnt\[13\]
+ _02053_ vssd1 vssd1 vccd1 vccd1 _02057_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09028_ _03698_ vssd1 vssd1 vccd1 vccd1 _03699_ sky130_fd_sc_hd__inv_2
XANTENNA__12452__D net222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold260 genblk2\[9\].wave_shpr.div.b1\[13\] vssd1 vssd1 vccd1 vccd1 net478 sky130_fd_sc_hd__dlygate4sd3_1
Xhold271 genblk2\[11\].wave_shpr.div.quo\[14\] vssd1 vssd1 vccd1 vccd1 net489 sky130_fd_sc_hd__dlygate4sd3_1
Xhold282 genblk2\[5\].wave_shpr.div.quo\[11\] vssd1 vssd1 vccd1 vccd1 net500 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09951__A0 _04250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold293 genblk2\[1\].wave_shpr.div.quo\[14\] vssd1 vssd1 vccd1 vccd1 net511 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08506__B2 _02468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12302__A2 _06009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12941_ clknet_leaf_111_clk _00270_ net136 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.fin_quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06517__B1 _01442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12872_ clknet_leaf_134_clk _00203_ net59 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.b1\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11823_ _05585_ _05668_ vssd1 vssd1 vccd1 vccd1 _05669_ sky130_fd_sc_hd__xnor2_1
XTAP_2454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_119_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_119_clk
+ sky130_fd_sc_hd__clkbuf_16
XTAP_1720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11754_ _05464_ genblk1\[9\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 _05625_
+ sky130_fd_sc_hd__and2_1
XTAP_1775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10705_ _04818_ _04819_ vssd1 vssd1 vccd1 vccd1 _04880_ sky130_fd_sc_hd__nor2_2
XTAP_1797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11685_ genblk2\[9\].wave_shpr.div.b1\[2\] genblk2\[9\].wave_shpr.div.acc\[2\] vssd1
+ vssd1 vccd1 vccd1 _05577_ sky130_fd_sc_hd__and2b_1
XFILLER_0_102_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13424_ clknet_leaf_87_clk _00743_ net179 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.acc\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10636_ _04845_ vssd1 vssd1 vccd1 vccd1 _00535_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_141_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09234__A2 _03841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13355_ clknet_leaf_4_clk _00676_ net45 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.acc\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10567_ _04773_ _04793_ _04794_ vssd1 vssd1 vccd1 vccd1 _04795_ sky130_fd_sc_hd__a21o_1
XFILLER_0_140_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12306_ net358 _06009_ _06010_ net397 vssd1 vssd1 vccd1 vccd1 _01040_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13286_ clknet_leaf_118_clk _00607_ net137 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.fin_quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10498_ genblk2\[4\].wave_shpr.div.acc\[18\] _04738_ vssd1 vssd1 vccd1 vccd1 _04739_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12237_ genblk2\[11\].wave_shpr.div.b1\[17\] genblk2\[11\].wave_shpr.div.acc\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05975_ sky130_fd_sc_hd__and2b_1
X_12168_ _05785_ _05899_ _05912_ vssd1 vssd1 vccd1 vccd1 _05913_ sky130_fd_sc_hd__o21ai_1
XANTENNA__07753__B _02459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11119_ _05177_ _05178_ vssd1 vssd1 vccd1 vccd1 _05179_ sky130_fd_sc_hd__nand2_1
X_12099_ genblk2\[10\].wave_shpr.div.acc\[6\] _05861_ _05787_ vssd1 vssd1 vccd1 vccd1
+ _05862_ sky130_fd_sc_hd__mux2_1
Xinput6 pb[14] vssd1 vssd1 vccd1 vccd1 net6 sky130_fd_sc_hd__clkbuf_1
XANTENNA__06508__B1 _01432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11501__B1 _05446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06369__B _01208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06660_ net1237 _01549_ _01552_ vssd1 vssd1 vccd1 vccd1 genblk1\[3\].osc.clkdiv_C.next_cnt\[15\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_36_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09460__S _00007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07720__A2 _01309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06591_ genblk1\[3\].osc.clkdiv_C.cnt\[2\] _01496_ _01498_ genblk1\[3\].osc.clkdiv_C.cnt\[14\]
+ vssd1 vssd1 vccd1 vccd1 _01499_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_143_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08330_ _02682_ _03035_ _03036_ vssd1 vssd1 vccd1 vccd1 _03037_ sky130_fd_sc_hd__o21ai_1
XANTENNA__06385__A _01326_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08261_ _02966_ _02965_ vssd1 vssd1 vccd1 vccd1 _02968_ sky130_fd_sc_hd__and2b_1
XFILLER_0_117_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07212_ _01308_ genblk1\[10\].osc.clkdiv_C.cnt\[2\] _01214_ _01993_ genblk1\[10\].osc.clkdiv_C.cnt\[17\]
+ vssd1 vssd1 vccd1 vccd1 _01994_ sky130_fd_sc_hd__a221o_1
X_08192_ _02897_ _02898_ vssd1 vssd1 vccd1 vccd1 _02899_ sky130_fd_sc_hd__or2_1
XFILLER_0_61_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09225__A2 _03836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_144_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_70_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07143_ genblk1\[9\].osc.clkdiv_C.cnt\[3\] _01514_ vssd1 vssd1 vccd1 vccd1 _01943_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_30_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07074_ _01879_ _01889_ vssd1 vssd1 vccd1 vccd1 _01890_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10354__B _01242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07976_ genblk2\[7\].wave_shpr.div.fin_quo\[5\] vssd1 vssd1 vccd1 vccd1 _02683_ sky130_fd_sc_hd__inv_2
X_09715_ genblk2\[2\].wave_shpr.div.b1\[11\] genblk2\[2\].wave_shpr.div.acc\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04195_ sky130_fd_sc_hd__and2b_1
XANTENNA__12296__A1 _03687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06927_ genblk1\[6\].osc.clkdiv_C.cnt\[8\] genblk1\[6\].osc.clkdiv_C.cnt\[7\] _01770_
+ vssd1 vssd1 vccd1 vccd1 _01773_ sky130_fd_sc_hd__and3_1
X_09646_ genblk2\[1\].wave_shpr.div.acc\[20\] _04133_ _04136_ vssd1 vssd1 vccd1 vccd1
+ _04137_ sky130_fd_sc_hd__a21o_1
X_06858_ genblk1\[5\].osc.clkdiv_C.cnt\[13\] genblk1\[5\].osc.clkdiv_C.cnt\[12\] _01714_
+ vssd1 vssd1 vccd1 vccd1 _01717_ sky130_fd_sc_hd__and3_1
XTAP_1005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09577_ _03978_ _03967_ vssd1 vssd1 vccd1 vccd1 _04084_ sky130_fd_sc_hd__nor2_1
XTAP_1027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06789_ genblk1\[5\].osc.clkdiv_C.cnt\[2\] _01660_ vssd1 vssd1 vccd1 vccd1 _01661_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__12297__A _03942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08528_ _03230_ _03234_ vssd1 vssd1 vccd1 vccd1 _03235_ sky130_fd_sc_hd__nor2_1
XFILLER_0_77_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08267__A3 _02350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08459_ genblk2\[6\].wave_shpr.div.fin_quo\[3\] _02734_ _02736_ _02261_ vssd1 vssd1
+ vccd1 vccd1 _03166_ sky130_fd_sc_hd__a31o_1
XFILLER_0_65_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_462 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11470_ net1187 _01946_ _05237_ vssd1 vssd1 vccd1 vccd1 _05432_ sky130_fd_sc_hd__mux2_1
XFILLER_0_80_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_404 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10421_ genblk2\[4\].wave_shpr.div.acc\[0\] _00012_ _04679_ net643 _04680_ vssd1
+ vssd1 vccd1 vccd1 _00485_ sky130_fd_sc_hd__o221a_1
XFILLER_0_61_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13140_ clknet_leaf_115_clk _00465_ net133 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10352_ net1279 _04643_ _04637_ vssd1 vssd1 vccd1 vccd1 _04644_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13071_ clknet_leaf_24_clk _00398_ net92 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.quo\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10283_ _04576_ _04593_ _04594_ vssd1 vssd1 vccd1 vccd1 _04595_ sky130_fd_sc_hd__a21o_1
X_12022_ _05815_ vssd1 vssd1 vccd1 vccd1 _05817_ sky130_fd_sc_hd__buf_4
XANTENNA__07950__A2 _01564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12924_ clknet_leaf_35_clk _00255_ net105 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.acc\[22\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_88_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09280__S _03804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12855_ clknet_leaf_91_clk _00186_ net146 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.fin_quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11806_ net1006 _05652_ _05653_ _05656_ vssd1 vssd1 vccd1 vccd1 _00894_ sky130_fd_sc_hd__a22o_1
XTAP_2284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12786_ clknet_leaf_43_clk _00119_ net124 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.b1\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11737_ _05621_ vssd1 vssd1 vccd1 vccd1 _00860_ sky130_fd_sc_hd__clkbuf_1
XTAP_1594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11668_ genblk2\[9\].wave_shpr.div.acc\[11\] genblk2\[9\].wave_shpr.div.b1\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05560_ sky130_fd_sc_hd__or2b_1
XFILLER_0_36_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13407_ clknet_leaf_90_clk _00726_ net144 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.quo\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_52_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10619_ _04835_ vssd1 vssd1 vccd1 vccd1 _00528_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07748__B _01576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11599_ net909 _05507_ _05484_ _05510_ vssd1 vssd1 vccd1 vccd1 _00833_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07769__A2 _01256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13338_ clknet_leaf_8_clk _00659_ net50 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.acc\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13188__D _00015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13269_ clknet_leaf_1_clk _00592_ net41 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.acc\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_110_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10525__A1 _04655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07830_ _02461_ _02463_ genblk2\[1\].wave_shpr.div.fin_quo\[4\] vssd1 vssd1 vccd1
+ vccd1 _02537_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_138_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07761_ _02467_ vssd1 vssd1 vccd1 vccd1 _02468_ sky130_fd_sc_hd__clkbuf_4
X_09500_ _03732_ net369 _03733_ vssd1 vssd1 vccd1 vccd1 _00204_ sky130_fd_sc_hd__o21a_1
X_06712_ _01601_ vssd1 vssd1 vccd1 vccd1 genblk1\[4\].osc.clkdiv_C.next_cnt\[0\] sky130_fd_sc_hd__clkbuf_1
X_07692_ genblk1\[10\].osc.clkdiv_C.cnt\[11\] _02011_ vssd1 vssd1 vccd1 vccd1 _02399_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_154_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09190__S _03822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09431_ _03959_ _03993_ _03994_ vssd1 vssd1 vccd1 vccd1 _03995_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06643_ net1145 _01538_ _01541_ vssd1 vssd1 vccd1 vccd1 genblk1\[3\].osc.clkdiv_C.next_cnt\[9\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_87_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09362_ _03802_ _03923_ vssd1 vssd1 vccd1 vccd1 _03934_ sky130_fd_sc_hd__nor2_1
X_06574_ _01452_ _01482_ vssd1 vssd1 vccd1 vccd1 genblk1\[2\].osc.clkdiv_C.next_cnt\[17\]
+ sky130_fd_sc_hd__nor2_1
X_08313_ _02406_ _02404_ _02408_ _02525_ vssd1 vssd1 vccd1 vccd1 _03020_ sky130_fd_sc_hd__o31a_1
XFILLER_0_75_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09293_ genblk2\[0\].wave_shpr.div.acc\[5\] _03882_ _03804_ vssd1 vssd1 vccd1 vccd1
+ _03883_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08244_ _02947_ _02948_ _02949_ _02950_ vssd1 vssd1 vccd1 vccd1 _02951_ sky130_fd_sc_hd__o211a_1
XFILLER_0_145_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08175_ _02872_ _02881_ _02877_ vssd1 vssd1 vccd1 vccd1 _02882_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07126_ genblk1\[9\].osc.clkdiv_C.cnt\[5\] _01925_ _01855_ genblk1\[9\].osc.clkdiv_C.cnt\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01926_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07057_ genblk1\[8\].osc.clkdiv_C.cnt\[14\] _01246_ genblk1\[8\].osc.clkdiv_C.cnt\[17\]
+ vssd1 vssd1 vccd1 vccd1 _01875_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_2_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07959_ genblk1\[7\].osc.clkdiv_C.cnt\[10\] _01311_ _01925_ genblk1\[7\].osc.clkdiv_C.cnt\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02666_ sky130_fd_sc_hd__a22o_1
Xmax_cap24 net1353 vssd1 vssd1 vccd1 vccd1 net24 sky130_fd_sc_hd__buf_1
X_10970_ _05059_ genblk1\[6\].osc.clkdiv_C.cnt\[9\] vssd1 vssd1 vccd1 vccd1 _05070_
+ sky130_fd_sc_hd__and2_1
XANTENNA__07145__B1 _01513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09629_ _04123_ _04001_ vssd1 vssd1 vccd1 vccd1 _04124_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_97_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12640_ clknet_leaf_15_clk genblk1\[5\].osc.clkdiv_C.next_cnt\[7\] net73 vssd1 vssd1
+ vccd1 vccd1 genblk1\[5\].osc.clkdiv_C.cnt\[7\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_78_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_155_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12571_ clknet_leaf_28_clk genblk1\[1\].osc.clkdiv_C.next_cnt\[10\] net89 vssd1 vssd1
+ vccd1 vccd1 genblk1\[1\].osc.clkdiv_C.cnt\[10\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_65_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_108_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_50_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_50_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_136_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11522_ net237 _05454_ _05449_ net312 _05457_ vssd1 vssd1 vccd1 vccd1 _00809_ sky130_fd_sc_hd__a221o_1
XFILLER_0_150_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11453_ _05423_ vssd1 vssd1 vccd1 vccd1 _00774_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_150_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_34_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10404_ genblk2\[4\].wave_shpr.div.quo\[19\] _04661_ _04663_ net255 _04670_ vssd1
+ vssd1 vccd1 vccd1 _00478_ sky130_fd_sc_hd__a221o_1
XFILLER_0_104_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11384_ genblk2\[8\].wave_shpr.div.acc\[15\] genblk2\[8\].wave_shpr.div.b1\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05360_ sky130_fd_sc_hd__or2b_1
XFILLER_0_150_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13123_ clknet_leaf_124_clk _00448_ net77 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.b1\[7\]
+ sky130_fd_sc_hd__dfrtp_2
X_10335_ _04635_ vssd1 vssd1 vccd1 vccd1 _00444_ sky130_fd_sc_hd__clkbuf_1
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13054_ clknet_leaf_113_clk net815 net128 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10266_ genblk2\[4\].wave_shpr.div.b1\[4\] genblk2\[4\].wave_shpr.div.acc\[4\] vssd1
+ vssd1 vccd1 vccd1 _04578_ sky130_fd_sc_hd__or2b_1
X_12005_ _05807_ vssd1 vssd1 vccd1 vccd1 _00942_ sky130_fd_sc_hd__clkbuf_1
X_10197_ _04407_ _04364_ vssd1 vssd1 vccd1 vccd1 _04526_ sky130_fd_sc_hd__or2b_1
XFILLER_0_88_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12907_ clknet_leaf_36_clk _00238_ net102 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.acc\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12838_ clknet_leaf_65_clk _00171_ net196 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.acc\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2070 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2081 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2092 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12769_ clknet_leaf_93_clk _00102_ net148 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.fin_quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_579 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_41_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_41_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08100__A2 _02805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06290_ genblk1\[0\].osc.clkdiv_C.cnt\[11\] _01251_ vssd1 vssd1 vccd1 vccd1 _01252_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_613 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_141_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold804 genblk2\[9\].wave_shpr.div.acc\[2\] vssd1 vssd1 vccd1 vccd1 net1022 sky130_fd_sc_hd__dlygate4sd3_1
Xhold815 genblk2\[0\].wave_shpr.div.acc\[4\] vssd1 vssd1 vccd1 vccd1 net1033 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold826 genblk2\[11\].wave_shpr.div.acc\[1\] vssd1 vssd1 vccd1 vccd1 net1044 sky130_fd_sc_hd__dlygate4sd3_1
Xhold837 genblk2\[3\].wave_shpr.div.acc\[20\] vssd1 vssd1 vccd1 vccd1 net1055 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold848 genblk2\[0\].wave_shpr.div.acc\[1\] vssd1 vssd1 vccd1 vccd1 net1066 sky130_fd_sc_hd__dlygate4sd3_1
X_09980_ _04374_ _04375_ vssd1 vssd1 vccd1 vccd1 _04376_ sky130_fd_sc_hd__nand2_1
XFILLER_0_110_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold859 genblk1\[3\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 net1077 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07494__A net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08931_ net1141 _02260_ _03626_ _03574_ vssd1 vssd1 vccd1 vccd1 _00049_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08862_ _03136_ _03224_ vssd1 vssd1 vccd1 vccd1 _03569_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08102__B _01574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07813_ _02424_ _02471_ _02519_ vssd1 vssd1 vccd1 vccd1 _02520_ sky130_fd_sc_hd__nor3_2
X_08793_ _03484_ _03498_ _03395_ _03499_ vssd1 vssd1 vccd1 vccd1 _03500_ sky130_fd_sc_hd__o211a_1
XANTENNA__11744__A _03693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07744_ genblk1\[1\].osc.clkdiv_C.cnt\[13\] _02425_ _01344_ genblk1\[1\].osc.clkdiv_C.cnt\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02451_ sky130_fd_sc_hd__o22ai_2
XANTENNA__07127__B1 _01923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09081__B1_N _03717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07675_ _02369_ _02370_ vssd1 vssd1 vccd1 vccd1 _02382_ sky130_fd_sc_hd__nand2_1
XFILLER_0_94_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09414_ genblk2\[1\].wave_shpr.div.b1\[4\] genblk2\[1\].wave_shpr.div.acc\[4\] vssd1
+ vssd1 vccd1 vccd1 _03978_ sky130_fd_sc_hd__and2b_1
XFILLER_0_149_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06626_ genblk1\[3\].osc.clkdiv_C.cnt\[3\] _01528_ vssd1 vssd1 vccd1 vccd1 _01531_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09345_ net604 _03903_ _03910_ _03922_ vssd1 vssd1 vccd1 vccd1 _00167_ sky130_fd_sc_hd__a22o_1
XFILLER_0_90_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06557_ net1213 _01468_ _01471_ vssd1 vssd1 vccd1 vccd1 genblk1\[2\].osc.clkdiv_C.next_cnt\[11\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_75_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_32_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_32_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__07669__A _01188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09276_ _03839_ _03867_ _03869_ _03841_ net1139 vssd1 vssd1 vccd1 vccd1 _00151_ sky130_fd_sc_hd__a32o_1
XFILLER_0_47_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06488_ genblk1\[2\].osc.clkdiv_C.cnt\[2\] vssd1 vssd1 vccd1 vccd1 _01414_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08227_ genblk2\[4\].wave_shpr.div.fin_quo\[5\] _02932_ _02842_ _02316_ vssd1 vssd1
+ vccd1 vccd1 _02934_ sky130_fd_sc_hd__a31o_1
XFILLER_0_118_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_105_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08158_ genblk1\[3\].osc.clkdiv_C.cnt\[7\] _01483_ _01858_ _01486_ _02864_ vssd1
+ vssd1 vccd1 vccd1 _02865_ sky130_fd_sc_hd__a221o_1
XFILLER_0_43_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07109_ _01886_ _01912_ vssd1 vssd1 vccd1 vccd1 _01913_ sky130_fd_sc_hd__nor2_1
X_08089_ genblk2\[5\].wave_shpr.div.fin_quo\[7\] _02309_ _02795_ _02527_ vssd1 vssd1
+ vccd1 vccd1 _02796_ sky130_fd_sc_hd__a22o_1
XFILLER_0_101_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_101_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10120_ _04465_ genblk1\[3\].osc.clkdiv_C.cnt\[10\] vssd1 vssd1 vccd1 vccd1 _04471_
+ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_99_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_99_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__08158__A2 _01483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10051_ _04434_ vssd1 vssd1 vccd1 vccd1 _00361_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12938__RESET_B net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09658__A2 _04048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13741_ clknet_leaf_46_clk _01052_ net121 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.quo\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10953_ net344 _05057_ _05055_ net477 _05060_ vssd1 vssd1 vccd1 vccd1 _00637_ sky130_fd_sc_hd__a221o_1
XFILLER_0_85_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_98_799 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13672_ clknet_leaf_40_clk _00985_ net117 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.acc\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10884_ genblk2\[6\].wave_shpr.div.fin_quo\[2\] net1338 _00017_ vssd1 vssd1 vccd1
+ vccd1 _05026_ sky130_fd_sc_hd__mux2_1
X_12623_ clknet_leaf_16_clk genblk1\[4\].osc.clkdiv_C.next_cnt\[8\] net74 vssd1 vssd1
+ vccd1 vccd1 genblk1\[4\].osc.clkdiv_C.cnt\[8\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_155_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06892__A2 _01675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_23_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_23_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_93_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12554_ clknet_leaf_55_clk genblk1\[0\].osc.clkdiv_C.next_cnt\[11\] net175 vssd1
+ vssd1 vccd1 vccd1 genblk1\[0\].osc.clkdiv_C.cnt\[11\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_54_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11505_ _05441_ vssd1 vssd1 vccd1 vccd1 _05447_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_108_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12485_ clknet_leaf_106_clk _00047_ net151 vssd1 vssd1 vccd1 vccd1 sig_norm.acc\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09794__A _04247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_908 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11436_ genblk2\[8\].wave_shpr.div.acc\[22\] _05411_ vssd1 vssd1 vccd1 vccd1 _05412_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_80_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08397__A2 _01209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11367_ net381 _05251_ _05248_ _05348_ vssd1 vssd1 vccd1 vccd1 _00763_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_0_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13106_ clknet_leaf_12_clk _00431_ net52 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.i\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10318_ genblk2\[4\].wave_shpr.div.fin_quo\[3\] genblk2\[4\].wave_shpr.div.quo\[2\]
+ _00013_ vssd1 vssd1 vccd1 vccd1 _04627_ sky130_fd_sc_hd__mux2_1
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11298_ net1009 _05279_ _05283_ _05297_ vssd1 vssd1 vccd1 vccd1 _00745_ sky130_fd_sc_hd__a22o_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13037_ clknet_leaf_125_clk _00364_ net72 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.b1\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10249_ genblk2\[3\].wave_shpr.div.i\[3\] _02168_ _04560_ vssd1 vssd1 vccd1 vccd1
+ _04563_ sky130_fd_sc_hd__and3_1
XFILLER_0_119_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10900__A1 _01991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_62_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10664__B1 _04857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07460_ genblk2\[7\].wave_shpr.div.busy _02191_ vssd1 vssd1 vccd1 vccd1 _02192_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06411_ _01354_ vssd1 vssd1 vccd1 vccd1 _01355_ sky130_fd_sc_hd__buf_4
XFILLER_0_57_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06883__A2 _01484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07391_ _02091_ _02138_ _02140_ vssd1 vssd1 vccd1 vccd1 _02141_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_151_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_14_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_14_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_146_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10416__B1 _04654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09130_ _03756_ _03776_ _03777_ vssd1 vssd1 vccd1 vccd1 _03778_ sky130_fd_sc_hd__a21o_1
XFILLER_0_57_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06342_ _01268_ _01291_ vssd1 vssd1 vccd1 vccd1 _01292_ sky130_fd_sc_hd__nor2_1
XANTENNA__07489__A _02147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06393__A _01336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_77_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09061_ _01193_ vssd1 vssd1 vccd1 vccd1 _03721_ sky130_fd_sc_hd__inv_2
X_06273_ _01231_ _01234_ vssd1 vssd1 vccd1 vccd1 _01235_ sky130_fd_sc_hd__nor2_4
XFILLER_0_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12169__B1 _05816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_120_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08012_ genblk1\[6\].osc.clkdiv_C.cnt\[4\] _01747_ vssd1 vssd1 vccd1 vccd1 _02719_
+ sky130_fd_sc_hd__or2_1
XANTENNA__07134__A1_N genblk1\[9\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold601 genblk2\[6\].wave_shpr.div.acc\[6\] vssd1 vssd1 vccd1 vccd1 net819 sky130_fd_sc_hd__dlygate4sd3_1
Xhold612 genblk2\[2\].wave_shpr.div.acc\[11\] vssd1 vssd1 vccd1 vccd1 net830 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold623 genblk2\[11\].wave_shpr.div.acc\[6\] vssd1 vssd1 vccd1 vccd1 net841 sky130_fd_sc_hd__dlygate4sd3_1
Xhold634 genblk2\[7\].wave_shpr.div.acc\[12\] vssd1 vssd1 vccd1 vccd1 net852 sky130_fd_sc_hd__dlygate4sd3_1
Xhold645 genblk2\[5\].wave_shpr.div.acc\[6\] vssd1 vssd1 vccd1 vccd1 net863 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout101_A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold656 genblk2\[1\].wave_shpr.div.acc\[20\] vssd1 vssd1 vccd1 vccd1 net874 sky130_fd_sc_hd__dlygate4sd3_1
Xhold667 genblk2\[5\].wave_shpr.div.acc\[5\] vssd1 vssd1 vccd1 vccd1 net885 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold678 genblk2\[5\].wave_shpr.div.acc\[19\] vssd1 vssd1 vccd1 vccd1 net896 sky130_fd_sc_hd__dlygate4sd3_1
X_09963_ net282 _04359_ _03855_ vssd1 vssd1 vccd1 vccd1 _04360_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_110_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_135_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold689 genblk2\[6\].wave_shpr.div.acc\[5\] vssd1 vssd1 vccd1 vccd1 net907 sky130_fd_sc_hd__dlygate4sd3_1
X_08914_ sig_norm.acc\[5\] _03611_ vssd1 vssd1 vccd1 vccd1 _03615_ sky130_fd_sc_hd__nand2_1
X_09894_ genblk2\[2\].wave_shpr.div.acc\[10\] _04310_ _04301_ vssd1 vssd1 vccd1 vccd1
+ _04311_ sky130_fd_sc_hd__mux2_1
XTAP_950 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_961 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_15_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12341__B1 _03941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_972 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08845_ _03533_ _03535_ vssd1 vssd1 vccd1 vccd1 _03552_ sky130_fd_sc_hd__and2b_1
XTAP_983 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_994 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08560__A2 _02362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08776_ _03298_ _03332_ _03331_ vssd1 vssd1 vccd1 vccd1 _03483_ sky130_fd_sc_hd__a21bo_1
XTAP_2806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07727_ genblk1\[1\].osc.clkdiv_C.cnt\[5\] _02433_ _01305_ genblk1\[1\].osc.clkdiv_C.cnt\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02434_ sky130_fd_sc_hd__o22ai_1
XTAP_2839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06287__B _01188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07658_ _02312_ vssd1 vssd1 vccd1 vccd1 _02365_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_67_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06323__A1 genblk1\[0\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06609_ genblk1\[3\].osc.clkdiv_C.cnt\[4\] _01514_ _01513_ genblk1\[3\].osc.clkdiv_C.cnt\[3\]
+ vssd1 vssd1 vccd1 vccd1 _01517_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_137_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_4_8_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_8_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_47_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07589_ _02282_ _02286_ _02292_ _02295_ vssd1 vssd1 vccd1 vccd1 _02296_ sky130_fd_sc_hd__o31a_1
X_09328_ net913 _03903_ _03877_ _03909_ vssd1 vssd1 vccd1 vccd1 _00163_ sky130_fd_sc_hd__a22o_1
XANTENNA__09812__A2 _04253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09259_ _03853_ genblk1\[0\].osc.clkdiv_C.cnt\[13\] vssd1 vssd1 vccd1 vccd1 _03859_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_7_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09025__B1 _03696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12270_ net1267 _04229_ _05994_ vssd1 vssd1 vccd1 vccd1 _05996_ sky130_fd_sc_hd__mux2_1
XANTENNA__11907__B1 _03855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11221_ genblk2\[7\].wave_shpr.div.quo\[4\] _05246_ _05250_ net331 vssd1 vssd1 vccd1
+ vccd1 _00715_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07587__B1 _01513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11152_ _05166_ _05210_ _05211_ vssd1 vssd1 vccd1 vccd1 _05212_ sky130_fd_sc_hd__a21oi_1
X_10103_ _04451_ vssd1 vssd1 vccd1 vccd1 _04461_ sky130_fd_sc_hd__buf_2
X_11083_ genblk2\[6\].wave_shpr.div.acc\[24\] _05057_ _05126_ _05150_ vssd1 vssd1
+ vccd1 vccd1 _00677_ sky130_fd_sc_hd__a22o_1
X_10034_ _04426_ vssd1 vssd1 vccd1 vccd1 _00352_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10894__A0 genblk2\[6\].wave_shpr.div.fin_quo\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11985_ _05797_ vssd1 vssd1 vccd1 vccd1 _00932_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__09500__A1 _03732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10936_ _05053_ vssd1 vssd1 vccd1 vccd1 _05054_ sky130_fd_sc_hd__clkbuf_4
X_13724_ clknet_leaf_96_clk _01035_ net160 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.quo\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13655_ clknet_leaf_41_clk _00968_ net116 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.quo\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10867_ _04969_ _05009_ _05010_ vssd1 vssd1 vccd1 vccd1 _05011_ sky130_fd_sc_hd__a21o_1
XFILLER_0_85_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12606_ clknet_leaf_22_clk genblk1\[3\].osc.clkdiv_C.next_cnt\[9\] net92 vssd1 vssd1
+ vccd1 vccd1 genblk1\[3\].osc.clkdiv_C.cnt\[9\] sky130_fd_sc_hd__dfrtp_2
XPHY_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13586_ clknet_leaf_72_clk _00901_ net215 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.acc\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09264__B1 _03838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10798_ genblk2\[5\].wave_shpr.div.acc\[23\] _04818_ vssd1 vssd1 vccd1 vccd1 _04950_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_38_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09803__A2 _04248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07102__A genblk1\[8\].osc.clkdiv_C.cnt\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12537_ clknet_leaf_41_clk _00089_ net123 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.b1\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12468_ clknet_leaf_34_clk smpl_rt_clkdiv.clkDiv_inst.next_cnt\[2\] net99 vssd1 vssd1
+ vccd1 vccd1 smpl_rt_clkdiv.clkDiv_inst.cnt\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11419_ _05365_ _05393_ _05394_ vssd1 vssd1 vccd1 vccd1 _05395_ sky130_fd_sc_hd__a21o_1
X_12399_ net949 _06039_ _06040_ _06071_ vssd1 vssd1 vccd1 vccd1 _01072_ sky130_fd_sc_hd__a22o_1
XANTENNA__07042__A2 _01436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06250__B1 _01210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06960_ genblk1\[7\].osc.clkdiv_C.cnt\[10\] genblk1\[7\].osc.clkdiv_C.cnt\[0\] _01514_
+ vssd1 vssd1 vccd1 vccd1 _01796_ sky130_fd_sc_hd__and3b_1
Xclkbuf_leaf_3_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_3_clk sky130_fd_sc_hd__clkbuf_16
X_06891_ genblk1\[6\].osc.clkdiv_C.cnt\[13\] _01666_ _01484_ genblk1\[6\].osc.clkdiv_C.cnt\[11\]
+ vssd1 vssd1 vccd1 vccd1 _01745_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__08542__A2 _02526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08630_ genblk2\[6\].wave_shpr.div.fin_quo\[2\] _02733_ _02735_ _02261_ vssd1 vssd1
+ vccd1 vccd1 _03337_ sky130_fd_sc_hd__a31o_1
XANTENNA__07491__B _02152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08561_ _03266_ _03267_ _02604_ vssd1 vssd1 vccd1 vccd1 _03268_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_77_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07512_ PWM.counter\[3\] vssd1 vssd1 vccd1 vccd1 _02232_ sky130_fd_sc_hd__inv_2
X_08492_ _03197_ _03198_ vssd1 vssd1 vccd1 vccd1 _03199_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07443_ genblk2\[5\].wave_shpr.div.i\[2\] genblk2\[5\].wave_shpr.div.i\[3\] genblk2\[5\].wave_shpr.div.i\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02179_ sky130_fd_sc_hd__nand3b_1
Xfanout39 net44 vssd1 vssd1 vccd1 vccd1 net39 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_92_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13648__RESET_B net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout149_A net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07374_ net1269 _02123_ _02127_ _02092_ vssd1 vssd1 vccd1 vccd1 genblk1\[11\].osc.clkdiv_C.next_cnt\[10\]
+ sky130_fd_sc_hd__o211a_1
XFILLER_0_45_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10357__B _01441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09113_ genblk2\[0\].wave_shpr.div.b1\[2\] vssd1 vssd1 vccd1 vccd1 _03761_ sky130_fd_sc_hd__inv_2
XFILLER_0_134_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06325_ genblk1\[0\].osc.clkdiv_C.cnt\[6\] _01279_ vssd1 vssd1 vccd1 vccd1 _01281_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_115_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_828 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09044_ _03710_ vssd1 vssd1 vccd1 vccd1 _00078_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06256_ genblk1\[0\].osc.clkdiv_C.cnt\[15\] _01210_ _01212_ _01217_ vssd1 vssd1 vccd1
+ vccd1 _01218_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_142_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold420 _00472_ vssd1 vssd1 vccd1 vccd1 net638 sky130_fd_sc_hd__dlygate4sd3_1
X_06187_ _01157_ vssd1 vssd1 vccd1 vccd1 _01158_ sky130_fd_sc_hd__inv_2
Xhold431 genblk2\[9\].wave_shpr.div.quo\[1\] vssd1 vssd1 vccd1 vccd1 net649 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold442 genblk2\[8\].wave_shpr.div.quo\[20\] vssd1 vssd1 vccd1 vccd1 net660 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold453 genblk2\[6\].wave_shpr.div.quo\[2\] vssd1 vssd1 vccd1 vccd1 net671 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold464 genblk2\[10\].wave_shpr.div.quo\[3\] vssd1 vssd1 vccd1 vccd1 net682 sky130_fd_sc_hd__dlygate4sd3_1
Xhold475 genblk2\[7\].wave_shpr.div.quo\[2\] vssd1 vssd1 vccd1 vccd1 net693 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08136__C_N _02837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold486 genblk2\[8\].wave_shpr.div.acc\[23\] vssd1 vssd1 vccd1 vccd1 net704 sky130_fd_sc_hd__dlygate4sd3_1
Xhold497 genblk2\[0\].wave_shpr.div.acc\[0\] vssd1 vssd1 vccd1 vccd1 net715 sky130_fd_sc_hd__dlygate4sd3_1
X_09946_ net1094 _04253_ _04251_ _04348_ vssd1 vssd1 vccd1 vccd1 _00342_ sky130_fd_sc_hd__a22o_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09877_ genblk2\[2\].wave_shpr.div.acc\[6\] _04297_ _04214_ vssd1 vssd1 vccd1 vccd1
+ _04298_ sky130_fd_sc_hd__mux2_1
Xhold1120 genblk2\[6\].wave_shpr.div.quo\[1\] vssd1 vssd1 vccd1 vccd1 net1338 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1131 genblk2\[6\].wave_shpr.div.quo\[6\] vssd1 vssd1 vccd1 vccd1 net1349 sky130_fd_sc_hd__dlygate4sd3_1
X_08828_ net8 _02744_ _03534_ vssd1 vssd1 vccd1 vccd1 _03535_ sky130_fd_sc_hd__and3_1
XTAP_2603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08759_ genblk2\[5\].wave_shpr.div.fin_quo\[0\] _02467_ _02791_ vssd1 vssd1 vccd1
+ vccd1 _03466_ sky130_fd_sc_hd__a21o_1
XTAP_2625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11770_ net304 _05628_ _05629_ net485 _05634_ vssd1 vssd1 vccd1 vccd1 _00880_ sky130_fd_sc_hd__a221o_1
XTAP_2669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10721_ genblk2\[5\].wave_shpr.div.acc\[3\] _04892_ _04821_ vssd1 vssd1 vccd1 vccd1
+ _04893_ sky130_fd_sc_hd__mux2_1
XTAP_1957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13440_ clknet_leaf_95_clk _00759_ net162 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.acc\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10652_ _02170_ genblk2\[5\].wave_shpr.div.busy _02180_ vssd1 vssd1 vccd1 vccd1 _04854_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_76_791 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08018__A _01739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13371_ clknet_leaf_117_clk _00690_ net140 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.fin_quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10583_ _04765_ _04809_ _04810_ vssd1 vssd1 vccd1 vccd1 _04811_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_36_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12322_ _05835_ genblk1\[11\].osc.clkdiv_C.cnt\[6\] vssd1 vssd1 vccd1 vccd1 _06019_
+ sky130_fd_sc_hd__and2_1
XANTENNA__10800__B1 _04858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_198 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11379__A _03690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12253_ genblk2\[11\].wave_shpr.div.fin_quo\[4\] genblk2\[11\].wave_shpr.div.quo\[3\]
+ _00005_ vssd1 vssd1 vccd1 vccd1 _05987_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11204_ _03727_ _01490_ _03687_ net1005 vssd1 vssd1 vccd1 vccd1 _00706_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_31_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12184_ _03690_ _05922_ _05923_ vssd1 vssd1 vccd1 vccd1 _01005_ sky130_fd_sc_hd__nor3_1
XFILLER_0_102_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11135_ genblk2\[7\].wave_shpr.div.b1\[7\] genblk2\[7\].wave_shpr.div.acc\[7\] vssd1
+ vssd1 vccd1 vccd1 _05195_ sky130_fd_sc_hd__and2b_1
XFILLER_0_101_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12305__B1 _06010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11066_ _05018_ net21 vssd1 vssd1 vccd1 vccd1 _05139_ sky130_fd_sc_hd__or2_1
X_10017_ genblk2\[3\].wave_shpr.div.b1\[17\] genblk2\[3\].wave_shpr.div.acc\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04413_ sky130_fd_sc_hd__and2b_1
XFILLER_0_86_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11968_ genblk2\[10\].wave_shpr.div.fin_quo\[1\] genblk2\[10\].wave_shpr.div.quo\[0\]
+ _00003_ vssd1 vssd1 vccd1 vccd1 _05789_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10095__A1 genblk2\[3\].wave_shpr.div.quo\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10095__B2 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13707_ clknet_leaf_37_clk _01018_ net104 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.b1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10919_ _05044_ vssd1 vssd1 vccd1 vccd1 _00619_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_27_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11899_ _03839_ _05723_ _05724_ _03841_ net1106 vssd1 vssd1 vccd1 vccd1 _00919_ sky130_fd_sc_hd__a32o_1
XFILLER_0_67_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13638_ clknet_leaf_94_clk net221 net159 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.quo\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_116_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09237__B1 _03839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13569_ clknet_leaf_55_clk _00884_ net182 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.quo\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07799__B1 _01577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_54_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09458__S _00007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_81_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06110_ net338 vssd1 vssd1 vccd1 vccd1 smpl_rt_clkdiv.clkDiv_inst.next_cnt\[0\] sky130_fd_sc_hd__inv_2
XFILLER_0_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_125_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07090_ genblk1\[8\].osc.clkdiv_C.cnt\[8\] genblk1\[8\].osc.clkdiv_C.cnt\[7\] _01897_
+ vssd1 vssd1 vccd1 vccd1 _01900_ sky130_fd_sc_hd__and3_1
XFILLER_0_42_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09800_ net812 _04248_ _04252_ net1054 vssd1 vssd1 vccd1 vccd1 _00292_ sky130_fd_sc_hd__a22o_1
Xfanout207 net208 vssd1 vssd1 vccd1 vccd1 net207 sky130_fd_sc_hd__clkbuf_4
Xfanout218 net16 vssd1 vssd1 vccd1 vccd1 net218 sky130_fd_sc_hd__clkbuf_4
X_07992_ genblk2\[6\].wave_shpr.div.fin_quo\[5\] vssd1 vssd1 vccd1 vccd1 _02699_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12623__RESET_B net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09731_ genblk2\[2\].wave_shpr.div.acc\[22\] genblk2\[2\].wave_shpr.div.acc\[21\]
+ genblk2\[2\].wave_shpr.div.acc\[20\] _04210_ vssd1 vssd1 vccd1 vccd1 _04211_ sky130_fd_sc_hd__or4_1
X_06943_ net28 _01783_ vssd1 vssd1 vccd1 vccd1 _01784_ sky130_fd_sc_hd__nor2_1
X_09662_ _04046_ _04042_ genblk2\[1\].wave_shpr.div.i\[0\] vssd1 vssd1 vccd1 vccd1
+ _04147_ sky130_fd_sc_hd__mux2_1
X_06874_ genblk1\[6\].osc.clkdiv_C.cnt\[16\] _01578_ vssd1 vssd1 vccd1 vccd1 _01728_
+ sky130_fd_sc_hd__xnor2_1
X_08613_ _03318_ _03319_ _02797_ vssd1 vssd1 vccd1 vccd1 _03320_ sky130_fd_sc_hd__a21bo_1
X_09593_ net827 _04076_ _04080_ _04096_ vssd1 vssd1 vccd1 vccd1 _00241_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_77_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08544_ _02603_ _03247_ _03248_ _03250_ vssd1 vssd1 vccd1 vccd1 _03251_ sky130_fd_sc_hd__and4_1
XFILLER_0_49_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11283__B1 _05283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08475_ _03180_ _03181_ _02797_ vssd1 vssd1 vccd1 vccd1 _03182_ sky130_fd_sc_hd__o21a_1
XANTENNA__06829__A2 genblk1\[5\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_432 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_419 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_49_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_343 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07426_ genblk2\[3\].wave_shpr.div.i\[2\] genblk2\[3\].wave_shpr.div.i\[3\] genblk2\[3\].wave_shpr.div.i\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02166_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_92_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07357_ _02092_ _02113_ _02114_ vssd1 vssd1 vccd1 vccd1 _02115_ sky130_fd_sc_hd__and3_1
XFILLER_0_73_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06308_ net1089 _01269_ vssd1 vssd1 vccd1 vccd1 genblk1\[0\].osc.clkdiv_C.next_cnt\[0\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_143_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07288_ genblk1\[10\].osc.clkdiv_C.cnt\[13\] _02053_ genblk1\[10\].osc.clkdiv_C.cnt\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02056_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09027_ genblk2\[9\].wave_shpr.div.i\[1\] genblk2\[9\].wave_shpr.div.i\[0\] genblk2\[9\].wave_shpr.div.i\[2\]
+ genblk2\[9\].wave_shpr.div.i\[3\] vssd1 vssd1 vccd1 vccd1 _03698_ sky130_fd_sc_hd__and4_1
XFILLER_0_60_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06239_ _01200_ vssd1 vssd1 vccd1 vccd1 _01201_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_14_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09559__B_N _04046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold250 _01044_ vssd1 vssd1 vccd1 vccd1 net468 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold261 genblk2\[11\].wave_shpr.div.quo\[9\] vssd1 vssd1 vccd1 vccd1 net479 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_376 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold272 genblk2\[3\].wave_shpr.div.quo\[23\] vssd1 vssd1 vccd1 vccd1 net490 sky130_fd_sc_hd__dlygate4sd3_1
Xhold283 _00555_ vssd1 vssd1 vccd1 vccd1 net501 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09951__A1 _04247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold294 _00222_ vssd1 vssd1 vccd1 vccd1 net512 sky130_fd_sc_hd__dlygate4sd3_1
X_09929_ _04336_ _04337_ vssd1 vssd1 vccd1 vccd1 _04338_ sky130_fd_sc_hd__nand2_1
X_12940_ clknet_leaf_110_clk _00269_ net136 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.fin_quo\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12871_ clknet_leaf_134_clk _00202_ net59 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.b1\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11822_ _05586_ _05564_ vssd1 vssd1 vccd1 vccd1 _05668_ sky130_fd_sc_hd__or2b_1
XTAP_2444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11753_ net526 _05623_ _05624_ net1085 vssd1 vssd1 vccd1 vccd1 _00873_ sky130_fd_sc_hd__a22o_1
XTAP_2499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10704_ _03819_ net493 _00014_ genblk2\[5\].wave_shpr.div.acc\[0\] _04879_ vssd1
+ vssd1 vccd1 vccd1 _00569_ sky130_fd_sc_hd__o221a_1
XTAP_1787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11684_ _05572_ genblk2\[9\].wave_shpr.div.acc\[1\] _05575_ vssd1 vssd1 vccd1 vccd1
+ _05576_ sky130_fd_sc_hd__a21o_1
XFILLER_0_138_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13423_ clknet_leaf_87_clk _00742_ net179 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.acc\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10635_ genblk2\[6\].wave_shpr.div.b1\[10\] _04844_ _04834_ vssd1 vssd1 vccd1 vccd1
+ _04845_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13354_ clknet_leaf_4_clk _00675_ net45 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.acc\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10566_ genblk2\[5\].wave_shpr.div.b1\[7\] genblk2\[5\].wave_shpr.div.acc\[7\] vssd1
+ vssd1 vccd1 vccd1 _04794_ sky130_fd_sc_hd__and2b_1
XFILLER_0_11_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_106_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12305_ net397 _06009_ _06010_ net731 vssd1 vssd1 vccd1 vccd1 _01039_ sky130_fd_sc_hd__a22o_1
X_13285_ clknet_leaf_117_clk _00606_ net137 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.fin_quo\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_10497_ _04617_ _04622_ vssd1 vssd1 vccd1 vccd1 _04738_ sky130_fd_sc_hd__nand2b_1
X_12236_ _05810_ genblk2\[11\].wave_shpr.div.acc\[16\] _05973_ vssd1 vssd1 vccd1 vccd1
+ _05974_ sky130_fd_sc_hd__a21o_1
X_12167_ genblk2\[10\].wave_shpr.div.acc\[24\] _05784_ vssd1 vssd1 vccd1 vccd1 _05912_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__07953__B1 _02656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11118_ genblk2\[7\].wave_shpr.div.acc\[4\] genblk2\[7\].wave_shpr.div.b1\[4\] vssd1
+ vssd1 vccd1 vccd1 _05178_ sky130_fd_sc_hd__or2b_1
X_12098_ _05757_ _05860_ vssd1 vssd1 vccd1 vccd1 _05861_ sky130_fd_sc_hd__xnor2_1
X_11049_ _05054_ vssd1 vssd1 vccd1 vccd1 _05126_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__06508__A1 _01201_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput7 pb[1] vssd1 vssd1 vccd1 vccd1 net7 sky130_fd_sc_hd__buf_4
XFILLER_0_79_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09741__S _00009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06590_ _01497_ vssd1 vssd1 vccd1 vccd1 _01498_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_47_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06385__B _01328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08260_ _02965_ _02966_ vssd1 vssd1 vccd1 vccd1 _02967_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_313 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07211_ genblk1\[10\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 _01993_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08191_ _02697_ _02747_ _02896_ vssd1 vssd1 vccd1 vccd1 _02898_ sky130_fd_sc_hd__and3_1
XFILLER_0_27_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07142_ genblk1\[9\].osc.clkdiv_C.cnt\[3\] _01514_ vssd1 vssd1 vccd1 vccd1 _01942_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_30_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07073_ _01862_ _01885_ _01888_ _01889_ vssd1 vssd1 vccd1 vccd1 genblk1\[8\].osc.clkdiv_C.next_cnt\[1\]
+ sky130_fd_sc_hd__o211a_1
XANTENNA__08105__B _01192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10651__A _02183_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07944__B1 _01514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09217__A _03838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07975_ _02681_ vssd1 vssd1 vccd1 vccd1 _02682_ sky130_fd_sc_hd__buf_2
X_09714_ _04163_ _04192_ _04193_ vssd1 vssd1 vccd1 vccd1 _04194_ sky130_fd_sc_hd__a21o_1
X_06926_ _01761_ _01772_ vssd1 vssd1 vccd1 vccd1 genblk1\[6\].osc.clkdiv_C.next_cnt\[7\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09645_ _04007_ _04129_ vssd1 vssd1 vccd1 vccd1 _04136_ sky130_fd_sc_hd__nor2_1
X_06857_ genblk1\[5\].osc.clkdiv_C.cnt\[12\] _01714_ _01716_ vssd1 vssd1 vccd1 vccd1
+ genblk1\[5\].osc.clkdiv_C.next_cnt\[12\] sky130_fd_sc_hd__o21a_1
XTAP_1006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09576_ net829 _04076_ _04080_ _04083_ vssd1 vssd1 vccd1 vccd1 _00237_ sky130_fd_sc_hd__a22o_1
XTAP_1017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06788_ _01179_ _01262_ vssd1 vssd1 vccd1 vccd1 _01660_ sky130_fd_sc_hd__nor2_1
XANTENNA__06576__A _01182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10059__A1 _01263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08527_ _03232_ _03233_ vssd1 vssd1 vccd1 vccd1 _03234_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08458_ _02734_ _02736_ genblk2\[6\].wave_shpr.div.fin_quo\[3\] vssd1 vssd1 vccd1
+ vccd1 _03165_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_53_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07409_ _02149_ _02153_ genblk2\[0\].wave_shpr.div.busy vssd1 vssd1 vccd1 vccd1 _02154_
+ sky130_fd_sc_hd__and3b_1
X_08389_ _03086_ _03095_ genblk1\[2\].osc.clkdiv_C.cnt\[7\] _02011_ vssd1 vssd1 vccd1
+ vccd1 _03096_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_107_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10420_ _03719_ genblk1\[4\].osc.clkdiv_C.cnt\[17\] vssd1 vssd1 vccd1 vccd1 _04680_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_150_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07200__A genblk1\[9\].osc.clkdiv_C.cnt\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10351_ _01355_ vssd1 vssd1 vccd1 vccd1 _04643_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10782__A2 _04880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13070_ clknet_leaf_24_clk _00397_ net92 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.quo\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10282_ genblk2\[4\].wave_shpr.div.b1\[6\] genblk2\[4\].wave_shpr.div.acc\[6\] vssd1
+ vssd1 vccd1 vccd1 _04594_ sky130_fd_sc_hd__and2b_1
X_12021_ genblk2\[10\].wave_shpr.div.quo\[0\] _05813_ _05787_ _05816_ vssd1 vssd1
+ vccd1 vccd1 _00949_ sky130_fd_sc_hd__a22o_1
XANTENNA__07935__B1 _02223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12923_ clknet_leaf_35_clk _00254_ net105 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.acc\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12854_ clknet_leaf_119_clk _00185_ net139 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.fin_quo\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11805_ genblk2\[9\].wave_shpr.div.acc\[2\] _05655_ _05613_ vssd1 vssd1 vccd1 vccd1
+ _05656_ sky130_fd_sc_hd__mux2_1
XTAP_2274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12785_ clknet_leaf_41_clk _00118_ net123 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.b1\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_28_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09797__A _04250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11736_ net1259 genblk2\[9\].wave_shpr.div.quo\[6\] _00023_ vssd1 vssd1 vccd1 vccd1
+ _05621_ sky130_fd_sc_hd__mux2_1
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11667_ genblk2\[9\].wave_shpr.div.acc\[12\] genblk2\[9\].wave_shpr.div.b1\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05559_ sky130_fd_sc_hd__or2b_1
XFILLER_0_142_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13406_ clknet_leaf_90_clk _00725_ net144 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.quo\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10618_ genblk2\[6\].wave_shpr.div.b1\[3\] _01758_ _04834_ vssd1 vssd1 vccd1 vccd1
+ _04835_ sky130_fd_sc_hd__mux2_1
XANTENNA__07218__A2 _01246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11598_ genblk2\[8\].wave_shpr.div.acc\[11\] _05509_ _05493_ vssd1 vssd1 vccd1 vccd1
+ _05510_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06426__B1 _01368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10549_ genblk2\[5\].wave_shpr.div.acc\[4\] genblk2\[5\].wave_shpr.div.b1\[4\] vssd1
+ vssd1 vccd1 vccd1 _04777_ sky130_fd_sc_hd__or2b_1
XFILLER_0_24_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13337_ clknet_leaf_8_clk _00658_ net49 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.acc\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_122_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13268_ clknet_leaf_1_clk _00591_ net44 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.acc\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12219_ genblk2\[11\].wave_shpr.div.b1\[8\] genblk2\[11\].wave_shpr.div.acc\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05957_ sky130_fd_sc_hd__and2b_1
X_13199_ clknet_leaf_114_clk _00522_ net134 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.fin_quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11722__A1 _05613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07760_ _02362_ vssd1 vssd1 vccd1 vccd1 _02467_ sky130_fd_sc_hd__clkbuf_4
X_06711_ genblk1\[4\].osc.clkdiv_C.cnt\[0\] _01600_ vssd1 vssd1 vccd1 vccd1 _01601_
+ sky130_fd_sc_hd__and2b_1
X_07691_ _02373_ _02384_ _02385_ _02397_ vssd1 vssd1 vccd1 vccd1 _02398_ sky130_fd_sc_hd__a211o_1
X_09430_ genblk2\[1\].wave_shpr.div.b1\[12\] genblk2\[1\].wave_shpr.div.acc\[12\]
+ vssd1 vssd1 vccd1 vccd1 _03994_ sky130_fd_sc_hd__and2b_1
X_06642_ _01523_ _01540_ vssd1 vssd1 vccd1 vccd1 _01541_ sky130_fd_sc_hd__nor2_1
XFILLER_0_154_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06396__A _01238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09361_ net653 _03841_ _03910_ _03933_ vssd1 vssd1 vccd1 vccd1 _00172_ sky130_fd_sc_hd__a22o_1
X_06573_ genblk1\[2\].osc.clkdiv_C.cnt\[17\] _01480_ vssd1 vssd1 vccd1 vccd1 _01482_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08312_ _02404_ _02408_ _02406_ vssd1 vssd1 vccd1 vccd1 _03019_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_118_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09292_ _03881_ _03772_ vssd1 vssd1 vccd1 vccd1 _03882_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08243_ _02225_ _02682_ vssd1 vssd1 vccd1 vccd1 _02950_ sky130_fd_sc_hd__nand2_1
XFILLER_0_117_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout131_A net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_55_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08174_ _02873_ _02874_ _02871_ vssd1 vssd1 vccd1 vccd1 _02881_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_144_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07125_ _01924_ vssd1 vssd1 vccd1 vccd1 _01925_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07056_ genblk1\[8\].osc.clkdiv_C.cnt\[3\] _01498_ vssd1 vssd1 vccd1 vccd1 _01874_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__10381__A _04477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07958_ _02655_ _02663_ _02664_ vssd1 vssd1 vccd1 vccd1 _02665_ sky130_fd_sc_hd__a21o_1
XFILLER_0_98_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06909_ genblk1\[6\].osc.clkdiv_C.cnt\[1\] net837 vssd1 vssd1 vccd1 vccd1 _01762_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__11477__B1 _04233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07889_ genblk2\[0\].wave_shpr.div.fin_quo\[6\] _02595_ vssd1 vssd1 vccd1 vccd1 _02596_
+ sky130_fd_sc_hd__xnor2_1
Xmax_cap36 _01423_ vssd1 vssd1 vccd1 vccd1 net36 sky130_fd_sc_hd__clkbuf_2
X_09628_ _04002_ _03955_ vssd1 vssd1 vccd1 vccd1 _04123_ sky130_fd_sc_hd__nor2_1
XANTENNA_fanout44_A net85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09559_ net588 _04046_ vssd1 vssd1 vccd1 vccd1 _04071_ sky130_fd_sc_hd__or2b_1
XFILLER_0_65_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_560 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12570_ clknet_leaf_28_clk genblk1\[1\].osc.clkdiv_C.next_cnt\[9\] net90 vssd1 vssd1
+ vccd1 vccd1 genblk1\[1\].osc.clkdiv_C.cnt\[9\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_66_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09842__B1 _04250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12441__A2 _03947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07999__A3 _01361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11521_ _05450_ genblk1\[8\].osc.clkdiv_C.cnt\[5\] vssd1 vssd1 vccd1 vccd1 _05457_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_108_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11452_ genblk2\[8\].wave_shpr.div.fin_quo\[5\] genblk2\[8\].wave_shpr.div.quo\[4\]
+ _00021_ vssd1 vssd1 vccd1 vccd1 _05423_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10403_ _04058_ _01588_ vssd1 vssd1 vccd1 vccd1 _04670_ sky130_fd_sc_hd__nor2_1
X_11383_ _05243_ genblk2\[8\].wave_shpr.div.acc\[16\] vssd1 vssd1 vccd1 vccd1 _05359_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_21_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_150_279 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13122_ clknet_leaf_136_clk _00447_ net43 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.b1\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10334_ net1212 _01240_ _04440_ vssd1 vssd1 vccd1 vccd1 _04635_ sky130_fd_sc_hd__mux2_1
XANTENNA__07865__A _02216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07620__A2 _01430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13053_ clknet_leaf_113_clk _00380_ net128 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10265_ genblk2\[4\].wave_shpr.div.acc\[5\] genblk2\[4\].wave_shpr.div.b1\[5\] vssd1
+ vssd1 vccd1 vccd1 _04577_ sky130_fd_sc_hd__or2b_1
X_12004_ genblk2\[11\].wave_shpr.div.b1\[11\] _01500_ _05802_ vssd1 vssd1 vccd1 vccd1
+ _05807_ sky130_fd_sc_hd__mux2_1
X_10196_ net862 _04518_ _04522_ _04525_ vssd1 vssd1 vccd1 vccd1 _00415_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08581__B1 _02525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12906_ clknet_leaf_36_clk _00237_ net104 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.acc\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07687__A2 _02011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10140__B1 _04457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2060 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12837_ clknet_leaf_65_clk _00170_ net196 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.acc\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2071 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2082 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2093 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12768_ clknet_leaf_93_clk _00101_ net148 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.fin_quo\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11719_ genblk2\[9\].wave_shpr.div.acc\[23\] genblk2\[9\].wave_shpr.div.acc\[25\]
+ genblk2\[9\].wave_shpr.div.acc\[24\] genblk2\[9\].wave_shpr.div.acc\[26\] vssd1
+ vssd1 vccd1 vccd1 _05611_ sky130_fd_sc_hd__or4_2
XFILLER_0_25_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12699_ clknet_leaf_54_clk genblk1\[8\].osc.clkdiv_C.next_cnt\[12\] net172 vssd1
+ vssd1 vccd1 vccd1 genblk1\[8\].osc.clkdiv_C.cnt\[12\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_116_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xinput10 pb[4] vssd1 vssd1 vccd1 vccd1 net10 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_625 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold805 genblk2\[9\].wave_shpr.div.acc\[19\] vssd1 vssd1 vccd1 vccd1 net1023 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold816 genblk2\[2\].wave_shpr.div.acc\[21\] vssd1 vssd1 vccd1 vccd1 net1034 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09466__S _03822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold827 genblk2\[9\].wave_shpr.div.acc\[25\] vssd1 vssd1 vccd1 vccd1 net1045 sky130_fd_sc_hd__dlygate4sd3_1
Xhold838 genblk2\[5\].wave_shpr.div.quo\[0\] vssd1 vssd1 vccd1 vccd1 net1056 sky130_fd_sc_hd__dlygate4sd3_1
Xhold849 genblk2\[3\].wave_shpr.div.acc\[1\] vssd1 vssd1 vccd1 vccd1 net1067 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07611__A2 _01437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08930_ sig_norm.acc\[10\] _03590_ _03625_ vssd1 vssd1 vccd1 vccd1 _03626_ sky130_fd_sc_hd__a21o_1
XANTENNA__09364__A2 _03841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08861_ _03565_ _03567_ _03519_ _03523_ vssd1 vssd1 vccd1 vccd1 _03568_ sky130_fd_sc_hd__or4_1
X_07812_ _02509_ _02516_ _02518_ vssd1 vssd1 vccd1 vccd1 _02519_ sky130_fd_sc_hd__o21ai_1
X_08792_ _03384_ _03394_ _03393_ vssd1 vssd1 vccd1 vccd1 _03499_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_74_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07743_ _02440_ _02443_ _02449_ vssd1 vssd1 vccd1 vccd1 _02450_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07127__A1 genblk1\[9\].osc.clkdiv_C.cnt\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07674_ _02378_ _02376_ _02380_ _02375_ vssd1 vssd1 vccd1 vccd1 _02381_ sky130_fd_sc_hd__or4b_1
XANTENNA__10131__B1 _04455_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06625_ genblk1\[3\].osc.clkdiv_C.cnt\[3\] _01528_ vssd1 vssd1 vccd1 vccd1 _01530_
+ sky130_fd_sc_hd__and2_1
X_09413_ _03968_ _03975_ _03976_ vssd1 vssd1 vccd1 vccd1 _03977_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06886__B1 _01739_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11760__A _02203_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09344_ genblk2\[0\].wave_shpr.div.acc\[17\] _03921_ _03803_ vssd1 vssd1 vccd1 vccd1
+ _03922_ sky130_fd_sc_hd__mux2_1
X_06556_ _01451_ _01470_ vssd1 vssd1 vccd1 vccd1 _01471_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12890__RESET_B net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09275_ _03804_ _03868_ vssd1 vssd1 vccd1 vccd1 _03869_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06487_ genblk1\[2\].osc.clkdiv_C.cnt\[12\] _01411_ _01412_ _01183_ vssd1 vssd1 vccd1
+ vccd1 _01413_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__07669__B _01440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08226_ _02932_ _02842_ genblk2\[4\].wave_shpr.div.fin_quo\[5\] vssd1 vssd1 vccd1
+ vccd1 _02933_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_133_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_105_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08157_ genblk1\[3\].osc.clkdiv_C.cnt\[14\] _01361_ _02851_ _02863_ vssd1 vssd1 vccd1
+ vccd1 _02864_ sky130_fd_sc_hd__a211o_1
XFILLER_0_16_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07108_ genblk1\[8\].osc.clkdiv_C.cnt\[14\] _01910_ vssd1 vssd1 vccd1 vccd1 _01912_
+ sky130_fd_sc_hd__and2_1
X_08088_ genblk2\[5\].wave_shpr.div.fin_quo\[6\] _02794_ vssd1 vssd1 vccd1 vccd1 _02795_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_101_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07039_ genblk1\[8\].osc.clkdiv_C.cnt\[5\] _01487_ vssd1 vssd1 vccd1 vccd1 _01857_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10050_ net1188 _01248_ _04238_ vssd1 vssd1 vccd1 vccd1 _04434_ sky130_fd_sc_hd__mux2_1
XFILLER_0_97_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10050__S _04238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13740_ clknet_leaf_46_clk _01051_ net121 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.quo\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10952_ _05059_ genblk1\[6\].osc.clkdiv_C.cnt\[1\] vssd1 vssd1 vccd1 vccd1 _05060_
+ sky130_fd_sc_hd__and2_1
X_13671_ clknet_leaf_40_clk _00984_ net118 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.acc\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10883_ _05025_ vssd1 vssd1 vccd1 vccd1 _00602_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12622_ clknet_leaf_17_clk genblk1\[4\].osc.clkdiv_C.next_cnt\[7\] net83 vssd1 vssd1
+ vccd1 vccd1 genblk1\[4\].osc.clkdiv_C.cnt\[7\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_39_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_155_349 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12553_ clknet_leaf_55_clk genblk1\[0\].osc.clkdiv_C.next_cnt\[10\] net176 vssd1
+ vssd1 vccd1 vccd1 genblk1\[0\].osc.clkdiv_C.cnt\[10\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__08094__A2 _01359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11504_ net404 _05442_ _05446_ net676 vssd1 vssd1 vccd1 vccd1 _00802_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12484_ clknet_leaf_107_clk _00046_ net151 vssd1 vssd1 vccd1 vccd1 sig_norm.acc\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09043__A1 _02002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11435_ genblk2\[8\].wave_shpr.div.acc\[21\] _05410_ vssd1 vssd1 vccd1 vccd1 _05411_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_110_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11366_ genblk2\[7\].wave_shpr.div.acc\[25\] _05346_ vssd1 vssd1 vccd1 vccd1 _05348_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_104_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13766__RESET_B net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10317_ _04626_ vssd1 vssd1 vccd1 vccd1 _00435_ sky130_fd_sc_hd__clkbuf_1
X_13105_ clknet_leaf_12_clk _00430_ net52 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.i\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11297_ net893 _05296_ _05222_ vssd1 vssd1 vccd1 vccd1 _05297_ sky130_fd_sc_hd__mux2_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13036_ clknet_leaf_123_clk _00363_ net76 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.b1\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10248_ _00010_ _04560_ net1148 vssd1 vssd1 vccd1 vccd1 _04562_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_119_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10179_ _04399_ _04368_ vssd1 vssd1 vccd1 vccd1 _04512_ sky130_fd_sc_hd__or2b_1
XANTENNA__06580__A2 _01344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10664__B2 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06410_ _01178_ _01176_ freq_div.state\[0\] vssd1 vssd1 vccd1 vccd1 _01354_ sky130_fd_sc_hd__mux2_2
XFILLER_0_29_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07390_ _02139_ vssd1 vssd1 vccd1 vccd1 _02140_ sky130_fd_sc_hd__inv_2
XANTENNA__09806__B1 _04252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09050__A _03708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06341_ genblk1\[0\].osc.clkdiv_C.cnt\[12\] _01290_ vssd1 vssd1 vccd1 vccd1 _01291_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_60_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06393__B _01226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09060_ _03720_ vssd1 vssd1 vccd1 vccd1 _00084_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06272_ _01229_ _01230_ _01233_ vssd1 vssd1 vccd1 vccd1 _01234_ sky130_fd_sc_hd__a21o_2
XFILLER_0_4_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08011_ genblk1\[6\].osc.clkdiv_C.cnt\[5\] _01367_ _01747_ genblk1\[6\].osc.clkdiv_C.cnt\[4\]
+ _02717_ vssd1 vssd1 vccd1 vccd1 _02718_ sky130_fd_sc_hd__a221o_1
XFILLER_0_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold602 genblk2\[3\].wave_shpr.div.quo\[6\] vssd1 vssd1 vccd1 vccd1 net820 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09196__S _03822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold613 PWM.counter\[2\] vssd1 vssd1 vccd1 vccd1 net831 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold624 genblk2\[4\].wave_shpr.div.acc\[4\] vssd1 vssd1 vccd1 vccd1 net842 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_40_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold635 _00749_ vssd1 vssd1 vccd1 vccd1 net853 sky130_fd_sc_hd__dlygate4sd3_1
Xhold646 genblk2\[8\].wave_shpr.div.b1\[0\] vssd1 vssd1 vccd1 vccd1 net864 sky130_fd_sc_hd__dlygate4sd3_1
Xhold657 genblk2\[11\].wave_shpr.div.acc\[12\] vssd1 vssd1 vccd1 vccd1 net875 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_96 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold668 genblk2\[9\].wave_shpr.div.acc\[4\] vssd1 vssd1 vccd1 vccd1 net886 sky130_fd_sc_hd__dlygate4sd3_1
Xhold679 genblk2\[11\].wave_shpr.div.acc\[15\] vssd1 vssd1 vccd1 vccd1 net897 sky130_fd_sc_hd__dlygate4sd3_1
X_09962_ _03690_ _04358_ _04359_ vssd1 vssd1 vccd1 vccd1 _00347_ sky130_fd_sc_hd__nor3_1
X_08913_ sig_norm.acc\[5\] _03611_ vssd1 vssd1 vccd1 vccd1 _03614_ sky130_fd_sc_hd__or2_1
X_09893_ _04192_ _04309_ vssd1 vssd1 vccd1 vccd1 _04310_ sky130_fd_sc_hd__xnor2_1
XTAP_940 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_962 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08844_ _03540_ _03550_ vssd1 vssd1 vccd1 vccd1 _03551_ sky130_fd_sc_hd__nand2_1
XTAP_984 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_995 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08775_ _03465_ _03480_ _03481_ vssd1 vssd1 vccd1 vccd1 _03482_ sky130_fd_sc_hd__nor3_2
XFILLER_0_79_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07726_ _01342_ _01241_ vssd1 vssd1 vccd1 vccd1 _02433_ sky130_fd_sc_hd__nor2_4
XTAP_2829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07657_ net136 vssd1 vssd1 vccd1 vccd1 _02364_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06608_ genblk1\[3\].osc.clkdiv_C.cnt\[9\] _01210_ vssd1 vssd1 vccd1 vccd1 _01516_
+ sky130_fd_sc_hd__xnor2_1
X_07588_ _02284_ _02283_ _02293_ _02294_ _02285_ vssd1 vssd1 vccd1 vccd1 _02295_ sky130_fd_sc_hd__o311a_1
XFILLER_0_137_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_36_826 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09327_ genblk2\[0\].wave_shpr.div.acc\[13\] _03908_ _03889_ vssd1 vssd1 vccd1 vccd1
+ _03909_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06539_ genblk1\[2\].osc.clkdiv_C.cnt\[4\] _01456_ genblk1\[2\].osc.clkdiv_C.cnt\[5\]
+ vssd1 vssd1 vccd1 vccd1 _01460_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_75_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08076__A2 _01678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_106_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09258_ net265 _03845_ _03847_ net636 _03858_ vssd1 vssd1 vccd1 vccd1 _00144_ sky130_fd_sc_hd__a221o_1
XFILLER_0_145_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08209_ _02910_ _02914_ _02915_ vssd1 vssd1 vccd1 vccd1 _02916_ sky130_fd_sc_hd__a21oi_1
X_09189_ _03701_ vssd1 vssd1 vccd1 vccd1 _03822_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_121_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11206__B1_N _03717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11220_ net331 _05246_ _05250_ net693 vssd1 vssd1 vccd1 vccd1 _00714_ sky130_fd_sc_hd__a22o_1
XANTENNA__07036__B1 _01578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11151_ genblk2\[7\].wave_shpr.div.b1\[15\] genblk2\[7\].wave_shpr.div.acc\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05211_ sky130_fd_sc_hd__and2b_1
X_10102_ net525 _04457_ _04454_ net631 _04460_ vssd1 vssd1 vccd1 vccd1 _00386_ sky130_fd_sc_hd__a221o_1
XFILLER_0_101_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11082_ genblk2\[6\].wave_shpr.div.acc\[23\] _05020_ _05149_ vssd1 vssd1 vccd1 vccd1
+ _05150_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10033_ genblk2\[3\].wave_shpr.div.fin_quo\[3\] genblk2\[3\].wave_shpr.div.quo\[2\]
+ _04422_ vssd1 vssd1 vccd1 vccd1 _04426_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11984_ genblk2\[11\].wave_shpr.div.b1\[1\] _03813_ _05433_ vssd1 vssd1 vccd1 vccd1
+ _05797_ sky130_fd_sc_hd__mux2_1
X_13723_ clknet_leaf_96_clk net431 net160 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.quo\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_726 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10935_ _02152_ genblk2\[6\].wave_shpr.div.busy _02186_ vssd1 vssd1 vccd1 vccd1 _05053_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_105_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13654_ clknet_leaf_41_clk _00967_ net116 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.quo\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10866_ genblk2\[6\].wave_shpr.div.b1\[14\] genblk2\[6\].wave_shpr.div.acc\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05010_ sky130_fd_sc_hd__and2b_1
XANTENNA__06494__A _01242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12605_ clknet_leaf_22_clk genblk1\[3\].osc.clkdiv_C.next_cnt\[8\] net94 vssd1 vssd1
+ vccd1 vccd1 genblk1\[3\].osc.clkdiv_C.cnt\[8\] sky130_fd_sc_hd__dfrtp_4
XPHY_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13585_ clknet_leaf_76_clk _00900_ net207 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.acc\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10797_ genblk2\[5\].wave_shpr.div.acc\[23\] _04818_ vssd1 vssd1 vccd1 vccd1 _04949_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_122 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12536_ clknet_leaf_44_clk _00088_ net123 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.b1\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07102__B genblk1\[8\].osc.clkdiv_C.cnt\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12467_ clknet_leaf_33_clk smpl_rt_clkdiv.clkDiv_inst.next_cnt\[1\] net99 vssd1 vssd1
+ vccd1 vccd1 smpl_rt_clkdiv.clkDiv_inst.cnt\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11418_ genblk2\[8\].wave_shpr.div.b1\[10\] genblk2\[8\].wave_shpr.div.acc\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05394_ sky130_fd_sc_hd__and2b_1
X_12398_ genblk2\[11\].wave_shpr.div.acc\[12\] _06070_ _06055_ vssd1 vssd1 vccd1 vccd1
+ _06071_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11349_ genblk2\[7\].wave_shpr.div.acc\[20\] _05334_ vssd1 vssd1 vccd1 vccd1 _05336_
+ sky130_fd_sc_hd__or2_1
XANTENNA__07042__A3 _01855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06250__B2 genblk1\[0\].osc.clkdiv_C.cnt\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13019_ clknet_leaf_123_clk _00346_ net76 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.i\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_06890_ genblk1\[6\].osc.clkdiv_C.cnt\[12\] _01519_ _01739_ genblk1\[6\].osc.clkdiv_C.cnt\[8\]
+ _01743_ vssd1 vssd1 vccd1 vccd1 _01744_ sky130_fd_sc_hd__a221o_1
XANTENNA__06669__A _01349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08560_ genblk2\[8\].wave_shpr.div.fin_quo\[2\] _02362_ _02636_ vssd1 vssd1 vccd1
+ vccd1 _03267_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07511_ _02230_ PWM.final_sample_in\[5\] vssd1 vssd1 vccd1 vccd1 _02231_ sky130_fd_sc_hd__and2_1
XANTENNA__10637__A1 _04223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08491_ _03066_ _03070_ vssd1 vssd1 vccd1 vccd1 _03198_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06305__A2 _01227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_42 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07442_ _02178_ vssd1 vssd1 vccd1 vccd1 _00013_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_76_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07373_ genblk1\[11\].osc.clkdiv_C.cnt\[10\] _02123_ vssd1 vssd1 vccd1 vccd1 _02127_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_128_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08058__A2 _01172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09112_ genblk2\[0\].wave_shpr.div.acc\[3\] genblk2\[0\].wave_shpr.div.b1\[3\] vssd1
+ vssd1 vccd1 vccd1 _03760_ sky130_fd_sc_hd__or2b_1
XANTENNA__10357__C _01367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06324_ _01269_ _01279_ _01280_ vssd1 vssd1 vccd1 vccd1 genblk1\[0\].osc.clkdiv_C.next_cnt\[5\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_72_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09043_ genblk2\[0\].wave_shpr.div.b1\[2\] _02002_ _03708_ vssd1 vssd1 vccd1 vccd1
+ _03710_ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06255_ genblk1\[0\].osc.clkdiv_C.cnt\[0\] _01211_ _01215_ genblk1\[0\].osc.clkdiv_C.cnt\[4\]
+ _01216_ vssd1 vssd1 vccd1 vccd1 _01217_ sky130_fd_sc_hd__a221o_1
XANTENNA__07947__B _01574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold410 genblk2\[7\].wave_shpr.div.acc\[18\] vssd1 vssd1 vccd1 vccd1 net628 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09558__A2 _04042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06186_ _01155_ _01150_ _01156_ vssd1 vssd1 vccd1 vccd1 _01157_ sky130_fd_sc_hd__a21oi_4
Xhold421 genblk2\[2\].wave_shpr.div.quo\[22\] vssd1 vssd1 vccd1 vccd1 net639 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold432 _00867_ vssd1 vssd1 vccd1 vccd1 net650 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07569__A1 genblk1\[9\].osc.clkdiv_C.cnt\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold443 genblk2\[7\].wave_shpr.div.quo\[4\] vssd1 vssd1 vccd1 vccd1 net661 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold454 genblk2\[4\].wave_shpr.div.quo\[10\] vssd1 vssd1 vccd1 vccd1 net672 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold465 _00953_ vssd1 vssd1 vccd1 vccd1 net683 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold476 genblk2\[4\].wave_shpr.div.acc\[20\] vssd1 vssd1 vccd1 vccd1 net694 sky130_fd_sc_hd__dlygate4sd3_1
Xhold487 genblk2\[10\].wave_shpr.div.acc\[20\] vssd1 vssd1 vccd1 vccd1 net705 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06241__A1 _01201_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold498 genblk2\[2\].wave_shpr.div.quo\[5\] vssd1 vssd1 vccd1 vccd1 net716 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09945_ _04346_ _04212_ genblk2\[2\].wave_shpr.div.acc\[24\] vssd1 vssd1 vccd1 vccd1
+ _04348_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09876_ _04184_ _04296_ vssd1 vssd1 vccd1 vccd1 _04297_ sky130_fd_sc_hd__xnor2_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1110 genblk2\[9\].wave_shpr.div.quo\[0\] vssd1 vssd1 vccd1 vccd1 net1328 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06579__A _01172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1121 sig_norm.quo\[4\] vssd1 vssd1 vccd1 vccd1 net1339 sky130_fd_sc_hd__dlygate4sd3_1
X_08827_ genblk2\[2\].wave_shpr.div.fin_quo\[0\] _02592_ _02468_ genblk2\[2\].wave_shpr.div.fin_quo\[1\]
+ _03114_ vssd1 vssd1 vccd1 vccd1 _03534_ sky130_fd_sc_hd__a221o_1
XANTENNA__07741__A1 genblk1\[1\].osc.clkdiv_C.cnt\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07741__B2 genblk1\[1\].osc.clkdiv_C.cnt\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08758_ _03258_ _03452_ _03464_ vssd1 vssd1 vccd1 vccd1 _03465_ sky130_fd_sc_hd__and3_1
XTAP_2626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10628__A1 _01189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07709_ _02415_ vssd1 vssd1 vccd1 vccd1 _02416_ sky130_fd_sc_hd__buf_2
XTAP_1903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08689_ _03366_ _03376_ vssd1 vssd1 vccd1 vccd1 _03396_ sky130_fd_sc_hd__and2b_1
XFILLER_0_67_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10720_ _04786_ _04891_ vssd1 vssd1 vccd1 vccd1 _04892_ sky130_fd_sc_hd__xnor2_1
XTAP_1947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07203__A genblk1\[9\].osc.clkdiv_C.cnt\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10651_ _02183_ vssd1 vssd1 vccd1 vccd1 _04853_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_153_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10582_ genblk2\[5\].wave_shpr.div.b1\[15\] genblk2\[5\].wave_shpr.div.acc\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04810_ sky130_fd_sc_hd__and2b_1
X_13370_ clknet_leaf_116_clk _00689_ net140 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.fin_quo\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_90_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12321_ genblk2\[11\].wave_shpr.div.quo\[14\] _06014_ _06015_ net342 _06018_ vssd1
+ vssd1 vccd1 vccd1 _01047_ sky130_fd_sc_hd__a221o_1
XFILLER_0_133_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12252_ _05986_ vssd1 vssd1 vccd1 vccd1 _01010_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11203_ _03726_ _01869_ _05242_ vssd1 vssd1 vccd1 vccd1 _00705_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_121_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12183_ genblk2\[10\].wave_shpr.div.i\[3\] _02207_ _05920_ vssd1 vssd1 vccd1 vccd1
+ _05923_ sky130_fd_sc_hd__and3_1
XFILLER_0_102_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_61_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11134_ _05175_ _05192_ _05193_ vssd1 vssd1 vccd1 vccd1 _05194_ sky130_fd_sc_hd__a21o_1
XANTENNA__12305__A1 net397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11065_ genblk2\[6\].wave_shpr.div.acc\[25\] genblk2\[6\].wave_shpr.div.acc\[24\]
+ genblk2\[6\].wave_shpr.div.acc\[26\] _05021_ vssd1 vssd1 vccd1 vccd1 _05138_ sky130_fd_sc_hd__nor4_1
X_10016_ _04362_ _04410_ _04411_ vssd1 vssd1 vccd1 vccd1 _04412_ sky130_fd_sc_hd__o21bai_1
XANTENNA_clkbuf_leaf_76_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12069__B1 _05815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11967_ _05788_ vssd1 vssd1 vccd1 vccd1 _00923_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10095__A2 _04452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13706_ clknet_leaf_37_clk _01017_ net114 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.b1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10918_ net1253 net34 _05042_ vssd1 vssd1 vccd1 vccd1 _05044_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11898_ genblk2\[0\].wave_shpr.div.i\[1\] genblk2\[0\].wave_shpr.div.i\[0\] vssd1
+ vssd1 vccd1 vccd1 _05724_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_134_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13637_ clknet_leaf_93_clk _00950_ net159 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.quo\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10849_ _04978_ _04991_ _04992_ vssd1 vssd1 vccd1 vccd1 _04993_ sky130_fd_sc_hd__a21o_1
XFILLER_0_143_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09739__S _00009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_14_clk_A clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13568_ clknet_leaf_55_clk _00883_ net176 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.quo\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_143_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07799__A1 genblk1\[0\].osc.clkdiv_C.cnt\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12519_ clknet_leaf_104_clk PWM.next_counter\[3\] net157 vssd1 vssd1 vccd1 vccd1
+ PWM.counter\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_140_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13499_ clknet_leaf_86_clk _00816_ net179 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.quo\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_29_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout208 net209 vssd1 vssd1 vccd1 vccd1 net208 sky130_fd_sc_hd__clkbuf_4
X_07991_ _02604_ _02645_ _02648_ _02696_ vssd1 vssd1 vccd1 vccd1 _02698_ sky130_fd_sc_hd__a22o_1
XANTENNA__07971__A1 _01201_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_7_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_7_0_clk sky130_fd_sc_hd__clkbuf_8
X_09730_ genblk2\[2\].wave_shpr.div.acc\[19\] _04209_ vssd1 vssd1 vccd1 vccd1 _04210_
+ sky130_fd_sc_hd__or2_1
X_06942_ genblk1\[6\].osc.clkdiv_C.cnt\[13\] genblk1\[6\].osc.clkdiv_C.cnt\[12\] _01779_
+ vssd1 vssd1 vccd1 vccd1 _01783_ sky130_fd_sc_hd__and3_1
X_09661_ net1107 _04048_ _04045_ _04146_ vssd1 vssd1 vccd1 vccd1 _00259_ sky130_fd_sc_hd__a22o_1
X_06873_ genblk1\[6\].osc.clkdiv_C.cnt\[10\] _01726_ genblk1\[6\].osc.clkdiv_C.cnt\[14\]
+ vssd1 vssd1 vccd1 vccd1 _01727_ sky130_fd_sc_hd__o21bai_1
X_08612_ genblk2\[5\].wave_shpr.div.fin_quo\[2\] _02521_ _02791_ vssd1 vssd1 vccd1
+ vccd1 _03319_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12663__RESET_B net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09592_ genblk2\[1\].wave_shpr.div.acc\[7\] _04094_ _04095_ vssd1 vssd1 vccd1 vccd1
+ _04096_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08543_ _02225_ _02682_ _03249_ vssd1 vssd1 vccd1 vccd1 _03250_ sky130_fd_sc_hd__a21o_1
XANTENNA__10649__A _02171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_70 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08474_ genblk2\[5\].wave_shpr.div.fin_quo\[4\] _02308_ _02791_ vssd1 vssd1 vccd1
+ vccd1 _03181_ sky130_fd_sc_hd__a21o_1
XFILLER_0_65_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_612 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07425_ _02165_ vssd1 vssd1 vccd1 vccd1 _00009_ sky130_fd_sc_hd__buf_4
XFILLER_0_9_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_9_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07356_ genblk1\[11\].osc.clkdiv_C.cnt\[6\] _02108_ vssd1 vssd1 vccd1 vccd1 _02114_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_33_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06307_ _01268_ vssd1 vssd1 vccd1 vccd1 _01269_ sky130_fd_sc_hd__clkbuf_4
X_07287_ genblk1\[10\].osc.clkdiv_C.cnt\[13\] _02053_ _02055_ vssd1 vssd1 vccd1 vccd1
+ genblk1\[10\].osc.clkdiv_C.next_cnt\[13\] sky130_fd_sc_hd__o21a_1
XFILLER_0_33_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09026_ genblk2\[9\].wave_shpr.div.i\[1\] genblk2\[9\].wave_shpr.div.i\[0\] genblk2\[9\].wave_shpr.div.i\[2\]
+ genblk2\[9\].wave_shpr.div.i\[3\] vssd1 vssd1 vccd1 vccd1 _03697_ sky130_fd_sc_hd__a31o_1
X_06238_ _01181_ vssd1 vssd1 vccd1 vccd1 _01200_ sky130_fd_sc_hd__buf_6
XFILLER_0_32_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_862 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06169_ _01129_ _01140_ vssd1 vssd1 vccd1 vccd1 _01141_ sky130_fd_sc_hd__nor2_1
Xhold240 _00305_ vssd1 vssd1 vccd1 vccd1 net458 sky130_fd_sc_hd__dlygate4sd3_1
Xhold251 genblk2\[8\].wave_shpr.div.quo\[10\] vssd1 vssd1 vccd1 vccd1 net469 sky130_fd_sc_hd__dlygate4sd3_1
Xhold262 genblk2\[2\].wave_shpr.div.quo\[14\] vssd1 vssd1 vccd1 vccd1 net480 sky130_fd_sc_hd__dlygate4sd3_1
Xhold273 _00399_ vssd1 vssd1 vccd1 vccd1 net491 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_388 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold284 genblk2\[8\].wave_shpr.div.quo\[16\] vssd1 vssd1 vccd1 vccd1 net502 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_580 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold295 genblk2\[9\].wave_shpr.div.quo\[18\] vssd1 vssd1 vccd1 vccd1 net513 sky130_fd_sc_hd__dlygate4sd3_1
X_09928_ _04208_ net22 genblk2\[2\].wave_shpr.div.acc\[18\] vssd1 vssd1 vccd1 vccd1
+ _04337_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12299__B1 _06010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout74_A net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07562__A2_N _01799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09859_ _04176_ _04283_ vssd1 vssd1 vccd1 vccd1 _04284_ sky130_fd_sc_hd__xnor2_1
X_12870_ clknet_leaf_134_clk _00201_ net59 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.b1\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11821_ net984 _05652_ _05653_ _05667_ vssd1 vssd1 vccd1 vccd1 _00898_ sky130_fd_sc_hd__a22o_1
XTAP_2434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11752_ genblk2\[9\].wave_shpr.div.quo\[7\] _05623_ _05624_ net267 vssd1 vssd1 vccd1
+ vccd1 _00872_ sky130_fd_sc_hd__a22o_1
XTAP_1744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10703_ genblk2\[5\].wave_shpr.div.acc_next\[0\] _04856_ vssd1 vssd1 vccd1 vccd1
+ _04879_ sky130_fd_sc_hd__or2b_1
XTAP_1777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11683_ genblk2\[9\].wave_shpr.div.b1\[0\] _05573_ _05574_ vssd1 vssd1 vccd1 vccd1
+ _05575_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_138_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13422_ clknet_leaf_92_clk _00741_ net149 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.acc\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10634_ _01742_ vssd1 vssd1 vccd1 vccd1 _04844_ sky130_fd_sc_hd__inv_2
XFILLER_0_11_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13353_ clknet_leaf_4_clk _00674_ net45 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.acc\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10565_ _04774_ _04791_ _04792_ vssd1 vssd1 vccd1 vccd1 _04793_ sky130_fd_sc_hd__a21o_1
XFILLER_0_106_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12304_ net731 _06009_ _06010_ net767 vssd1 vssd1 vccd1 vccd1 _01038_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13284_ clknet_leaf_117_clk _00605_ net137 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.fin_quo\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_10496_ net1074 _04715_ _04722_ _04737_ vssd1 vssd1 vccd1 vccd1 _00503_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12235_ _05926_ _05972_ vssd1 vssd1 vccd1 vccd1 _05973_ sky130_fd_sc_hd__and2b_1
X_12166_ _05816_ _05910_ _05911_ _05818_ net536 vssd1 vssd1 vccd1 vccd1 _00999_ sky130_fd_sc_hd__a32o_1
X_11117_ genblk2\[7\].wave_shpr.div.b1\[4\] genblk2\[7\].wave_shpr.div.acc\[4\] vssd1
+ vssd1 vccd1 vccd1 _05177_ sky130_fd_sc_hd__or2b_1
X_12097_ genblk2\[10\].wave_shpr.div.b1\[6\] genblk2\[10\].wave_shpr.div.acc\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05860_ sky130_fd_sc_hd__xor2_1
XANTENNA__12014__A _02171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07108__A genblk1\[8\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11048_ net921 _05119_ _05093_ _05125_ vssd1 vssd1 vccd1 vccd1 _00667_ sky130_fd_sc_hd__a22o_1
Xinput8 pb[2] vssd1 vssd1 vccd1 vccd1 net8 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_127_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12999_ clknet_leaf_132_clk _00328_ net60 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.acc\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_98_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11265__A1 _03819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09469__S _03822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07210_ _01359_ _01224_ _01241_ vssd1 vssd1 vccd1 vccd1 _01992_ sky130_fd_sc_hd__a21o_1
XFILLER_0_144_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08190_ _02697_ _02747_ _02896_ vssd1 vssd1 vccd1 vccd1 _02897_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_859 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07141_ _01935_ _01939_ _01940_ vssd1 vssd1 vccd1 vccd1 _01941_ sky130_fd_sc_hd__and3_1
XFILLER_0_54_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07072_ genblk1\[8\].osc.clkdiv_C.cnt\[1\] genblk1\[8\].osc.clkdiv_C.cnt\[0\] vssd1
+ vssd1 vccd1 vccd1 _01889_ sky130_fd_sc_hd__nand2_2
XFILLER_0_140_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08105__C _01208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__12844__RESET_B net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10143__S _04420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07974_ _02676_ _02679_ _02680_ vssd1 vssd1 vccd1 vccd1 _02681_ sky130_fd_sc_hd__o21ai_2
X_09713_ genblk2\[2\].wave_shpr.div.b1\[10\] genblk2\[2\].wave_shpr.div.acc\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04193_ sky130_fd_sc_hd__and2b_1
X_06925_ genblk1\[6\].osc.clkdiv_C.cnt\[7\] _01770_ vssd1 vssd1 vccd1 vccd1 _01772_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_93_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09644_ net874 _04109_ _04113_ _04135_ vssd1 vssd1 vccd1 vccd1 _00253_ sky130_fd_sc_hd__a22o_1
XFILLER_0_93_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06856_ _01693_ _01715_ vssd1 vssd1 vccd1 vccd1 _01716_ sky130_fd_sc_hd__nor2_1
XANTENNA__10700__B1 _04856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09575_ genblk2\[1\].wave_shpr.div.acc\[3\] _04082_ _04011_ vssd1 vssd1 vccd1 vccd1
+ _04083_ sky130_fd_sc_hd__mux2_1
XTAP_1007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06787_ genblk1\[5\].osc.clkdiv_C.cnt\[10\] _01658_ vssd1 vssd1 vccd1 vccd1 _01659_
+ sky130_fd_sc_hd__xor2_1
XTAP_1018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06576__B _01302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08526_ _03227_ _03229_ vssd1 vssd1 vccd1 vccd1 _03233_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08457_ _02648_ _03162_ _03158_ vssd1 vssd1 vccd1 vccd1 _03164_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_147_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_857 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_740 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13632__RESET_B net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07408_ _02152_ vssd1 vssd1 vccd1 vccd1 _02153_ sky130_fd_sc_hd__buf_6
XFILLER_0_80_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08388_ _03090_ _03092_ _03094_ vssd1 vssd1 vccd1 vccd1 _03095_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_61_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07339_ _02100_ vssd1 vssd1 vccd1 vccd1 genblk1\[11\].osc.clkdiv_C.next_cnt\[2\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_103_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07200__B genblk1\[9\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10350_ _04642_ vssd1 vssd1 vccd1 vccd1 _00452_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_60_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_670 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06986__A2 _01227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09009_ _03684_ vssd1 vssd1 vccd1 vccd1 _00069_ sky130_fd_sc_hd__clkbuf_1
X_10281_ _04577_ _04591_ _04592_ vssd1 vssd1 vccd1 vccd1 _04593_ sky130_fd_sc_hd__a21o_1
XFILLER_0_130_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12020_ _05815_ vssd1 vssd1 vccd1 vccd1 _05816_ sky130_fd_sc_hd__buf_4
X_12922_ clknet_leaf_35_clk _00253_ net105 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.acc\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_12853_ clknet_leaf_119_clk _00184_ net139 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.fin_quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11804_ _05576_ _05654_ vssd1 vssd1 vccd1 vccd1 _05655_ sky130_fd_sc_hd__xnor2_1
XTAP_2264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12784_ clknet_leaf_40_clk _00117_ net123 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.b1\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08982__A _01097_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11735_ _05620_ vssd1 vssd1 vccd1 vccd1 _00859_ sky130_fd_sc_hd__clkbuf_1
XTAP_1574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08663__A2 _02521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09289__S _03804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11666_ genblk2\[9\].wave_shpr.div.acc\[13\] genblk2\[9\].wave_shpr.div.b1\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05558_ sky130_fd_sc_hd__or2b_1
X_13405_ clknet_leaf_90_clk _00724_ net143 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.quo\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_592 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10617_ _03701_ vssd1 vssd1 vccd1 vccd1 _04834_ sky130_fd_sc_hd__buf_4
XFILLER_0_3_306 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11597_ _05395_ _05508_ vssd1 vssd1 vccd1 vccd1 _05509_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06426__A1 _01197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13336_ clknet_leaf_6_clk _00657_ net48 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.acc\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06426__B2 genblk1\[1\].osc.clkdiv_C.cnt\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10548_ genblk2\[5\].wave_shpr.div.b1\[4\] genblk2\[5\].wave_shpr.div.acc\[4\] vssd1
+ vssd1 vccd1 vccd1 _04776_ sky130_fd_sc_hd__or2b_1
XFILLER_0_122_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13267_ clknet_leaf_1_clk _00590_ net38 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.acc\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10479_ genblk2\[4\].wave_shpr.div.acc\[13\] _04724_ _04704_ vssd1 vssd1 vccd1 vccd1
+ _04725_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12218_ _05935_ _05954_ _05955_ vssd1 vssd1 vccd1 vccd1 _05956_ sky130_fd_sc_hd__a21o_1
X_13198_ clknet_leaf_114_clk _00521_ net134 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.fin_quo\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_12149_ _05782_ _05899_ vssd1 vssd1 vccd1 vccd1 _05900_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10930__B1 _03736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09752__S _04039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06710_ _01599_ vssd1 vssd1 vccd1 vccd1 _01600_ sky130_fd_sc_hd__buf_2
XFILLER_0_79_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11486__A1 _03831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07690_ _02003_ _01991_ _02393_ _02396_ vssd1 vssd1 vccd1 vccd1 _02397_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_79_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06641_ genblk1\[3\].osc.clkdiv_C.cnt\[9\] _01538_ vssd1 vssd1 vccd1 vccd1 _01540_
+ sky130_fd_sc_hd__and2_1
XANTENNA__06396__B _01262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09360_ genblk2\[0\].wave_shpr.div.acc\[22\] _03931_ vssd1 vssd1 vccd1 vccd1 _03933_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06572_ genblk1\[2\].osc.clkdiv_C.cnt\[16\] _01478_ _01481_ vssd1 vssd1 vccd1 vccd1
+ genblk1\[2\].osc.clkdiv_C.next_cnt\[16\] sky130_fd_sc_hd__o21a_1
XFILLER_0_87_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08311_ _02366_ _03017_ vssd1 vssd1 vccd1 vccd1 _03018_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09291_ _03773_ _03758_ vssd1 vssd1 vccd1 vccd1 _03881_ sky130_fd_sc_hd__or2b_1
XANTENNA__09199__S _03822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_879 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08242_ genblk2\[7\].wave_shpr.div.fin_quo\[6\] _02309_ vssd1 vssd1 vccd1 vccd1 _02949_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__07862__B1 _02361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08173_ _01486_ _01858_ vssd1 vssd1 vccd1 vccd1 _02880_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07124_ _01336_ _01355_ vssd1 vssd1 vccd1 vccd1 _01924_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_42_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06968__A2 _01801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07055_ genblk1\[8\].osc.clkdiv_C.cnt\[8\] _01430_ vssd1 vssd1 vccd1 vccd1 _01873_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_112_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07917__A1 genblk1\[8\].osc.clkdiv_C.cnt\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06601__A2_N _01507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07957_ genblk1\[7\].osc.clkdiv_C.cnt\[8\] _01920_ _01947_ genblk1\[7\].osc.clkdiv_C.cnt\[7\]
+ vssd1 vssd1 vccd1 vccd1 _02664_ sky130_fd_sc_hd__a22o_1
XANTENNA__11493__A _02152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06908_ net837 _01761_ vssd1 vssd1 vccd1 vccd1 genblk1\[6\].osc.clkdiv_C.next_cnt\[0\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__11477__A1 _03704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07888_ _02513_ genblk2\[0\].wave_shpr.div.fin_quo\[5\] _02510_ vssd1 vssd1 vccd1
+ vccd1 _02595_ sky130_fd_sc_hd__or3b_1
Xmax_cap26 _03602_ vssd1 vssd1 vccd1 vccd1 net26 sky130_fd_sc_hd__buf_1
XANTENNA__07145__A2 _01514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap37 _01320_ vssd1 vssd1 vccd1 vccd1 net37 sky130_fd_sc_hd__buf_4
X_09627_ net774 _04109_ _04113_ _04122_ vssd1 vssd1 vccd1 vccd1 _00249_ sky130_fd_sc_hd__a22o_1
X_06839_ genblk1\[5\].osc.clkdiv_C.cnt\[6\] _01703_ vssd1 vssd1 vccd1 vccd1 _01705_
+ sky130_fd_sc_hd__and2_1
X_09558_ net588 _04042_ _04046_ genblk2\[1\].wave_shpr.div.quo\[24\] _04070_ vssd1
+ vssd1 vccd1 vccd1 _00232_ sky130_fd_sc_hd__a221o_1
XFILLER_0_155_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08509_ _03208_ _03215_ vssd1 vssd1 vccd1 vccd1 _03216_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_136_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09489_ _01420_ vssd1 vssd1 vccd1 vccd1 _04034_ sky130_fd_sc_hd__inv_2
XFILLER_0_148_572 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_65_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11520_ net312 _05454_ _05449_ net482 _05456_ vssd1 vssd1 vccd1 vccd1 _00808_ sky130_fd_sc_hd__a221o_1
XFILLER_0_135_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11451_ _05422_ vssd1 vssd1 vccd1 vccd1 _00773_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10048__S _04238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10402_ net255 _04661_ _04663_ net531 _04669_ vssd1 vssd1 vccd1 vccd1 _00477_ sky130_fd_sc_hd__a221o_1
XFILLER_0_61_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11382_ genblk2\[8\].wave_shpr.div.acc\[17\] genblk2\[8\].wave_shpr.div.b1\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05358_ sky130_fd_sc_hd__or2b_1
XFILLER_0_150_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13121_ clknet_leaf_136_clk _00446_ net43 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.b1\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10333_ _03714_ net692 _01262_ _03705_ vssd1 vssd1 vccd1 vccd1 _00443_ sky130_fd_sc_hd__o22a_1
XANTENNA__12263__S _05802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13052_ clknet_leaf_113_clk net780 net131 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.quo\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10264_ genblk2\[4\].wave_shpr.div.acc\[6\] genblk2\[4\].wave_shpr.div.b1\[6\] vssd1
+ vssd1 vccd1 vccd1 _04576_ sky130_fd_sc_hd__or2b_1
XANTENNA__12762__SET_B net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12003_ _05806_ vssd1 vssd1 vccd1 vccd1 _00941_ sky130_fd_sc_hd__clkbuf_1
X_10195_ genblk2\[3\].wave_shpr.div.acc\[13\] _04524_ _04507_ vssd1 vssd1 vccd1 vccd1
+ _04525_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11468__A1 _01811_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12905_ clknet_leaf_37_clk _00236_ net104 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.acc\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10140__A1 _04454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12836_ clknet_leaf_64_clk _00169_ net196 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.acc\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07105__B genblk1\[8\].osc.clkdiv_C.cnt\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2050 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2061 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2072 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2083 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_output18_A net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2094 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12767_ clknet_leaf_93_clk _00100_ net148 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.fin_quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11718_ genblk2\[9\].wave_shpr.div.acc\[22\] _05609_ vssd1 vssd1 vccd1 vccd1 _05610_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_126_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12698_ clknet_leaf_54_clk genblk1\[8\].osc.clkdiv_C.next_cnt\[11\] net172 vssd1
+ vssd1 vccd1 vccd1 genblk1\[8\].osc.clkdiv_C.cnt\[11\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_127_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11649_ _05545_ vssd1 vssd1 vccd1 vccd1 _00848_ sky130_fd_sc_hd__clkbuf_1
Xinput11 pb[5] vssd1 vssd1 vccd1 vccd1 net11 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_142_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09747__S _00009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_52_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold806 genblk2\[4\].wave_shpr.div.acc\[10\] vssd1 vssd1 vccd1 vccd1 net1024 sky130_fd_sc_hd__dlygate4sd3_1
Xhold817 genblk2\[10\].wave_shpr.div.acc\[9\] vssd1 vssd1 vccd1 vccd1 net1035 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13319_ clknet_leaf_26_clk net621 net87 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.quo\[13\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold828 genblk2\[9\].wave_shpr.div.acc\[12\] vssd1 vssd1 vccd1 vccd1 net1046 sky130_fd_sc_hd__dlygate4sd3_1
Xhold839 genblk2\[3\].wave_shpr.div.acc\[3\] vssd1 vssd1 vccd1 vccd1 net1057 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_150_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08860_ _03507_ _03451_ _03506_ _03566_ vssd1 vssd1 vccd1 vccd1 _03567_ sky130_fd_sc_hd__or4_1
X_07811_ _02517_ vssd1 vssd1 vccd1 vccd1 _02518_ sky130_fd_sc_hd__buf_2
XANTENNA__08572__B2 _02362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08791_ _03484_ _03485_ _03497_ vssd1 vssd1 vccd1 vccd1 _03498_ sky130_fd_sc_hd__nor3b_2
X_07742_ _02445_ _02446_ _02447_ _02448_ vssd1 vssd1 vccd1 vccd1 _02449_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_74_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09521__B1 _04045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07673_ genblk1\[10\].osc.clkdiv_C.cnt\[0\] _02001_ _02379_ _02013_ genblk1\[10\].osc.clkdiv_C.cnt\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02380_ sky130_fd_sc_hd__a32o_1
XANTENNA__13295__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09412_ genblk2\[1\].wave_shpr.div.b1\[3\] genblk2\[1\].wave_shpr.div.acc\[3\] vssd1
+ vssd1 vccd1 vccd1 _03976_ sky130_fd_sc_hd__and2b_1
X_06624_ _01523_ _01528_ _01529_ vssd1 vssd1 vccd1 vccd1 genblk1\[3\].osc.clkdiv_C.next_cnt\[2\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_48_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09343_ _03796_ _03920_ vssd1 vssd1 vccd1 vccd1 _03921_ sky130_fd_sc_hd__xnor2_1
X_06555_ genblk1\[2\].osc.clkdiv_C.cnt\[11\] _01468_ vssd1 vssd1 vccd1 vccd1 _01470_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_118_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09274_ _03764_ _03765_ vssd1 vssd1 vccd1 vccd1 _03868_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_145_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06486_ genblk1\[2\].osc.clkdiv_C.cnt\[8\] vssd1 vssd1 vccd1 vccd1 _01412_ sky130_fd_sc_hd__inv_2
XFILLER_0_118_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_56_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08225_ _02837_ vssd1 vssd1 vccd1 vccd1 _02932_ sky130_fd_sc_hd__buf_2
XFILLER_0_118_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_486 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08156_ genblk1\[3\].osc.clkdiv_C.cnt\[14\] _01361_ _01576_ genblk1\[3\].osc.clkdiv_C.cnt\[15\]
+ vssd1 vssd1 vccd1 vccd1 _02863_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_31_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07063__A1 _01441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07107_ net1182 _01908_ _01911_ vssd1 vssd1 vccd1 vccd1 genblk1\[8\].osc.clkdiv_C.next_cnt\[13\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_141_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08087_ genblk2\[5\].wave_shpr.div.fin_quo\[5\] _02789_ _02793_ vssd1 vssd1 vccd1
+ vccd1 _02794_ sky130_fd_sc_hd__or3b_1
XFILLER_0_30_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07038_ _01436_ _01855_ genblk1\[8\].osc.clkdiv_C.cnt\[1\] vssd1 vssd1 vccd1 vccd1
+ _01856_ sky130_fd_sc_hd__a21oi_1
X_08989_ sig_norm.quo\[9\] _03672_ _01155_ vssd1 vssd1 vccd1 vccd1 _03673_ sky130_fd_sc_hd__mux2_1
XANTENNA__10370__B2 _04655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10331__S _03689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09512__B1 _04047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10951_ _04268_ vssd1 vssd1 vccd1 vccd1 _05059_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_98_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08866__A2 _02248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13670_ clknet_leaf_40_clk _00983_ net117 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.acc\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10882_ genblk2\[6\].wave_shpr.div.fin_quo\[1\] genblk2\[6\].wave_shpr.div.quo\[0\]
+ _00017_ vssd1 vssd1 vccd1 vccd1 _05025_ sky130_fd_sc_hd__mux2_1
X_12621_ clknet_leaf_17_clk genblk1\[4\].osc.clkdiv_C.next_cnt\[6\] net80 vssd1 vssd1
+ vccd1 vccd1 genblk1\[4\].osc.clkdiv_C.cnt\[6\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_78_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12552_ clknet_leaf_60_clk genblk1\[0\].osc.clkdiv_C.next_cnt\[9\] net186 vssd1 vssd1
+ vccd1 vccd1 genblk1\[0\].osc.clkdiv_C.cnt\[9\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_65_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08037__A _02364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11503_ net676 _05442_ _05446_ net751 vssd1 vssd1 vccd1 vccd1 _00801_ sky130_fd_sc_hd__a22o_1
XFILLER_0_124_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12483_ clknet_leaf_108_clk _00045_ net151 vssd1 vssd1 vccd1 vccd1 sig_norm.acc\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11434_ genblk2\[8\].wave_shpr.div.acc\[20\] genblk2\[8\].wave_shpr.div.acc\[18\]
+ genblk2\[8\].wave_shpr.div.acc\[19\] _05409_ vssd1 vssd1 vccd1 vccd1 _05410_ sky130_fd_sc_hd__or4_1
XANTENNA__07054__A1 genblk1\[8\].osc.clkdiv_C.cnt\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_100_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_100_clk
+ sky130_fd_sc_hd__clkbuf_16
X_11365_ net1053 _05251_ _05248_ _05347_ vssd1 vssd1 vccd1 vccd1 _00762_ sky130_fd_sc_hd__a22o_1
X_13104_ clknet_leaf_13_clk _00429_ net52 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.i\[1\]
+ sky130_fd_sc_hd__dfrtp_2
X_10316_ genblk2\[4\].wave_shpr.div.fin_quo\[2\] genblk2\[4\].wave_shpr.div.quo\[1\]
+ _00013_ vssd1 vssd1 vccd1 vccd1 _04626_ sky130_fd_sc_hd__mux2_1
XFILLER_0_21_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06801__B2 _01436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11296_ _05194_ _05295_ vssd1 vssd1 vccd1 vccd1 _05296_ sky130_fd_sc_hd__xnor2_1
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_119_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13035_ clknet_leaf_122_clk _00362_ net76 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.b1\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10247_ _04454_ _04559_ _04561_ _04457_ net725 vssd1 vssd1 vccd1 vccd1 _00430_ sky130_fd_sc_hd__a32o_1
X_10178_ net790 _04486_ _04490_ _04511_ vssd1 vssd1 vccd1 vccd1 _00411_ sky130_fd_sc_hd__a22o_1
XANTENNA__12022__A _05815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09503__B1 _03736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10664__A2 _04853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12819_ clknet_leaf_66_clk _00152_ net196 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.acc\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08609__A2 _02789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_816 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10416__A2 _04651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06340_ _01269_ _01289_ _01290_ vssd1 vssd1 vccd1 vccd1 genblk1\[0\].osc.clkdiv_C.next_cnt\[11\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_151_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12688__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06271_ _01232_ vssd1 vssd1 vccd1 vccd1 _01233_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_60_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12169__A2 _05818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08010_ genblk1\[6\].osc.clkdiv_C.cnt\[5\] _01365_ genblk1\[6\].osc.clkdiv_C.cnt\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02717_ sky130_fd_sc_hd__o21a_1
XFILLER_0_115_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_4_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_4_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold603 genblk2\[0\].wave_shpr.div.acc\[26\] vssd1 vssd1 vccd1 vccd1 net821 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold614 _01160_ vssd1 vssd1 vccd1 vccd1 net832 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold625 _00489_ vssd1 vssd1 vccd1 vccd1 net843 sky130_fd_sc_hd__dlygate4sd3_1
Xhold636 genblk2\[0\].wave_shpr.div.acc\[3\] vssd1 vssd1 vccd1 vccd1 net854 sky130_fd_sc_hd__dlygate4sd3_1
Xhold647 genblk2\[1\].wave_shpr.div.acc\[13\] vssd1 vssd1 vccd1 vccd1 net865 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11101__A _03690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold658 genblk2\[11\].wave_shpr.div.acc\[8\] vssd1 vssd1 vccd1 vccd1 net876 sky130_fd_sc_hd__dlygate4sd3_1
X_09961_ genblk2\[2\].wave_shpr.div.i\[3\] _02163_ _04356_ vssd1 vssd1 vccd1 vccd1
+ _04359_ sky130_fd_sc_hd__and3_1
Xhold669 genblk2\[2\].wave_shpr.div.acc\[6\] vssd1 vssd1 vccd1 vccd1 net887 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_100_94 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08912_ net1027 _02260_ _03613_ _03574_ vssd1 vssd1 vccd1 vccd1 _00043_ sky130_fd_sc_hd__a22o_1
XFILLER_0_0_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_110_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09892_ _04193_ _04163_ vssd1 vssd1 vccd1 vccd1 _04309_ sky130_fd_sc_hd__or2b_1
XTAP_930 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_952 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12341__A2 _03942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08843_ _03529_ _03547_ _03549_ vssd1 vssd1 vccd1 vccd1 _03550_ sky130_fd_sc_hd__and3_1
XTAP_963 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09506__A _02170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_974 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout191_A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_985 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10352__A1 _04643_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_996 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08774_ _03258_ _03452_ _03464_ vssd1 vssd1 vccd1 vccd1 _03481_ sky130_fd_sc_hd__a21oi_1
XTAP_2808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07725_ genblk1\[1\].osc.clkdiv_C.cnt\[4\] _01305_ _01313_ genblk1\[1\].osc.clkdiv_C.cnt\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02432_ sky130_fd_sc_hd__a22o_1
XTAP_2819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_149_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07656_ genblk2\[11\].wave_shpr.div.fin_quo\[7\] _02362_ vssd1 vssd1 vccd1 vccd1
+ _02363_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_138_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06607_ genblk1\[3\].osc.clkdiv_C.cnt\[3\] _01513_ _01514_ genblk1\[3\].osc.clkdiv_C.cnt\[4\]
+ vssd1 vssd1 vccd1 vccd1 _01515_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__12078__S _05787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10387__A _04651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07587_ genblk1\[9\].osc.clkdiv_C.cnt\[7\] _01234_ _01513_ genblk1\[9\].osc.clkdiv_C.cnt\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02294_ sky130_fd_sc_hd__a211o_1
XFILLER_0_36_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_48_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09326_ _03788_ _03907_ vssd1 vssd1 vccd1 vccd1 _03908_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06538_ genblk1\[2\].osc.clkdiv_C.cnt\[5\] genblk1\[2\].osc.clkdiv_C.cnt\[4\] _01456_
+ vssd1 vssd1 vccd1 vccd1 _01459_ sky130_fd_sc_hd__and3_1
XANTENNA__07808__B1 _02224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_36_838 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11080__A2 _05057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09257_ _03853_ genblk1\[0\].osc.clkdiv_C.cnt\[12\] vssd1 vssd1 vccd1 vccd1 _03858_
+ sky130_fd_sc_hd__and2_1
X_06469_ genblk1\[1\].osc.clkdiv_C.cnt\[12\] _01398_ _01400_ vssd1 vssd1 vccd1 vccd1
+ genblk1\[1\].osc.clkdiv_C.next_cnt\[12\] sky130_fd_sc_hd__o21a_1
XFILLER_0_133_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08208_ _02901_ _02419_ _02905_ _02909_ vssd1 vssd1 vccd1 vccd1 _02915_ sky130_fd_sc_hd__and4_1
XFILLER_0_105_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09188_ _03714_ _03821_ _03705_ vssd1 vssd1 vccd1 vccd1 _00111_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11368__A0 _05249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09025__A2 _03694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07036__A1 genblk1\[8\].osc.clkdiv_C.cnt\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08139_ net10 _02364_ _02365_ vssd1 vssd1 vccd1 vccd1 _02846_ sky130_fd_sc_hd__and3_2
XFILLER_0_121_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07587__A2 _01234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11150_ _05167_ _05208_ _05209_ vssd1 vssd1 vccd1 vccd1 _05210_ sky130_fd_sc_hd__a21o_1
X_10101_ _04269_ genblk1\[3\].osc.clkdiv_C.cnt\[2\] vssd1 vssd1 vccd1 vccd1 _04460_
+ sky130_fd_sc_hd__and2_1
X_11081_ _05021_ _05138_ vssd1 vssd1 vccd1 vccd1 _05149_ sky130_fd_sc_hd__nor2_1
XFILLER_0_101_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10032_ _04425_ vssd1 vssd1 vccd1 vccd1 _00351_ sky130_fd_sc_hd__clkbuf_1
X_11983_ _03732_ net1007 _05796_ vssd1 vssd1 vccd1 vccd1 _00931_ sky130_fd_sc_hd__o21a_1
XFILLER_0_98_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13722_ clknet_leaf_97_clk _01033_ net161 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.quo\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10934_ _05051_ vssd1 vssd1 vccd1 vccd1 _05052_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_738 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13653_ clknet_leaf_41_clk net354 net116 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.quo\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10865_ _04970_ _05007_ _05008_ vssd1 vssd1 vccd1 vccd1 _05009_ sky130_fd_sc_hd__a21o_1
XFILLER_0_85_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06494__B _01223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12604_ clknet_leaf_21_clk genblk1\[3\].osc.clkdiv_C.next_cnt\[7\] net97 vssd1 vssd1
+ vccd1 vccd1 genblk1\[3\].osc.clkdiv_C.cnt\[7\] sky130_fd_sc_hd__dfrtp_4
XPHY_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13584_ clknet_leaf_75_clk _00899_ net207 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.acc\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10796_ net1012 _04858_ _04922_ _04948_ vssd1 vssd1 vccd1 vccd1 _00592_ sky130_fd_sc_hd__a22o_1
XPHY_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12535_ clknet_leaf_45_clk _00087_ net186 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.b1\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08472__B1 _02526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09297__S _03804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12466_ clknet_leaf_33_clk smpl_rt_clkdiv.clkDiv_inst.next_cnt\[0\] net101 vssd1
+ vssd1 vccd1 vccd1 smpl_rt_clkdiv.clkDiv_inst.cnt\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11417_ _05366_ _05391_ _05392_ vssd1 vssd1 vccd1 vccd1 _05393_ sky130_fd_sc_hd__a21o_1
X_12397_ _05964_ _06069_ vssd1 vssd1 vccd1 vccd1 _06070_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_111_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11348_ net923 _05311_ _05315_ _05335_ vssd1 vssd1 vccd1 vccd1 _00757_ sky130_fd_sc_hd__a22o_1
XANTENNA__06250__A2 _01211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10760__A _04856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11279_ _05249_ vssd1 vssd1 vccd1 vccd1 _05283_ sky130_fd_sc_hd__clkbuf_4
X_13018_ clknet_leaf_123_clk _00345_ net76 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.i\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10334__A1 _01240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06669__B _01180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07510_ PWM.counter\[5\] vssd1 vssd1 vccd1 vccd1 _02230_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10098__B1 _04454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08490_ _03164_ _03169_ _03163_ vssd1 vssd1 vccd1 vccd1 _03197_ sky130_fd_sc_hd__a21bo_1
X_07441_ _02175_ _02153_ genblk2\[4\].wave_shpr.div.busy vssd1 vssd1 vccd1 vccd1 _02178_
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_71_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_900 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07372_ _02126_ vssd1 vssd1 vccd1 vccd1 genblk1\[11\].osc.clkdiv_C.next_cnt\[9\]
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08058__A3 _01180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09111_ genblk2\[0\].wave_shpr.div.acc\[4\] genblk2\[0\].wave_shpr.div.b1\[4\] vssd1
+ vssd1 vccd1 vccd1 _03759_ sky130_fd_sc_hd__or2b_1
XFILLER_0_44_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06323_ genblk1\[0\].osc.clkdiv_C.cnt\[4\] _01276_ genblk1\[0\].osc.clkdiv_C.cnt\[5\]
+ vssd1 vssd1 vccd1 vccd1 _01280_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10935__A _02152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_142_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12451__RESET_B net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09042_ _03709_ vssd1 vssd1 vccd1 vccd1 _00077_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_754 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06254_ genblk1\[0\].osc.clkdiv_C.cnt\[4\] _01215_ _01193_ genblk1\[0\].osc.clkdiv_C.cnt\[9\]
+ vssd1 vssd1 vccd1 vccd1 _01216_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_143_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12011__A1 _03687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold400 _00814_ vssd1 vssd1 vccd1 vccd1 net618 sky130_fd_sc_hd__dlygate4sd3_1
X_06185_ _01152_ _01097_ sig_norm.busy vssd1 vssd1 vccd1 vccd1 _01156_ sky130_fd_sc_hd__and3b_1
Xhold411 sig_norm.acc\[1\] vssd1 vssd1 vccd1 vccd1 net629 sky130_fd_sc_hd__dlygate4sd3_1
Xhold422 genblk2\[7\].wave_shpr.div.quo\[13\] vssd1 vssd1 vccd1 vccd1 net640 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout204_A net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07569__A2 _01577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold433 genblk2\[10\].wave_shpr.div.b1\[5\] vssd1 vssd1 vccd1 vccd1 net651 sky130_fd_sc_hd__dlygate4sd3_1
Xhold444 _00716_ vssd1 vssd1 vccd1 vccd1 net662 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09963__B1 _03855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold455 _00469_ vssd1 vssd1 vccd1 vccd1 net673 sky130_fd_sc_hd__dlygate4sd3_1
Xhold466 genblk2\[1\].wave_shpr.div.quo\[1\] vssd1 vssd1 vccd1 vccd1 net684 sky130_fd_sc_hd__dlygate4sd3_1
Xhold477 genblk1\[10\].osc.clkdiv_C.cnt\[17\] vssd1 vssd1 vccd1 vccd1 net695 sky130_fd_sc_hd__dlygate4sd3_1
X_09944_ genblk2\[2\].wave_shpr.div.acc\[24\] _04253_ _04322_ _04347_ vssd1 vssd1
+ vccd1 vccd1 _00341_ sky130_fd_sc_hd__a22o_1
Xhold488 genblk2\[7\].wave_shpr.div.acc\[22\] vssd1 vssd1 vccd1 vccd1 net706 sky130_fd_sc_hd__dlygate4sd3_1
Xhold499 sig_norm.acc\[9\] vssd1 vssd1 vccd1 vccd1 net717 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12361__S _05982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09875_ _04185_ _04167_ vssd1 vssd1 vccd1 vccd1 _04296_ sky130_fd_sc_hd__or2b_1
Xhold1100 genblk2\[7\].wave_shpr.div.quo\[3\] vssd1 vssd1 vccd1 vccd1 net1318 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11522__B1 _05449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06579__B _01182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1111 genblk2\[2\].wave_shpr.div.quo\[2\] vssd1 vssd1 vccd1 vccd1 net1329 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1122 genblk2\[4\].wave_shpr.div.acc\[7\] vssd1 vssd1 vccd1 vccd1 net1340 sky130_fd_sc_hd__dlygate4sd3_1
X_08826_ _02575_ _03532_ vssd1 vssd1 vccd1 vccd1 _03533_ sky130_fd_sc_hd__xor2_2
XANTENNA__07741__A2 _01337_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08757_ _03461_ _03463_ vssd1 vssd1 vccd1 vccd1 _03464_ sky130_fd_sc_hd__and2_1
XTAP_2605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10089__B1 _04456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07708_ _02225_ _02403_ vssd1 vssd1 vccd1 vccd1 _02415_ sky130_fd_sc_hd__and2_1
XTAP_2649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08688_ _03384_ _03393_ _03394_ vssd1 vssd1 vccd1 vccd1 _03395_ sky130_fd_sc_hd__or3_2
XTAP_1915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07639_ _02333_ _02334_ vssd1 vssd1 vccd1 vccd1 _02346_ sky130_fd_sc_hd__or2b_1
XTAP_1959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11006__A _05054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10650_ _04852_ vssd1 vssd1 vccd1 vccd1 _00542_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_137_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09309_ _03780_ _03894_ vssd1 vssd1 vccd1 vccd1 _03895_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_134_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10581_ _04766_ _04807_ _04808_ vssd1 vssd1 vccd1 vccd1 _04809_ sky130_fd_sc_hd__a21o_1
XFILLER_0_146_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12320_ _05835_ genblk1\[11\].osc.clkdiv_C.cnt\[5\] vssd1 vssd1 vccd1 vccd1 _06018_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_106_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10800__A2 _04855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12002__A1 _02002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12251_ genblk2\[11\].wave_shpr.div.fin_quo\[3\] net402 _00005_ vssd1 vssd1 vccd1
+ vccd1 _05986_ sky130_fd_sc_hd__mux2_1
X_11202_ _03702_ net1147 vssd1 vssd1 vccd1 vccd1 _05242_ sky130_fd_sc_hd__nor2_1
X_12182_ _00002_ _05920_ net1153 vssd1 vssd1 vccd1 vccd1 _05922_ sky130_fd_sc_hd__a21oi_1
X_11133_ genblk2\[7\].wave_shpr.div.b1\[6\] genblk2\[7\].wave_shpr.div.acc\[6\] vssd1
+ vssd1 vccd1 vccd1 _05193_ sky130_fd_sc_hd__and2b_1
XANTENNA__12305__A2 _06009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11064_ net560 _05119_ _05126_ _05137_ vssd1 vssd1 vccd1 vccd1 _00671_ sky130_fd_sc_hd__a22o_1
XANTENNA__11513__B1 _05449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09182__A1 _01214_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10015_ _04245_ genblk2\[3\].wave_shpr.div.acc\[16\] vssd1 vssd1 vccd1 vccd1 _04411_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_99_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07732__A2 _02433_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11966_ genblk2\[10\].wave_shpr.div.fin_quo\[0\] _05787_ _00003_ vssd1 vssd1 vccd1
+ vccd1 _05788_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10917_ _05043_ vssd1 vssd1 vccd1 vccd1 _00618_ sky130_fd_sc_hd__clkbuf_1
X_13705_ clknet_leaf_37_clk _01016_ net113 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.b1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_11897_ genblk2\[0\].wave_shpr.div.i\[1\] genblk2\[0\].wave_shpr.div.i\[0\] vssd1
+ vssd1 vccd1 vccd1 _05723_ sky130_fd_sc_hd__or2_1
XFILLER_0_129_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_132_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13636_ clknet_leaf_68_clk _00949_ net195 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.quo\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_27_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10848_ genblk2\[6\].wave_shpr.div.b1\[5\] genblk2\[6\].wave_shpr.div.acc\[5\] vssd1
+ vssd1 vccd1 vccd1 _04992_ sky130_fd_sc_hd__and2b_1
XFILLER_0_73_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13567_ clknet_leaf_55_clk net350 net176 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.quo\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10779_ genblk2\[5\].wave_shpr.div.acc\[17\] _04936_ _04907_ vssd1 vssd1 vccd1 vccd1
+ _04937_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10755__A _02183_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_156 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07799__A2 _01349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12518_ clknet_leaf_105_clk PWM.next_counter\[2\] net155 vssd1 vssd1 vccd1 vccd1
+ PWM.counter\[2\] sky130_fd_sc_hd__dfrtp_1
XANTENNA__08225__A _02837_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_329 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13498_ clknet_leaf_86_clk _00815_ net178 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.quo\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12449_ clknet_leaf_106_clk net766 net153 vssd1 vssd1 vccd1 vccd1 sig_norm.i\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09755__S _04039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11752__B1 _05624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07990_ _02604_ _02645_ _02648_ _02696_ vssd1 vssd1 vccd1 vccd1 _02697_ sky130_fd_sc_hd__nand4_2
Xfanout209 net210 vssd1 vssd1 vccd1 vccd1 net209 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_5_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06941_ genblk1\[6\].osc.clkdiv_C.cnt\[12\] _01779_ _01782_ vssd1 vssd1 vccd1 vccd1
+ genblk1\[6\].osc.clkdiv_C.next_cnt\[12\] sky130_fd_sc_hd__o21a_1
XANTENNA__11504__B1 _05446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09660_ genblk2\[1\].wave_shpr.div.acc\[25\] _04009_ _04145_ vssd1 vssd1 vccd1 vccd1
+ _04146_ sky130_fd_sc_hd__a21bo_1
X_06872_ _01441_ _01366_ vssd1 vssd1 vccd1 vccd1 _01726_ sky130_fd_sc_hd__nor2_1
X_08611_ _03316_ _02223_ _03317_ vssd1 vssd1 vccd1 vccd1 _03318_ sky130_fd_sc_hd__or3b_1
XANTENNA__07723__A2 _01323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09591_ _04010_ vssd1 vssd1 vccd1 vccd1 _04095_ sky130_fd_sc_hd__buf_4
X_08542_ genblk2\[7\].wave_shpr.div.fin_quo\[0\] _02526_ _02308_ genblk2\[7\].wave_shpr.div.fin_quo\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03249_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11205__B1_N _03728_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08473_ genblk2\[5\].wave_shpr.div.fin_quo\[3\] _03178_ _03179_ vssd1 vssd1 vccd1
+ vccd1 _03180_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11283__A2 _05279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07424_ _02162_ _02153_ genblk2\[2\].wave_shpr.div.busy vssd1 vssd1 vccd1 vccd1 _02165_
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_64_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12632__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_147_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07355_ _02112_ vssd1 vssd1 vccd1 vccd1 _02113_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10243__B1 _04457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06306_ _01169_ _01185_ _01219_ _01267_ vssd1 vssd1 vccd1 vccd1 _01268_ sky130_fd_sc_hd__o211a_2
XFILLER_0_122_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07286_ genblk1\[10\].osc.clkdiv_C.cnt\[13\] _02053_ _02027_ vssd1 vssd1 vccd1 vccd1
+ _02055_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_115 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09025_ _03691_ _03694_ _03695_ _03696_ net1149 vssd1 vssd1 vccd1 vccd1 _00073_ sky130_fd_sc_hd__a32o_1
X_06237_ genblk1\[0\].osc.clkdiv_C.cnt\[17\] _01197_ _01198_ vssd1 vssd1 vccd1 vccd1
+ _01199_ sky130_fd_sc_hd__a21o_1
Xhold230 genblk2\[1\].wave_shpr.div.acc\[24\] vssd1 vssd1 vccd1 vccd1 net448 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_896 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06168_ _01133_ _01137_ _01139_ vssd1 vssd1 vccd1 vccd1 _01140_ sky130_fd_sc_hd__a21oi_1
Xhold241 genblk2\[5\].wave_shpr.div.quo\[23\] vssd1 vssd1 vccd1 vccd1 net459 sky130_fd_sc_hd__dlygate4sd3_1
Xhold252 _00806_ vssd1 vssd1 vccd1 vccd1 net470 sky130_fd_sc_hd__dlygate4sd3_1
Xhold263 genblk2\[9\].wave_shpr.div.quo\[11\] vssd1 vssd1 vccd1 vccd1 net481 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12091__S _05787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold274 genblk2\[7\].wave_shpr.div.quo\[8\] vssd1 vssd1 vccd1 vccd1 net492 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10604__S _00015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold285 genblk2\[5\].wave_shpr.div.quo\[20\] vssd1 vssd1 vccd1 vccd1 net503 sky130_fd_sc_hd__dlygate4sd3_1
Xhold296 genblk2\[3\].wave_shpr.div.quo\[15\] vssd1 vssd1 vccd1 vccd1 net514 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09927_ _04209_ net22 vssd1 vssd1 vccd1 vccd1 _04336_ sky130_fd_sc_hd__or2_1
XANTENNA__12299__B2 _05982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09858_ genblk2\[2\].wave_shpr.div.b1\[2\] genblk2\[2\].wave_shpr.div.acc\[2\] vssd1
+ vssd1 vccd1 vccd1 _04283_ sky130_fd_sc_hd__xor2_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout67_A net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08809_ _03513_ _03514_ _03511_ _03515_ vssd1 vssd1 vccd1 vccd1 _03516_ sky130_fd_sc_hd__a211o_1
X_09789_ net730 vssd1 vssd1 vccd1 vccd1 _04245_ sky130_fd_sc_hd__inv_2
XTAP_2402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11820_ genblk2\[9\].wave_shpr.div.acc\[6\] _05666_ _05613_ vssd1 vssd1 vccd1 vccd1
+ _05667_ sky130_fd_sc_hd__mux2_1
XTAP_2424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07214__A _01181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11751_ net267 _05623_ _05624_ net712 vssd1 vssd1 vccd1 vccd1 _00871_ sky130_fd_sc_hd__a22o_1
XTAP_1734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_80_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_80_clk sky130_fd_sc_hd__clkbuf_16
XTAP_1756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10702_ genblk2\[5\].wave_shpr.div.acc_next\[0\] _02183_ _04856_ net324 _04878_ vssd1
+ vssd1 vccd1 vccd1 _00568_ sky130_fd_sc_hd__a221o_1
XTAP_1767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11682_ genblk2\[9\].wave_shpr.div.b1\[1\] genblk2\[9\].wave_shpr.div.acc\[1\] vssd1
+ vssd1 vccd1 vccd1 _05574_ sky130_fd_sc_hd__xor2_1
XTAP_1789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13421_ clknet_leaf_92_clk _00740_ net147 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.acc\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10633_ _04843_ vssd1 vssd1 vccd1 vccd1 _00534_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13352_ clknet_leaf_4_clk _00673_ net45 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.acc\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_118_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10564_ genblk2\[5\].wave_shpr.div.b1\[6\] genblk2\[5\].wave_shpr.div.acc\[6\] vssd1
+ vssd1 vccd1 vccd1 _04792_ sky130_fd_sc_hd__and2b_1
XFILLER_0_140_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_649 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12303_ net767 _06009_ _06010_ net776 vssd1 vssd1 vccd1 vccd1 _01037_ sky130_fd_sc_hd__a22o_1
XANTENNA__11982__B1 _03702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13283_ clknet_leaf_117_clk _00604_ net137 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.fin_quo\[3\]
+ sky130_fd_sc_hd__dfrtp_2
X_10495_ genblk2\[4\].wave_shpr.div.acc\[17\] _04736_ _04622_ vssd1 vssd1 vccd1 vccd1
+ _04737_ sky130_fd_sc_hd__mux2_1
XANTENNA__09575__S _04011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12234_ _05927_ _05970_ _05971_ vssd1 vssd1 vccd1 vccd1 _05972_ sky130_fd_sc_hd__a21o_1
XFILLER_0_20_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12165_ genblk2\[10\].wave_shpr.div.acc\[22\] _05908_ genblk2\[10\].wave_shpr.div.acc\[23\]
+ vssd1 vssd1 vccd1 vccd1 _05911_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_20_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11116_ genblk2\[7\].wave_shpr.div.acc\[5\] genblk2\[7\].wave_shpr.div.b1\[5\] vssd1
+ vssd1 vccd1 vccd1 _05176_ sky130_fd_sc_hd__or2b_1
XANTENNA__07953__A2 _01732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12096_ net1241 _05844_ _05850_ _05859_ vssd1 vssd1 vccd1 vccd1 _00981_ sky130_fd_sc_hd__a22o_1
XFILLER_0_127_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11047_ genblk2\[6\].wave_shpr.div.acc\[13\] _05124_ _05105_ vssd1 vssd1 vccd1 vccd1
+ _05125_ sky130_fd_sc_hd__mux2_1
Xinput9 pb[3] vssd1 vssd1 vccd1 vccd1 net9 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_98_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12998_ clknet_leaf_131_clk _00327_ net64 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.acc\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07124__A _01336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08666__B1 _02316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11949_ _05736_ _05769_ _05770_ vssd1 vssd1 vccd1 vccd1 _05771_ sky130_fd_sc_hd__a21o_1
XFILLER_0_143_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_71_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_71_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_86_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_74_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13619_ clknet_leaf_68_clk _00932_ net211 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.b1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_144_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07140_ genblk1\[9\].osc.clkdiv_C.cnt\[6\] _01334_ _01328_ genblk1\[9\].osc.clkdiv_C.cnt\[13\]
+ vssd1 vssd1 vccd1 vccd1 _01940_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_109_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07071_ genblk1\[8\].osc.clkdiv_C.cnt\[1\] genblk1\[8\].osc.clkdiv_C.cnt\[0\] vssd1
+ vssd1 vccd1 vccd1 _01888_ sky130_fd_sc_hd__or2_1
XFILLER_0_112_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_11_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07973_ genblk1\[7\].osc.clkdiv_C.cnt\[16\] genblk1\[7\].osc.clkdiv_C.cnt\[17\] vssd1
+ vssd1 vccd1 vccd1 _02680_ sky130_fd_sc_hd__nor2_1
X_09712_ _04164_ _04190_ _04191_ vssd1 vssd1 vccd1 vccd1 _04192_ sky130_fd_sc_hd__a21o_1
X_06924_ _01761_ _01770_ _01771_ vssd1 vssd1 vccd1 vccd1 genblk1\[6\].osc.clkdiv_C.next_cnt\[6\]
+ sky130_fd_sc_hd__nor3_1
X_09643_ _04133_ _04134_ vssd1 vssd1 vccd1 vccd1 _04135_ sky130_fd_sc_hd__nand2_1
X_06855_ genblk1\[5\].osc.clkdiv_C.cnt\[12\] _01714_ vssd1 vssd1 vccd1 vccd1 _01715_
+ sky130_fd_sc_hd__and2_1
X_09574_ _03975_ _04081_ vssd1 vssd1 vccd1 vccd1 _04082_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06786_ _01489_ net37 vssd1 vssd1 vccd1 vccd1 _01658_ sky130_fd_sc_hd__nand2_2
XTAP_1008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08525_ _02310_ _03231_ _02314_ vssd1 vssd1 vccd1 vccd1 _03232_ sky130_fd_sc_hd__o21a_1
XANTENNA__07034__A genblk1\[8\].osc.clkdiv_C.cnt\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_62_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_62_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__08121__A2 _01439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_60_clk_A clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08456_ _02946_ _03158_ _03162_ vssd1 vssd1 vccd1 vccd1 _03163_ sky130_fd_sc_hd__or3b_2
XFILLER_0_65_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07407_ genblk2\[0\].wave_shpr.div.start vssd1 vssd1 vccd1 vccd1 _02152_ sky130_fd_sc_hd__inv_6
XFILLER_0_46_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08387_ genblk1\[2\].osc.clkdiv_C.cnt\[6\] _01433_ _03093_ vssd1 vssd1 vccd1 vccd1
+ _03094_ sky130_fd_sc_hd__o21a_1
XANTENNA__10395__A _04477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06592__B _01437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07338_ _02092_ _02098_ _02099_ vssd1 vssd1 vccd1 vccd1 _02100_ sky130_fd_sc_hd__and3_1
XANTENNA_clkbuf_leaf_75_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07269_ genblk1\[10\].osc.clkdiv_C.cnt\[7\] _02041_ vssd1 vssd1 vccd1 vccd1 _02044_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_6_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09008_ net1132 sig_norm.quo\[5\] _01154_ vssd1 vssd1 vccd1 vccd1 _03684_ sky130_fd_sc_hd__mux2_1
XANTENNA__07132__A1_N genblk1\[9\].osc.clkdiv_C.cnt\[16\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_103_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10280_ genblk2\[4\].wave_shpr.div.b1\[5\] genblk2\[4\].wave_shpr.div.acc\[5\] vssd1
+ vssd1 vccd1 vccd1 _04592_ sky130_fd_sc_hd__and2b_1
XFILLER_0_103_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10334__S _04440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07209__A _01556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_133_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_13_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12921_ clknet_leaf_35_clk _00252_ net105 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.acc\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12852_ clknet_leaf_118_clk _00183_ net138 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.fin_quo\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_2221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold915_A genblk1\[0\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06371__B2 genblk1\[1\].osc.clkdiv_C.cnt\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11803_ _05577_ _05571_ vssd1 vssd1 vccd1 vccd1 _05654_ sky130_fd_sc_hd__or2b_1
XTAP_2254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12783_ clknet_leaf_40_clk _00116_ net117 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.b1\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_28_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_53_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_53_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_96_674 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11734_ genblk2\[9\].wave_shpr.div.fin_quo\[6\] genblk2\[9\].wave_shpr.div.quo\[5\]
+ _00023_ vssd1 vssd1 vccd1 vccd1 _05620_ sky130_fd_sc_hd__mux2_1
XTAP_2298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_113_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11665_ genblk2\[9\].wave_shpr.div.acc\[14\] genblk2\[9\].wave_shpr.div.b1\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05557_ sky130_fd_sc_hd__or2b_1
Xclkbuf_4_6_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_6_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_154_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10616_ _04833_ vssd1 vssd1 vccd1 vccd1 _00527_ sky130_fd_sc_hd__clkbuf_1
X_13404_ clknet_leaf_90_clk net371 net143 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.quo\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11596_ _05396_ _05364_ vssd1 vssd1 vccd1 vccd1 _05508_ sky130_fd_sc_hd__or2b_1
XFILLER_0_51_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_141_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13335_ clknet_leaf_6_clk _00656_ net48 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.acc\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10547_ genblk2\[5\].wave_shpr.div.acc\[5\] genblk2\[5\].wave_shpr.div.b1\[5\] vssd1
+ vssd1 vccd1 vccd1 _04775_ sky130_fd_sc_hd__or2b_1
XFILLER_0_40_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13266_ clknet_leaf_0_clk _00589_ net38 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.acc\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10478_ _04607_ _04723_ vssd1 vssd1 vccd1 vccd1 _04724_ sky130_fd_sc_hd__xnor2_1
X_12217_ genblk2\[11\].wave_shpr.div.b1\[7\] genblk2\[11\].wave_shpr.div.acc\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05955_ sky130_fd_sc_hd__and2b_1
X_13197_ clknet_leaf_113_clk _00520_ net134 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.fin_quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11183__A1 _04242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12148_ genblk2\[10\].wave_shpr.div.acc\[25\] genblk2\[10\].wave_shpr.div.acc\[26\]
+ _05785_ vssd1 vssd1 vccd1 vccd1 _05899_ sky130_fd_sc_hd__nor3_2
XANTENNA__10930__A1 _03726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12079_ net989 _05844_ _05817_ _05846_ vssd1 vssd1 vccd1 vccd1 _00977_ sky130_fd_sc_hd__a22o_1
XANTENNA__07139__B1 _01196_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06677__B _01565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10694__B1 _04856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06640_ _01523_ _01538_ _01539_ vssd1 vssd1 vccd1 vccd1 genblk1\[3\].osc.clkdiv_C.next_cnt\[8\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_78_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08639__B1 _02526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06571_ _01451_ _01480_ vssd1 vssd1 vccd1 vccd1 _01481_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_44_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_44_clk sky130_fd_sc_hd__clkbuf_16
X_08310_ _03014_ _03015_ _03016_ _02360_ vssd1 vssd1 vccd1 vccd1 _03017_ sky130_fd_sc_hd__o211a_1
X_09290_ net823 _03870_ _03877_ _03880_ vssd1 vssd1 vccd1 vccd1 _00154_ sky130_fd_sc_hd__a22o_1
XFILLER_0_74_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07311__B1 _01262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08241_ _02683_ _02682_ _02689_ _02527_ vssd1 vssd1 vccd1 vccd1 _02948_ sky130_fd_sc_hd__o31ai_1
XANTENNA__07862__A1 _02525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08172_ genblk1\[3\].osc.clkdiv_C.cnt\[13\] _01498_ _02867_ vssd1 vssd1 vccd1 vccd1
+ _02879_ sky130_fd_sc_hd__a21o_1
XANTENNA__07301__B _01595_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07123_ _01432_ _01344_ vssd1 vssd1 vccd1 vccd1 _01923_ sky130_fd_sc_hd__nand2_4
XFILLER_0_132_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07614__A1 _01171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07054_ genblk1\[8\].osc.clkdiv_C.cnt\[15\] _01436_ _01864_ _01868_ _01871_ vssd1
+ vssd1 vccd1 vccd1 _01872_ sky130_fd_sc_hd__a2111o_1
XANTENNA__11758__B genblk1\[9\].osc.clkdiv_C.cnt\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_112_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07917__A2 _01858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07956_ genblk1\[7\].osc.clkdiv_C.cnt\[3\] _02656_ _02659_ _02660_ _02662_ vssd1
+ vssd1 vccd1 vccd1 _02663_ sky130_fd_sc_hd__a221o_1
X_06907_ net28 vssd1 vssd1 vccd1 vccd1 _01761_ sky130_fd_sc_hd__clkbuf_4
X_07887_ _02469_ _02593_ vssd1 vssd1 vccd1 vccd1 _02594_ sky130_fd_sc_hd__or2_1
XFILLER_0_97_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06587__B _01494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09626_ genblk2\[1\].wave_shpr.div.acc\[15\] _04121_ _04095_ vssd1 vssd1 vccd1 vccd1
+ _04122_ sky130_fd_sc_hd__mux2_1
X_06838_ _01693_ _01703_ _01704_ vssd1 vssd1 vccd1 vccd1 genblk1\[5\].osc.clkdiv_C.next_cnt\[5\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_97_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09557_ _04069_ genblk1\[1\].osc.clkdiv_C.cnt\[16\] vssd1 vssd1 vccd1 vccd1 _04070_
+ sky130_fd_sc_hd__and2_1
X_06769_ _01644_ _01642_ _01645_ _01600_ vssd1 vssd1 vccd1 vccd1 genblk1\[4\].osc.clkdiv_C.next_cnt\[13\]
+ sky130_fd_sc_hd__o211a_1
Xclkbuf_leaf_35_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_35_clk sky130_fd_sc_hd__clkbuf_16
X_08508_ _03210_ _03214_ vssd1 vssd1 vccd1 vccd1 _03215_ sky130_fd_sc_hd__xnor2_1
X_09488_ _04033_ vssd1 vssd1 vccd1 vccd1 _00199_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07302__B1 _02064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09842__A2 _04247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08439_ _02404_ _02407_ genblk2\[10\].wave_shpr.div.fin_quo\[2\] vssd1 vssd1 vccd1
+ vccd1 _03146_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_93_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11450_ genblk2\[8\].wave_shpr.div.fin_quo\[4\] net1321 _00021_ vssd1 vssd1 vccd1
+ vccd1 _05422_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10401_ _04477_ genblk1\[4\].osc.clkdiv_C.cnt\[9\] vssd1 vssd1 vccd1 vccd1 _04669_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_104_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06408__A2 _01323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11381_ net328 _05356_ _05357_ vssd1 vssd1 vccd1 vccd1 _00768_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13120_ clknet_leaf_136_clk _00445_ net43 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.b1\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10332_ _03717_ _04634_ vssd1 vssd1 vccd1 vccd1 _00442_ sky130_fd_sc_hd__nand2_1
XFILLER_0_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13051_ clknet_leaf_113_clk net738 net128 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10064__S _04440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10263_ genblk2\[4\].wave_shpr.div.acc\[7\] genblk2\[4\].wave_shpr.div.b1\[7\] vssd1
+ vssd1 vccd1 vccd1 _04575_ sky130_fd_sc_hd__or2b_1
XFILLER_0_103_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08042__B _01359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12002_ net1204 _02002_ _05802_ vssd1 vssd1 vccd1 vccd1 _05806_ sky130_fd_sc_hd__mux2_1
X_10194_ _04404_ _04523_ vssd1 vssd1 vccd1 vccd1 _04524_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12904_ clknet_leaf_37_clk _00235_ net104 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.acc\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2040 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12835_ clknet_leaf_64_clk net689 net196 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.acc\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2051 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_124_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_26_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_26_clk sky130_fd_sc_hd__clkbuf_16
XTAP_2062 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2073 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2084 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2095 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12766_ clknet_leaf_91_clk _00099_ net146 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.fin_quo\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_584 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11717_ genblk2\[9\].wave_shpr.div.acc\[21\] genblk2\[9\].wave_shpr.div.acc\[20\]
+ genblk2\[9\].wave_shpr.div.acc\[19\] _05608_ vssd1 vssd1 vccd1 vccd1 _05609_ sky130_fd_sc_hd__or4_1
X_12697_ clknet_leaf_54_clk genblk1\[8\].osc.clkdiv_C.next_cnt\[10\] net172 vssd1
+ vssd1 vccd1 vccd1 genblk1\[8\].osc.clkdiv_C.cnt\[10\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_127_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11648_ _05444_ _05441_ genblk2\[8\].wave_shpr.div.i\[0\] vssd1 vssd1 vccd1 vccd1
+ _05545_ sky130_fd_sc_hd__mux2_1
Xinput12 pb[6] vssd1 vssd1 vccd1 vccd1 net12 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_154_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11579_ _05388_ _05368_ vssd1 vssd1 vccd1 vccd1 _05495_ sky130_fd_sc_hd__or2b_1
XFILLER_0_3_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold807 genblk2\[2\].wave_shpr.div.b1\[16\] vssd1 vssd1 vccd1 vccd1 net1025 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09329__A _03838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold818 genblk2\[2\].wave_shpr.div.acc\[15\] vssd1 vssd1 vccd1 vccd1 net1036 sky130_fd_sc_hd__dlygate4sd3_1
X_13318_ clknet_leaf_25_clk net624 net86 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.quo\[12\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold829 genblk2\[2\].wave_shpr.div.b1\[2\] vssd1 vssd1 vccd1 vccd1 net1047 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13249_ clknet_leaf_2_clk _00572_ net52 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.acc\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07810_ net1 net150 _02312_ vssd1 vssd1 vccd1 vccd1 _02517_ sky130_fd_sc_hd__and3_1
XANTENNA__07791__B _01263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08790_ _03489_ _03496_ vssd1 vssd1 vccd1 vccd1 _03497_ sky130_fd_sc_hd__xor2_1
XANTENNA__06688__A _01577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07780__B1 _01215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07741_ genblk1\[1\].osc.clkdiv_C.cnt\[11\] _01337_ _01312_ genblk1\[1\].osc.clkdiv_C.cnt\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02448_ sky130_fd_sc_hd__o22a_1
XANTENNA__10667__B1 _04855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07672_ _01308_ genblk1\[10\].osc.clkdiv_C.cnt\[1\] vssd1 vssd1 vccd1 vccd1 _02379_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_79_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10131__A2 _04451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09411_ _03969_ _03973_ _03974_ vssd1 vssd1 vccd1 vccd1 _03975_ sky130_fd_sc_hd__a21o_1
X_06623_ genblk1\[3\].osc.clkdiv_C.cnt\[1\] genblk1\[3\].osc.clkdiv_C.cnt\[0\] genblk1\[3\].osc.clkdiv_C.cnt\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01529_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06886__A2 _01738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_17_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_17_clk sky130_fd_sc_hd__clkbuf_16
X_09342_ _03797_ _03746_ vssd1 vssd1 vccd1 vccd1 _03920_ sky130_fd_sc_hd__or2b_1
X_06554_ net1159 _01466_ _01469_ vssd1 vssd1 vccd1 vccd1 genblk1\[2\].osc.clkdiv_C.next_cnt\[10\]
+ sky130_fd_sc_hd__o21a_1
XANTENNA__09285__B1 _03840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09273_ genblk2\[0\].wave_shpr.div.acc\[1\] _03803_ vssd1 vssd1 vccd1 vccd1 _03867_
+ sky130_fd_sc_hd__or2_1
X_06485_ _01241_ _01337_ vssd1 vssd1 vccd1 vccd1 _01411_ sky130_fd_sc_hd__or2_2
XFILLER_0_117_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08224_ _02527_ _02928_ _02929_ _02930_ vssd1 vssd1 vccd1 vccd1 _02931_ sky130_fd_sc_hd__a31o_1
XANTENNA__13264__RESET_B net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_7_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08155_ genblk1\[3\].osc.clkdiv_C.cnt\[7\] _01483_ _01494_ genblk1\[3\].osc.clkdiv_C.cnt\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02862_ sky130_fd_sc_hd__o22a_1
X_07106_ _01886_ _01910_ vssd1 vssd1 vccd1 vccd1 _01911_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_287 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08086_ genblk2\[5\].wave_shpr.div.fin_quo\[4\] _02792_ vssd1 vssd1 vccd1 vccd1 _02793_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_141_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07037_ _01230_ _01564_ vssd1 vssd1 vccd1 vccd1 _01855_ sky130_fd_sc_hd__nand2_4
X_08988_ _03670_ _03671_ vssd1 vssd1 vccd1 vccd1 _03672_ sky130_fd_sc_hd__xnor2_1
X_07939_ _02217_ _02553_ vssd1 vssd1 vccd1 vccd1 _02646_ sky130_fd_sc_hd__nor2_1
XANTENNA__10658__B1 _04857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10950_ net477 _05057_ _05055_ net515 _05058_ vssd1 vssd1 vccd1 vccd1 _00636_ sky130_fd_sc_hd__a221o_1
X_09609_ genblk2\[1\].wave_shpr.div.acc\[12\] _04076_ _04080_ _04108_ vssd1 vssd1
+ vccd1 vccd1 _00245_ sky130_fd_sc_hd__a22o_1
X_10881_ _05024_ vssd1 vssd1 vccd1 vccd1 _00601_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_38_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12620_ clknet_leaf_17_clk genblk1\[4\].osc.clkdiv_C.next_cnt\[5\] net83 vssd1 vssd1
+ vccd1 vccd1 genblk1\[4\].osc.clkdiv_C.cnt\[5\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__09276__B1 _03841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12551_ clknet_leaf_60_clk genblk1\[0\].osc.clkdiv_C.next_cnt\[8\] net187 vssd1 vssd1
+ vccd1 vccd1 genblk1\[0\].osc.clkdiv_C.cnt\[8\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__10059__S _04238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11502_ net751 _05442_ _05446_ net795 vssd1 vssd1 vccd1 vccd1 _00800_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12482_ clknet_leaf_108_clk _00044_ net151 vssd1 vssd1 vccd1 vccd1 sig_norm.acc\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11433_ _05358_ _05407_ _05408_ vssd1 vssd1 vccd1 vccd1 _05409_ sky130_fd_sc_hd__a21o_1
XFILLER_0_110_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11364_ _05345_ _05342_ _05346_ vssd1 vssd1 vccd1 vccd1 _05347_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11398__B genblk2\[8\].wave_shpr.div.b1\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07054__A2 _01436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10315_ _04625_ vssd1 vssd1 vccd1 vccd1 _00434_ sky130_fd_sc_hd__clkbuf_1
X_13103_ clknet_leaf_12_clk _00428_ net51 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.i\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__06262__B1 _01223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11295_ _05195_ _05174_ vssd1 vssd1 vccd1 vccd1 _05295_ sky130_fd_sc_hd__or2b_1
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09583__S _04011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13034_ clknet_leaf_127_clk _00361_ net66 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.b1\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10246_ _04560_ vssd1 vssd1 vccd1 vccd1 _04561_ sky130_fd_sc_hd__inv_2
XFILLER_0_119_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10177_ genblk2\[3\].wave_shpr.div.acc\[9\] _04510_ _04507_ vssd1 vssd1 vccd1 vccd1
+ _04511_ sky130_fd_sc_hd__mux2_1
XANTENNA__06301__A _01238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09503__A1 _03714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_76_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12818_ clknet_leaf_67_clk _00151_ net193 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.acc\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_57_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09806__A2 _04248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12749_ clknet_leaf_46_clk genblk1\[11\].osc.clkdiv_C.next_cnt\[8\] net119 vssd1
+ vssd1 vccd1 vccd1 genblk1\[11\].osc.clkdiv_C.cnt\[8\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_151_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09758__S _04039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06270_ freq_div.state\[0\] freq_div.state\[1\] vssd1 vssd1 vccd1 vccd1 _01232_ sky130_fd_sc_hd__and2_1
XFILLER_0_115_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold604 genblk2\[7\].wave_shpr.div.quo\[0\] vssd1 vssd1 vccd1 vccd1 net822 sky130_fd_sc_hd__dlygate4sd3_1
Xhold615 genblk2\[8\].wave_shpr.div.acc\[13\] vssd1 vssd1 vccd1 vccd1 net833 sky130_fd_sc_hd__dlygate4sd3_1
Xhold626 genblk2\[10\].wave_shpr.div.acc\[11\] vssd1 vssd1 vccd1 vccd1 net844 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold637 genblk2\[5\].wave_shpr.div.i\[4\] vssd1 vssd1 vccd1 vccd1 net855 sky130_fd_sc_hd__dlygate4sd3_1
Xhold648 genblk2\[0\].wave_shpr.div.acc\[6\] vssd1 vssd1 vccd1 vccd1 net866 sky130_fd_sc_hd__dlygate4sd3_1
X_09960_ _00008_ _04356_ net1123 vssd1 vssd1 vccd1 vccd1 _04358_ sky130_fd_sc_hd__a21oi_1
Xhold659 genblk2\[7\].wave_shpr.div.acc\[4\] vssd1 vssd1 vccd1 vccd1 net877 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_6_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_6_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_122_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08911_ _03611_ _03612_ vssd1 vssd1 vccd1 vccd1 _03613_ sky130_fd_sc_hd__nand2_1
XTAP_920 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09891_ net952 _04282_ _04289_ _04308_ vssd1 vssd1 vccd1 vccd1 _00327_ sky130_fd_sc_hd__a22o_1
XTAP_931 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_953 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08842_ _03545_ _03548_ vssd1 vssd1 vccd1 vccd1 _03549_ sky130_fd_sc_hd__and2b_1
XTAP_964 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_986 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_997 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08773_ _03474_ _03479_ vssd1 vssd1 vccd1 vccd1 _03480_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_109_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout184_A net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07724_ genblk1\[1\].osc.clkdiv_C.cnt\[2\] _01323_ _01313_ genblk1\[1\].osc.clkdiv_C.cnt\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02431_ sky130_fd_sc_hd__o22a_1
XTAP_2809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07505__B1 _02225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09522__A _03853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07655_ _02361_ vssd1 vssd1 vccd1 vccd1 _02362_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_79_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10668__A _04672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06606_ _01234_ vssd1 vssd1 vccd1 vccd1 _01514_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_125_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_149_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07586_ _02278_ _02279_ _02281_ vssd1 vssd1 vccd1 vccd1 _02293_ sky130_fd_sc_hd__a21o_1
X_09325_ _03789_ _03750_ vssd1 vssd1 vccd1 vccd1 _03907_ sky130_fd_sc_hd__or2b_1
X_06537_ _01452_ _01458_ vssd1 vssd1 vccd1 vccd1 genblk1\[2\].osc.clkdiv_C.next_cnt\[4\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09256_ genblk2\[0\].wave_shpr.div.quo\[20\] _03845_ _03847_ net298 _03857_ vssd1
+ vssd1 vccd1 vccd1 _00143_ sky130_fd_sc_hd__a221o_1
X_06468_ _01373_ _01399_ vssd1 vssd1 vccd1 vccd1 _01400_ sky130_fd_sc_hd__nor2_1
XANTENNA__06881__A _01189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_16_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_796 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08207_ _02310_ _02913_ _02314_ vssd1 vssd1 vccd1 vccd1 _02914_ sky130_fd_sc_hd__o21a_1
XFILLER_0_106_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09187_ net1173 vssd1 vssd1 vccd1 vccd1 _03821_ sky130_fd_sc_hd__inv_2
X_06399_ _01173_ _01175_ vssd1 vssd1 vccd1 vccd1 _01343_ sky130_fd_sc_hd__or2_1
XANTENNA__11368__A1 _05245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08138_ genblk2\[4\].wave_shpr.div.fin_quo\[7\] _02309_ _02844_ _02527_ vssd1 vssd1
+ vccd1 vccd1 _02845_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08069_ genblk1\[5\].osc.clkdiv_C.cnt\[2\] _01592_ _02775_ vssd1 vssd1 vccd1 vccd1
+ _02776_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10100_ net631 _04457_ _04454_ net538 _04459_ vssd1 vssd1 vccd1 vccd1 _00385_ sky130_fd_sc_hd__a221o_1
XANTENNA_fanout97_A net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11080_ net659 _05057_ _05126_ _05148_ vssd1 vssd1 vccd1 vccd1 _00676_ sky130_fd_sc_hd__a22o_1
X_10031_ genblk2\[3\].wave_shpr.div.fin_quo\[2\] net326 _04422_ vssd1 vssd1 vccd1
+ vccd1 _04425_ sky130_fd_sc_hd__mux2_1
XANTENNA__10342__S _04637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07744__B1 _01344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12096__A2 _05844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11982_ _01441_ _01320_ _03702_ vssd1 vssd1 vccd1 vccd1 _05796_ sky130_fd_sc_hd__o21ai_4
X_13721_ clknet_leaf_40_clk _01032_ net118 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.b1\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10933_ _02188_ vssd1 vssd1 vccd1 vccd1 _05051_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13652_ clknet_leaf_40_clk _00965_ net116 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.quo\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10864_ genblk2\[6\].wave_shpr.div.b1\[13\] genblk2\[6\].wave_shpr.div.acc\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05008_ sky130_fd_sc_hd__and2b_1
XFILLER_0_39_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12603_ clknet_leaf_21_clk genblk1\[3\].osc.clkdiv_C.next_cnt\[6\] net97 vssd1 vssd1
+ vccd1 vccd1 genblk1\[3\].osc.clkdiv_C.cnt\[6\] sky130_fd_sc_hd__dfrtp_4
XPHY_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10795_ genblk2\[5\].wave_shpr.div.acc\[22\] _04817_ _04947_ vssd1 vssd1 vccd1 vccd1
+ _04948_ sky130_fd_sc_hd__a21o_1
X_13583_ clknet_leaf_76_clk _00898_ net207 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.acc\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_27_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12534_ clknet_leaf_45_clk _00086_ net186 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.b1\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_30_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12465_ clknet_leaf_31_clk smpl_rt_clkdiv.clkDiv_inst.next_hzX net99 vssd1 vssd1
+ vccd1 vccd1 genblk2\[0\].wave_shpr.div.start sky130_fd_sc_hd__dfrtp_4
XFILLER_0_34_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_124_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11202__A _03702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08224__A1 _02527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11416_ genblk2\[8\].wave_shpr.div.b1\[9\] genblk2\[8\].wave_shpr.div.acc\[9\] vssd1
+ vssd1 vccd1 vccd1 _05392_ sky130_fd_sc_hd__and2b_1
X_12396_ _05965_ _05930_ vssd1 vssd1 vccd1 vccd1 _06069_ sky130_fd_sc_hd__or2b_1
XFILLER_0_1_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11347_ genblk2\[7\].wave_shpr.div.acc\[19\] _05217_ _05334_ vssd1 vssd1 vccd1 vccd1
+ _05335_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_120_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11278_ net992 _05279_ _05250_ _05282_ vssd1 vssd1 vccd1 vccd1 _00740_ sky130_fd_sc_hd__a22o_1
X_10229_ genblk2\[3\].wave_shpr.div.acc\[23\] _04417_ vssd1 vssd1 vccd1 vccd1 _04549_
+ sky130_fd_sc_hd__nor2_1
X_13017_ clknet_leaf_124_clk _00344_ net76 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.i\[0\]
+ sky130_fd_sc_hd__dfrtp_2
Xhold1 PWM.pwm_out vssd1 vssd1 vccd1 vccd1 net219 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06966__A _01192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10098__B2 genblk2\[3\].wave_shpr.div.quo\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07440_ _02177_ vssd1 vssd1 vccd1 vccd1 _00012_ sky130_fd_sc_hd__inv_2
XFILLER_0_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07371_ _02091_ _02124_ _02125_ vssd1 vssd1 vccd1 vccd1 _02126_ sky130_fd_sc_hd__and3_1
X_09110_ genblk2\[0\].wave_shpr.div.acc\[5\] genblk2\[0\].wave_shpr.div.b1\[5\] vssd1
+ vssd1 vccd1 vccd1 _03758_ sky130_fd_sc_hd__or2b_1
X_06322_ genblk1\[0\].osc.clkdiv_C.cnt\[5\] genblk1\[0\].osc.clkdiv_C.cnt\[4\] _01276_
+ vssd1 vssd1 vccd1 vccd1 _01279_ sky130_fd_sc_hd__and3_1
XFILLER_0_33_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_143_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09041_ net1243 _03706_ _03708_ vssd1 vssd1 vccd1 vccd1 _03709_ sky130_fd_sc_hd__mux2_1
X_06253_ _01213_ _01214_ vssd1 vssd1 vccd1 vccd1 _01215_ sky130_fd_sc_hd__nand2_2
XFILLER_0_115_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_766 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06184_ _01094_ _01095_ _01096_ vssd1 vssd1 vccd1 vccd1 _01155_ sky130_fd_sc_hd__or3_4
Xhold401 genblk2\[11\].wave_shpr.div.acc\[23\] vssd1 vssd1 vccd1 vccd1 net619 sky130_fd_sc_hd__dlygate4sd3_1
Xhold412 genblk2\[5\].wave_shpr.div.acc\[18\] vssd1 vssd1 vccd1 vccd1 net630 sky130_fd_sc_hd__dlygate4sd3_1
Xhold423 genblk2\[11\].wave_shpr.div.acc\[19\] vssd1 vssd1 vccd1 vccd1 net641 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold434 genblk2\[0\].wave_shpr.div.quo\[5\] vssd1 vssd1 vccd1 vccd1 net652 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12491__RESET_B net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold445 sig_norm.acc\[10\] vssd1 vssd1 vccd1 vccd1 net663 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10951__A _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold456 genblk2\[10\].wave_shpr.div.b1\[15\] vssd1 vssd1 vccd1 vccd1 net674 sky130_fd_sc_hd__dlygate4sd3_1
Xhold467 _00209_ vssd1 vssd1 vccd1 vccd1 net685 sky130_fd_sc_hd__dlygate4sd3_1
Xhold478 genblk2\[2\].wave_shpr.div.quo\[4\] vssd1 vssd1 vccd1 vccd1 net696 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09943_ genblk2\[2\].wave_shpr.div.acc\[23\] _04211_ _04346_ vssd1 vssd1 vccd1 vccd1
+ _04347_ sky130_fd_sc_hd__a21o_1
Xhold489 genblk2\[2\].wave_shpr.div.acc\[23\] vssd1 vssd1 vccd1 vccd1 net707 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09874_ net887 _04282_ _04289_ _04295_ vssd1 vssd1 vccd1 vccd1 _00323_ sky130_fd_sc_hd__a22o_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1101 genblk2\[6\].wave_shpr.div.quo\[3\] vssd1 vssd1 vccd1 vccd1 net1319 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1112 genblk2\[5\].wave_shpr.div.quo\[4\] vssd1 vssd1 vccd1 vccd1 net1330 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08825_ _02581_ _02580_ vssd1 vssd1 vccd1 vccd1 _03532_ sky130_fd_sc_hd__or2b_1
Xhold1123 genblk2\[11\].wave_shpr.div.quo\[6\] vssd1 vssd1 vccd1 vccd1 net1341 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08756_ _03234_ _03462_ vssd1 vssd1 vccd1 vccd1 _03463_ sky130_fd_sc_hd__nor2_1
XTAP_2606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06876__A _01336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09252__A _03719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07707_ _02316_ _02411_ _02413_ vssd1 vssd1 vccd1 vccd1 _02414_ sky130_fd_sc_hd__or3_1
XANTENNA__11286__B1 _05283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08687_ _03381_ _03382_ _03298_ _03333_ vssd1 vssd1 vccd1 vccd1 _03394_ sky130_fd_sc_hd__o211a_1
XTAP_1905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08151__B1 _01514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07638_ _01229_ _02081_ _02085_ vssd1 vssd1 vccd1 vccd1 _02345_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_137_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07569_ genblk1\[9\].osc.clkdiv_C.cnt\[15\] _01577_ _02274_ _02275_ vssd1 vssd1 vccd1
+ vccd1 _02276_ sky130_fd_sc_hd__a211o_1
XFILLER_0_48_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_75_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09308_ _03781_ _03754_ vssd1 vssd1 vccd1 vccd1 _03894_ sky130_fd_sc_hd__or2b_1
X_10580_ genblk2\[5\].wave_shpr.div.b1\[14\] genblk2\[5\].wave_shpr.div.acc\[14\]
+ vssd1 vssd1 vccd1 vccd1 _04808_ sky130_fd_sc_hd__and2b_1
XFILLER_0_106_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09239_ _03725_ genblk1\[0\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 _03848_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_133_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12250_ _05985_ vssd1 vssd1 vccd1 vccd1 _01009_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08206__B2 _02362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11201_ _05241_ vssd1 vssd1 vccd1 vccd1 _00704_ sky130_fd_sc_hd__clkbuf_1
X_12181_ _05816_ _05919_ _05921_ _05818_ net748 vssd1 vssd1 vccd1 vccd1 _01004_ sky130_fd_sc_hd__a32o_1
XANTENNA__07965__B1 _01675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11132_ _05176_ _05190_ _05191_ vssd1 vssd1 vccd1 vccd1 _05192_ sky130_fd_sc_hd__a21o_1
Xhold990 genblk2\[9\].wave_shpr.div.b1\[5\] vssd1 vssd1 vccd1 vccd1 net1208 sky130_fd_sc_hd__dlygate4sd3_1
X_11063_ genblk2\[6\].wave_shpr.div.acc\[17\] _05136_ _05022_ vssd1 vssd1 vccd1 vccd1
+ _05137_ sky130_fd_sc_hd__mux2_1
XANTENNA__08050__B _01355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10014_ _04363_ _04408_ _04409_ vssd1 vssd1 vccd1 vccd1 _04410_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08390__B1 _02011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_25_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06786__A _01489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11965_ _05786_ vssd1 vssd1 vccd1 vccd1 _05787_ sky130_fd_sc_hd__clkbuf_8
X_13704_ clknet_leaf_37_clk _01015_ net113 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.b1\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10916_ net1286 _01797_ _05042_ vssd1 vssd1 vccd1 vccd1 _05043_ sky130_fd_sc_hd__mux2_1
XANTENNA__10101__A _04269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11896_ _05722_ vssd1 vssd1 vccd1 vccd1 _00918_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13635_ clknet_leaf_69_clk _00948_ net212 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.b1\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_132_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10847_ _04979_ _04989_ _04990_ vssd1 vssd1 vccd1 vccd1 _04991_ sky130_fd_sc_hd__a21o_1
XFILLER_0_66_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13566_ clknet_leaf_56_clk net305 net182 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.quo\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10778_ _04813_ _04935_ vssd1 vssd1 vccd1 vccd1 _04936_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_26_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07410__A _02154_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_630 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_168 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12517_ clknet_leaf_105_clk PWM.next_counter\[1\] net155 vssd1 vssd1 vccd1 vccd1
+ PWM.counter\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_136_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13497_ clknet_leaf_86_clk net618 net178 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.quo\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12448_ clknet_leaf_105_clk _00027_ net153 vssd1 vssd1 vccd1 vccd1 sig_norm.i\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_22_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_140_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12379_ net876 _06039_ _06040_ _06056_ vssd1 vssd1 vccd1 vccd1 _01067_ sky130_fd_sc_hd__a22o_1
XFILLER_0_10_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06940_ net28 _01781_ vssd1 vssd1 vccd1 vccd1 _01782_ sky130_fd_sc_hd__nor2_1
XANTENNA__07971__A3 _01362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06871_ net493 _01724_ vssd1 vssd1 vccd1 vccd1 genblk1\[5\].osc.clkdiv_C.next_cnt\[17\]
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__08381__B1 _02336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08610_ _03314_ _03315_ _02789_ vssd1 vssd1 vccd1 vccd1 _03317_ sky130_fd_sc_hd__or3_1
X_09590_ _03983_ _04093_ vssd1 vssd1 vccd1 vccd1 _04094_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07222__A2_N _02001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08541_ genblk2\[8\].wave_shpr.div.fin_quo\[0\] _02526_ _02308_ genblk2\[8\].wave_shpr.div.fin_quo\[1\]
+ _02636_ vssd1 vssd1 vccd1 vccd1 _03248_ sky130_fd_sc_hd__a221o_1
XFILLER_0_49_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08472_ genblk2\[5\].wave_shpr.div.fin_quo\[3\] _03178_ _02526_ vssd1 vssd1 vccd1
+ vccd1 _03179_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07423_ _02164_ vssd1 vssd1 vccd1 vccd1 _00008_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout147_A net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07354_ genblk1\[11\].osc.clkdiv_C.cnt\[6\] _02108_ vssd1 vssd1 vccd1 vccd1 _02112_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_116_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10243__A1 _04454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06305_ genblk1\[0\].osc.clkdiv_C.cnt\[3\] _01227_ _01236_ _01266_ vssd1 vssd1 vccd1
+ vccd1 _01267_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07285_ net1119 _02052_ _02054_ vssd1 vssd1 vccd1 vccd1 genblk1\[10\].osc.clkdiv_C.next_cnt\[12\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_5_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_127 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09024_ _02203_ vssd1 vssd1 vccd1 vccd1 _03696_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_131_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06236_ _01174_ genblk1\[0\].osc.clkdiv_C.cnt\[6\] vssd1 vssd1 vccd1 vccd1 _01198_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_115_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11777__A _04676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold220 genblk2\[11\].wave_shpr.div.quo\[22\] vssd1 vssd1 vccd1 vccd1 net438 sky130_fd_sc_hd__dlygate4sd3_1
X_06167_ _01129_ _01138_ vssd1 vssd1 vccd1 vccd1 _01139_ sky130_fd_sc_hd__or2_1
Xhold231 genblk2\[2\].wave_shpr.div.quo\[6\] vssd1 vssd1 vccd1 vccd1 net449 sky130_fd_sc_hd__dlygate4sd3_1
Xhold242 genblk2\[1\].wave_shpr.div.quo\[8\] vssd1 vssd1 vccd1 vccd1 net460 sky130_fd_sc_hd__dlygate4sd3_1
Xhold253 genblk2\[5\].wave_shpr.div.quo\[22\] vssd1 vssd1 vccd1 vccd1 net471 sky130_fd_sc_hd__dlygate4sd3_1
Xhold264 genblk2\[8\].wave_shpr.div.quo\[12\] vssd1 vssd1 vccd1 vccd1 net482 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold275 genblk1\[5\].osc.clkdiv_C.cnt\[17\] vssd1 vssd1 vccd1 vccd1 net493 sky130_fd_sc_hd__dlygate4sd3_1
Xhold286 genblk2\[11\].wave_shpr.div.quo\[21\] vssd1 vssd1 vccd1 vccd1 net504 sky130_fd_sc_hd__dlygate4sd3_1
Xhold297 genblk2\[6\].wave_shpr.div.quo\[8\] vssd1 vssd1 vccd1 vccd1 net515 sky130_fd_sc_hd__dlygate4sd3_1
X_09926_ genblk2\[2\].wave_shpr.div.acc\[25\] genblk2\[2\].wave_shpr.div.acc\[24\]
+ genblk2\[2\].wave_shpr.div.acc\[26\] _04212_ vssd1 vssd1 vccd1 vccd1 _04335_ sky130_fd_sc_hd__nor4_1
XANTENNA__12299__A2 _06009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09857_ _04247_ vssd1 vssd1 vccd1 vccd1 _04282_ sky130_fd_sc_hd__clkbuf_4
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08808_ _03217_ _03510_ _03442_ _03443_ vssd1 vssd1 vccd1 vccd1 _03515_ sky130_fd_sc_hd__o211a_1
X_09788_ _04244_ vssd1 vssd1 vccd1 vccd1 _00288_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12401__A _03941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11259__B1 _05249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08739_ _03443_ _03444_ _03428_ _03420_ vssd1 vssd1 vccd1 vccd1 _03446_ sky130_fd_sc_hd__a211oi_2
XTAP_2425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08124__B1 _01304_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11750_ genblk2\[9\].wave_shpr.div.quo\[5\] _05623_ _05624_ net586 vssd1 vssd1 vccd1
+ vccd1 _00870_ sky130_fd_sc_hd__a22o_1
XTAP_1724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10701_ _04869_ genblk1\[5\].osc.clkdiv_C.cnt\[16\] vssd1 vssd1 vccd1 vccd1 _04878_
+ sky130_fd_sc_hd__and2_1
XTAP_1757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11681_ genblk2\[9\].wave_shpr.div.acc\[0\] vssd1 vssd1 vccd1 vccd1 _05573_ sky130_fd_sc_hd__inv_2
XFILLER_0_154_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13420_ clknet_leaf_91_clk _00739_ net147 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.acc\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10632_ genblk2\[6\].wave_shpr.div.b1\[9\] _01923_ _04834_ vssd1 vssd1 vccd1 vccd1
+ _04843_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_153_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10563_ _04775_ _04789_ _04790_ vssd1 vssd1 vccd1 vccd1 _04791_ sky130_fd_sc_hd__a21o_1
X_13351_ clknet_leaf_5_clk _00672_ net47 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.acc\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_855 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11982__A1 _01441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_691 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12302_ genblk2\[11\].wave_shpr.div.quo\[3\] _06009_ _06010_ net402 vssd1 vssd1 vccd1
+ vccd1 _01036_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10494_ _04615_ _04735_ vssd1 vssd1 vccd1 vccd1 _04736_ sky130_fd_sc_hd__xnor2_1
X_13282_ clknet_leaf_117_clk _00603_ net137 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.fin_quo\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_122_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12233_ genblk2\[11\].wave_shpr.div.b1\[15\] genblk2\[11\].wave_shpr.div.acc\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05971_ sky130_fd_sc_hd__and2b_1
XFILLER_0_32_683 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12164_ genblk2\[10\].wave_shpr.div.acc\[22\] _05908_ genblk2\[10\].wave_shpr.div.acc\[23\]
+ vssd1 vssd1 vccd1 vccd1 _05910_ sky130_fd_sc_hd__or3b_1
X_11115_ genblk2\[7\].wave_shpr.div.acc\[6\] genblk2\[7\].wave_shpr.div.b1\[6\] vssd1
+ vssd1 vccd1 vccd1 _05175_ sky130_fd_sc_hd__or2b_1
XANTENNA__13548__RESET_B net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12095_ genblk2\[10\].wave_shpr.div.acc\[5\] _05858_ _05787_ vssd1 vssd1 vccd1 vccd1
+ _05859_ sky130_fd_sc_hd__mux2_1
X_11046_ _05007_ _05123_ vssd1 vssd1 vccd1 vccd1 _05124_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11498__B1 _05446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07405__A _02147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12997_ clknet_leaf_132_clk _00326_ net60 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.acc\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07124__B _01355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11948_ genblk2\[10\].wave_shpr.div.b1\[12\] genblk2\[10\].wave_shpr.div.acc\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05770_ sky130_fd_sc_hd__and2b_1
X_11879_ net556 _05684_ _05685_ _05711_ vssd1 vssd1 vccd1 vccd1 _00912_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13618_ clknet_leaf_84_clk _00931_ net204 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.b1\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08236__A net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_403 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13549_ clknet_leaf_110_clk _00864_ net152 vssd1 vssd1 vccd1 vccd1 sig_norm.b1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07070_ net1092 _01887_ vssd1 vssd1 vccd1 vccd1 genblk1\[8\].osc.clkdiv_C.next_cnt\[0\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_140_611 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_11_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09067__A _02155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06601__B1 _01508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07972_ _02672_ _02673_ _02678_ vssd1 vssd1 vccd1 vccd1 _02679_ sky130_fd_sc_hd__o21ai_2
X_09711_ genblk2\[2\].wave_shpr.div.b1\[9\] genblk2\[2\].wave_shpr.div.acc\[9\] vssd1
+ vssd1 vccd1 vccd1 _04191_ sky130_fd_sc_hd__and2b_1
X_06923_ genblk1\[6\].osc.clkdiv_C.cnt\[6\] _01768_ vssd1 vssd1 vccd1 vccd1 _01771_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__06227__B1_N _01188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09642_ genblk2\[1\].wave_shpr.div.acc\[19\] _04130_ vssd1 vssd1 vccd1 vccd1 _04134_
+ sky130_fd_sc_hd__nand2_1
X_06854_ _01693_ _01713_ _01714_ vssd1 vssd1 vccd1 vccd1 genblk1\[5\].osc.clkdiv_C.next_cnt\[11\]
+ sky130_fd_sc_hd__nor3_1
XANTENNA__10700__A2 _02183_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06785_ genblk1\[5\].osc.clkdiv_C.cnt\[4\] _01483_ vssd1 vssd1 vccd1 vccd1 _01657_
+ sky130_fd_sc_hd__xnor2_1
X_09573_ _03976_ _03968_ vssd1 vssd1 vccd1 vccd1 _04081_ sky130_fd_sc_hd__or2b_1
XTAP_1009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08524_ _02216_ _02552_ genblk2\[9\].wave_shpr.div.fin_quo\[0\] vssd1 vssd1 vccd1
+ vccd1 _03231_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07034__B _01359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09530__A _03707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08455_ _03159_ _03160_ _03161_ _02694_ vssd1 vssd1 vccd1 vccd1 _03162_ sky130_fd_sc_hd__a211o_1
XANTENNA__10676__A _04672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07406_ _02151_ vssd1 vssd1 vccd1 vccd1 _00000_ sky130_fd_sc_hd__inv_2
X_08386_ _01200_ genblk1\[2\].osc.clkdiv_C.cnt\[4\] genblk1\[2\].osc.clkdiv_C.cnt\[5\]
+ _01441_ vssd1 vssd1 vccd1 vccd1 _03093_ sky130_fd_sc_hd__a211o_1
XFILLER_0_133_92 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07337_ genblk1\[11\].osc.clkdiv_C.cnt\[1\] genblk1\[11\].osc.clkdiv_C.cnt\[0\] genblk1\[11\].osc.clkdiv_C.cnt\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02099_ sky130_fd_sc_hd__a21o_1
XFILLER_0_151_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_33_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07268_ genblk1\[10\].osc.clkdiv_C.cnt\[7\] _02041_ vssd1 vssd1 vccd1 vccd1 _02043_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07632__A2 _01262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09007_ _03683_ vssd1 vssd1 vccd1 vccd1 _00068_ sky130_fd_sc_hd__clkbuf_1
X_06219_ _01174_ vssd1 vssd1 vccd1 vccd1 _01181_ sky130_fd_sc_hd__buf_6
XFILLER_0_104_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10615__S _04637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07199_ genblk1\[9\].osc.clkdiv_C.cnt\[14\] _01981_ _01984_ vssd1 vssd1 vccd1 vccd1
+ genblk1\[9\].osc.clkdiv_C.next_cnt\[14\] sky130_fd_sc_hd__o21a_1
XFILLER_0_60_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08593__B1 _02361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07209__B _01564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09909_ _04250_ vssd1 vssd1 vccd1 vccd1 _04322_ sky130_fd_sc_hd__clkbuf_4
X_12920_ clknet_leaf_35_clk _00251_ net118 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.acc\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12851_ clknet_leaf_118_clk _00182_ net138 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.fin_quo\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_2211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06371__A2 _01311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11802_ _03693_ vssd1 vssd1 vccd1 vccd1 _05653_ sky130_fd_sc_hd__clkbuf_4
XTAP_2244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12782_ clknet_leaf_40_clk _00115_ net117 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.b1\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_68_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11733_ _05619_ vssd1 vssd1 vccd1 vccd1 _00858_ sky130_fd_sc_hd__clkbuf_1
XTAP_1554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11652__B1 _05448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_22_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11664_ genblk2\[9\].wave_shpr.div.acc\[15\] genblk2\[9\].wave_shpr.div.b1\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05556_ sky130_fd_sc_hd__or2b_1
XFILLER_0_52_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13403_ clknet_leaf_92_clk _00722_ net147 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.quo\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10615_ genblk2\[6\].wave_shpr.div.b1\[2\] _01684_ _04637_ vssd1 vssd1 vccd1 vccd1
+ _04833_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_4_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11595_ _05441_ vssd1 vssd1 vccd1 vccd1 _05507_ sky130_fd_sc_hd__clkbuf_4
X_13334_ clknet_leaf_6_clk _00655_ net48 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.acc\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10546_ genblk2\[5\].wave_shpr.div.acc\[6\] genblk2\[5\].wave_shpr.div.b1\[6\] vssd1
+ vssd1 vccd1 vccd1 _04774_ sky130_fd_sc_hd__or2b_1
XFILLER_0_51_266 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_121_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13265_ clknet_leaf_0_clk _00588_ net38 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.acc\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10477_ _04608_ _04569_ vssd1 vssd1 vccd1 vccd1 _04723_ sky130_fd_sc_hd__or2b_1
XFILLER_0_20_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12216_ _05936_ _05952_ _05953_ vssd1 vssd1 vccd1 vccd1 _05954_ sky130_fd_sc_hd__a21o_1
XFILLER_0_122_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13196_ clknet_leaf_114_clk _00519_ net134 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.fin_quo\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_103_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_138_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12147_ net590 _05876_ _05883_ _05898_ vssd1 vssd1 vccd1 vccd1 _00993_ sky130_fd_sc_hd__a22o_1
XANTENNA__07119__B _01227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09615__A _04046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07139__A1 genblk1\[9\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12078_ genblk2\[10\].wave_shpr.div.acc\[1\] _05845_ _05787_ vssd1 vssd1 vccd1 vccd1
+ _05846_ sky130_fd_sc_hd__mux2_1
X_11029_ _04999_ _05110_ vssd1 vssd1 vccd1 vccd1 _05111_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07899__A1_N _01181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06570_ genblk1\[2\].osc.clkdiv_C.cnt\[16\] _01478_ vssd1 vssd1 vccd1 vccd1 _01480_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_86_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07789__B _01263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09851__A3 _04214_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08240_ _02682_ _02689_ _02683_ vssd1 vssd1 vccd1 vccd1 _02947_ sky130_fd_sc_hd__o21a_1
XFILLER_0_117_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_144_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08171_ _02861_ _02862_ _02865_ _02876_ _02877_ vssd1 vssd1 vccd1 vccd1 _02878_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_133_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07122_ genblk1\[9\].osc.clkdiv_C.cnt\[6\] _01334_ _01328_ genblk1\[9\].osc.clkdiv_C.cnt\[13\]
+ _01921_ vssd1 vssd1 vccd1 vccd1 _01922_ sky130_fd_sc_hd__o221a_1
XANTENNA__07614__A2 _01192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_789 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07053_ genblk1\[8\].osc.clkdiv_C.cnt\[12\] _01869_ _01870_ genblk1\[8\].osc.clkdiv_C.cnt\[11\]
+ vssd1 vssd1 vccd1 vccd1 _01871_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_3_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_113_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10382__B1 _04655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07955_ _02661_ _02653_ _02652_ vssd1 vssd1 vccd1 vccd1 _02662_ sky130_fd_sc_hd__or3b_1
X_06906_ _01675_ _01727_ _01737_ _01756_ _01759_ vssd1 vssd1 vccd1 vccd1 _01760_ sky130_fd_sc_hd__a2111oi_1
XANTENNA__10134__B1 _04455_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07886_ genblk2\[1\].wave_shpr.div.fin_quo\[7\] _02539_ _02591_ _02592_ vssd1 vssd1
+ vccd1 vccd1 _02593_ sky130_fd_sc_hd__a22o_1
X_09625_ _03999_ _04120_ vssd1 vssd1 vccd1 vccd1 _04121_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06837_ genblk1\[5\].osc.clkdiv_C.cnt\[4\] _01700_ genblk1\[5\].osc.clkdiv_C.cnt\[5\]
+ vssd1 vssd1 vccd1 vccd1 _01704_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_78_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09556_ _03707_ vssd1 vssd1 vccd1 vccd1 _04069_ sky130_fd_sc_hd__clkbuf_4
X_06768_ genblk1\[4\].osc.clkdiv_C.cnt\[13\] _01641_ vssd1 vssd1 vccd1 vccd1 _01645_
+ sky130_fd_sc_hd__or2_1
XANTENNA__06884__A _01241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08507_ _03114_ _03213_ _03122_ vssd1 vssd1 vccd1 vccd1 _03214_ sky130_fd_sc_hd__o21a_1
XFILLER_0_93_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09487_ net1304 _04032_ _04024_ vssd1 vssd1 vccd1 vccd1 _04033_ sky130_fd_sc_hd__mux2_1
X_06699_ _01320_ _01321_ vssd1 vssd1 vccd1 vccd1 _01589_ sky130_fd_sc_hd__nand2_4
X_08438_ _03141_ _03144_ _02901_ vssd1 vssd1 vccd1 vccd1 _03145_ sky130_fd_sc_hd__o21a_1
XFILLER_0_108_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09055__A1 _03704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08369_ _03052_ _03053_ _03030_ _03051_ vssd1 vssd1 vccd1 vccd1 _03076_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_150_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10400_ net531 _04661_ _04663_ genblk2\[4\].wave_shpr.div.quo\[16\] _04668_ vssd1
+ vssd1 vccd1 vccd1 _00476_ sky130_fd_sc_hd__a221o_1
XANTENNA__07066__B1 _01870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11380_ net328 _05356_ _03855_ vssd1 vssd1 vccd1 vccd1 _05357_ sky130_fd_sc_hd__o21ai_1
XANTENNA__08604__A _02261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07053__A2_N _01869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10331_ _04633_ _01304_ _03689_ vssd1 vssd1 vccd1 vccd1 _04634_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10345__S _04637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10262_ genblk2\[4\].wave_shpr.div.acc\[8\] genblk2\[4\].wave_shpr.div.b1\[8\] vssd1
+ vssd1 vccd1 vccd1 _04574_ sky130_fd_sc_hd__or2b_1
X_13050_ clknet_leaf_113_clk net327 net128 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.quo\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12001_ _05805_ vssd1 vssd1 vccd1 vccd1 _00940_ sky130_fd_sc_hd__clkbuf_1
X_10193_ _04405_ _04365_ vssd1 vssd1 vccd1 vccd1 _04523_ sky130_fd_sc_hd__or2b_1
XANTENNA__11190__B1_N _04241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12903_ clknet_leaf_37_clk net753 net104 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.acc\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12834_ clknet_leaf_64_clk _00167_ net196 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.acc\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2030 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06794__A _01440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2041 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2052 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2063 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2074 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12765_ clknet_leaf_93_clk _00098_ net146 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.fin_quo\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_2085 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2096 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11716_ genblk2\[9\].wave_shpr.div.acc\[18\] _05607_ vssd1 vssd1 vccd1 vccd1 _05608_
+ sky130_fd_sc_hd__or2_1
XTAP_1395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_596 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12696_ clknet_leaf_54_clk genblk1\[8\].osc.clkdiv_C.next_cnt\[9\] net172 vssd1 vssd1
+ vccd1 vccd1 genblk1\[8\].osc.clkdiv_C.cnt\[9\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_154_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11647_ net615 _05448_ _05445_ _05544_ vssd1 vssd1 vccd1 vccd1 _00847_ sky130_fd_sc_hd__a22o_1
Xinput13 pb[7] vssd1 vssd1 vccd1 vccd1 net13 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_141_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_13_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11578_ net950 _05447_ _05484_ _05494_ vssd1 vssd1 vccd1 vccd1 _00828_ sky130_fd_sc_hd__a22o_1
XFILLER_0_107_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06960__C _01514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13317_ clknet_leaf_24_clk net345 net88 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.quo\[11\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold808 genblk2\[9\].wave_shpr.div.acc\[24\] vssd1 vssd1 vccd1 vccd1 net1026 sky130_fd_sc_hd__dlygate4sd3_1
Xhold819 genblk2\[5\].wave_shpr.div.acc\[7\] vssd1 vssd1 vccd1 vccd1 net1037 sky130_fd_sc_hd__dlygate4sd3_1
X_10529_ _04655_ _04757_ _04759_ _04657_ net734 vssd1 vssd1 vccd1 vccd1 _00514_ sky130_fd_sc_hd__a32o_1
XANTENNA__08233__B _02885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13248_ clknet_leaf_13_clk net911 net52 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.acc\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_149_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08557__B1 genblk2\[8\].wave_shpr.div.fin_quo\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13179_ clknet_leaf_131_clk _00504_ net65 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.acc\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08021__A2 _01577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06969__A _01179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07740_ genblk1\[1\].osc.clkdiv_C.cnt\[9\] _01334_ _01356_ genblk1\[1\].osc.clkdiv_C.cnt\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02447_ sky130_fd_sc_hd__o22a_1
XANTENNA_clkbuf_leaf_74_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09521__A2 _04048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07671_ _01308_ genblk1\[10\].osc.clkdiv_C.cnt\[1\] vssd1 vssd1 vccd1 vccd1 _02378_
+ sky130_fd_sc_hd__and2_1
X_09410_ genblk2\[1\].wave_shpr.div.b1\[2\] genblk2\[1\].wave_shpr.div.acc\[2\] vssd1
+ vssd1 vccd1 vccd1 _03974_ sky130_fd_sc_hd__and2b_1
X_06622_ genblk1\[3\].osc.clkdiv_C.cnt\[2\] genblk1\[3\].osc.clkdiv_C.cnt\[1\] genblk1\[3\].osc.clkdiv_C.cnt\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01528_ sky130_fd_sc_hd__and3_1
X_09341_ net786 _03903_ _03910_ _03919_ vssd1 vssd1 vccd1 vccd1 _00166_ sky130_fd_sc_hd__a22o_1
X_06553_ _01451_ _01468_ vssd1 vssd1 vccd1 vccd1 _01469_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_8_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_89_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06484_ genblk1\[2\].osc.clkdiv_C.cnt\[3\] vssd1 vssd1 vccd1 vccd1 _01410_ sky130_fd_sc_hd__inv_2
XFILLER_0_75_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09272_ _03865_ _03866_ net1066 _03836_ vssd1 vssd1 vccd1 vccd1 _00150_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_23_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_132_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08223_ genblk2\[5\].wave_shpr.div.fin_quo\[6\] _02308_ _02791_ vssd1 vssd1 vccd1
+ vccd1 _02930_ sky130_fd_sc_hd__a21o_1
XFILLER_0_117_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09037__A1 _03704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10954__A _04676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07048__B1 _01336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12041__B1 _05816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_12_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08154_ _02858_ _02859_ _02860_ vssd1 vssd1 vccd1 vccd1 _02861_ sky130_fd_sc_hd__a21o_1
XFILLER_0_132_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_244 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07105_ genblk1\[8\].osc.clkdiv_C.cnt\[13\] genblk1\[8\].osc.clkdiv_C.cnt\[12\] _01906_
+ vssd1 vssd1 vccd1 vccd1 _01910_ sky130_fd_sc_hd__and3_1
XFILLER_0_125_290 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08085_ genblk2\[5\].wave_shpr.div.fin_quo\[0\] genblk2\[5\].wave_shpr.div.fin_quo\[1\]
+ genblk2\[5\].wave_shpr.div.fin_quo\[2\] genblk2\[5\].wave_shpr.div.fin_quo\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02792_ sky130_fd_sc_hd__or4_1
XANTENNA__09239__B genblk1\[0\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07036_ genblk1\[8\].osc.clkdiv_C.cnt\[16\] _01853_ _01578_ vssd1 vssd1 vccd1 vccd1
+ _01854_ sky130_fd_sc_hd__o21a_1
XFILLER_0_113_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_27_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09255__A _03853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08987_ _03134_ _03135_ vssd1 vssd1 vccd1 vccd1 _03671_ sky130_fd_sc_hd__nor2_1
XANTENNA__06598__B _01197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_4_5_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_5_0_clk sky130_fd_sc_hd__clkbuf_8
X_07938_ genblk2\[8\].wave_shpr.div.fin_quo\[7\] _02539_ _02636_ _02644_ vssd1 vssd1
+ vccd1 vccd1 _02645_ sky130_fd_sc_hd__a211o_1
XANTENNA__09512__A2 _04043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07869_ genblk2\[0\].wave_shpr.div.fin_quo\[0\] _02524_ _02307_ genblk2\[0\].wave_shpr.div.fin_quo\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02576_ sky130_fd_sc_hd__a22o_1
XANTENNA__11724__S _00023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09608_ net366 _04107_ _04095_ vssd1 vssd1 vccd1 vccd1 _04108_ sky130_fd_sc_hd__mux2_1
X_10880_ genblk2\[6\].wave_shpr.div.fin_quo\[0\] _05023_ _00017_ vssd1 vssd1 vccd1
+ vccd1 _05024_ sky130_fd_sc_hd__mux2_1
XANTENNA__07503__A _02223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09539_ net462 _04052_ _04053_ genblk2\[1\].wave_shpr.div.quo\[15\] _04060_ vssd1
+ vssd1 vccd1 vccd1 _00223_ sky130_fd_sc_hd__a221o_1
XANTENNA__08079__A2 _01355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09276__A1 _03839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12550_ clknet_leaf_60_clk genblk1\[0\].osc.clkdiv_C.next_cnt\[7\] net186 vssd1 vssd1
+ vccd1 vccd1 genblk1\[0\].osc.clkdiv_C.cnt\[7\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_136_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11501_ genblk2\[8\].wave_shpr.div.quo\[4\] _05442_ _05446_ net346 vssd1 vssd1 vccd1
+ vccd1 _00799_ sky130_fd_sc_hd__a22o_1
X_12481_ clknet_leaf_108_clk net1028 net151 vssd1 vssd1 vccd1 vccd1 sig_norm.acc\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11432_ genblk2\[8\].wave_shpr.div.b1\[17\] genblk2\[8\].wave_shpr.div.acc\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05408_ sky130_fd_sc_hd__and2b_1
XFILLER_0_80_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_21_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10075__S _04440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11363_ genblk2\[7\].wave_shpr.div.acc\[24\] _05273_ _05342_ vssd1 vssd1 vccd1 vccd1
+ _05346_ sky130_fd_sc_hd__or3b_1
XFILLER_0_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09864__S _04214_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13102_ clknet_leaf_118_clk _00013_ net139 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.done
+ sky130_fd_sc_hd__dfrtp_1
X_10314_ genblk2\[4\].wave_shpr.div.fin_quo\[1\] net1309 _00013_ vssd1 vssd1 vccd1
+ vccd1 _04625_ sky130_fd_sc_hd__mux2_1
X_11294_ net893 _05279_ _05283_ _05294_ vssd1 vssd1 vccd1 vccd1 _00744_ sky130_fd_sc_hd__a22o_1
XFILLER_0_131_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13033_ clknet_leaf_123_clk _00360_ net79 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.b1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_30_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10245_ genblk2\[3\].wave_shpr.div.i\[1\] genblk2\[3\].wave_shpr.div.i\[0\] genblk2\[3\].wave_shpr.div.i\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04560_ sky130_fd_sc_hd__and3_1
XANTENNA__08003__A2 _01666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10176_ _04396_ _04509_ vssd1 vssd1 vccd1 vccd1 _04510_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07762__A1 _02458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10104__A _04455_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout190 net198 vssd1 vssd1 vccd1 vccd1 net190 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06301__B _01262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12817_ clknet_leaf_59_clk _00150_ net193 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.acc\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_139_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12748_ clknet_leaf_50_clk genblk1\[11\].osc.clkdiv_C.next_cnt\[7\] net111 vssd1
+ vssd1 vccd1 vccd1 genblk1\[11\].osc.clkdiv_C.cnt\[7\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_29_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_44_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12679_ clknet_leaf_120_clk genblk1\[7\].osc.clkdiv_C.next_cnt\[10\] net82 vssd1
+ vssd1 vccd1 vccd1 genblk1\[7\].osc.clkdiv_C.cnt\[10\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_154_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12023__B1 _05817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold605 genblk2\[0\].wave_shpr.div.acc\[5\] vssd1 vssd1 vccd1 vccd1 net823 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold616 genblk2\[5\].wave_shpr.div.b1\[16\] vssd1 vssd1 vccd1 vccd1 net834 sky130_fd_sc_hd__dlygate4sd3_1
Xhold627 genblk2\[2\].wave_shpr.div.acc\[16\] vssd1 vssd1 vccd1 vccd1 net845 sky130_fd_sc_hd__dlygate4sd3_1
Xhold638 _04964_ vssd1 vssd1 vccd1 vccd1 net856 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_69_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold649 genblk2\[6\].wave_shpr.div.acc\[8\] vssd1 vssd1 vccd1 vccd1 net867 sky130_fd_sc_hd__dlygate4sd3_1
X_08910_ _03586_ net26 sig_norm.acc\[4\] vssd1 vssd1 vccd1 vccd1 _03612_ sky130_fd_sc_hd__o21ai_1
XANTENNA__11809__S _05613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_910 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09890_ genblk2\[2\].wave_shpr.div.acc\[9\] _04307_ _04301_ vssd1 vssd1 vccd1 vccd1
+ _04308_ sky130_fd_sc_hd__mux2_1
XTAP_921 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08841_ _03542_ _03544_ vssd1 vssd1 vccd1 vccd1 _03548_ sky130_fd_sc_hd__or2_1
XTAP_943 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_954 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_976 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_987 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08772_ _03477_ _03478_ vssd1 vssd1 vccd1 vccd1 _03479_ sky130_fd_sc_hd__xnor2_1
XTAP_998 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12626__RESET_B net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07307__B _01223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07723_ genblk1\[1\].osc.clkdiv_C.cnt\[2\] _01323_ _02429_ genblk1\[1\].osc.clkdiv_C.cnt\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02430_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07654_ _02307_ vssd1 vssd1 vccd1 vccd1 _02361_ sky130_fd_sc_hd__buf_4
XFILLER_0_149_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_94_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_88_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06605_ _01512_ vssd1 vssd1 vccd1 vccd1 _01513_ sky130_fd_sc_hd__clkbuf_4
X_07585_ genblk1\[9\].osc.clkdiv_C.cnt\[3\] _01311_ _02290_ _02291_ vssd1 vssd1 vccd1
+ vccd1 _02292_ sky130_fd_sc_hd__a22o_1
X_09324_ net920 _03903_ _03877_ _03906_ vssd1 vssd1 vccd1 vccd1 _00162_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06536_ genblk1\[2\].osc.clkdiv_C.cnt\[4\] _01456_ vssd1 vssd1 vccd1 vccd1 _01458_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_118_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09255_ _03853_ genblk1\[0\].osc.clkdiv_C.cnt\[11\] vssd1 vssd1 vccd1 vccd1 _03857_
+ sky130_fd_sc_hd__and2_1
XANTENNA__10684__A _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06467_ genblk1\[1\].osc.clkdiv_C.cnt\[12\] _01398_ vssd1 vssd1 vccd1 vccd1 _01399_
+ sky130_fd_sc_hd__and2_1
XANTENNA__06881__B _01678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08206_ _02911_ _02912_ genblk2\[9\].wave_shpr.div.fin_quo\[6\] _02362_ vssd1 vssd1
+ vccd1 vccd1 _02913_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_145_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09186_ _03704_ net651 _03820_ vssd1 vssd1 vccd1 vccd1 _00110_ sky130_fd_sc_hd__a21o_1
X_06398_ _01188_ vssd1 vssd1 vccd1 vccd1 _01342_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_31_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08137_ genblk2\[4\].wave_shpr.div.fin_quo\[6\] _02843_ vssd1 vssd1 vccd1 vccd1 _02844_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08068_ _01196_ _01254_ genblk1\[5\].osc.clkdiv_C.cnt\[3\] vssd1 vssd1 vccd1 vccd1
+ _02775_ sky130_fd_sc_hd__o21a_1
XFILLER_0_12_770 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07019_ _01822_ _01842_ vssd1 vssd1 vccd1 vccd1 _01843_ sky130_fd_sc_hd__nor2_1
X_10030_ _04424_ vssd1 vssd1 vccd1 vccd1 _00350_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07744__A1 genblk1\[1\].osc.clkdiv_C.cnt\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11540__A2 _05441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07744__B2 genblk1\[1\].osc.clkdiv_C.cnt\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11981_ _05795_ vssd1 vssd1 vccd1 vccd1 _00930_ sky130_fd_sc_hd__clkbuf_1
X_13720_ clknet_leaf_39_clk _01031_ net115 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.b1\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10932_ _05050_ vssd1 vssd1 vccd1 vccd1 _00626_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_98_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13651_ clknet_leaf_41_clk _00964_ net116 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.quo\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_79_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10863_ _04971_ _05005_ _05006_ vssd1 vssd1 vccd1 vccd1 _05007_ sky130_fd_sc_hd__a21o_1
XFILLER_0_128_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12602_ clknet_leaf_21_clk genblk1\[3\].osc.clkdiv_C.next_cnt\[5\] net95 vssd1 vssd1
+ vccd1 vccd1 genblk1\[3\].osc.clkdiv_C.cnt\[5\] sky130_fd_sc_hd__dfrtp_4
XPHY_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13582_ clknet_leaf_76_clk _00897_ net207 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.acc\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10794_ _04818_ _04819_ vssd1 vssd1 vccd1 vccd1 _04947_ sky130_fd_sc_hd__and2b_1
XPHY_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12533_ clknet_leaf_61_clk _00085_ net186 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.b1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06791__B _01578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12464_ clknet_leaf_103_clk _00037_ net156 vssd1 vssd1 vccd1 vccd1 PWM.final_sample_in\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11415_ _05367_ _05389_ _05390_ vssd1 vssd1 vccd1 vccd1 _05391_ sky130_fd_sc_hd__a21o_1
X_12395_ net875 _06039_ _06040_ _06068_ vssd1 vssd1 vccd1 vccd1 _01071_ sky130_fd_sc_hd__a22o_1
XFILLER_0_50_843 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_417 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11346_ genblk2\[7\].wave_shpr.div.acc\[19\] _05331_ vssd1 vssd1 vccd1 vccd1 _05334_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_120_720 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11277_ genblk2\[7\].wave_shpr.div.acc\[2\] _05281_ _05222_ vssd1 vssd1 vccd1 vccd1
+ _05282_ sky130_fd_sc_hd__mux2_1
XANTENNA__12314__A _03942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09185__B1 _03819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13016_ clknet_leaf_121_clk _00011_ net77 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.done
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07408__A _02152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10228_ net1000 _04457_ _04522_ _04548_ vssd1 vssd1 vccd1 vccd1 _00424_ sky130_fd_sc_hd__a22o_1
XFILLER_0_146_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10159_ _04496_ _04388_ vssd1 vssd1 vccd1 vccd1 _04497_ sky130_fd_sc_hd__xnor2_1
Xhold2 genblk2\[10\].wave_shpr.div.quo\[1\] vssd1 vssd1 vccd1 vccd1 net220 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_89_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10098__A2 _04457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07143__A genblk1\[9\].osc.clkdiv_C.cnt\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07370_ genblk1\[11\].osc.clkdiv_C.cnt\[9\] _02119_ vssd1 vssd1 vccd1 vccd1 _02125_
+ sky130_fd_sc_hd__or2_1
X_06321_ net1133 _01276_ _01278_ vssd1 vssd1 vccd1 vccd1 genblk1\[0\].osc.clkdiv_C.next_cnt\[4\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_127_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06252_ _01187_ _01188_ vssd1 vssd1 vccd1 vccd1 _01214_ sky130_fd_sc_hd__nand2b_4
X_09040_ _03707_ vssd1 vssd1 vccd1 vccd1 _03708_ sky130_fd_sc_hd__buf_8
XFILLER_0_60_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06183_ _01099_ _01150_ _01154_ vssd1 vssd1 vccd1 vccd1 _00025_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_143_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold402 genblk2\[6\].wave_shpr.div.quo\[13\] vssd1 vssd1 vccd1 vccd1 net620 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold413 genblk2\[3\].wave_shpr.div.quo\[10\] vssd1 vssd1 vccd1 vccd1 net631 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold424 PWM.counter\[1\] vssd1 vssd1 vccd1 vccd1 net642 sky130_fd_sc_hd__dlygate4sd3_1
Xhold435 genblk2\[0\].wave_shpr.div.acc\[23\] vssd1 vssd1 vccd1 vccd1 net653 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_887 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold446 genblk2\[1\].wave_shpr.div.acc\[18\] vssd1 vssd1 vccd1 vccd1 net664 sky130_fd_sc_hd__dlygate4sd3_1
Xhold457 genblk2\[4\].wave_shpr.div.quo\[12\] vssd1 vssd1 vccd1 vccd1 net675 sky130_fd_sc_hd__dlygate4sd3_1
Xhold468 genblk2\[9\].wave_shpr.div.quo\[2\] vssd1 vssd1 vccd1 vccd1 net686 sky130_fd_sc_hd__dlygate4sd3_1
X_09942_ _04212_ _04335_ vssd1 vssd1 vccd1 vccd1 _04346_ sky130_fd_sc_hd__nor2_1
Xhold479 _00296_ vssd1 vssd1 vccd1 vccd1 net697 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_461 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09873_ genblk2\[2\].wave_shpr.div.acc\[5\] _04294_ _04214_ vssd1 vssd1 vccd1 vccd1
+ _04295_ sky130_fd_sc_hd__mux2_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08824_ _03482_ _03529_ _03530_ vssd1 vssd1 vccd1 vccd1 _03531_ sky130_fd_sc_hd__or3_1
Xhold1102 genblk2\[6\].wave_shpr.div.quo\[2\] vssd1 vssd1 vccd1 vccd1 net1320 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1113 genblk2\[8\].wave_shpr.div.quo\[0\] vssd1 vssd1 vccd1 vccd1 net1331 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07037__B _01564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1124 genblk2\[5\].wave_shpr.div.quo\[0\] vssd1 vssd1 vccd1 vccd1 net1342 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08755_ _03232_ _03233_ vssd1 vssd1 vccd1 vccd1 _03462_ sky130_fd_sc_hd__nor2_1
XANTENNA__06876__B net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10089__A2 _04452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07706_ genblk2\[10\].wave_shpr.div.fin_quo\[4\] genblk2\[10\].wave_shpr.div.fin_quo\[5\]
+ _02404_ _02409_ _02412_ vssd1 vssd1 vccd1 vccd1 _02413_ sky130_fd_sc_hd__o41a_1
XTAP_2629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08686_ _03386_ _03392_ vssd1 vssd1 vccd1 vccd1 _03393_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_67_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07637_ _02338_ _02340_ _02341_ _02342_ vssd1 vssd1 vccd1 vccd1 _02344_ sky130_fd_sc_hd__o2bb2a_1
XTAP_1939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_138_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07568_ genblk1\[9\].osc.clkdiv_C.cnt\[14\] _01349_ _01246_ genblk1\[9\].osc.clkdiv_C.cnt\[13\]
+ vssd1 vssd1 vccd1 vccd1 _02275_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_0_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09307_ net956 _03870_ _03877_ _03893_ vssd1 vssd1 vccd1 vccd1 _00158_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06519_ genblk1\[2\].osc.clkdiv_C.cnt\[7\] _01433_ _01418_ genblk1\[2\].osc.clkdiv_C.cnt\[4\]
+ vssd1 vssd1 vccd1 vccd1 _01445_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_119_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10618__S _04834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07499_ net18 net17 vssd1 vssd1 vccd1 vccd1 _02220_ sky130_fd_sc_hd__or2b_1
XFILLER_0_63_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09238_ _03838_ vssd1 vssd1 vccd1 vccd1 _03847_ sky130_fd_sc_hd__buf_2
XFILLER_0_35_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_134_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_44_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09169_ genblk2\[0\].wave_shpr.div.fin_quo\[6\] net652 _00001_ vssd1 vssd1 vccd1
+ vccd1 _03811_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11200_ genblk2\[8\].wave_shpr.div.b1\[11\] _01565_ _05237_ vssd1 vssd1 vccd1 vccd1
+ _05241_ sky130_fd_sc_hd__mux2_1
X_12180_ _05920_ vssd1 vssd1 vccd1 vccd1 _05921_ sky130_fd_sc_hd__inv_2
XFILLER_0_102_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_102_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11131_ genblk2\[7\].wave_shpr.div.b1\[5\] genblk2\[7\].wave_shpr.div.acc\[5\] vssd1
+ vssd1 vccd1 vccd1 _05191_ sky130_fd_sc_hd__and2b_1
Xhold980 _04222_ vssd1 vssd1 vccd1 vccd1 net1198 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_8_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold991 genblk2\[9\].wave_shpr.div.acc\[0\] vssd1 vssd1 vccd1 vccd1 net1209 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11062_ _05015_ _05135_ vssd1 vssd1 vccd1 vccd1 _05136_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06132__A net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11513__A2 _05448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10013_ genblk2\[3\].wave_shpr.div.b1\[15\] genblk2\[3\].wave_shpr.div.acc\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04409_ sky130_fd_sc_hd__and2b_1
XFILLER_0_99_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06786__B net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11964_ genblk2\[10\].wave_shpr.div.acc\[25\] genblk2\[10\].wave_shpr.div.acc\[26\]
+ _05785_ vssd1 vssd1 vccd1 vccd1 _05786_ sky130_fd_sc_hd__or3_2
XFILLER_0_59_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_217 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13703_ clknet_leaf_96_clk _01014_ net161 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.fin_quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10915_ _03707_ vssd1 vssd1 vccd1 vccd1 _05042_ sky130_fd_sc_hd__buf_4
XFILLER_0_58_239 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11895_ _03838_ _03835_ genblk2\[0\].wave_shpr.div.i\[0\] vssd1 vssd1 vccd1 vccd1
+ _05722_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13634_ clknet_leaf_69_clk _00947_ net211 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.b1\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10846_ genblk2\[6\].wave_shpr.div.b1\[4\] genblk2\[6\].wave_shpr.div.acc\[4\] vssd1
+ vssd1 vccd1 vccd1 _04990_ sky130_fd_sc_hd__and2b_1
XFILLER_0_41_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13565_ clknet_leaf_57_clk _00880_ net182 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.quo\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10777_ _04814_ _04763_ vssd1 vssd1 vccd1 vccd1 _04935_ sky130_fd_sc_hd__or2b_1
XFILLER_0_81_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_743 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11213__A _02170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12516_ clknet_leaf_105_clk PWM.next_counter\[0\] net155 vssd1 vssd1 vccd1 vccd1
+ PWM.counter\[0\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07653__B1 _02221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13496_ clknet_leaf_86_clk net264 net178 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.quo\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12447_ clknet_leaf_106_clk net940 net153 vssd1 vssd1 vccd1 vccd1 sig_norm.i\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_128 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12378_ genblk2\[11\].wave_shpr.div.acc\[7\] _06054_ _06055_ vssd1 vssd1 vccd1 vccd1
+ _06056_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11752__A2 _05623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11329_ net809 _05311_ _05315_ _05321_ vssd1 vssd1 vccd1 vccd1 _00752_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_66_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08905__B1 _02248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06870_ _01725_ vssd1 vssd1 vccd1 vccd1 genblk1\[5\].osc.clkdiv_C.next_cnt\[16\]
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10712__B1 _04857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08540_ _02647_ vssd1 vssd1 vccd1 vccd1 _03247_ sky130_fd_sc_hd__inv_2
X_08471_ _03176_ _03177_ _02789_ vssd1 vssd1 vccd1 vccd1 _03178_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07422_ _02147_ _02163_ vssd1 vssd1 vccd1 vccd1 _02164_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_18_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07353_ _02111_ vssd1 vssd1 vccd1 vccd1 genblk1\[11\].osc.clkdiv_C.next_cnt\[5\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06304_ genblk1\[0\].osc.clkdiv_C.cnt\[1\] _01235_ _01253_ _01260_ _01265_ vssd1
+ vssd1 vccd1 vccd1 _01266_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_61_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_491 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07284_ _02026_ _02053_ vssd1 vssd1 vccd1 vccd1 _02054_ sky130_fd_sc_hd__nor2_1
XFILLER_0_33_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09023_ genblk2\[9\].wave_shpr.div.i\[1\] genblk2\[9\].wave_shpr.div.i\[0\] genblk2\[9\].wave_shpr.div.i\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03695_ sky130_fd_sc_hd__nand3_1
XFILLER_0_142_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06235_ _01196_ vssd1 vssd1 vccd1 vccd1 _01197_ sky130_fd_sc_hd__buf_4
XFILLER_0_86_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_575 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold210 sig_norm.acc_next\[0\] vssd1 vssd1 vccd1 vccd1 net428 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09528__A _03853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06166_ _01128_ _01113_ _01117_ vssd1 vssd1 vccd1 vccd1 _01138_ sky130_fd_sc_hd__and3_1
Xhold221 _01056_ vssd1 vssd1 vccd1 vccd1 net439 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_41_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold232 genblk2\[8\].wave_shpr.div.quo\[8\] vssd1 vssd1 vccd1 vccd1 net450 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold243 _00215_ vssd1 vssd1 vccd1 vccd1 net461 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10173__S _04507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold254 genblk2\[4\].wave_shpr.div.acc\[21\] vssd1 vssd1 vccd1 vccd1 net472 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold265 genblk2\[11\].wave_shpr.div.quo\[19\] vssd1 vssd1 vccd1 vccd1 net483 sky130_fd_sc_hd__dlygate4sd3_1
Xhold276 _00569_ vssd1 vssd1 vccd1 vccd1 net494 sky130_fd_sc_hd__dlygate4sd3_1
Xhold287 genblk2\[8\].wave_shpr.div.quo\[23\] vssd1 vssd1 vccd1 vccd1 net505 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09925_ net580 _04315_ _04322_ _04334_ vssd1 vssd1 vccd1 vccd1 _00335_ sky130_fd_sc_hd__a22o_1
Xhold298 _00636_ vssd1 vssd1 vccd1 vccd1 net516 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09856_ _04251_ _04279_ _04281_ _04253_ net1137 vssd1 vssd1 vccd1 vccd1 _00319_ sky130_fd_sc_hd__a32o_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08807_ _03431_ _03438_ vssd1 vssd1 vccd1 vccd1 _03514_ sky130_fd_sc_hd__nand2_1
XANTENNA__09263__A _03853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09787_ genblk2\[3\].wave_shpr.div.b1\[15\] _01365_ _04238_ vssd1 vssd1 vccd1 vccd1
+ _04244_ sky130_fd_sc_hd__mux2_1
X_06999_ genblk1\[7\].osc.clkdiv_C.cnt\[5\] genblk1\[7\].osc.clkdiv_C.cnt\[4\] _01827_
+ vssd1 vssd1 vccd1 vccd1 _01830_ sky130_fd_sc_hd__and3_1
XTAP_2404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08738_ _03428_ _03420_ _03443_ _03444_ vssd1 vssd1 vccd1 vccd1 _03445_ sky130_fd_sc_hd__o211a_2
XTAP_2415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_537 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08669_ _03371_ _03375_ vssd1 vssd1 vccd1 vccd1 _03376_ sky130_fd_sc_hd__xnor2_1
XTAP_1725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11732__S _00023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10700_ net324 _02183_ _04856_ net459 _04877_ vssd1 vssd1 vccd1 vccd1 _00567_ sky130_fd_sc_hd__a221o_1
XTAP_1747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11680_ genblk2\[9\].wave_shpr.div.b1\[1\] vssd1 vssd1 vccd1 vccd1 _05572_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10631_ _04842_ vssd1 vssd1 vccd1 vccd1 _00533_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_812 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_63_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13350_ clknet_leaf_5_clk _00671_ net45 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.acc\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07635__B1 _01235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07230__B _01432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10562_ genblk2\[5\].wave_shpr.div.b1\[5\] genblk2\[5\].wave_shpr.div.acc\[5\] vssd1
+ vssd1 vccd1 vccd1 _04790_ sky130_fd_sc_hd__and2b_1
XFILLER_0_63_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12301_ net402 _06009_ _06010_ net769 vssd1 vssd1 vccd1 vccd1 _01035_ sky130_fd_sc_hd__a22o_1
XFILLER_0_51_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13281_ clknet_leaf_122_clk _00602_ net79 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.fin_quo\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_16_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10493_ _04616_ _04565_ vssd1 vssd1 vccd1 vccd1 _04735_ sky130_fd_sc_hd__or2b_1
XFILLER_0_32_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09388__B1 _03819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12232_ _05928_ _05968_ _05969_ vssd1 vssd1 vccd1 vccd1 _05970_ sky130_fd_sc_hd__a21o_1
X_12163_ net906 _05818_ _05883_ _05909_ vssd1 vssd1 vccd1 vccd1 _00998_ sky130_fd_sc_hd__a22o_1
XANTENNA__10942__B1 _05056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11114_ genblk2\[7\].wave_shpr.div.acc\[7\] genblk2\[7\].wave_shpr.div.b1\[7\] vssd1
+ vssd1 vccd1 vccd1 _05174_ sky130_fd_sc_hd__or2b_1
X_12094_ _05857_ _05755_ vssd1 vssd1 vccd1 vccd1 _05858_ sky130_fd_sc_hd__xnor2_1
X_11045_ _05008_ _04970_ vssd1 vssd1 vccd1 vccd1 _05123_ sky130_fd_sc_hd__or2b_1
XFILLER_0_36_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09173__A _01342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13517__RESET_B net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12996_ clknet_leaf_132_clk _00325_ net60 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.acc\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08115__A1 _01172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11947_ _05737_ _05767_ _05768_ vssd1 vssd1 vccd1 vccd1 _05769_ sky130_fd_sc_hd__a21o_1
XFILLER_0_143_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_52_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13170__RESET_B net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_58 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_129_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11878_ _05709_ _05710_ vssd1 vssd1 vccd1 vccd1 _05711_ sky130_fd_sc_hd__nand2_1
X_13617_ clknet_leaf_94_clk _00930_ net160 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.fin_quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10829_ genblk2\[6\].wave_shpr.div.acc\[10\] genblk2\[6\].wave_shpr.div.b1\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04973_ sky130_fd_sc_hd__or2b_1
XFILLER_0_43_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13548_ clknet_leaf_110_clk _00863_ net152 vssd1 vssd1 vccd1 vccd1 sig_norm.b1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_501 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13479_ clknet_leaf_99_clk net744 net168 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.quo\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_140_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_2_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07971_ _01201_ genblk1\[7\].osc.clkdiv_C.cnt\[15\] _01362_ _02677_ vssd1 vssd1 vccd1
+ vccd1 _02678_ sky130_fd_sc_hd__o31a_1
X_09710_ _04165_ _04188_ _04189_ vssd1 vssd1 vccd1 vccd1 _04190_ sky130_fd_sc_hd__a21o_1
X_06922_ genblk1\[6\].osc.clkdiv_C.cnt\[6\] _01768_ vssd1 vssd1 vccd1 vccd1 _01770_
+ sky130_fd_sc_hd__and2_1
XANTENNA__10721__S _04821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09551__B1 _04046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09083__A _02170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09641_ genblk2\[1\].wave_shpr.div.acc\[19\] _04130_ vssd1 vssd1 vccd1 vccd1 _04133_
+ sky130_fd_sc_hd__or2_1
X_06853_ genblk1\[5\].osc.clkdiv_C.cnt\[11\] genblk1\[5\].osc.clkdiv_C.cnt\[10\] _01710_
+ vssd1 vssd1 vccd1 vccd1 _01714_ sky130_fd_sc_hd__and3_1
X_09572_ _04046_ vssd1 vssd1 vccd1 vccd1 _04080_ sky130_fd_sc_hd__clkbuf_4
X_06784_ _01436_ _01304_ genblk1\[5\].osc.clkdiv_C.cnt\[1\] vssd1 vssd1 vccd1 vccd1
+ _01656_ sky130_fd_sc_hd__a21oi_1
X_08523_ _03227_ _03229_ vssd1 vssd1 vccd1 vccd1 _03230_ sky130_fd_sc_hd__and2b_1
XANTENNA__09811__A _04069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08454_ _02216_ _02553_ genblk2\[7\].wave_shpr.div.fin_quo\[4\] vssd1 vssd1 vccd1
+ vccd1 _03161_ sky130_fd_sc_hd__and3_1
XFILLER_0_147_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_46_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07405_ _02147_ _02150_ vssd1 vssd1 vccd1 vccd1 _02151_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10168__S _04420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08385_ genblk1\[2\].osc.clkdiv_C.cnt\[4\] _01439_ _01418_ genblk1\[2\].osc.clkdiv_C.cnt\[3\]
+ _03091_ vssd1 vssd1 vccd1 vccd1 _03092_ sky130_fd_sc_hd__a221o_1
XFILLER_0_34_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07617__B1 _02064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07336_ _02097_ vssd1 vssd1 vccd1 vccd1 _02098_ sky130_fd_sc_hd__inv_2
XFILLER_0_116_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12893__RESET_B net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07267_ _02027_ _02041_ _02042_ vssd1 vssd1 vccd1 vccd1 genblk1\[10\].osc.clkdiv_C.next_cnt\[6\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_103_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09006_ net1168 net1170 _01154_ vssd1 vssd1 vccd1 vccd1 _03683_ sky130_fd_sc_hd__mux2_1
X_06218_ _01174_ _01177_ _01179_ vssd1 vssd1 vccd1 vccd1 _01180_ sky130_fd_sc_hd__a21o_2
XFILLER_0_104_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07198_ _01952_ _01983_ vssd1 vssd1 vccd1 vccd1 _01984_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06149_ _01119_ _01120_ vssd1 vssd1 vccd1 vccd1 _01121_ sky130_fd_sc_hd__nor2_1
XFILLER_0_130_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09790__B1 _03736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09908_ net1002 _04315_ _04289_ _04321_ vssd1 vssd1 vccd1 vccd1 _00331_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout72_A net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09839_ _04269_ genblk1\[2\].osc.clkdiv_C.cnt\[13\] vssd1 vssd1 vccd1 vccd1 _04271_
+ sky130_fd_sc_hd__and2_1
X_12850_ clknet_leaf_118_clk _00181_ net138 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.fin_quo\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_2201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11801_ _02203_ vssd1 vssd1 vccd1 vccd1 _05652_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_68_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12781_ clknet_leaf_40_clk _00114_ net115 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.b1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11732_ genblk2\[9\].wave_shpr.div.fin_quo\[5\] net1317 _00023_ vssd1 vssd1 vccd1
+ vccd1 _05619_ sky130_fd_sc_hd__mux2_1
XTAP_1544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11652__A1 _05449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07320__A2 _01513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11663_ _05439_ genblk2\[9\].wave_shpr.div.acc\[16\] vssd1 vssd1 vccd1 vccd1 _05555_
+ sky130_fd_sc_hd__nor2_1
XTAP_1599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_154_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13402_ clknet_leaf_90_clk net303 net147 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.quo\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10614_ _04832_ vssd1 vssd1 vccd1 vccd1 _00526_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11594_ net917 _05447_ _05484_ _05506_ vssd1 vssd1 vccd1 vccd1 _00832_ sky130_fd_sc_hd__a22o_1
X_13333_ clknet_leaf_9_clk _00654_ net54 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.acc\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10545_ genblk2\[5\].wave_shpr.div.acc\[7\] genblk2\[5\].wave_shpr.div.b1\[7\] vssd1
+ vssd1 vccd1 vccd1 _04773_ sky130_fd_sc_hd__or2b_1
XFILLER_0_52_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_130_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_130_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_107_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13264_ clknet_leaf_1_clk _00587_ net38 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.acc\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10476_ _04654_ vssd1 vssd1 vccd1 vccd1 _04722_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12215_ genblk2\[11\].wave_shpr.div.b1\[6\] genblk2\[11\].wave_shpr.div.acc\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05953_ sky130_fd_sc_hd__and2b_1
XFILLER_0_20_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13195_ clknet_leaf_128_clk _00518_ net132 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.fin_quo\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__10107__A _04269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12146_ genblk2\[10\].wave_shpr.div.acc\[17\] _05897_ _05786_ vssd1 vssd1 vccd1 vccd1
+ _05898_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_676 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13769__RESET_B net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07236__A2_N _02001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12077_ _05746_ _05747_ vssd1 vssd1 vccd1 vccd1 _05845_ sky130_fd_sc_hd__xor2_1
XANTENNA__07139__A2 _01246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11028_ _05000_ _04974_ vssd1 vssd1 vccd1 vccd1 _05110_ sky130_fd_sc_hd__or2b_1
XFILLER_0_154_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10694__A2 _02183_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12979_ clknet_leaf_124_clk _00308_ net72 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.quo\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_86_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06974__B _01675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_75_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08170_ genblk1\[3\].osc.clkdiv_C.cnt\[10\] _01508_ _01507_ genblk1\[3\].osc.clkdiv_C.cnt\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02877_ sky130_fd_sc_hd__a22o_1
X_07121_ genblk1\[9\].osc.clkdiv_C.cnt\[2\] _01920_ _01855_ genblk1\[9\].osc.clkdiv_C.cnt\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01921_ sky130_fd_sc_hd__o22a_1
XFILLER_0_132_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10716__S _04821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_121_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_121_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__07614__A3 _01208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07052_ _01441_ _01226_ vssd1 vssd1 vccd1 vccd1 _01870_ sky130_fd_sc_hd__nor2_4
XANTENNA__09078__A _03702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_140_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_10_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07954_ genblk1\[7\].osc.clkdiv_C.cnt\[4\] _01805_ vssd1 vssd1 vccd1 vccd1 _02661_
+ sky130_fd_sc_hd__and2_1
X_06905_ genblk1\[6\].osc.clkdiv_C.cnt\[3\] _01758_ vssd1 vssd1 vccd1 vccd1 _01759_
+ sky130_fd_sc_hd__xor2_1
X_07885_ _02526_ vssd1 vssd1 vccd1 vccd1 _02592_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_128_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_98_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09624_ _04000_ _03956_ vssd1 vssd1 vccd1 vccd1 _04120_ sky130_fd_sc_hd__or2b_1
X_06836_ genblk1\[5\].osc.clkdiv_C.cnt\[5\] genblk1\[5\].osc.clkdiv_C.cnt\[4\] _01700_
+ vssd1 vssd1 vccd1 vccd1 _01703_ sky130_fd_sc_hd__and3_1
XANTENNA__07045__B _01430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap29 _01372_ vssd1 vssd1 vccd1 vccd1 net29 sky130_fd_sc_hd__dlymetal6s2s_1
X_09555_ net632 _04042_ _04046_ genblk2\[1\].wave_shpr.div.quo\[23\] _04068_ vssd1
+ vssd1 vccd1 vccd1 _00231_ sky130_fd_sc_hd__a221o_1
X_06767_ genblk1\[4\].osc.clkdiv_C.cnt\[13\] vssd1 vssd1 vccd1 vccd1 _01644_ sky130_fd_sc_hd__inv_2
XANTENNA__11282__S _05222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08506_ _03211_ _03212_ genblk2\[2\].wave_shpr.div.fin_quo\[6\] _02468_ vssd1 vssd1
+ vccd1 vccd1 _03213_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_148_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09486_ _01431_ vssd1 vssd1 vccd1 vccd1 _04032_ sky130_fd_sc_hd__inv_2
X_06698_ genblk1\[4\].osc.clkdiv_C.cnt\[10\] vssd1 vssd1 vccd1 vccd1 _01588_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07302__A2 _01256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08437_ _02525_ _03142_ _03143_ _02361_ genblk2\[11\].wave_shpr.div.fin_quo\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03144_ sky130_fd_sc_hd__a32o_1
XFILLER_0_65_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08368_ _03071_ _03074_ vssd1 vssd1 vccd1 vccd1 _03075_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_746 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07066__A1 genblk1\[8\].osc.clkdiv_C.cnt\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07319_ _02080_ _01242_ _01423_ _02081_ _02082_ vssd1 vssd1 vccd1 vccd1 _02083_ sky130_fd_sc_hd__o221a_1
XFILLER_0_34_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10626__S _04834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07066__B2 genblk1\[8\].osc.clkdiv_C.cnt\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_112_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_112_clk
+ sky130_fd_sc_hd__clkbuf_16
X_08299_ _02897_ _02925_ _02926_ vssd1 vssd1 vccd1 vccd1 _03006_ sky130_fd_sc_hd__or3_1
XFILLER_0_21_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10330_ genblk2\[5\].wave_shpr.div.b1\[1\] vssd1 vssd1 vccd1 vccd1 _04633_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_33_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06405__A _01172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10261_ genblk2\[4\].wave_shpr.div.acc\[9\] genblk2\[4\].wave_shpr.div.b1\[9\] vssd1
+ vssd1 vccd1 vccd1 _04573_ sky130_fd_sc_hd__or2b_1
XANTENNA_hold586_A genblk2\[0\].wave_shpr.div.quo\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12000_ net1217 _03706_ _05802_ vssd1 vssd1 vccd1 vccd1 _05805_ sky130_fd_sc_hd__mux2_1
X_10192_ _04455_ vssd1 vssd1 vccd1 vccd1 _04522_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__06585__A1_N _01490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_884 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09515__B1 _04047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11484__A2_N _01490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12902_ clknet_leaf_30_clk _00233_ net104 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.acc\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12833_ clknet_leaf_64_clk _00166_ net196 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.acc\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2020 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2031 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2042 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06794__B _01171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2053 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2064 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12764_ clknet_leaf_92_clk _00097_ net148 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.fin_quo\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_2075 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2086 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2097 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_68_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11715_ _05554_ _05605_ _05606_ vssd1 vssd1 vccd1 vccd1 _05607_ sky130_fd_sc_hd__a21o_1
XTAP_1374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12695_ clknet_leaf_54_clk genblk1\[8\].osc.clkdiv_C.next_cnt\[8\] net172 vssd1 vssd1
+ vccd1 vccd1 genblk1\[8\].osc.clkdiv_C.cnt\[8\] sky130_fd_sc_hd__dfrtp_4
XTAP_1396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11646_ genblk2\[8\].wave_shpr.div.acc\[25\] _05414_ _05543_ vssd1 vssd1 vccd1 vccd1
+ _05544_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_37_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_24_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput14 pb[8] vssd1 vssd1 vccd1 vccd1 net14 sky130_fd_sc_hd__clkbuf_2
XANTENNA__07057__A1 genblk1\[8\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_589 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08254__B1 _02261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_leaf_103_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_103_clk
+ sky130_fd_sc_hd__clkbuf_16
X_11577_ genblk2\[8\].wave_shpr.div.acc\[6\] _05492_ _05493_ vssd1 vssd1 vccd1 vccd1
+ _05494_ sky130_fd_sc_hd__mux2_1
XFILLER_0_107_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13316_ clknet_leaf_9_clk _00637_ net50 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.quo\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10528_ _04758_ vssd1 vssd1 vccd1 vccd1 _04759_ sky130_fd_sc_hd__inv_2
Xhold809 sig_norm.acc\[5\] vssd1 vssd1 vccd1 vccd1 net1027 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13247_ clknet_leaf_2_clk _00570_ net52 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.acc\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08006__B1 _01738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10459_ _04600_ _04573_ vssd1 vssd1 vccd1 vccd1 _04709_ sky130_fd_sc_hd__or2b_1
XFILLER_0_58_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08557__A1 genblk2\[8\].wave_shpr.div.fin_quo\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_13178_ clknet_leaf_131_clk _00503_ net65 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.acc\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_12129_ _05771_ _05884_ vssd1 vssd1 vccd1 vccd1 _05885_ sky130_fd_sc_hd__xnor2_1
XANTENNA__12105__A2 _05844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07146__A _01336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10667__A2 _04858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07670_ _02375_ _02376_ vssd1 vssd1 vccd1 vccd1 _02377_ sky130_fd_sc_hd__or2_1
X_06621_ _01527_ vssd1 vssd1 vccd1 vccd1 genblk1\[3\].osc.clkdiv_C.next_cnt\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09340_ genblk2\[0\].wave_shpr.div.acc\[16\] _03918_ _03889_ vssd1 vssd1 vccd1 vccd1
+ _03919_ sky130_fd_sc_hd__mux2_1
X_06552_ genblk1\[2\].osc.clkdiv_C.cnt\[10\] genblk1\[2\].osc.clkdiv_C.cnt\[9\] _01464_
+ vssd1 vssd1 vccd1 vccd1 _01468_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09271_ genblk2\[0\].wave_shpr.div.b1\[0\] genblk2\[0\].wave_shpr.div.acc\[0\] _03804_
+ _03863_ vssd1 vssd1 vccd1 vccd1 _03866_ sky130_fd_sc_hd__a31o_1
X_06483_ genblk1\[1\].osc.clkdiv_C.cnt\[17\] _01407_ _01409_ _01374_ vssd1 vssd1 vccd1
+ vccd1 genblk1\[1\].osc.clkdiv_C.next_cnt\[17\] sky130_fd_sc_hd__o211a_1
XFILLER_0_117_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08222_ _02789_ _02793_ genblk2\[5\].wave_shpr.div.fin_quo\[5\] vssd1 vssd1 vccd1
+ vccd1 _02929_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_117_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_31 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07048__A1 _01174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08153_ genblk1\[3\].osc.clkdiv_C.cnt\[5\] _01500_ _01494_ genblk1\[3\].osc.clkdiv_C.cnt\[6\]
+ vssd1 vssd1 vccd1 vccd1 _02860_ sky130_fd_sc_hd__a22o_1
XFILLER_0_133_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_16_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_71_852 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout122_A net126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07104_ genblk1\[8\].osc.clkdiv_C.cnt\[12\] _01906_ _01909_ vssd1 vssd1 vccd1 vccd1
+ genblk1\[8\].osc.clkdiv_C.next_cnt\[12\] sky130_fd_sc_hd__o21a_1
XFILLER_0_15_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08084_ _02790_ vssd1 vssd1 vccd1 vccd1 _02791_ sky130_fd_sc_hd__buf_2
XFILLER_0_43_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_130_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07035_ genblk1\[8\].osc.clkdiv_C.cnt\[10\] _01852_ _01248_ vssd1 vssd1 vccd1 vccd1
+ _01853_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_101_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09536__A _04058_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11785__B genblk1\[9\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10355__A1 _04645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11277__S _05222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10181__S _04507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08986_ _03225_ _03570_ vssd1 vssd1 vccd1 vccd1 _03670_ sky130_fd_sc_hd__nor2_1
XANTENNA__07056__A genblk1\[8\].osc.clkdiv_C.cnt\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07937_ _02642_ _02643_ vssd1 vssd1 vccd1 vccd1 _02644_ sky130_fd_sc_hd__and2b_1
XANTENNA__10658__A2 _04853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07868_ _02509_ _02572_ _02574_ _02517_ vssd1 vssd1 vccd1 vccd1 _02575_ sky130_fd_sc_hd__o211a_1
XFILLER_0_3_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09607_ _03991_ _04106_ vssd1 vssd1 vccd1 vccd1 _04107_ sky130_fd_sc_hd__xnor2_1
X_06819_ _01665_ _01668_ _01673_ _01690_ vssd1 vssd1 vccd1 vccd1 _01691_ sky130_fd_sc_hd__or4b_1
X_07799_ genblk1\[0\].osc.clkdiv_C.cnt\[15\] _01349_ _01577_ genblk1\[0\].osc.clkdiv_C.cnt\[16\]
+ _02505_ vssd1 vssd1 vccd1 vccd1 _02506_ sky130_fd_sc_hd__o221a_1
XFILLER_0_39_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09538_ _04055_ genblk1\[1\].osc.clkdiv_C.cnt\[7\] vssd1 vssd1 vccd1 vccd1 _04060_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_39_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08484__B1 _02885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09469_ genblk2\[2\].wave_shpr.div.b1\[3\] _01231_ _03822_ vssd1 vssd1 vccd1 vccd1
+ _04022_ sky130_fd_sc_hd__mux2_1
XANTENNA__11083__A2 _05057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11500_ net346 _05442_ _05446_ net709 vssd1 vssd1 vccd1 vccd1 _00798_ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12480_ clknet_leaf_108_clk _00042_ net152 vssd1 vssd1 vccd1 vccd1 sig_norm.acc\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11431_ _05359_ _05405_ _05406_ vssd1 vssd1 vccd1 vccd1 _05407_ sky130_fd_sc_hd__a21o_1
XFILLER_0_151_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10043__B1 _03733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08787__B2 _02468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11362_ genblk2\[7\].wave_shpr.div.acc\[24\] vssd1 vssd1 vccd1 vccd1 _05345_ sky130_fd_sc_hd__inv_2
XANTENNA__06135__A net11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10594__A1 _04821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13101_ clknet_leaf_122_clk _00012_ net78 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.busy
+ sky130_fd_sc_hd__dfrtp_1
X_10313_ _04624_ vssd1 vssd1 vccd1 vccd1 _00433_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07898__A1_N genblk1\[8\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__06262__A2 _01221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11293_ genblk2\[7\].wave_shpr.div.acc\[6\] _05293_ _05222_ vssd1 vssd1 vccd1 vccd1
+ _05294_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_104_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13032_ clknet_leaf_121_clk _00359_ net78 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.b1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10244_ genblk2\[3\].wave_shpr.div.i\[1\] genblk2\[3\].wave_shpr.div.i\[0\] genblk2\[3\].wave_shpr.div.i\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04559_ sky130_fd_sc_hd__a21o_1
XFILLER_0_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10175_ _04397_ _04369_ vssd1 vssd1 vccd1 vccd1 _04509_ sky130_fd_sc_hd__or2b_1
XANTENNA__07762__A2 _02459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout180 net185 vssd1 vssd1 vccd1 vccd1 net180 sky130_fd_sc_hd__buf_2
XANTENNA__06970__B1 _01801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout191 net198 vssd1 vssd1 vccd1 vccd1 net191 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_135_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12816_ clknet_leaf_58_clk _00149_ net192 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.acc\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_97_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_69_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12747_ clknet_leaf_49_clk genblk1\[11\].osc.clkdiv_C.next_cnt\[6\] net108 vssd1
+ vssd1 vccd1 vccd1 genblk1\[11\].osc.clkdiv_C.cnt\[6\] sky130_fd_sc_hd__dfrtp_4
XTAP_1182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12678_ clknet_leaf_120_clk genblk1\[7\].osc.clkdiv_C.next_cnt\[9\] net142 vssd1
+ vssd1 vccd1 vccd1 genblk1\[7\].osc.clkdiv_C.cnt\[9\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_37_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08227__B1 _02316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11629_ _05471_ _05532_ net690 _05442_ vssd1 vssd1 vccd1 vccd1 _00841_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_115_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_13_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold606 _00154_ vssd1 vssd1 vccd1 vccd1 net824 sky130_fd_sc_hd__dlygate4sd3_1
Xhold617 genblk2\[5\].wave_shpr.div.acc\[15\] vssd1 vssd1 vccd1 vccd1 net835 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold628 genblk2\[8\].wave_shpr.div.acc\[14\] vssd1 vssd1 vccd1 vccd1 net846 sky130_fd_sc_hd__dlygate4sd3_1
Xhold639 genblk2\[2\].wave_shpr.div.acc\[12\] vssd1 vssd1 vccd1 vccd1 net857 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_900 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08840_ _03464_ _03526_ _03528_ vssd1 vssd1 vccd1 vccd1 _03547_ sky130_fd_sc_hd__o21ai_1
XTAP_933 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07202__A1 genblk1\[9\].osc.clkdiv_C.cnt\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_944 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_977 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08771_ _03304_ _03306_ vssd1 vssd1 vccd1 vccd1 _03478_ sky130_fd_sc_hd__xnor2_1
XTAP_988 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_109_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_999 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07307__C _01678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07722_ _01330_ _01262_ _01591_ _01172_ vssd1 vssd1 vccd1 vccd1 _02429_ sky130_fd_sc_hd__o211ai_1
XANTENNA_clkbuf_4_7_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09091__A _01201_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07653_ _02349_ _02351_ _02221_ vssd1 vssd1 vccd1 vccd1 _02360_ sky130_fd_sc_hd__a21o_1
XANTENNA__12666__RESET_B net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07910__C1 _01238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_76_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06604_ _01171_ _01192_ _01208_ vssd1 vssd1 vccd1 vccd1 _01512_ sky130_fd_sc_hd__and3_1
X_07584_ genblk1\[9\].osc.clkdiv_C.cnt\[2\] _01234_ _01310_ genblk1\[9\].osc.clkdiv_C.cnt\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02291_ sky130_fd_sc_hd__o22a_1
XFILLER_0_149_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09323_ genblk2\[0\].wave_shpr.div.acc\[12\] _03905_ _03889_ vssd1 vssd1 vccd1 vccd1
+ _03906_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06535_ _01452_ _01456_ _01457_ vssd1 vssd1 vccd1 vccd1 genblk1\[2\].osc.clkdiv_C.next_cnt\[3\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_47_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09254_ net298 _03845_ _03847_ net466 _03856_ vssd1 vssd1 vccd1 vccd1 _00142_ sky130_fd_sc_hd__a221o_1
XFILLER_0_35_318 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06466_ _01373_ _01397_ _01398_ vssd1 vssd1 vccd1 vccd1 genblk1\[1\].osc.clkdiv_C.next_cnt\[11\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_29_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08205_ genblk2\[9\].wave_shpr.div.fin_quo\[5\] _02303_ _02265_ _02316_ vssd1 vssd1
+ vccd1 vccd1 _02912_ sky130_fd_sc_hd__a31o_1
XFILLER_0_106_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09185_ _01430_ _01344_ _03819_ vssd1 vssd1 vccd1 vccd1 _03820_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_141_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06397_ genblk1\[1\].osc.clkdiv_C.cnt\[17\] vssd1 vssd1 vccd1 vccd1 _01341_ sky130_fd_sc_hd__inv_2
XFILLER_0_105_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08136_ _02842_ genblk2\[4\].wave_shpr.div.fin_quo\[5\] _02837_ vssd1 vssd1 vccd1
+ vccd1 _02843_ sky130_fd_sc_hd__or3b_1
XFILLER_0_43_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06244__A2 _01190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08067_ _01660_ _02773_ genblk1\[5\].osc.clkdiv_C.cnt\[1\] vssd1 vssd1 vccd1 vccd1
+ _02774_ sky130_fd_sc_hd__o21a_1
XANTENNA__10904__S _04848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_481 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07018_ genblk1\[7\].osc.clkdiv_C.cnt\[12\] _01841_ vssd1 vssd1 vccd1 vccd1 _01842_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_12_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10328__A1 _01735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09194__A1 _01991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07744__A2 _02425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08969_ _03565_ _03567_ _03508_ vssd1 vssd1 vccd1 vccd1 _03656_ sky130_fd_sc_hd__o21a_1
X_11980_ genblk2\[10\].wave_shpr.div.fin_quo\[7\] genblk2\[10\].wave_shpr.div.quo\[6\]
+ _00003_ vssd1 vssd1 vccd1 vccd1 _05795_ sky130_fd_sc_hd__mux2_1
XFILLER_0_98_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06891__A2_N _01666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10931_ _02171_ net1234 vssd1 vssd1 vccd1 vccd1 _05050_ sky130_fd_sc_hd__and2_1
XFILLER_0_98_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13650_ clknet_leaf_38_clk _00963_ net116 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.quo\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10862_ genblk2\[6\].wave_shpr.div.b1\[12\] genblk2\[6\].wave_shpr.div.acc\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05006_ sky130_fd_sc_hd__and2b_1
XFILLER_0_14_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_66_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12601_ clknet_leaf_21_clk genblk1\[3\].osc.clkdiv_C.next_cnt\[4\] net97 vssd1 vssd1
+ vccd1 vccd1 genblk1\[3\].osc.clkdiv_C.cnt\[4\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_94_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13581_ clknet_leaf_76_clk _00896_ net207 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.acc\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10793_ net654 _04918_ _04922_ _04946_ vssd1 vssd1 vccd1 vccd1 _00591_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12532_ clknet_leaf_61_clk _00084_ net186 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.b1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12463_ clknet_leaf_103_clk _00036_ net156 vssd1 vssd1 vccd1 vccd1 PWM.final_sample_in\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_34_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11414_ genblk2\[8\].wave_shpr.div.b1\[8\] genblk2\[8\].wave_shpr.div.acc\[8\] vssd1
+ vssd1 vccd1 vccd1 _05390_ sky130_fd_sc_hd__and2b_1
X_12394_ genblk2\[11\].wave_shpr.div.acc\[11\] _06067_ _06055_ vssd1 vssd1 vccd1 vccd1
+ _06068_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_leaf_73_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_429 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11345_ net1048 _05311_ _05315_ _05333_ vssd1 vssd1 vccd1 vccd1 _00756_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_120_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11276_ _05185_ _05280_ vssd1 vssd1 vccd1 vccd1 _05281_ sky130_fd_sc_hd__xnor2_1
X_13015_ clknet_leaf_12_clk _00010_ net52 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.busy
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09185__A1 _01430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10227_ genblk2\[3\].wave_shpr.div.acc\[22\] _04416_ _04547_ vssd1 vssd1 vccd1 vccd1
+ _04548_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_88_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07735__A2 _02433_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10158_ _04389_ _04373_ vssd1 vssd1 vccd1 vccd1 _04496_ sky130_fd_sc_hd__or2b_1
XANTENNA_clkbuf_leaf_131_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold3 _00951_ vssd1 vssd1 vccd1 vccd1 net221 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10089_ genblk2\[3\].wave_shpr.div.quo\[2\] _04452_ _04456_ net326 vssd1 vssd1 vccd1
+ vccd1 _00377_ sky130_fd_sc_hd__a22o_1
XANTENNA__12330__A _03689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_11_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08145__C1 _01362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07143__B _01514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08954__S _02248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08448__B1 genblk2\[8\].wave_shpr.div.fin_quo\[3\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_26_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06320_ genblk1\[0\].osc.clkdiv_C.cnt\[4\] _01276_ _01270_ vssd1 vssd1 vccd1 vccd1
+ _01278_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_29_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_84_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_57_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06251_ _01174_ _01187_ vssd1 vssd1 vccd1 vccd1 _01213_ sky130_fd_sc_hd__nand2_2
Xclkbuf_4_4_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_4_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_60_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09785__S _04238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06182_ _01153_ vssd1 vssd1 vccd1 vccd1 _01154_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__11755__B1 _03694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold403 _00640_ vssd1 vssd1 vccd1 vccd1 net621 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold414 genblk2\[1\].wave_shpr.div.quo\[24\] vssd1 vssd1 vccd1 vccd1 net632 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10724__S _04821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold425 genblk2\[4\].wave_shpr.div.acc_next\[0\] vssd1 vssd1 vccd1 vccd1 net643 sky130_fd_sc_hd__dlygate4sd3_1
Xhold436 genblk2\[5\].wave_shpr.div.acc\[22\] vssd1 vssd1 vccd1 vccd1 net654 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold447 genblk2\[4\].wave_shpr.div.quo\[22\] vssd1 vssd1 vccd1 vccd1 net665 sky130_fd_sc_hd__dlygate4sd3_1
Xhold458 genblk2\[8\].wave_shpr.div.quo\[6\] vssd1 vssd1 vccd1 vccd1 net676 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09086__A modein.delay_octave_down_in\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09941_ net707 _04253_ _04322_ _04345_ vssd1 vssd1 vccd1 vccd1 _00340_ sky130_fd_sc_hd__a22o_1
Xhold469 _00868_ vssd1 vssd1 vccd1 vccd1 net687 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09176__A1 _01368_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07318__B _01262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09872_ _04293_ _04182_ vssd1 vssd1 vccd1 vccd1 _04294_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10025__A _02170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08823_ _03465_ _03481_ _03480_ vssd1 vssd1 vccd1 vccd1 _03530_ sky130_fd_sc_hd__o21a_1
Xhold1103 genblk2\[8\].wave_shpr.div.quo\[3\] vssd1 vssd1 vccd1 vccd1 net1321 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1114 genblk2\[11\].wave_shpr.div.quo\[5\] vssd1 vssd1 vccd1 vccd1 net1332 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_31_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1125 genblk2\[2\].wave_shpr.div.quo\[1\] vssd1 vssd1 vccd1 vccd1 net1343 sky130_fd_sc_hd__dlygate4sd3_1
X_08754_ _03454_ _03460_ vssd1 vssd1 vccd1 vccd1 _03461_ sky130_fd_sc_hd__xnor2_1
XTAP_2608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07705_ genblk2\[10\].wave_shpr.div.fin_quo\[6\] vssd1 vssd1 vccd1 vccd1 _02412_
+ sky130_fd_sc_hd__inv_2
XTAP_2619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08685_ _03387_ _03391_ vssd1 vssd1 vccd1 vccd1 _03392_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11286__A2 _05279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_92_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_92_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_95_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08149__B _01513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08151__A2 _01250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07636_ _02337_ _02341_ _02342_ vssd1 vssd1 vccd1 vccd1 _02343_ sky130_fd_sc_hd__or3b_1
XTAP_1929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07567_ genblk1\[9\].osc.clkdiv_C.cnt\[14\] _01936_ _01349_ vssd1 vssd1 vccd1 vccd1
+ _02274_ sky130_fd_sc_hd__o21a_1
X_09306_ genblk2\[0\].wave_shpr.div.acc\[8\] _03892_ _03889_ vssd1 vssd1 vccd1 vccd1
+ _03893_ sky130_fd_sc_hd__mux2_1
X_06518_ genblk1\[2\].osc.clkdiv_C.cnt\[9\] _01442_ _01439_ genblk1\[2\].osc.clkdiv_C.cnt\[5\]
+ vssd1 vssd1 vccd1 vccd1 _01444_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_8_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07498_ _02218_ _02219_ vssd1 vssd1 vccd1 vccd1 FSM.next_mode\[0\] sky130_fd_sc_hd__nand2_1
XFILLER_0_118_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09237_ net584 _03845_ _03839_ net599 _03846_ vssd1 vssd1 vccd1 vccd1 _00135_ sky130_fd_sc_hd__a221o_1
XFILLER_0_145_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06449_ genblk1\[1\].osc.clkdiv_C.cnt\[6\] _01385_ vssd1 vssd1 vccd1 vccd1 _01387_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_16_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_50_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_32_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09168_ _03810_ vssd1 vssd1 vccd1 vccd1 _00102_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11746__B1 _05624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08119_ _02822_ _02823_ _02824_ _02825_ vssd1 vssd1 vccd1 vccd1 _02826_ sky130_fd_sc_hd__o31a_1
XFILLER_0_32_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09099_ genblk2\[0\].wave_shpr.div.acc\[16\] genblk2\[0\].wave_shpr.div.b1\[16\]
+ vssd1 vssd1 vccd1 vccd1 _03747_ sky130_fd_sc_hd__or2b_1
XFILLER_0_102_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07965__A2 _01577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11130_ _05179_ _05189_ _05177_ vssd1 vssd1 vccd1 vccd1 _05190_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_101_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold970 genblk2\[4\].wave_shpr.div.b1\[4\] vssd1 vssd1 vccd1 vccd1 net1188 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06413__A genblk1\[1\].osc.clkdiv_C.cnt\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold981 genblk2\[10\].wave_shpr.div.b1\[12\] vssd1 vssd1 vccd1 vccd1 net1199 sky130_fd_sc_hd__dlygate4sd3_1
X_11061_ _05016_ _04966_ vssd1 vssd1 vccd1 vccd1 _05135_ sky130_fd_sc_hd__or2b_1
Xhold992 _00891_ vssd1 vssd1 vccd1 vccd1 net1210 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06132__B net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10012_ _04364_ _04406_ _04407_ vssd1 vssd1 vccd1 vccd1 _04408_ sky130_fd_sc_hd__a21o_1
XANTENNA__08390__A2 _01442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11963_ genblk2\[10\].wave_shpr.div.acc\[24\] _05784_ vssd1 vssd1 vccd1 vccd1 _05785_
+ sky130_fd_sc_hd__or2_2
XFILLER_0_25_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_83_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_83_clk sky130_fd_sc_hd__clkbuf_16
X_13702_ clknet_leaf_97_clk _01013_ net167 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.fin_quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10914_ _05041_ vssd1 vssd1 vccd1 vccd1 _00617_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__06153__A1 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11894_ net348 _03696_ _03694_ _05721_ vssd1 vssd1 vccd1 vccd1 _00917_ sky130_fd_sc_hd__a22o_1
X_13633_ clknet_leaf_69_clk _00946_ net213 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.b1\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10845_ _04980_ _04987_ _04988_ vssd1 vssd1 vccd1 vccd1 _04989_ sky130_fd_sc_hd__a21o_1
XFILLER_0_132_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_38 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10776_ net828 _04918_ _04922_ _04934_ vssd1 vssd1 vccd1 vccd1 _00586_ sky130_fd_sc_hd__a22o_1
XFILLER_0_109_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13564_ clknet_leaf_57_clk _00879_ net182 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.quo\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_12515_ clknet_leaf_106_clk _00024_ net154 vssd1 vssd1 vccd1 vccd1 sig_norm.busy
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_695 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13495_ clknet_leaf_88_clk _00812_ net178 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.quo\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12446_ clknet_leaf_99_clk net219 net168 vssd1 vssd1 vccd1 vccd1 net19 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12377_ _05981_ vssd1 vssd1 vccd1 vccd1 _06055_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07956__A2 _02656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11328_ genblk2\[7\].wave_shpr.div.acc\[14\] _05320_ _05300_ vssd1 vssd1 vccd1 vccd1
+ _05321_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11259_ genblk2\[7\].wave_shpr.div.quo\[23\] _05245_ _05249_ net487 _05269_ vssd1
+ vssd1 vccd1 vccd1 _00734_ sky130_fd_sc_hd__a221o_1
XANTENNA__12940__RESET_B net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08381__A2 _01209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11268__A2 _05222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_74_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_74_clk sky130_fd_sc_hd__clkbuf_16
X_08470_ genblk2\[5\].wave_shpr.div.fin_quo\[0\] genblk2\[5\].wave_shpr.div.fin_quo\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03177_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_148_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07421_ genblk2\[2\].wave_shpr.div.busy _02162_ vssd1 vssd1 vccd1 vccd1 _02163_ sky130_fd_sc_hd__and2_1
XFILLER_0_46_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_73_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07352_ _02092_ _02109_ _02110_ vssd1 vssd1 vccd1 vccd1 _02111_ sky130_fd_sc_hd__and3_1
XFILLER_0_134_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06303_ genblk1\[0\].osc.clkdiv_C.cnt\[14\] _01256_ _01258_ genblk1\[0\].osc.clkdiv_C.cnt\[5\]
+ _01264_ vssd1 vssd1 vccd1 vccd1 _01265_ sky130_fd_sc_hd__a221o_1
XFILLER_0_127_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07283_ genblk1\[10\].osc.clkdiv_C.cnt\[12\] _02052_ vssd1 vssd1 vccd1 vccd1 _02053_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_73_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09022_ _03693_ vssd1 vssd1 vccd1 vccd1 _03694_ sky130_fd_sc_hd__clkbuf_4
X_06234_ _01195_ vssd1 vssd1 vccd1 vccd1 _01196_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_115_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09809__A _04069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_827 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_587 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_130_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold200 genblk2\[4\].wave_shpr.div.quo\[0\] vssd1 vssd1 vccd1 vccd1 net418 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_131_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold211 _00062_ vssd1 vssd1 vccd1 vccd1 net429 sky130_fd_sc_hd__dlygate4sd3_1
X_06165_ _01134_ _01136_ vssd1 vssd1 vccd1 vccd1 _01137_ sky130_fd_sc_hd__or2_1
XFILLER_0_142_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold222 genblk2\[10\].wave_shpr.div.quo\[19\] vssd1 vssd1 vccd1 vccd1 net440 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold233 genblk2\[3\].wave_shpr.div.quo\[18\] vssd1 vssd1 vccd1 vccd1 net451 sky130_fd_sc_hd__dlygate4sd3_1
Xhold244 genblk2\[1\].wave_shpr.div.quo\[16\] vssd1 vssd1 vccd1 vccd1 net462 sky130_fd_sc_hd__dlygate4sd3_1
Xhold255 _00507_ vssd1 vssd1 vccd1 vccd1 net473 sky130_fd_sc_hd__dlygate4sd3_1
Xhold266 genblk2\[7\].wave_shpr.div.b1\[14\] vssd1 vssd1 vccd1 vccd1 net484 sky130_fd_sc_hd__dlygate4sd3_1
Xhold277 genblk2\[0\].wave_shpr.div.quo\[13\] vssd1 vssd1 vccd1 vccd1 net495 sky130_fd_sc_hd__dlygate4sd3_1
Xhold288 genblk2\[8\].wave_shpr.div.quo\[11\] vssd1 vssd1 vccd1 vccd1 net506 sky130_fd_sc_hd__dlygate4sd3_1
X_09924_ genblk2\[2\].wave_shpr.div.acc\[17\] _04333_ _04213_ vssd1 vssd1 vccd1 vccd1
+ _04334_ sky130_fd_sc_hd__mux2_1
Xhold299 genblk2\[1\].wave_shpr.div.quo\[9\] vssd1 vssd1 vccd1 vccd1 net517 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09855_ _04214_ _04280_ vssd1 vssd1 vccd1 vccd1 _04281_ sky130_fd_sc_hd__nand2_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11285__S _05222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08806_ _03433_ _03437_ vssd1 vssd1 vccd1 vccd1 _03513_ sky130_fd_sc_hd__or2b_1
XANTENNA__09263__B genblk1\[0\].osc.clkdiv_C.cnt\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09786_ _04243_ vssd1 vssd1 vccd1 vccd1 _00287_ sky130_fd_sc_hd__clkbuf_1
X_06998_ _01823_ _01829_ vssd1 vssd1 vccd1 vccd1 genblk1\[7\].osc.clkdiv_C.next_cnt\[4\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__07580__B1 genblk1\[9\].osc.clkdiv_C.cnt\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08737_ _03442_ _03441_ _03439_ vssd1 vssd1 vccd1 vccd1 _03444_ sky130_fd_sc_hd__a21bo_1
XANTENNA__11259__A2 _05245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_65_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_65_clk sky130_fd_sc_hd__clkbuf_16
XTAP_2427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08124__A2 _01340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08668_ _02838_ _03374_ _02846_ vssd1 vssd1 vccd1 vccd1 _03375_ sky130_fd_sc_hd__o21a_1
XTAP_1704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07619_ genblk1\[11\].osc.clkdiv_C.cnt\[5\] _01595_ _02323_ _02324_ _02325_ vssd1
+ vssd1 vccd1 vccd1 _02326_ sky130_fd_sc_hd__o221a_1
X_08599_ net9 _02744_ _03305_ vssd1 vssd1 vccd1 vccd1 _03306_ sky130_fd_sc_hd__and3_1
XTAP_1759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10630_ net1308 _02725_ _04834_ vssd1 vssd1 vccd1 vccd1 _04842_ sky130_fd_sc_hd__mux2_1
XANTENNA__09085__B1 _03736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_882 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_824 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10561_ _04778_ _04788_ _04776_ vssd1 vssd1 vccd1 vccd1 _04789_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_63_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_632 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_619 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_799 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12300_ genblk2\[11\].wave_shpr.div.quo\[1\] _06009_ _06010_ net430 vssd1 vssd1 vccd1
+ vccd1 _01034_ sky130_fd_sc_hd__a22o_1
X_13280_ clknet_leaf_122_clk _00601_ net79 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.fin_quo\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_51_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10492_ net926 _04715_ _04722_ _04734_ vssd1 vssd1 vccd1 vccd1 _00502_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12231_ genblk2\[11\].wave_shpr.div.b1\[14\] genblk2\[11\].wave_shpr.div.acc\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05969_ sky130_fd_sc_hd__and2b_1
XFILLER_0_122_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11195__A1 _05236_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07938__A2 _02539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12162_ genblk2\[10\].wave_shpr.div.acc\[22\] _05908_ vssd1 vssd1 vccd1 vccd1 _05909_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_31_173 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06143__A net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11113_ genblk2\[7\].wave_shpr.div.acc\[8\] genblk2\[7\].wave_shpr.div.b1\[8\] vssd1
+ vssd1 vccd1 vccd1 _05173_ sky130_fd_sc_hd__or2b_1
X_12093_ _05756_ _05742_ vssd1 vssd1 vccd1 vccd1 _05857_ sky130_fd_sc_hd__nor2_1
XANTENNA__06610__A2 _01231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_4_15_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11044_ net883 _05119_ _05093_ _05122_ vssd1 vssd1 vccd1 vccd1 _00666_ sky130_fd_sc_hd__a22o_1
XANTENNA__08899__B1 _01157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09560__A1 _03819_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09173__B _01441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06374__B2 genblk1\[1\].osc.clkdiv_C.cnt\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12995_ clknet_leaf_131_clk _00324_ net64 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.acc\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_56_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_56_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__08115__A2 _01180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11946_ genblk2\[10\].wave_shpr.div.b1\[11\] genblk2\[10\].wave_shpr.div.acc\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05768_ sky130_fd_sc_hd__and2b_1
XFILLER_0_98_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08520__C1 _02364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11877_ genblk2\[9\].wave_shpr.div.acc\[20\] _05707_ vssd1 vssd1 vccd1 vccd1 _05710_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_55_700 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13616_ clknet_leaf_94_clk _00929_ net160 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.fin_quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_55_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10828_ genblk2\[6\].wave_shpr.div.acc\[11\] genblk2\[6\].wave_shpr.div.b1\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04972_ sky130_fd_sc_hd__or2b_1
XFILLER_0_82_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08236__C _02365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13547_ clknet_leaf_109_clk _00862_ net152 vssd1 vssd1 vccd1 vccd1 sig_norm.b1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10759_ net981 _04918_ _04890_ _04921_ vssd1 vssd1 vccd1 vccd1 _00582_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13478_ clknet_leaf_99_clk _00795_ net168 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.quo\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_2_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12429_ genblk2\[11\].wave_shpr.div.acc\[20\] _06092_ vssd1 vssd1 vccd1 vccd1 _06094_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_124_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11186__A1 _01508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_23_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07970_ genblk1\[7\].osc.clkdiv_C.cnt\[15\] _01577_ _02668_ vssd1 vssd1 vccd1 vccd1
+ _02677_ sky130_fd_sc_hd__a21o_1
XFILLER_0_77_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06921_ _01761_ _01768_ _01769_ vssd1 vssd1 vccd1 vccd1 genblk1\[6\].osc.clkdiv_C.next_cnt\[5\]
+ sky130_fd_sc_hd__nor3_1
X_09640_ net983 _04109_ _04113_ _04132_ vssd1 vssd1 vccd1 vccd1 _00252_ sky130_fd_sc_hd__a22o_1
X_06852_ genblk1\[5\].osc.clkdiv_C.cnt\[10\] _01710_ genblk1\[5\].osc.clkdiv_C.cnt\[11\]
+ vssd1 vssd1 vccd1 vccd1 _01713_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09083__B _01201_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_93_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09571_ net965 _04076_ _04047_ _04079_ vssd1 vssd1 vccd1 vccd1 _00236_ sky130_fd_sc_hd__a22o_1
X_06783_ net851 _01654_ vssd1 vssd1 vccd1 vccd1 genblk1\[4\].osc.clkdiv_C.next_cnt\[17\]
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_47_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_47_clk sky130_fd_sc_hd__clkbuf_16
X_08522_ _02416_ _03228_ net2 _02364_ vssd1 vssd1 vccd1 vccd1 _03229_ sky130_fd_sc_hd__o211a_1
XFILLER_0_77_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07314__B1 genblk1\[11\].osc.clkdiv_C.cnt\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08453_ _02684_ _02681_ _02687_ _02526_ vssd1 vssd1 vccd1 vccd1 _03160_ sky130_fd_sc_hd__o31a_1
XFILLER_0_147_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout152_A net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_148_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07404_ genblk2\[0\].wave_shpr.div.busy _02149_ vssd1 vssd1 vccd1 vccd1 _02150_ sky130_fd_sc_hd__and2_1
X_08384_ _01437_ genblk1\[2\].osc.clkdiv_C.cnt\[5\] vssd1 vssd1 vccd1 vccd1 _03091_
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_18_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07335_ genblk1\[11\].osc.clkdiv_C.cnt\[2\] genblk1\[11\].osc.clkdiv_C.cnt\[1\] genblk1\[11\].osc.clkdiv_C.cnt\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02097_ sky130_fd_sc_hd__and3_1
XFILLER_0_34_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_33_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07266_ genblk1\[10\].osc.clkdiv_C.cnt\[6\] _02039_ vssd1 vssd1 vccd1 vccd1 _02042_
+ sky130_fd_sc_hd__nor2_1
X_09005_ net1151 vssd1 vssd1 vccd1 vccd1 _00067_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_115_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06217_ _01178_ _01176_ vssd1 vssd1 vccd1 vccd1 _01179_ sky130_fd_sc_hd__nor2_4
XFILLER_0_103_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07197_ genblk1\[9\].osc.clkdiv_C.cnt\[14\] _01981_ vssd1 vssd1 vccd1 vccd1 _01983_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_103_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06148_ _01118_ _01108_ vssd1 vssd1 vccd1 vccd1 _01120_ sky130_fd_sc_hd__and2b_1
XANTENNA__10924__A1 _02374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08593__A2 _02526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09790__A1 _03714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09907_ genblk2\[2\].wave_shpr.div.acc\[13\] _04320_ _04301_ vssd1 vssd1 vccd1 vccd1
+ _04321_ sky130_fd_sc_hd__mux2_1
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09838_ net261 _04257_ _04259_ net656 _04270_ vssd1 vssd1 vccd1 vccd1 _00312_ sky130_fd_sc_hd__a221o_1
XANTENNA__06356__A1 genblk1\[0\].osc.clkdiv_C.cnt\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout65_A net68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09769_ _04234_ vssd1 vssd1 vccd1 vccd1 _00279_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_38_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_38_clk sky130_fd_sc_hd__clkbuf_16
XTAP_2202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11800_ net1022 _05623_ _05624_ _05651_ vssd1 vssd1 vccd1 vccd1 _00893_ sky130_fd_sc_hd__a22o_1
XTAP_2224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12780_ clknet_leaf_40_clk _00113_ net116 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.b1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11731_ _05618_ vssd1 vssd1 vccd1 vccd1 _00857_ sky130_fd_sc_hd__clkbuf_1
XTAP_1534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10359__S _04637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_22_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11662_ genblk2\[9\].wave_shpr.div.acc\[17\] genblk2\[9\].wave_shpr.div.b1\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05554_ sky130_fd_sc_hd__or2b_1
X_13401_ clknet_leaf_92_clk _00720_ net143 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.quo\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10613_ genblk2\[6\].wave_shpr.div.b1\[1\] _04831_ _04637_ vssd1 vssd1 vccd1 vccd1
+ _04832_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_37_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11593_ genblk2\[8\].wave_shpr.div.acc\[10\] _05505_ _05493_ vssd1 vssd1 vccd1 vccd1
+ _05506_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_714 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10544_ genblk2\[5\].wave_shpr.div.acc\[8\] genblk2\[5\].wave_shpr.div.b1\[8\] vssd1
+ vssd1 vccd1 vccd1 _04772_ sky130_fd_sc_hd__or2b_1
X_13332_ clknet_leaf_9_clk net284 net54 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.acc\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13263_ clknet_leaf_0_clk _00586_ net38 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.acc\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10475_ net901 _04715_ _04690_ _04721_ vssd1 vssd1 vccd1 vccd1 _00498_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12214_ _05937_ _05950_ _05951_ vssd1 vssd1 vccd1 vccd1 _05952_ sky130_fd_sc_hd__a21o_1
X_13194_ clknet_leaf_127_clk _00517_ net67 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.fin_quo\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__09230__B1 _03839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12145_ _05779_ _05896_ vssd1 vssd1 vccd1 vccd1 _05897_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09184__A _03719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12076_ _05812_ vssd1 vssd1 vccd1 vccd1 _05844_ sky130_fd_sc_hd__clkbuf_4
X_11027_ net806 _05086_ _05093_ _05109_ vssd1 vssd1 vccd1 vccd1 _00662_ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06898__A2 _01367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_29_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_29_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_86_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12978_ clknet_leaf_124_clk net316 net72 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.quo\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07432__A _02170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11929_ _05745_ _05749_ _05750_ vssd1 vssd1 vccd1 vccd1 _05751_ sky130_fd_sc_hd__a21o_1
XFILLER_0_87_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_27_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_67_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_703 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_872 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_788 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07120_ _01432_ _01221_ vssd1 vssd1 vccd1 vccd1 _01920_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07051_ _01336_ _01183_ vssd1 vssd1 vccd1 vccd1 _01869_ sky130_fd_sc_hd__nor2_2
XFILLER_0_140_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12356__B1 _06010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_23_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09221__B1 _03840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09772__A1 _01256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10732__S _04821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10382__A2 _04657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09094__A _01367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07953_ genblk1\[7\].osc.clkdiv_C.cnt\[2\] _01732_ _02656_ genblk1\[7\].osc.clkdiv_C.cnt\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02660_ sky130_fd_sc_hd__o22a_1
XANTENNA__08327__A2 _02467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06904_ _01576_ _01757_ vssd1 vssd1 vccd1 vccd1 _01758_ sky130_fd_sc_hd__nand2_2
X_07884_ genblk2\[1\].wave_shpr.div.fin_quo\[6\] _02590_ vssd1 vssd1 vccd1 vccd1 _02591_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__10134__A2 _04451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07535__B1 _01099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09623_ net905 _04109_ _04113_ _04119_ vssd1 vssd1 vccd1 vccd1 _00248_ sky130_fd_sc_hd__a22o_1
X_06835_ net1105 _01700_ _01702_ vssd1 vssd1 vccd1 vccd1 genblk1\[5\].osc.clkdiv_C.next_cnt\[4\]
+ sky130_fd_sc_hd__a21oi_1
XANTENNA__11563__S _05417_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06766_ _01643_ vssd1 vssd1 vccd1 vccd1 genblk1\[4\].osc.clkdiv_C.next_cnt\[12\]
+ sky130_fd_sc_hd__clkbuf_1
X_09554_ _04055_ genblk1\[1\].osc.clkdiv_C.cnt\[15\] vssd1 vssd1 vccd1 vccd1 _04068_
+ sky130_fd_sc_hd__and2_1
X_08505_ genblk2\[2\].wave_shpr.div.fin_quo\[5\] _03113_ _03118_ _02224_ vssd1 vssd1
+ vccd1 vccd1 _03212_ sky130_fd_sc_hd__a31o_1
XFILLER_0_78_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09485_ _04031_ vssd1 vssd1 vccd1 vccd1 _00198_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06697_ genblk1\[4\].osc.clkdiv_C.cnt\[1\] _01436_ _01304_ genblk1\[4\].osc.clkdiv_C.cnt\[7\]
+ _01586_ vssd1 vssd1 vccd1 vccd1 _01587_ sky130_fd_sc_hd__a221o_1
XFILLER_0_53_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08436_ genblk2\[11\].wave_shpr.div.fin_quo\[2\] _02349_ _02351_ _02352_ vssd1 vssd1
+ vccd1 vccd1 _03143_ sky130_fd_sc_hd__nand4_1
XFILLER_0_65_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08367_ _03072_ _03073_ vssd1 vssd1 vccd1 vccd1 _03074_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10907__S _04848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07318_ genblk1\[11\].osc.clkdiv_C.cnt\[11\] _01262_ vssd1 vssd1 vccd1 vccd1 _02082_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__07066__A2 _01578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08298_ _02969_ _03003_ _03004_ vssd1 vssd1 vccd1 vccd1 _03005_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06274__B1 _01235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07249_ genblk1\[10\].osc.clkdiv_C.cnt\[1\] genblk1\[10\].osc.clkdiv_C.cnt\[0\] vssd1
+ vssd1 vccd1 vccd1 _02030_ sky130_fd_sc_hd__nand2_1
XFILLER_0_143_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10260_ genblk2\[4\].wave_shpr.div.acc\[10\] genblk2\[4\].wave_shpr.div.b1\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04572_ sky130_fd_sc_hd__or2b_1
XFILLER_0_103_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10191_ net1017 _04518_ _04490_ _04521_ vssd1 vssd1 vccd1 vccd1 _00414_ sky130_fd_sc_hd__a22o_1
XANTENNA__10642__S _04848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06421__A _01336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_896 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07526__B1 _01099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12901_ clknet_leaf_30_clk net589 net102 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.acc_next\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2010 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12832_ clknet_leaf_64_clk _00165_ net189 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.acc\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2021 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2032 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2043 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2054 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2065 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12763_ clknet_leaf_20_clk _00096_ net108 vssd1 vssd1 vccd1 vccd1 freq_div.state\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_96_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2076 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2087 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2098 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11714_ genblk2\[9\].wave_shpr.div.b1\[17\] genblk2\[9\].wave_shpr.div.acc\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05606_ sky130_fd_sc_hd__and2b_1
XTAP_1375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12694_ clknet_leaf_54_clk genblk1\[8\].osc.clkdiv_C.next_cnt\[7\] net172 vssd1 vssd1
+ vccd1 vccd1 genblk1\[8\].osc.clkdiv_C.cnt\[7\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_84_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11645_ _05414_ genblk2\[8\].wave_shpr.div.acc\[25\] genblk2\[8\].wave_shpr.div.acc\[26\]
+ vssd1 vssd1 vccd1 vccd1 _05543_ sky130_fd_sc_hd__or3b_1
XFILLER_0_140_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_154_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07057__A2 _01246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput15 pb[9] vssd1 vssd1 vccd1 vccd1 net15 sky130_fd_sc_hd__buf_4
XANTENNA__08083__A _02225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11576_ _05416_ vssd1 vssd1 vccd1 vccd1 _05493_ sky130_fd_sc_hd__clkbuf_4
X_13315_ clknet_leaf_9_clk net516 net48 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.quo\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10527_ genblk2\[4\].wave_shpr.div.i\[1\] genblk2\[4\].wave_shpr.div.i\[0\] genblk2\[4\].wave_shpr.div.i\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04758_ sky130_fd_sc_hd__and3_1
XANTENNA__06804__A2 _01362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10458_ net928 _04683_ _04690_ _04708_ vssd1 vssd1 vccd1 vccd1 _00494_ sky130_fd_sc_hd__a22o_1
X_13246_ clknet_leaf_11_clk net494 net56 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.acc\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_149_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13177_ clknet_leaf_130_clk _00502_ net65 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.acc\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10389_ net675 _04661_ _04655_ net602 _04662_ vssd1 vssd1 vccd1 vccd1 _00471_ sky130_fd_sc_hd__a221o_1
XANTENNA__07765__B1 _01208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12128_ _05772_ _05735_ vssd1 vssd1 vccd1 vccd1 _05884_ sky130_fd_sc_hd__or2b_1
X_12059_ _03833_ _02023_ vssd1 vssd1 vccd1 vccd1 _05834_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06620_ _01524_ _01525_ _01526_ vssd1 vssd1 vccd1 vccd1 _01527_ sky130_fd_sc_hd__and3_1
X_06551_ _01451_ _01466_ _01467_ vssd1 vssd1 vccd1 vccd1 genblk1\[2\].osc.clkdiv_C.next_cnt\[9\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_59_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09270_ genblk2\[0\].wave_shpr.div.b1\[0\] _03804_ genblk2\[0\].wave_shpr.div.acc\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03865_ sky130_fd_sc_hd__a21oi_1
X_06482_ genblk1\[1\].osc.clkdiv_C.cnt\[17\] _01407_ vssd1 vssd1 vccd1 vccd1 _01409_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_90_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08221_ _02793_ _02789_ genblk2\[5\].wave_shpr.div.fin_quo\[5\] vssd1 vssd1 vccd1
+ vccd1 _02928_ sky130_fd_sc_hd__or3b_1
XFILLER_0_7_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_894 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08152_ genblk1\[3\].osc.clkdiv_C.cnt\[5\] _01500_ _01250_ genblk1\[3\].osc.clkdiv_C.cnt\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02859_ sky130_fd_sc_hd__o22a_1
XANTENNA__07048__A2 _01182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_911 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10052__A1 _01870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07103_ _01887_ _01908_ vssd1 vssd1 vccd1 vccd1 _01909_ sky130_fd_sc_hd__nor2_1
XANTENNA_clkbuf_4_3_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08083_ _02225_ _02789_ vssd1 vssd1 vccd1 vccd1 _02790_ sky130_fd_sc_hd__and2_1
XFILLER_0_125_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_9_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_9_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_113_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_641 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07034_ genblk1\[8\].osc.clkdiv_C.cnt\[15\] _01359_ vssd1 vssd1 vccd1 vccd1 _01852_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_130_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_3_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11001__B1 _05056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08440__B _02403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08985_ _03669_ vssd1 vssd1 vccd1 vccd1 _00060_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07936_ _02637_ _02638_ _02641_ genblk2\[8\].wave_shpr.div.fin_quo\[6\] vssd1 vssd1
+ vccd1 vccd1 _02643_ sky130_fd_sc_hd__a31o_1
XANTENNA__07056__B _01498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07867_ _02469_ _02573_ _02529_ vssd1 vssd1 vccd1 vccd1 _02574_ sky130_fd_sc_hd__o21a_1
XANTENNA__11293__S _05222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06895__B _01362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09606_ _03992_ _03960_ vssd1 vssd1 vccd1 vccd1 _04106_ sky130_fd_sc_hd__or2b_1
XFILLER_0_3_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06818_ _01669_ _01559_ _01675_ genblk1\[5\].osc.clkdiv_C.cnt\[14\] _01689_ vssd1
+ vssd1 vccd1 vccd1 _01690_ sky130_fd_sc_hd__o221a_1
X_07798_ genblk1\[0\].osc.clkdiv_C.cnt\[15\] genblk1\[0\].osc.clkdiv_C.cnt\[14\] _01209_
+ vssd1 vssd1 vccd1 vccd1 _02505_ sky130_fd_sc_hd__or3_1
XFILLER_0_78_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09537_ genblk2\[1\].wave_shpr.div.quo\[15\] _04052_ _04053_ net511 _04059_ vssd1
+ vssd1 vccd1 vccd1 _00222_ sky130_fd_sc_hd__a221o_1
XFILLER_0_149_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06749_ _01630_ vssd1 vssd1 vccd1 vccd1 genblk1\[4\].osc.clkdiv_C.next_cnt\[8\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09468_ _03732_ net1047 _03733_ vssd1 vssd1 vccd1 vccd1 _00191_ sky130_fd_sc_hd__o21a_1
XFILLER_0_109_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08419_ _03001_ _03078_ _03055_ _03077_ vssd1 vssd1 vccd1 vccd1 _03126_ sky130_fd_sc_hd__o211a_1
XFILLER_0_93_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10637__S _04834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09399_ genblk2\[1\].wave_shpr.div.acc\[8\] genblk2\[1\].wave_shpr.div.b1\[8\] vssd1
+ vssd1 vccd1 vccd1 _03963_ sky130_fd_sc_hd__or2b_1
XFILLER_0_34_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11430_ _05243_ genblk2\[8\].wave_shpr.div.acc\[16\] vssd1 vssd1 vccd1 vccd1 _05406_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_117_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06416__A _01359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10043__A1 _03732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11361_ _05220_ _05248_ _05344_ _05251_ net1029 vssd1 vssd1 vccd1 vccd1 _00761_ sky130_fd_sc_hd__a32o_1
XFILLER_0_104_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_22_739 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10312_ genblk2\[4\].wave_shpr.div.fin_quo\[0\] _04623_ _00013_ vssd1 vssd1 vccd1
+ vccd1 _04624_ sky130_fd_sc_hd__mux2_1
X_13100_ clknet_leaf_136_clk _00427_ net42 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.acc\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_104_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11292_ _05192_ _05292_ vssd1 vssd1 vccd1 vccd1 _05293_ sky130_fd_sc_hd__xnor2_1
X_13031_ clknet_leaf_122_clk _00358_ net79 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.b1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10243_ _04454_ _04557_ _04558_ _04457_ net1079 vssd1 vssd1 vccd1 vccd1 _00429_ sky130_fd_sc_hd__a32o_1
X_10174_ net796 _04486_ _04490_ _04508_ vssd1 vssd1 vccd1 vccd1 _00410_ sky130_fd_sc_hd__a22o_1
Xfanout170 net171 vssd1 vssd1 vccd1 vccd1 net170 sky130_fd_sc_hd__buf_2
Xfanout181 net185 vssd1 vssd1 vccd1 vccd1 net181 sky130_fd_sc_hd__clkbuf_4
Xfanout192 net193 vssd1 vssd1 vccd1 vccd1 net192 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10401__A _04477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12815_ clknet_leaf_58_clk net579 net192 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.acc_next\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10806__B1 _04855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12746_ clknet_leaf_49_clk genblk1\[11\].osc.clkdiv_C.next_cnt\[5\] net108 vssd1
+ vssd1 vccd1 vccd1 genblk1\[11\].osc.clkdiv_C.cnt\[5\] sky130_fd_sc_hd__dfrtp_4
XTAP_1161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_151_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12677_ clknet_leaf_120_clk genblk1\[7\].osc.clkdiv_C.next_cnt\[8\] net142 vssd1
+ vssd1 vccd1 vccd1 genblk1\[7\].osc.clkdiv_C.cnt\[8\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__12328__A _03689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11628_ genblk2\[8\].wave_shpr.div.acc\[19\] _05531_ vssd1 vssd1 vccd1 vccd1 _05532_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__12023__A2 _05813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11559_ genblk2\[8\].wave_shpr.div.acc\[2\] _05479_ _05417_ vssd1 vssd1 vccd1 vccd1
+ _05480_ sky130_fd_sc_hd__mux2_1
Xhold607 genblk2\[1\].wave_shpr.div.acc\[5\] vssd1 vssd1 vccd1 vccd1 net825 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07986__B1 _02527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold618 genblk2\[2\].wave_shpr.div.acc\[7\] vssd1 vssd1 vccd1 vccd1 net836 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_52_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold629 genblk2\[1\].wave_shpr.div.acc\[9\] vssd1 vssd1 vccd1 vccd1 net847 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_122_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13229_ clknet_leaf_15_clk _00552_ net56 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.quo\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_901 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_912 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_923 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07157__A genblk1\[9\].osc.clkdiv_C.cnt\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_934 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_978 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08770_ _03454_ _03475_ _03476_ vssd1 vssd1 vccd1 vccd1 _03477_ sky130_fd_sc_hd__o21ai_2
XTAP_989 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11298__B1 _05283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07721_ genblk1\[1\].osc.clkdiv_C.cnt\[13\] _02425_ _02426_ _02427_ vssd1 vssd1 vccd1
+ vccd1 _02428_ sky130_fd_sc_hd__a211oi_2
XFILLER_0_18_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_79_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12002__S _05802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07652_ _02316_ _02357_ _02358_ vssd1 vssd1 vccd1 vccd1 _02359_ sky130_fd_sc_hd__or3b_1
XFILLER_0_79_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06603_ _01486_ _01487_ _01492_ _01504_ _01510_ vssd1 vssd1 vccd1 vccd1 _01511_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_125_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07583_ genblk1\[9\].osc.clkdiv_C.cnt\[2\] _01234_ _02287_ _02288_ _02289_ vssd1
+ vssd1 vccd1 vccd1 _02290_ sky130_fd_sc_hd__a221o_1
XFILLER_0_149_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09322_ _03786_ _03904_ vssd1 vssd1 vccd1 vccd1 _03905_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06534_ genblk1\[2\].osc.clkdiv_C.cnt\[3\] _01454_ vssd1 vssd1 vccd1 vccd1 _01457_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_146_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_861 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06465_ genblk1\[1\].osc.clkdiv_C.cnt\[11\] genblk1\[1\].osc.clkdiv_C.cnt\[10\] _01394_
+ vssd1 vssd1 vccd1 vccd1 _01398_ sky130_fd_sc_hd__and3_1
X_09253_ _03855_ _01169_ vssd1 vssd1 vccd1 vccd1 _03856_ sky130_fd_sc_hd__nor2_1
XANTENNA__10457__S _04704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12635__RESET_B net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_243 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08204_ _02303_ _02265_ genblk2\[9\].wave_shpr.div.fin_quo\[5\] vssd1 vssd1 vccd1
+ vccd1 _02911_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_56_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09184_ _03719_ vssd1 vssd1 vccd1 vccd1 _03819_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_133_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06396_ _01238_ _01262_ vssd1 vssd1 vccd1 vccd1 _01340_ sky130_fd_sc_hd__nor2_4
XFILLER_0_90_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06236__A _01174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_538 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08135_ genblk2\[4\].wave_shpr.div.fin_quo\[4\] _02841_ vssd1 vssd1 vccd1 vccd1 _02842_
+ sky130_fd_sc_hd__or2_1
XANTENNA__11222__B1 _05250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_886 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10981__A _05074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08066_ _01179_ _01222_ _01254_ _01171_ genblk1\[5\].osc.clkdiv_C.cnt\[0\] vssd1
+ vssd1 vccd1 vccd1 _02773_ sky130_fd_sc_hd__o311a_1
X_07017_ _01822_ _01840_ _01841_ vssd1 vssd1 vccd1 vccd1 genblk1\[7\].osc.clkdiv_C.next_cnt\[11\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_3_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06401__B1 _01344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10920__S _05042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08968_ _03655_ vssd1 vssd1 vccd1 vccd1 _00057_ sky130_fd_sc_hd__clkbuf_1
X_07919_ genblk1\[8\].osc.clkdiv_C.cnt\[7\] _01430_ _01858_ genblk1\[8\].osc.clkdiv_C.cnt\[5\]
+ _02625_ vssd1 vssd1 vccd1 vccd1 _02626_ sky130_fd_sc_hd__a221o_1
X_08899_ _03574_ _03600_ _03603_ _01157_ net1069 vssd1 vssd1 vccd1 vccd1 _00040_ sky130_fd_sc_hd__a32o_1
X_10930_ _03726_ _05049_ _03736_ vssd1 vssd1 vccd1 vccd1 _00625_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_98_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07901__B1 _01328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10861_ _04972_ _05003_ _05004_ vssd1 vssd1 vccd1 vccd1 _05005_ sky130_fd_sc_hd__a21o_1
XFILLER_0_94_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12600_ clknet_leaf_21_clk genblk1\[3\].osc.clkdiv_C.next_cnt\[3\] net97 vssd1 vssd1
+ vccd1 vccd1 genblk1\[3\].osc.clkdiv_C.cnt\[3\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_149_660 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13580_ clknet_leaf_76_clk _00895_ net207 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.acc\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10792_ _04817_ _04880_ _04943_ genblk2\[5\].wave_shpr.div.acc\[21\] vssd1 vssd1
+ vccd1 vccd1 _04946_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_66_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12531_ clknet_leaf_61_clk _00083_ net186 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.b1\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XPHY_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12462_ clknet_leaf_104_clk _00035_ net155 vssd1 vssd1 vccd1 vccd1 PWM.final_sample_in\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11413_ _05368_ _05387_ _05388_ vssd1 vssd1 vccd1 vccd1 _05389_ sky130_fd_sc_hd__a21o_1
XFILLER_0_152_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12393_ _05962_ _06066_ vssd1 vssd1 vccd1 vccd1 _06067_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11344_ _05331_ _05332_ vssd1 vssd1 vccd1 vccd1 _05333_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11275_ _05186_ _05181_ vssd1 vssd1 vccd1 vccd1 _05280_ sky130_fd_sc_hd__or2b_1
XFILLER_0_30_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13014_ clknet_leaf_132_clk _00343_ net60 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.acc\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09185__A2 _01344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10226_ _04417_ _04418_ vssd1 vssd1 vccd1 vccd1 _04547_ sky130_fd_sc_hd__and2b_1
XANTENNA__07196__A1 genblk1\[9\].osc.clkdiv_C.cnt\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10157_ net963 _04486_ _04490_ _04495_ vssd1 vssd1 vccd1 vccd1 _00406_ sky130_fd_sc_hd__a22o_1
Xhold4 modein.delay_in\[0\] vssd1 vssd1 vccd1 vccd1 net222 sky130_fd_sc_hd__clkbuf_2
X_10088_ net326 _04452_ _04456_ net794 vssd1 vssd1 vccd1 vccd1 _00376_ sky130_fd_sc_hd__a22o_1
XANTENNA__11227__A _05074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07424__B _02153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12729_ clknet_leaf_38_clk genblk1\[10\].osc.clkdiv_C.next_cnt\[6\] net115 vssd1
+ vssd1 vccd1 vccd1 genblk1\[10\].osc.clkdiv_C.cnt\[6\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_155_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06250_ genblk1\[0\].osc.clkdiv_C.cnt\[0\] _01211_ _01210_ genblk1\[0\].osc.clkdiv_C.cnt\[15\]
+ vssd1 vssd1 vccd1 vccd1 _01212_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_115_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11204__B1 _03687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06181_ sig_norm.busy _01152_ _01098_ vssd1 vssd1 vccd1 vccd1 _01153_ sky130_fd_sc_hd__and3_1
XFILLER_0_41_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07959__B1 _01925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold404 genblk2\[6\].wave_shpr.div.acc\[19\] vssd1 vssd1 vccd1 vccd1 net622 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11755__B2 net526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold415 _00231_ vssd1 vssd1 vccd1 vccd1 net633 sky130_fd_sc_hd__dlygate4sd3_1
Xhold426 _00484_ vssd1 vssd1 vccd1 vccd1 net644 sky130_fd_sc_hd__dlygate4sd3_1
Xhold437 genblk2\[0\].wave_shpr.div.quo\[1\] vssd1 vssd1 vccd1 vccd1 net655 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold448 _00481_ vssd1 vssd1 vccd1 vccd1 net666 sky130_fd_sc_hd__dlygate4sd3_1
X_09940_ genblk2\[2\].wave_shpr.div.acc\[22\] _04343_ vssd1 vssd1 vccd1 vccd1 _04345_
+ sky130_fd_sc_hd__xnor2_1
Xhold459 genblk2\[8\].wave_shpr.div.quo\[19\] vssd1 vssd1 vccd1 vccd1 net677 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09871_ _04183_ _04168_ vssd1 vssd1 vccd1 vccd1 _04293_ sky130_fd_sc_hd__or2b_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_110_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08822_ _03464_ _03526_ _03528_ vssd1 vssd1 vccd1 vccd1 _03529_ sky130_fd_sc_hd__or3_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1104 genblk2\[0\].wave_shpr.div.quo\[1\] vssd1 vssd1 vccd1 vccd1 net1322 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1115 genblk2\[4\].wave_shpr.div.quo\[3\] vssd1 vssd1 vccd1 vccd1 net1333 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1126 genblk2\[5\].wave_shpr.div.quo\[6\] vssd1 vssd1 vccd1 vccd1 net1344 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08753_ _03457_ _03459_ vssd1 vssd1 vccd1 vccd1 _03460_ sky130_fd_sc_hd__xnor2_1
XANTENNA_fanout182_A net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_24_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07704_ _02404_ _02405_ genblk2\[10\].wave_shpr.div.fin_quo\[6\] _02410_ vssd1 vssd1
+ vccd1 vccd1 _02411_ sky130_fd_sc_hd__and4b_1
XTAP_2609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08684_ _03114_ _03390_ _03122_ vssd1 vssd1 vccd1 vccd1 _03391_ sky130_fd_sc_hd__o21a_1
XFILLER_0_136_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07635_ genblk1\[11\].osc.clkdiv_C.cnt\[9\] _01190_ _01235_ genblk1\[11\].osc.clkdiv_C.cnt\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02342_ sky130_fd_sc_hd__o22a_1
XTAP_1919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07566_ _02269_ _02271_ _02272_ vssd1 vssd1 vccd1 vccd1 _02273_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09041__S _03708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09305_ _03778_ _03891_ vssd1 vssd1 vccd1 vccd1 _03892_ sky130_fd_sc_hd__xnor2_1
X_06517_ genblk1\[2\].osc.clkdiv_C.cnt\[5\] _01439_ _01442_ genblk1\[2\].osc.clkdiv_C.cnt\[9\]
+ vssd1 vssd1 vccd1 vccd1 _01443_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_36_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07497_ _02217_ _02215_ net760 vssd1 vssd1 vccd1 vccd1 _02219_ sky130_fd_sc_hd__or3_1
XANTENNA__08165__B _01508_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_118_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09236_ _03725_ genblk1\[0\].osc.clkdiv_C.cnt\[3\] vssd1 vssd1 vccd1 vccd1 _03846_
+ sky130_fd_sc_hd__and2_1
X_06448_ _01373_ _01385_ _01386_ vssd1 vssd1 vccd1 vccd1 genblk1\[1\].osc.clkdiv_C.next_cnt\[5\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_106_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_847 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09167_ genblk2\[0\].wave_shpr.div.fin_quo\[5\] net1334 _00001_ vssd1 vssd1 vccd1
+ vccd1 _03810_ sky130_fd_sc_hd__mux2_1
X_06379_ _01322_ vssd1 vssd1 vccd1 vccd1 _01323_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_32_834 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08118_ genblk1\[4\].osc.clkdiv_C.cnt\[2\] _01326_ _01213_ genblk1\[4\].osc.clkdiv_C.cnt\[3\]
+ vssd1 vssd1 vccd1 vccd1 _02825_ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09098_ _03734_ genblk2\[0\].wave_shpr.div.acc\[17\] vssd1 vssd1 vccd1 vccd1 _03746_
+ sky130_fd_sc_hd__or2_1
X_08049_ genblk1\[5\].osc.clkdiv_C.cnt\[11\] _01355_ vssd1 vssd1 vccd1 vccd1 _02756_
+ sky130_fd_sc_hd__nor2_1
Xhold960 genblk2\[4\].wave_shpr.div.b1\[6\] vssd1 vssd1 vccd1 vccd1 net1178 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06413__B _01356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold971 genblk1\[7\].osc.clkdiv_C.cnt\[12\] vssd1 vssd1 vccd1 vccd1 net1189 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout95_A net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11060_ net899 _05119_ _05126_ _05134_ vssd1 vssd1 vccd1 vccd1 _00670_ sky130_fd_sc_hd__a22o_1
Xhold982 genblk2\[7\].wave_shpr.div.b1\[4\] vssd1 vssd1 vccd1 vccd1 net1200 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold993 genblk2\[6\].wave_shpr.div.b1\[7\] vssd1 vssd1 vccd1 vccd1 net1211 sky130_fd_sc_hd__dlygate4sd3_1
X_10011_ genblk2\[3\].wave_shpr.div.b1\[14\] genblk2\[3\].wave_shpr.div.acc\[14\]
+ vssd1 vssd1 vccd1 vccd1 _04407_ sky130_fd_sc_hd__and2b_1
XFILLER_0_101_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11962_ genblk2\[10\].wave_shpr.div.acc\[23\] genblk2\[10\].wave_shpr.div.acc\[22\]
+ genblk2\[10\].wave_shpr.div.acc\[21\] _05783_ vssd1 vssd1 vccd1 vccd1 _05784_ sky130_fd_sc_hd__or4_1
XFILLER_0_99_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13701_ clknet_leaf_99_clk _01012_ net166 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.fin_quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06689__B1 _01578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10913_ net1201 _01819_ _04848_ vssd1 vssd1 vccd1 vccd1 _05041_ sky130_fd_sc_hd__mux2_1
X_11893_ genblk2\[9\].wave_shpr.div.acc\[25\] _05719_ vssd1 vssd1 vccd1 vccd1 _05721_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_79_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13632_ clknet_leaf_69_clk _00945_ net213 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.b1\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10844_ genblk2\[6\].wave_shpr.div.b1\[3\] genblk2\[6\].wave_shpr.div.acc\[3\] vssd1
+ vssd1 vccd1 vccd1 _04988_ sky130_fd_sc_hd__and2b_1
XFILLER_0_82_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_11_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13563_ clknet_leaf_57_clk net244 net184 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.quo\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10775_ genblk2\[5\].wave_shpr.div.acc\[16\] _04933_ _04907_ vssd1 vssd1 vccd1 vccd1
+ _04934_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12514_ clknet_leaf_106_clk _00025_ net153 vssd1 vssd1 vccd1 vccd1 PWM.start sky130_fd_sc_hd__dfrtp_4
XFILLER_0_54_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13494_ clknet_leaf_86_clk _00811_ net178 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.quo\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_136_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12445_ net960 _03947_ _03944_ _06104_ vssd1 vssd1 vccd1 vccd1 _01085_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12376_ _05954_ _06053_ vssd1 vssd1 vccd1 vccd1 _06054_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06604__A _01171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11327_ _05208_ _05319_ vssd1 vssd1 vccd1 vccd1 _05320_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11258_ _05260_ genblk1\[7\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 _05269_
+ sky130_fd_sc_hd__and2_1
X_10209_ _04413_ _04361_ vssd1 vssd1 vccd1 vccd1 _04535_ sky130_fd_sc_hd__or2b_1
X_11189_ _05234_ vssd1 vssd1 vccd1 vccd1 _00699_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10712__A2 _04853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08118__B1 _01213_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07420_ genblk2\[2\].wave_shpr.div.i\[1\] _02161_ genblk2\[2\].wave_shpr.div.i\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02162_ sky130_fd_sc_hd__or3b_1
XFILLER_0_147_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07170__A genblk1\[9\].osc.clkdiv_C.cnt\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07351_ genblk1\[11\].osc.clkdiv_C.cnt\[4\] genblk1\[11\].osc.clkdiv_C.cnt\[3\] _02097_
+ genblk1\[11\].osc.clkdiv_C.cnt\[5\] vssd1 vssd1 vccd1 vccd1 _02110_ sky130_fd_sc_hd__a31o_1
XFILLER_0_17_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_803 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06302_ genblk1\[0\].osc.clkdiv_C.cnt\[12\] _01263_ vssd1 vssd1 vccd1 vccd1 _01264_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_122_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07282_ _02027_ _02051_ _02052_ vssd1 vssd1 vccd1 vccd1 genblk1\[10\].osc.clkdiv_C.next_cnt\[11\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_17_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_14_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06233_ _01194_ _01175_ _01191_ vssd1 vssd1 vccd1 vccd1 _01195_ sky130_fd_sc_hd__nor3_1
X_09021_ _03692_ vssd1 vssd1 vccd1 vccd1 _03693_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_142_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06164_ _01133_ _01135_ vssd1 vssd1 vccd1 vccd1 _01136_ sky130_fd_sc_hd__nand2_1
Xhold201 _00460_ vssd1 vssd1 vccd1 vccd1 net419 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_14_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_599 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold212 genblk2\[11\].wave_shpr.div.quo\[0\] vssd1 vssd1 vccd1 vccd1 net430 sky130_fd_sc_hd__dlygate4sd3_1
Xhold223 genblk2\[2\].wave_shpr.div.quo\[10\] vssd1 vssd1 vccd1 vccd1 net441 sky130_fd_sc_hd__dlygate4sd3_1
Xhold234 _00393_ vssd1 vssd1 vccd1 vccd1 net452 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07801__C1 genblk1\[0\].osc.clkdiv_C.cnt\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold245 _00223_ vssd1 vssd1 vccd1 vccd1 net463 sky130_fd_sc_hd__dlygate4sd3_1
Xhold256 genblk2\[10\].wave_shpr.div.quo\[22\] vssd1 vssd1 vccd1 vccd1 net474 sky130_fd_sc_hd__dlygate4sd3_1
Xhold267 genblk2\[9\].wave_shpr.div.quo\[14\] vssd1 vssd1 vccd1 vccd1 net485 sky130_fd_sc_hd__dlygate4sd3_1
Xhold278 _00137_ vssd1 vssd1 vccd1 vccd1 net496 sky130_fd_sc_hd__dlygate4sd3_1
X_09923_ _04206_ _04332_ vssd1 vssd1 vccd1 vccd1 _04333_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09825__A _04069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold289 genblk2\[5\].wave_shpr.div.quo\[18\] vssd1 vssd1 vccd1 vccd1 net507 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10470__S _04704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09854_ _04174_ _04175_ vssd1 vssd1 vccd1 vccd1 _04280_ sky130_fd_sc_hd__xnor2_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09544__B genblk1\[1\].osc.clkdiv_C.cnt\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08805_ _03511_ vssd1 vssd1 vccd1 vccd1 _03512_ sky130_fd_sc_hd__inv_2
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09785_ genblk2\[3\].wave_shpr.div.b1\[14\] _04242_ _04238_ vssd1 vssd1 vccd1 vccd1
+ _04243_ sky130_fd_sc_hd__mux2_1
XFILLER_0_147_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06997_ genblk1\[7\].osc.clkdiv_C.cnt\[4\] _01827_ vssd1 vssd1 vccd1 vccd1 _01829_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__07580__A1 _01432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08736_ _03439_ _03441_ _03442_ vssd1 vssd1 vccd1 vccd1 _03443_ sky130_fd_sc_hd__nand3b_2
XTAP_2406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_72_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08667_ _03372_ _03373_ genblk2\[4\].wave_shpr.div.fin_quo\[3\] _02362_ vssd1 vssd1
+ vccd1 vccd1 _03374_ sky130_fd_sc_hd__a2bb2o_1
XTAP_1705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07618_ genblk1\[11\].osc.clkdiv_C.cnt\[4\] _02064_ vssd1 vssd1 vccd1 vccd1 _02325_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_138_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08598_ genblk2\[3\].wave_shpr.div.fin_quo\[0\] _02592_ _02467_ genblk2\[3\].wave_shpr.div.fin_quo\[1\]
+ _02939_ vssd1 vssd1 vccd1 vccd1 _03305_ sky130_fd_sc_hd__a221o_1
XFILLER_0_49_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09085__A1 _03714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07549_ net1157 net1132 PWM.start vssd1 vssd1 vccd1 vccd1 _02258_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_87_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10560_ _04779_ _04786_ _04787_ vssd1 vssd1 vccd1 vccd1 _04788_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07635__A2 _01190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_119_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_836 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_130_clk_A clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09219_ _03838_ vssd1 vssd1 vccd1 vccd1 _03840_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__10645__S _04848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10491_ genblk2\[4\].wave_shpr.div.acc\[16\] _04733_ _04704_ vssd1 vssd1 vccd1 vccd1
+ _04734_ sky130_fd_sc_hd__mux2_1
XFILLER_0_122_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12230_ _05929_ _05966_ _05967_ vssd1 vssd1 vccd1 vccd1 _05968_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_10_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06424__A _01365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12161_ genblk2\[10\].wave_shpr.div.acc\[21\] _05783_ _05899_ vssd1 vssd1 vccd1 vccd1
+ _05908_ sky130_fd_sc_hd__or3_1
XANTENNA__07239__B _01215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10942__A2 _05052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11112_ genblk2\[7\].wave_shpr.div.acc\[9\] genblk2\[7\].wave_shpr.div.b1\[9\] vssd1
+ vssd1 vccd1 vccd1 _05172_ sky130_fd_sc_hd__or2b_1
XANTENNA__10047__A1_N _03727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12092_ net977 _05844_ _05850_ _05856_ vssd1 vssd1 vccd1 vccd1 _00980_ sky130_fd_sc_hd__a22o_1
Xhold790 genblk2\[4\].wave_shpr.div.acc\[11\] vssd1 vssd1 vccd1 vccd1 net1008 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_leaf_25_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11043_ genblk2\[6\].wave_shpr.div.acc\[12\] _05121_ _05105_ vssd1 vssd1 vccd1 vccd1
+ _05122_ sky130_fd_sc_hd__mux2_1
Xclkbuf_4_3_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_3_0_clk sky130_fd_sc_hd__clkbuf_8
XANTENNA__06374__A2 _01311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12994_ clknet_leaf_131_clk _00323_ net64 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.acc\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11945_ _05738_ _05765_ _05766_ vssd1 vssd1 vccd1 vccd1 _05767_ sky130_fd_sc_hd__a21o_1
XFILLER_0_86_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08520__B1 net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11505__A _05441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11876_ genblk2\[9\].wave_shpr.div.acc\[20\] _05707_ vssd1 vssd1 vccd1 vccd1 _05709_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_28_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13615_ clknet_leaf_94_clk _00928_ net160 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.fin_quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_145_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09076__A1 _01483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10827_ genblk2\[6\].wave_shpr.div.acc\[12\] genblk2\[6\].wave_shpr.div.b1\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04971_ sky130_fd_sc_hd__or2b_1
XFILLER_0_67_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13546_ clknet_leaf_109_clk _00861_ net152 vssd1 vssd1 vccd1 vccd1 sig_norm.b1\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10758_ genblk2\[5\].wave_shpr.div.acc\[12\] _04920_ _04907_ vssd1 vssd1 vccd1 vccd1
+ _04921_ sky130_fd_sc_hd__mux2_1
XANTENNA__07626__A2 _01241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13597__RESET_B net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13477_ clknet_leaf_72_clk _00794_ net216 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.b1\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10689_ _04869_ genblk1\[5\].osc.clkdiv_C.cnt\[10\] vssd1 vssd1 vccd1 vccd1 _04872_
+ sky130_fd_sc_hd__and2_1
XANTENNA__12336__A _03689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12428_ net1203 _06072_ _06073_ _06093_ vssd1 vssd1 vccd1 vccd1 _01079_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_2_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12359_ _05947_ _05939_ vssd1 vssd1 vccd1 vccd1 _06041_ sky130_fd_sc_hd__or2b_1
XFILLER_0_77_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06920_ genblk1\[6\].osc.clkdiv_C.cnt\[4\] _01765_ genblk1\[6\].osc.clkdiv_C.cnt\[5\]
+ vssd1 vssd1 vccd1 vccd1 _01769_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12071__A _03719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06851_ genblk1\[5\].osc.clkdiv_C.cnt\[10\] _01710_ _01712_ _01694_ vssd1 vssd1 vccd1
+ vccd1 genblk1\[5\].osc.clkdiv_C.next_cnt\[10\] sky130_fd_sc_hd__o211a_1
XANTENNA__11894__B1 _03694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09551__A2 _04042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09083__C _01363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12479__RESET_B net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06500__C net35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09570_ genblk2\[1\].wave_shpr.div.acc\[2\] _04078_ _04011_ vssd1 vssd1 vccd1 vccd1
+ _04079_ sky130_fd_sc_hd__mux2_1
X_06782_ _01655_ vssd1 vssd1 vccd1 vccd1 genblk1\[4\].osc.clkdiv_C.next_cnt\[16\]
+ sky130_fd_sc_hd__clkbuf_1
X_08521_ _02216_ _02552_ genblk2\[10\].wave_shpr.div.fin_quo\[0\] vssd1 vssd1 vccd1
+ vccd1 _03228_ sky130_fd_sc_hd__and3_1
XFILLER_0_26_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_77_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08452_ _02682_ _02687_ _02684_ vssd1 vssd1 vccd1 vccd1 _03159_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07403_ genblk2\[0\].wave_shpr.div.i\[1\] _02148_ genblk2\[0\].wave_shpr.div.i\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02149_ sky130_fd_sc_hd__or3b_1
XFILLER_0_148_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_92_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_46_723 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08383_ _03087_ _03088_ _03089_ vssd1 vssd1 vccd1 vccd1 _03090_ sky130_fd_sc_hd__o21a_1
XFILLER_0_58_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout145_A net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06228__B _01189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07334_ _02096_ vssd1 vssd1 vccd1 vccd1 genblk1\[11\].osc.clkdiv_C.next_cnt\[1\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07617__A2 _01513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07265_ genblk1\[10\].osc.clkdiv_C.cnt\[6\] _02039_ vssd1 vssd1 vccd1 vccd1 _02041_
+ sky130_fd_sc_hd__and2_1
XANTENNA__10465__S _04704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13267__RESET_B net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09004_ net1150 sig_norm.quo\[3\] _01154_ vssd1 vssd1 vccd1 vccd1 _03682_ sky130_fd_sc_hd__mux2_1
X_06216_ freq_div.state\[1\] vssd1 vssd1 vccd1 vccd1 _01178_ sky130_fd_sc_hd__buf_4
X_07196_ genblk1\[9\].osc.clkdiv_C.cnt\[13\] _01979_ _01982_ vssd1 vssd1 vccd1 vccd1
+ genblk1\[9\].osc.clkdiv_C.next_cnt\[13\] sky130_fd_sc_hd__o21a_1
X_06147_ net1 net7 _01118_ vssd1 vssd1 vccd1 vccd1 _01119_ sky130_fd_sc_hd__and3_1
XFILLER_0_41_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09906_ _04198_ _04319_ vssd1 vssd1 vccd1 vccd1 _04320_ sky130_fd_sc_hd__xnor2_1
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09837_ _04269_ genblk1\[2\].osc.clkdiv_C.cnt\[12\] vssd1 vssd1 vccd1 vccd1 _04270_
+ sky130_fd_sc_hd__and2_1
XANTENNA__10213__B _04480_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09768_ genblk2\[3\].wave_shpr.div.b1\[6\] _01262_ _04039_ vssd1 vssd1 vccd1 vccd1
+ _04234_ sky130_fd_sc_hd__mux2_1
XTAP_2203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout58_A net85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08719_ _03420_ _03421_ _03383_ _03395_ vssd1 vssd1 vccd1 vccd1 _03426_ sky130_fd_sc_hd__o211a_1
XANTENNA__07803__A net31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09699_ genblk2\[2\].wave_shpr.div.b1\[3\] genblk2\[2\].wave_shpr.div.acc\[3\] vssd1
+ vssd1 vccd1 vccd1 _04179_ sky130_fd_sc_hd__and2b_1
XFILLER_0_69_848 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_68_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11730_ genblk2\[9\].wave_shpr.div.fin_quo\[4\] genblk2\[9\].wave_shpr.div.quo\[3\]
+ _00023_ vssd1 vssd1 vccd1 vccd1 _05618_ sky130_fd_sc_hd__mux2_1
XTAP_1524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07856__A2 net31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06419__A _01362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11661_ net319 _05552_ _05553_ vssd1 vssd1 vccd1 vccd1 _00852_ sky130_fd_sc_hd__a21oi_1
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13400_ clknet_leaf_119_clk net422 net143 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.quo\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10612_ _01738_ vssd1 vssd1 vccd1 vccd1 _04831_ sky130_fd_sc_hd__inv_2
XFILLER_0_107_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_9_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11592_ _05393_ _05504_ vssd1 vssd1 vccd1 vccd1 _05505_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_153_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13331_ clknet_leaf_24_clk _00652_ net92 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.acc_next\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_106_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10543_ genblk2\[5\].wave_shpr.div.acc\[9\] genblk2\[5\].wave_shpr.div.b1\[9\] vssd1
+ vssd1 vccd1 vccd1 _04771_ sky130_fd_sc_hd__or2b_1
XFILLER_0_107_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08281__A2 _02521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13262_ clknet_leaf_0_clk _00585_ net38 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.acc\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10474_ genblk2\[4\].wave_shpr.div.acc\[12\] _04720_ _04704_ vssd1 vssd1 vccd1 vccd1
+ _04721_ sky130_fd_sc_hd__mux2_1
X_12213_ genblk2\[11\].wave_shpr.div.b1\[5\] genblk2\[11\].wave_shpr.div.acc\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05951_ sky130_fd_sc_hd__and2b_1
XFILLER_0_20_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13193_ clknet_leaf_118_clk _00516_ net138 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.i\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_12144_ _05780_ _05731_ vssd1 vssd1 vccd1 vccd1 _05896_ sky130_fd_sc_hd__or2b_1
XFILLER_0_138_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06595__A2 _01363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07792__A1 _01246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12075_ _05842_ _05843_ net1118 _05813_ vssd1 vssd1 vccd1 vccd1 _00976_ sky130_fd_sc_hd__a2bb2o_1
X_11026_ genblk2\[6\].wave_shpr.div.acc\[8\] _05108_ _05105_ vssd1 vssd1 vccd1 vccd1
+ _05109_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12977_ clknet_leaf_123_clk _00306_ net72 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.quo\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11235__A _05074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_656 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11928_ genblk2\[10\].wave_shpr.div.b1\[2\] genblk2\[10\].wave_shpr.div.acc\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05750_ sky130_fd_sc_hd__and2b_1
XFILLER_0_75_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11859_ genblk2\[9\].wave_shpr.div.acc\[15\] _05696_ _05673_ vssd1 vssd1 vccd1 vccd1
+ _05697_ sky130_fd_sc_hd__mux2_1
XFILLER_0_145_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_7_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_715 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13529_ clknet_leaf_98_clk _00846_ net169 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.acc\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11800__B1 _05624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_12_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_153_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07050_ genblk1\[8\].osc.clkdiv_C.cnt\[9\] _01865_ _01867_ vssd1 vssd1 vccd1 vccd1
+ _01868_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_112_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_11_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_10_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__07232__B1 _02013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07783__A1 _01200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07952_ genblk1\[7\].osc.clkdiv_C.cnt\[0\] _01801_ _02657_ _02658_ vssd1 vssd1 vccd1
+ vccd1 _02659_ sky130_fd_sc_hd__a31o_1
X_06903_ _01325_ _01327_ vssd1 vssd1 vccd1 vccd1 _01757_ sky130_fd_sc_hd__nor2_2
X_07883_ _02464_ genblk2\[1\].wave_shpr.div.fin_quo\[5\] _02461_ vssd1 vssd1 vccd1
+ vccd1 _02590_ sky130_fd_sc_hd__or3b_1
X_09622_ genblk2\[1\].wave_shpr.div.acc\[14\] _04118_ _04095_ vssd1 vssd1 vccd1 vccd1
+ _04119_ sky130_fd_sc_hd__mux2_1
X_06834_ genblk1\[5\].osc.clkdiv_C.cnt\[4\] _01700_ _01694_ vssd1 vssd1 vccd1 vccd1
+ _01702_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_37_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09553_ genblk2\[1\].wave_shpr.div.quo\[23\] _04042_ _04046_ net340 _04067_ vssd1
+ vssd1 vccd1 vccd1 _00230_ sky130_fd_sc_hd__a221o_1
X_06765_ _01599_ _01640_ _01642_ vssd1 vssd1 vccd1 vccd1 _01643_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08504_ _03113_ _03118_ genblk2\[2\].wave_shpr.div.fin_quo\[5\] vssd1 vssd1 vccd1
+ vccd1 _03211_ sky130_fd_sc_hd__a21oi_1
X_09484_ genblk2\[2\].wave_shpr.div.b1\[9\] _01302_ _04024_ vssd1 vssd1 vccd1 vccd1
+ _04031_ sky130_fd_sc_hd__mux2_1
XANTENNA__07838__A2 _02539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06239__A _01200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06696_ genblk1\[4\].osc.clkdiv_C.cnt\[3\] _01326_ _01574_ genblk1\[4\].osc.clkdiv_C.cnt\[12\]
+ vssd1 vssd1 vccd1 vccd1 _01586_ sky130_fd_sc_hd__a22o_1
XFILLER_0_148_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08435_ net33 _02350_ _02352_ genblk2\[11\].wave_shpr.div.fin_quo\[2\] vssd1 vssd1
+ vccd1 vccd1 _03142_ sky130_fd_sc_hd__a31o_1
XFILLER_0_92_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_59_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_108_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08366_ _02938_ _02944_ vssd1 vssd1 vccd1 vccd1 _03073_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08454__A _02216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07317_ genblk1\[11\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 _02081_ sky130_fd_sc_hd__inv_2
XANTENNA__10195__S _04507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08297_ _03002_ _02970_ vssd1 vssd1 vccd1 vccd1 _03004_ sky130_fd_sc_hd__and2b_1
XFILLER_0_33_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08173__B _01858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_104_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07248_ genblk1\[10\].osc.clkdiv_C.cnt\[1\] genblk1\[10\].osc.clkdiv_C.cnt\[0\] vssd1
+ vssd1 vccd1 vccd1 _02029_ sky130_fd_sc_hd__or2_1
XFILLER_0_103_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_5_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10358__B1 _04647_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07179_ _01971_ vssd1 vssd1 vccd1 vccd1 genblk1\[9\].osc.clkdiv_C.next_cnt\[7\] sky130_fd_sc_hd__clkbuf_1
XANTENNA__07223__B1 _01196_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10190_ genblk2\[3\].wave_shpr.div.acc\[12\] _04520_ _04507_ vssd1 vssd1 vccd1 vccd1
+ _04521_ sky130_fd_sc_hd__mux2_1
XANTENNA__06702__A _01171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09515__A2 _04043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12900_ clknet_leaf_30_clk net633 net102 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.quo\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07533__A _02248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12831_ clknet_leaf_64_clk _00164_ net189 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.acc\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2000 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2011 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2022 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2033 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2044 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12762_ clknet_leaf_20_clk _00095_ net109 vssd1 vssd1 vccd1 vccd1 freq_div.state\[1\]
+ sky130_fd_sc_hd__dfstp_2
XTAP_2055 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2066 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2077 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2088 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11713_ _05555_ _05603_ _05604_ vssd1 vssd1 vccd1 vccd1 _05605_ sky130_fd_sc_hd__o21bai_2
XTAP_2099 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12693_ clknet_leaf_54_clk genblk1\[8\].osc.clkdiv_C.next_cnt\[6\] net172 vssd1 vssd1
+ vccd1 vccd1 genblk1\[8\].osc.clkdiv_C.cnt\[6\] sky130_fd_sc_hd__dfrtp_4
XTAP_1376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11644_ net1052 _05448_ _05445_ _05542_ vssd1 vssd1 vccd1 vccd1 _00846_ sky130_fd_sc_hd__a22o_1
XFILLER_0_83_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xinput16 reset vssd1 vssd1 vccd1 vccd1 net16 sky130_fd_sc_hd__clkbuf_8
XANTENNA__08254__A2 _02733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11575_ _05385_ _05491_ vssd1 vssd1 vccd1 vccd1 _05492_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08083__B _02789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13314_ clknet_leaf_12_clk _00635_ net54 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.quo\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10526_ genblk2\[4\].wave_shpr.div.i\[1\] genblk2\[4\].wave_shpr.div.i\[0\] genblk2\[4\].wave_shpr.div.i\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04757_ sky130_fd_sc_hd__a21o_1
XFILLER_0_52_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13245_ clknet_leaf_11_clk net325 net54 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.acc_next\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09203__A1 _01302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10457_ genblk2\[4\].wave_shpr.div.acc\[8\] _04707_ _04704_ vssd1 vssd1 vccd1 vccd1
+ _04708_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08006__A2 _01735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07708__A _02225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13176_ clknet_leaf_130_clk _00501_ net65 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.acc\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10388_ _04477_ genblk1\[4\].osc.clkdiv_C.cnt\[3\] vssd1 vssd1 vccd1 vccd1 _04662_
+ sky130_fd_sc_hd__and2_1
XANTENNA__07765__A1 genblk1\[0\].osc.clkdiv_C.cnt\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07765__B2 genblk1\[0\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12127_ _05815_ vssd1 vssd1 vccd1 vccd1 _05883_ sky130_fd_sc_hd__clkbuf_4
X_12058_ net383 _05823_ _05825_ net440 _05833_ vssd1 vssd1 vccd1 vccd1 _00969_ sky130_fd_sc_hd__a221o_1
X_11009_ genblk2\[6\].wave_shpr.div.acc\[4\] _05095_ _05023_ vssd1 vssd1 vccd1 vccd1
+ _05096_ sky130_fd_sc_hd__mux2_1
XANTENNA__10521__A0 _04654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06689__A2_N _01574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06550_ genblk1\[2\].osc.clkdiv_C.cnt\[9\] _01464_ vssd1 vssd1 vccd1 vccd1 _01467_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_48_818 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_59_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06481_ genblk1\[1\].osc.clkdiv_C.cnt\[16\] _01405_ _01408_ vssd1 vssd1 vccd1 vccd1
+ genblk1\[1\].osc.clkdiv_C.next_cnt\[16\] sky130_fd_sc_hd__o21a_1
XFILLER_0_114_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08220_ _02925_ _02926_ _02897_ vssd1 vssd1 vccd1 vccd1 _02927_ sky130_fd_sc_hd__o21ai_1
XANTENNA__12026__B1 _05817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_28_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_71_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08151_ genblk1\[3\].osc.clkdiv_C.cnt\[4\] _01250_ _01514_ genblk1\[3\].osc.clkdiv_C.cnt\[3\]
+ _02857_ vssd1 vssd1 vccd1 vccd1 _02858_ sky130_fd_sc_hd__a221o_1
XFILLER_0_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07102_ genblk1\[8\].osc.clkdiv_C.cnt\[12\] genblk1\[8\].osc.clkdiv_C.cnt\[11\] _01904_
+ vssd1 vssd1 vccd1 vccd1 _01908_ sky130_fd_sc_hd__and3_1
XANTENNA__06256__A1 genblk1\[0\].osc.clkdiv_C.cnt\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08082_ _02784_ _02788_ genblk1\[5\].osc.clkdiv_C.cnt\[16\] genblk1\[5\].osc.clkdiv_C.cnt\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02789_ sky130_fd_sc_hd__a211o_4
XFILLER_0_31_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_99_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_3_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07033_ net848 _01850_ vssd1 vssd1 vccd1 vccd1 genblk1\[7\].osc.clkdiv_C.next_cnt\[17\]
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_2_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_11_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout108_A net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08984_ net1156 _03668_ _01158_ vssd1 vssd1 vccd1 vccd1 _03669_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09833__A _04069_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07935_ _02637_ genblk2\[8\].wave_shpr.div.fin_quo\[6\] _02638_ _02641_ _02223_ vssd1
+ vssd1 vccd1 vccd1 _02642_ sky130_fd_sc_hd__a41o_1
XANTENNA__10979__A _05074_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09552__B genblk1\[1\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07866_ net17 _02552_ genblk2\[1\].wave_shpr.div.fin_quo\[0\] vssd1 vssd1 vccd1 vccd1
+ _02573_ sky130_fd_sc_hd__and3_1
X_09605_ net366 _04076_ _04080_ _04105_ vssd1 vssd1 vccd1 vccd1 _00244_ sky130_fd_sc_hd__a22o_1
X_06817_ _01681_ _01686_ _01687_ _01688_ vssd1 vssd1 vccd1 vccd1 _01689_ sky130_fd_sc_hd__and4bb_1
X_07797_ _02493_ _02500_ _02502_ _02498_ _02503_ vssd1 vssd1 vccd1 vccd1 _02504_ sky130_fd_sc_hd__a32oi_1
XANTENNA__07072__B genblk1\[8\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09536_ _04058_ _01307_ vssd1 vssd1 vccd1 vccd1 _04059_ sky130_fd_sc_hd__nor2_1
X_06748_ _01599_ _01628_ _01629_ vssd1 vssd1 vccd1 vccd1 _01630_ sky130_fd_sc_hd__and3_1
XFILLER_0_149_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09467_ _04021_ vssd1 vssd1 vccd1 vccd1 _00190_ sky130_fd_sc_hd__clkbuf_1
X_06679_ genblk1\[4\].osc.clkdiv_C.cnt\[15\] _01363_ _01242_ _01568_ genblk1\[4\].osc.clkdiv_C.cnt\[17\]
+ vssd1 vssd1 vccd1 vccd1 _01569_ sky130_fd_sc_hd__a221o_1
XANTENNA__10918__S _05042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08418_ _03083_ _03124_ vssd1 vssd1 vccd1 vccd1 _03125_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_19_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09398_ genblk2\[1\].wave_shpr.div.acc\[9\] genblk2\[1\].wave_shpr.div.b1\[9\] vssd1
+ vssd1 vccd1 vccd1 _03962_ sky130_fd_sc_hd__or2b_1
XANTENNA__08184__A _02225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08349_ _02789_ _02792_ vssd1 vssd1 vccd1 vccd1 _03056_ sky130_fd_sc_hd__and2b_1
XFILLER_0_46_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_123_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_567 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11360_ _05342_ _05343_ vssd1 vssd1 vccd1 vccd1 _05344_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10311_ _04622_ vssd1 vssd1 vccd1 vccd1 _04623_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_132_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11291_ _05193_ _05175_ vssd1 vssd1 vccd1 vccd1 _05292_ sky130_fd_sc_hd__or2b_1
XFILLER_0_104_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13030_ clknet_leaf_122_clk _00357_ net79 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.b1\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10242_ genblk2\[3\].wave_shpr.div.i\[1\] genblk2\[3\].wave_shpr.div.i\[0\] vssd1
+ vssd1 vccd1 vccd1 _04558_ sky130_fd_sc_hd__nand2_1
XFILLER_0_131_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10173_ genblk2\[3\].wave_shpr.div.acc\[8\] _04506_ _04507_ vssd1 vssd1 vccd1 vccd1
+ _04508_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout160 net162 vssd1 vssd1 vccd1 vccd1 net160 sky130_fd_sc_hd__clkbuf_4
Xfanout171 net16 vssd1 vssd1 vccd1 vccd1 net171 sky130_fd_sc_hd__buf_4
Xfanout182 net185 vssd1 vssd1 vccd1 vccd1 net182 sky130_fd_sc_hd__buf_2
Xfanout193 net195 vssd1 vssd1 vccd1 vccd1 net193 sky130_fd_sc_hd__buf_2
XFILLER_0_97_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12814_ clknet_leaf_58_clk net455 net192 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.quo\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12745_ clknet_leaf_50_clk genblk1\[11\].osc.clkdiv_C.next_cnt\[4\] net108 vssd1
+ vssd1 vccd1 vccd1 genblk1\[11\].osc.clkdiv_C.cnt\[4\] sky130_fd_sc_hd__dfrtp_4
XTAP_1151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12676_ clknet_leaf_120_clk genblk1\[7\].osc.clkdiv_C.next_cnt\[7\] net82 vssd1 vssd1
+ vccd1 vccd1 genblk1\[7\].osc.clkdiv_C.cnt\[7\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_72_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11627_ genblk2\[8\].wave_shpr.div.acc\[18\] _05529_ vssd1 vssd1 vccd1 vccd1 _05531_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_127_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_52_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11558_ _05377_ _05478_ vssd1 vssd1 vccd1 vccd1 _05479_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold608 genblk2\[6\].wave_shpr.div.acc\[7\] vssd1 vssd1 vccd1 vccd1 net826 sky130_fd_sc_hd__dlygate4sd3_1
X_10509_ genblk2\[4\].wave_shpr.div.acc\[22\] _04657_ _04722_ _04746_ vssd1 vssd1
+ vccd1 vccd1 _00507_ sky130_fd_sc_hd__a22o_1
Xhold619 genblk1\[6\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 net837 sky130_fd_sc_hd__buf_1
XFILLER_0_111_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12344__A genblk2\[11\].wave_shpr.div.acc_next\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_11489_ _02171_ net1239 vssd1 vssd1 vccd1 vccd1 _05440_ sky130_fd_sc_hd__and2_1
XANTENNA__09188__B1 _03705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13228_ clknet_leaf_125_clk net309 net69 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.quo\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_21_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_902 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13159_ clknet_leaf_121_clk net644 net78 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.acc_next\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07157__B genblk1\[9\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_935 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_968 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_979 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07720_ genblk1\[1\].osc.clkdiv_C.cnt\[15\] _01309_ _01208_ genblk1\[1\].osc.clkdiv_C.cnt\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02427_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07651_ _02349_ _02351_ _02356_ genblk2\[11\].wave_shpr.div.fin_quo\[6\] vssd1 vssd1
+ vccd1 vccd1 _02358_ sky130_fd_sc_hd__a31o_1
XFILLER_0_79_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06602_ genblk1\[3\].osc.clkdiv_C.cnt\[0\] _01484_ _01505_ _01506_ _01509_ vssd1
+ vssd1 vccd1 vccd1 _01510_ sky130_fd_sc_hd__a221o_1
X_07582_ genblk1\[9\].osc.clkdiv_C.cnt\[1\] _01230_ _01221_ vssd1 vssd1 vccd1 vccd1
+ _02289_ sky130_fd_sc_hd__and3_1
XFILLER_0_149_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09321_ _03787_ _03751_ vssd1 vssd1 vccd1 vccd1 _03904_ sky130_fd_sc_hd__or2b_1
XFILLER_0_48_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06533_ genblk1\[2\].osc.clkdiv_C.cnt\[3\] _01454_ vssd1 vssd1 vccd1 vccd1 _01456_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_8_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11470__A1 _01946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09252_ _03719_ vssd1 vssd1 vccd1 vccd1 _03855_ sky130_fd_sc_hd__buf_6
X_06464_ genblk1\[1\].osc.clkdiv_C.cnt\[10\] _01394_ genblk1\[1\].osc.clkdiv_C.cnt\[11\]
+ vssd1 vssd1 vccd1 vccd1 _01397_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_35_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_29_873 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08203_ _02901_ _02905_ _02909_ _02419_ vssd1 vssd1 vccd1 vccd1 _02910_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09183_ _03818_ vssd1 vssd1 vccd1 vccd1 _00109_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_255 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06395_ genblk1\[1\].osc.clkdiv_C.cnt\[15\] _01210_ _01337_ genblk1\[1\].osc.clkdiv_C.cnt\[12\]
+ vssd1 vssd1 vccd1 vccd1 _01339_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_180 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08134_ genblk2\[4\].wave_shpr.div.fin_quo\[3\] _02840_ vssd1 vssd1 vccd1 vccd1 _02841_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_71_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08065_ _02770_ _02771_ vssd1 vssd1 vccd1 vccd1 _02772_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_12_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07016_ genblk1\[7\].osc.clkdiv_C.cnt\[11\] genblk1\[7\].osc.clkdiv_C.cnt\[10\] _01837_
+ vssd1 vssd1 vccd1 vccd1 _01841_ sky130_fd_sc_hd__and3_1
XFILLER_0_101_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07729__A1 _01360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06401__A1 _01342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06401__B2 genblk1\[1\].osc.clkdiv_C.cnt\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08967_ sig_norm.quo\[6\] _03654_ _00024_ vssd1 vssd1 vccd1 vccd1 _03655_ sky130_fd_sc_hd__mux2_1
X_07918_ _01489_ genblk1\[8\].osc.clkdiv_C.cnt\[6\] vssd1 vssd1 vccd1 vccd1 _02625_
+ sky130_fd_sc_hd__xor2_1
X_08898_ _03581_ _03601_ net26 vssd1 vssd1 vccd1 vccd1 _03603_ sky130_fd_sc_hd__a21o_1
X_07849_ _02461_ _02462_ genblk2\[1\].wave_shpr.div.fin_quo\[2\] vssd1 vssd1 vccd1
+ vccd1 _02556_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07901__B2 genblk1\[8\].osc.clkdiv_C.cnt\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10860_ genblk2\[6\].wave_shpr.div.b1\[11\] genblk2\[6\].wave_shpr.div.acc\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05004_ sky130_fd_sc_hd__and2b_1
XANTENNA_fanout40_A net44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09519_ _04042_ vssd1 vssd1 vccd1 vccd1 _04048_ sky130_fd_sc_hd__clkbuf_4
XPHY_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10791_ net566 _04918_ _04922_ _04945_ vssd1 vssd1 vccd1 vccd1 _00590_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12530_ clknet_leaf_61_clk _00082_ net188 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.b1\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_94_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_137_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12461_ clknet_leaf_104_clk _00034_ net155 vssd1 vssd1 vccd1 vccd1 PWM.final_sample_in\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_124_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11412_ genblk2\[8\].wave_shpr.div.b1\[7\] genblk2\[8\].wave_shpr.div.acc\[7\] vssd1
+ vssd1 vccd1 vccd1 _05388_ sky130_fd_sc_hd__and2b_1
X_12392_ _05963_ _05931_ vssd1 vssd1 vccd1 vccd1 _06066_ sky130_fd_sc_hd__or2b_1
XFILLER_0_50_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11343_ _05216_ _05273_ genblk2\[7\].wave_shpr.div.acc\[18\] vssd1 vssd1 vccd1 vccd1
+ _05332_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_105_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06162__A net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11274_ _05245_ vssd1 vssd1 vccd1 vccd1 _05279_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_39_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13013_ clknet_leaf_133_clk _00342_ net60 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.acc\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10225_ net710 _04518_ _04522_ _04546_ vssd1 vssd1 vccd1 vccd1 _00423_ sky130_fd_sc_hd__a22o_1
X_10156_ genblk2\[3\].wave_shpr.div.acc\[4\] _04494_ _04420_ vssd1 vssd1 vccd1 vccd1
+ _04495_ sky130_fd_sc_hd__mux2_1
XFILLER_0_146_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11508__A _05444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold5 genblk2\[10\].wave_shpr.div.quo\[11\] vssd1 vssd1 vccd1 vccd1 net223 sky130_fd_sc_hd__dlygate4sd3_1
X_10087_ _04455_ vssd1 vssd1 vccd1 vccd1 _04456_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__10412__A _04672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08145__A1 _01201_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_69_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10989_ genblk2\[6\].wave_shpr.div.acc\[0\] _00016_ _05079_ net283 _05080_ vssd1
+ vssd1 vccd1 vccd1 _00653_ sky130_fd_sc_hd__o221a_1
XFILLER_0_57_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12728_ clknet_leaf_38_clk genblk1\[10\].osc.clkdiv_C.next_cnt\[5\] net113 vssd1
+ vssd1 vccd1 vccd1 genblk1\[10\].osc.clkdiv_C.cnt\[5\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12659_ clknet_leaf_27_clk genblk1\[6\].osc.clkdiv_C.next_cnt\[8\] net90 vssd1 vssd1
+ vccd1 vccd1 genblk1\[6\].osc.clkdiv_C.cnt\[8\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_155_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06180_ sig_norm.i\[1\] sig_norm.i\[0\] sig_norm.i\[3\] _01151_ vssd1 vssd1 vccd1
+ vccd1 _01152_ sky130_fd_sc_hd__and4_1
XFILLER_0_25_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_25_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_20_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11755__A2 _03696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold405 genblk2\[6\].wave_shpr.div.quo\[11\] vssd1 vssd1 vccd1 vccd1 net623 sky130_fd_sc_hd__dlygate4sd3_1
Xhold416 genblk2\[3\].wave_shpr.div.quo\[14\] vssd1 vssd1 vccd1 vccd1 net634 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold427 genblk2\[1\].wave_shpr.div.quo\[11\] vssd1 vssd1 vccd1 vccd1 net645 sky130_fd_sc_hd__dlygate4sd3_1
Xhold438 genblk2\[2\].wave_shpr.div.quo\[20\] vssd1 vssd1 vccd1 vccd1 net656 sky130_fd_sc_hd__dlygate4sd3_1
Xhold449 genblk2\[4\].wave_shpr.div.b1\[16\] vssd1 vssd1 vccd1 vccd1 net667 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_110_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09870_ net919 _04282_ _04289_ _04292_ vssd1 vssd1 vccd1 vccd1 _00322_ sky130_fd_sc_hd__a22o_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08821_ _03473_ _03527_ vssd1 vssd1 vccd1 vccd1 _03528_ sky130_fd_sc_hd__or2_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1105 genblk2\[10\].wave_shpr.div.quo\[3\] vssd1 vssd1 vccd1 vccd1 net1323 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06395__B1 _01337_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1116 genblk2\[0\].wave_shpr.div.quo\[4\] vssd1 vssd1 vccd1 vccd1 net1334 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1127 genblk2\[5\].wave_shpr.div.acc\[20\] vssd1 vssd1 vccd1 vccd1 net1345 sky130_fd_sc_hd__dlygate4sd3_1
X_08752_ _02950_ _03458_ _02647_ vssd1 vssd1 vccd1 vccd1 _03459_ sky130_fd_sc_hd__a21oi_1
X_07703_ genblk2\[10\].wave_shpr.div.fin_quo\[4\] _02409_ vssd1 vssd1 vccd1 vccd1
+ _02410_ sky130_fd_sc_hd__nor2_1
X_08683_ _03388_ _03389_ genblk2\[2\].wave_shpr.div.fin_quo\[3\] _02468_ vssd1 vssd1
+ vccd1 vccd1 _03390_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_45_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_17_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07634_ genblk1\[11\].osc.clkdiv_C.cnt\[9\] _01190_ _02339_ _02340_ vssd1 vssd1 vccd1
+ vccd1 _02341_ sky130_fd_sc_hd__a211o_1
XTAP_1909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07565_ genblk1\[9\].osc.clkdiv_C.cnt\[12\] _01328_ _01799_ genblk1\[9\].osc.clkdiv_C.cnt\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02272_ sky130_fd_sc_hd__a22oi_1
X_09304_ _03779_ _03755_ vssd1 vssd1 vccd1 vccd1 _03891_ sky130_fd_sc_hd__or2b_1
X_06516_ _01200_ _01441_ vssd1 vssd1 vccd1 vccd1 _01442_ sky130_fd_sc_hd__nand2_4
XFILLER_0_152_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07496_ _02215_ net760 _02217_ vssd1 vssd1 vccd1 vccd1 _02218_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_76_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06247__A _01208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_810 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09235_ _03835_ vssd1 vssd1 vccd1 vccd1 _03845_ sky130_fd_sc_hd__clkbuf_4
X_06447_ genblk1\[1\].osc.clkdiv_C.cnt\[4\] _01380_ genblk1\[1\].osc.clkdiv_C.cnt\[5\]
+ vssd1 vssd1 vccd1 vccd1 _01386_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_91_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_106_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_859 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_16_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09166_ _03809_ vssd1 vssd1 vccd1 vccd1 _00101_ sky130_fd_sc_hd__clkbuf_1
X_06378_ net37 _01321_ vssd1 vssd1 vccd1 vccd1 _01322_ sky130_fd_sc_hd__and2_1
XFILLER_0_16_375 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11746__A2 _05623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08117_ genblk1\[4\].osc.clkdiv_C.cnt\[2\] _01326_ vssd1 vssd1 vccd1 vccd1 _02824_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_32_846 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09097_ _03745_ vssd1 vssd1 vccd1 vccd1 _00096_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_142_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08181__B _02885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07078__A genblk1\[8\].osc.clkdiv_C.cnt\[3\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08048_ _02752_ _02754_ vssd1 vssd1 vccd1 vccd1 _02755_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold950 PWM.final_in\[5\] vssd1 vssd1 vccd1 vccd1 net1168 sky130_fd_sc_hd__dlygate4sd3_1
Xhold961 smpl_rt_clkdiv.clkDiv_inst.cnt\[6\] vssd1 vssd1 vccd1 vccd1 net1179 sky130_fd_sc_hd__dlygate4sd3_1
Xhold972 genblk2\[3\].wave_shpr.div.b1\[17\] vssd1 vssd1 vccd1 vccd1 net1190 sky130_fd_sc_hd__dlygate4sd3_1
Xhold983 genblk2\[7\].wave_shpr.div.b1\[8\] vssd1 vssd1 vccd1 vccd1 net1201 sky130_fd_sc_hd__dlygate4sd3_1
Xhold994 genblk2\[5\].wave_shpr.div.b1\[3\] vssd1 vssd1 vccd1 vccd1 net1212 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10010_ _04365_ _04404_ _04405_ vssd1 vssd1 vccd1 vccd1 _04406_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout88_A net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07499__B_N net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09999_ genblk2\[3\].wave_shpr.div.b1\[8\] genblk2\[3\].wave_shpr.div.acc\[8\] vssd1
+ vssd1 vccd1 vccd1 _04395_ sky130_fd_sc_hd__and2b_1
X_11961_ genblk2\[10\].wave_shpr.div.acc\[20\] genblk2\[10\].wave_shpr.div.acc\[19\]
+ _05782_ vssd1 vssd1 vccd1 vccd1 _05783_ sky130_fd_sc_hd__or3_1
X_13700_ clknet_leaf_97_clk _01011_ net166 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.fin_quo\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10912_ _05040_ vssd1 vssd1 vccd1 vccd1 _00616_ sky130_fd_sc_hd__clkbuf_1
X_11892_ net1045 _03696_ _03694_ _05720_ vssd1 vssd1 vccd1 vccd1 _00916_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13631_ clknet_leaf_66_clk _00944_ net197 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.b1\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10843_ _04981_ genblk2\[6\].wave_shpr.div.acc\[2\] _04986_ vssd1 vssd1 vccd1 vccd1
+ _04987_ sky130_fd_sc_hd__a21o_1
XANTENNA__09088__C1 _03738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_119 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_456 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13562_ clknet_leaf_85_clk _00877_ net184 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.quo\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10774_ _04932_ _04811_ vssd1 vssd1 vccd1 vccd1 _04933_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_66_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12513_ clknet_leaf_84_clk _00075_ net202 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.i\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13493_ clknet_leaf_86_clk net238 net177 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.quo\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_151_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12444_ _06102_ _06103_ vssd1 vssd1 vccd1 vccd1 _06104_ sky130_fd_sc_hd__nand2_1
XFILLER_0_152_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11510__B genblk1\[8\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12375_ _05955_ _05935_ vssd1 vssd1 vccd1 vccd1 _06053_ sky130_fd_sc_hd__or2b_1
XFILLER_0_23_868 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10407__A _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10945__B1 _05056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06604__B _01192_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11326_ _05209_ _05167_ vssd1 vssd1 vccd1 vccd1 _05319_ sky130_fd_sc_hd__or2b_1
XFILLER_0_10_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11257_ net487 _05245_ _05249_ net542 _05268_ vssd1 vssd1 vccd1 vccd1 _00733_ sky130_fd_sc_hd__a221o_1
X_10208_ net948 _04518_ _04522_ _04534_ vssd1 vssd1 vccd1 vccd1 _00418_ sky130_fd_sc_hd__a22o_1
XANTENNA__09563__B1 _04048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11188_ genblk2\[8\].wave_shpr.div.b1\[6\] _01507_ _05042_ vssd1 vssd1 vccd1 vccd1
+ _05234_ sky130_fd_sc_hd__mux2_1
X_10139_ genblk2\[3\].wave_shpr.div.b1\[0\] _04420_ genblk2\[3\].wave_shpr.div.acc\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04482_ sky130_fd_sc_hd__a21o_1
XFILLER_0_89_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_57_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10228__A2 _04457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07170__B genblk1\[9\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07350_ _02108_ vssd1 vssd1 vccd1 vccd1 _02109_ sky130_fd_sc_hd__inv_2
X_06301_ _01238_ _01262_ vssd1 vssd1 vccd1 vccd1 _01263_ sky130_fd_sc_hd__or2_4
XFILLER_0_128_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07281_ genblk1\[10\].osc.clkdiv_C.cnt\[11\] genblk1\[10\].osc.clkdiv_C.cnt\[10\]
+ _02048_ vssd1 vssd1 vccd1 vccd1 _02052_ sky130_fd_sc_hd__and3_1
XFILLER_0_122_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_155_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09020_ _02152_ genblk2\[9\].wave_shpr.div.busy _02201_ vssd1 vssd1 vccd1 vccd1 _03692_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_115_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06232_ freq_div.state\[0\] vssd1 vssd1 vccd1 vccd1 _01194_ sky130_fd_sc_hd__buf_2
XFILLER_0_127_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_142_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06163_ _01130_ _01132_ vssd1 vssd1 vccd1 vccd1 _01135_ sky130_fd_sc_hd__nand2_1
XFILLER_0_142_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12008__S _05802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold202 genblk2\[11\].wave_shpr.div.b1\[8\] vssd1 vssd1 vccd1 vccd1 net420 sky130_fd_sc_hd__dlygate4sd3_1
Xhold213 _01034_ vssd1 vssd1 vccd1 vccd1 net431 sky130_fd_sc_hd__dlygate4sd3_1
Xhold224 _00302_ vssd1 vssd1 vccd1 vccd1 net442 sky130_fd_sc_hd__dlygate4sd3_1
Xhold235 genblk2\[5\].wave_shpr.div.quo\[12\] vssd1 vssd1 vccd1 vccd1 net453 sky130_fd_sc_hd__dlygate4sd3_1
Xhold246 genblk2\[4\].wave_shpr.div.quo\[1\] vssd1 vssd1 vccd1 vccd1 net464 sky130_fd_sc_hd__dlygate4sd3_1
Xhold257 _00972_ vssd1 vssd1 vccd1 vccd1 net475 sky130_fd_sc_hd__dlygate4sd3_1
Xhold268 genblk2\[6\].wave_shpr.div.quo\[18\] vssd1 vssd1 vccd1 vccd1 net486 sky130_fd_sc_hd__dlygate4sd3_1
Xhold279 sig_norm.b1\[1\] vssd1 vssd1 vccd1 vccd1 net497 sky130_fd_sc_hd__dlygate4sd3_1
X_09922_ _04207_ _04156_ vssd1 vssd1 vccd1 vccd1 _04332_ sky130_fd_sc_hd__or2b_1
X_09853_ genblk2\[2\].wave_shpr.div.acc\[1\] _04213_ vssd1 vssd1 vccd1 vccd1 _04279_
+ sky130_fd_sc_hd__or2_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08804_ _03442_ _03443_ _03217_ _03510_ vssd1 vssd1 vccd1 vccd1 _03511_ sky130_fd_sc_hd__a211oi_2
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09784_ _01490_ _01233_ vssd1 vssd1 vccd1 vccd1 _04242_ sky130_fd_sc_hd__nor2_4
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06996_ _01823_ _01827_ _01828_ vssd1 vssd1 vccd1 vccd1 genblk1\[7\].osc.clkdiv_C.next_cnt\[3\]
+ sky130_fd_sc_hd__nor3_1
XANTENNA__07580__A2 _01221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08735_ _03405_ _03406_ _03202_ _03440_ vssd1 vssd1 vccd1 vccd1 _03442_ sky130_fd_sc_hd__a211o_1
XANTENNA__09841__A _04269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10987__A _05054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08666_ genblk2\[4\].wave_shpr.div.fin_quo\[2\] _02932_ _02839_ _02316_ vssd1 vssd1
+ vccd1 vccd1 _03373_ sky130_fd_sc_hd__a31o_1
XFILLER_0_68_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07617_ genblk1\[11\].osc.clkdiv_C.cnt\[3\] _01513_ _02064_ genblk1\[11\].osc.clkdiv_C.cnt\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02324_ sky130_fd_sc_hd__a22o_1
X_08597_ _03302_ _03303_ vssd1 vssd1 vccd1 vccd1 _03304_ sky130_fd_sc_hd__nor2_1
XTAP_1739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_95_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07548_ net1169 vssd1 vssd1 vccd1 vccd1 _00035_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07479_ genblk2\[10\].wave_shpr.div.i\[2\] genblk2\[10\].wave_shpr.div.i\[3\] genblk2\[10\].wave_shpr.div.i\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02205_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_146_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09218_ net804 _03836_ _03804_ _03839_ vssd1 vssd1 vccd1 vccd1 _00123_ sky130_fd_sc_hd__a22o_1
XFILLER_0_134_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10490_ _04732_ _04613_ vssd1 vssd1 vccd1 vccd1 _04733_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06705__A _01489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_106_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09149_ _03734_ genblk2\[0\].wave_shpr.div.acc\[17\] vssd1 vssd1 vccd1 vccd1 _03797_
+ sky130_fd_sc_hd__and2_1
XANTENNA__06424__B _01367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12160_ net1257 _05818_ _05883_ _05907_ vssd1 vssd1 vccd1 vccd1 _00997_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11111_ genblk2\[7\].wave_shpr.div.acc\[10\] genblk2\[7\].wave_shpr.div.b1\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05171_ sky130_fd_sc_hd__or2b_1
X_12091_ genblk2\[10\].wave_shpr.div.acc\[4\] _05855_ _05787_ vssd1 vssd1 vccd1 vccd1
+ _05856_ sky130_fd_sc_hd__mux2_1
Xhold780 genblk2\[4\].wave_shpr.div.acc\[6\] vssd1 vssd1 vccd1 vccd1 net998 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_6_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold791 genblk2\[7\].wave_shpr.div.acc\[8\] vssd1 vssd1 vccd1 vccd1 net1009 sky130_fd_sc_hd__dlygate4sd3_1
X_11042_ _05005_ _05120_ vssd1 vssd1 vccd1 vccd1 _05121_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09751__A _01211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12993_ clknet_leaf_131_clk _00322_ net64 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.acc\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_11944_ genblk2\[10\].wave_shpr.div.b1\[10\] genblk2\[10\].wave_shpr.div.acc\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05766_ sky130_fd_sc_hd__and2b_1
XFILLER_0_86_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11875_ net935 _05684_ _05685_ _05708_ vssd1 vssd1 vccd1 vccd1 _00911_ sky130_fd_sc_hd__a22o_1
XFILLER_0_28_916 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10826_ genblk2\[6\].wave_shpr.div.acc\[13\] genblk2\[6\].wave_shpr.div.b1\[13\]
+ vssd1 vssd1 vccd1 vccd1 _04970_ sky130_fd_sc_hd__or2b_1
X_13614_ clknet_leaf_94_clk _00927_ net159 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.fin_quo\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_95_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10757_ _04803_ _04919_ vssd1 vssd1 vccd1 vccd1 _04920_ sky130_fd_sc_hd__xnor2_1
X_13545_ clknet_leaf_101_clk _00860_ net165 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.fin_quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_133_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_133_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_55_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10091__B1 _04456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13476_ clknet_leaf_72_clk _00793_ net216 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.b1\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10688_ genblk2\[5\].wave_shpr.div.quo\[18\] _04861_ _04862_ net235 _04871_ vssd1
+ vssd1 vccd1 vccd1 _00561_ sky130_fd_sc_hd__a221o_1
XFILLER_0_124_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12427_ genblk2\[11\].wave_shpr.div.acc\[19\] _06089_ _06092_ vssd1 vssd1 vccd1 vccd1
+ _06093_ sky130_fd_sc_hd__a21o_1
XFILLER_0_152_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12358_ _03941_ vssd1 vssd1 vccd1 vccd1 _06040_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_10_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11309_ _05200_ _05305_ vssd1 vssd1 vccd1 vccd1 _05306_ sky130_fd_sc_hd__xnor2_1
X_12289_ _06006_ vssd1 vssd1 vccd1 vccd1 _01027_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07446__A _02147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06850_ genblk1\[5\].osc.clkdiv_C.cnt\[10\] _01710_ vssd1 vssd1 vccd1 vccd1 _01712_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_93_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06781_ _01599_ _01653_ _01654_ vssd1 vssd1 vccd1 vccd1 _01655_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08520_ _03141_ _03226_ net3 _02364_ vssd1 vssd1 vccd1 vccd1 _03227_ sky130_fd_sc_hd__o211ai_2
XANTENNA__07314__A2 _02077_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08451_ _02636_ _03157_ _02604_ vssd1 vssd1 vccd1 vccd1 _03158_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_77_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_77_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07402_ genblk2\[0\].wave_shpr.div.i\[2\] genblk2\[0\].wave_shpr.div.i\[3\] genblk2\[0\].wave_shpr.div.i\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02148_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_9_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08382_ genblk1\[2\].osc.clkdiv_C.cnt\[2\] _02336_ _01418_ genblk1\[2\].osc.clkdiv_C.cnt\[3\]
+ vssd1 vssd1 vccd1 vccd1 _03089_ sky130_fd_sc_hd__o22a_1
XFILLER_0_85_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09600__S _04095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_521 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07333_ _02092_ _02094_ _02095_ vssd1 vssd1 vccd1 vccd1 _02096_ sky130_fd_sc_hd__and3_1
XFILLER_0_116_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_124_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_124_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA_fanout138_A net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07264_ _02027_ _02039_ _02040_ vssd1 vssd1 vccd1 vccd1 genblk1\[10\].osc.clkdiv_C.next_cnt\[5\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_45_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09003_ _03681_ vssd1 vssd1 vccd1 vccd1 _00066_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06215_ _01175_ _01176_ vssd1 vssd1 vccd1 vccd1 _01177_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_115_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07195_ _01953_ _01981_ vssd1 vssd1 vccd1 vccd1 _01982_ sky130_fd_sc_hd__nor2_1
XFILLER_0_103_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_14_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06146_ net11 _01105_ _01104_ vssd1 vssd1 vccd1 vccd1 _01118_ sky130_fd_sc_hd__a21bo_1
XANTENNA__09836__A _04268_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__13236__RESET_B net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09905_ _04199_ _04160_ vssd1 vssd1 vccd1 vccd1 _04319_ sky130_fd_sc_hd__or2b_1
XFILLER_0_6_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09836_ _04268_ vssd1 vssd1 vccd1 vccd1 _04269_ sky130_fd_sc_hd__buf_2
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09767_ _03704_ net1099 _04233_ vssd1 vssd1 vccd1 vccd1 _00278_ sky130_fd_sc_hd__a21o_1
X_06979_ genblk1\[7\].osc.clkdiv_C.cnt\[15\] _01363_ _01196_ _01813_ _01814_ vssd1
+ vssd1 vccd1 vccd1 _01815_ sky130_fd_sc_hd__o221a_1
XFILLER_0_69_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08718_ _03383_ _03395_ _03420_ _03421_ vssd1 vssd1 vccd1 vccd1 _03425_ sky130_fd_sc_hd__a211oi_2
XTAP_2215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09698_ _04171_ genblk2\[2\].wave_shpr.div.acc\[2\] _04177_ vssd1 vssd1 vccd1 vccd1
+ _04178_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08649_ _03353_ _03355_ vssd1 vssd1 vccd1 vccd1 _03356_ sky130_fd_sc_hd__xnor2_1
XTAP_1514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_2259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11660_ net319 _05552_ _03855_ vssd1 vssd1 vccd1 vccd1 _05553_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_138_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10611_ _04830_ vssd1 vssd1 vccd1 vccd1 _00525_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_leaf_115_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_115_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_9_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11591_ _05394_ _05365_ vssd1 vssd1 vccd1 vccd1 _05504_ sky130_fd_sc_hd__or2b_1
XFILLER_0_36_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13330_ clknet_leaf_24_clk net386 net91 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.quo\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10542_ genblk2\[5\].wave_shpr.div.acc\[10\] genblk2\[5\].wave_shpr.div.b1\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04770_ sky130_fd_sc_hd__or2b_1
XFILLER_0_52_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13261_ clknet_leaf_0_clk _00584_ net38 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.acc\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10473_ _04605_ _04719_ vssd1 vssd1 vccd1 vccd1 _04720_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_121_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12212_ _05938_ _05948_ _05949_ vssd1 vssd1 vccd1 vccd1 _05950_ sky130_fd_sc_hd__a21o_1
X_13192_ clknet_leaf_122_clk _00515_ net79 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.i\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09230__A2 _03841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12143_ net859 _05876_ _05883_ _05895_ vssd1 vssd1 vccd1 vccd1 _00992_ sky130_fd_sc_hd__a22o_1
XFILLER_0_103_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12117__A2 _05844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09518__B1 _04047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07792__A2 _01439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12074_ genblk2\[10\].wave_shpr.div.b1\[0\] genblk2\[10\].wave_shpr.div.acc\[0\]
+ _05787_ _05840_ vssd1 vssd1 vccd1 vccd1 _05843_ sky130_fd_sc_hd__a31o_1
X_11025_ _04997_ _05107_ vssd1 vssd1 vccd1 vccd1 _05108_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07633__A2_N _01262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11516__A _05441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10420__A _03719_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12976_ clknet_leaf_123_clk net458 net71 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.quo\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11927_ _05746_ _05747_ _05748_ vssd1 vssd1 vccd1 vccd1 _05749_ sky130_fd_sc_hd__a21o_1
XTAP_2760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11858_ _05601_ _05695_ vssd1 vssd1 vccd1 vccd1 _05696_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_145_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_106_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_106_clk
+ sky130_fd_sc_hd__clkbuf_16
X_10809_ genblk2\[5\].wave_shpr.div.i\[1\] genblk2\[5\].wave_shpr.div.i\[0\] vssd1
+ vssd1 vccd1 vccd1 _04957_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11789_ _05631_ genblk1\[9\].osc.clkdiv_C.cnt\[16\] vssd1 vssd1 vccd1 vccd1 _05644_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_55_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_12_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13528_ clknet_leaf_98_clk _00845_ net169 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.acc\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_113_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13459_ clknet_leaf_99_clk _00776_ net166 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.fin_quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12356__A2 _06009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_71_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09221__A2 _03836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11564__B1 _05446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08980__A1 _01157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07951_ genblk1\[7\].osc.clkdiv_C.cnt\[1\] _01556_ _01564_ _01732_ genblk1\[7\].osc.clkdiv_C.cnt\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02658_ sky130_fd_sc_hd__a32o_1
XFILLER_0_10_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06902_ _01741_ _01744_ _01746_ _01755_ vssd1 vssd1 vccd1 vccd1 _01756_ sky130_fd_sc_hd__or4_1
XFILLER_0_128_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07882_ _02547_ _02586_ _02520_ _02587_ _02588_ vssd1 vssd1 vccd1 vccd1 _02589_ sky130_fd_sc_hd__a2111oi_1
XANTENNA_clkbuf_leaf_86_clk_A clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09621_ _03997_ _04117_ vssd1 vssd1 vccd1 vccd1 _04118_ sky130_fd_sc_hd__xnor2_1
X_06833_ _01693_ _01700_ _01701_ vssd1 vssd1 vccd1 vccd1 genblk1\[5\].osc.clkdiv_C.next_cnt\[3\]
+ sky130_fd_sc_hd__nor3_1
XANTENNA__07904__A genblk1\[8\].osc.clkdiv_C.cnt\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09552_ _04055_ genblk1\[1\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 _04067_
+ sky130_fd_sc_hd__and2_1
X_06764_ _01641_ vssd1 vssd1 vccd1 vccd1 _01642_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08503_ _03196_ _03199_ _03209_ vssd1 vssd1 vccd1 vccd1 _03210_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12292__A1 _01327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09483_ _04030_ vssd1 vssd1 vccd1 vccd1 _00197_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06695_ genblk1\[4\].osc.clkdiv_C.cnt\[10\] _01323_ vssd1 vssd1 vccd1 vccd1 _01585_
+ sky130_fd_sc_hd__nor2_1
X_08434_ _02349_ _02351_ _02221_ vssd1 vssd1 vccd1 vccd1 _03141_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_148_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_148_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08365_ _03042_ _03047_ _03041_ vssd1 vssd1 vccd1 vccd1 _03072_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_117_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_135_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_24_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07316_ genblk1\[11\].osc.clkdiv_C.cnt\[15\] vssd1 vssd1 vccd1 vccd1 _02080_ sky130_fd_sc_hd__inv_2
X_08296_ _02970_ _03002_ vssd1 vssd1 vccd1 vccd1 _03003_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_6_640 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06274__A2 _01227_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07247_ _02026_ vssd1 vssd1 vccd1 vccd1 _02028_ sky130_fd_sc_hd__inv_2
XFILLER_0_143_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xclkbuf_4_2_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_2_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_5_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12347__A2 _05982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_39_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07178_ _01954_ _01969_ _01970_ vssd1 vssd1 vccd1 vccd1 _01971_ sky130_fd_sc_hd__and3_1
XANTENNA__10358__A1 _03704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_478 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06129_ net13 net15 vssd1 vssd1 vccd1 vccd1 _01101_ sky130_fd_sc_hd__nand2_1
XANTENNA__07223__A1 _01174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06702__B _01591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07086__A genblk1\[8\].osc.clkdiv_C.cnt\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11307__B1 _05283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_876 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout70_A net75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07814__A _02308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09819_ _04069_ genblk1\[2\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 _04260_
+ sky130_fd_sc_hd__and2_1
X_12830_ clknet_leaf_62_clk _00163_ net189 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.acc\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2001 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2012 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2023 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2034 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2045 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12761_ clknet_leaf_20_clk _00094_ net108 vssd1 vssd1 vccd1 vccd1 freq_div.state\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_2056 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12283__A1 _01946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2067 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2078 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2089 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11712_ _05439_ genblk2\[9\].wave_shpr.div.acc\[16\] vssd1 vssd1 vccd1 vccd1 _05604_
+ sky130_fd_sc_hd__and2_1
XTAP_1355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12692_ clknet_leaf_53_clk genblk1\[8\].osc.clkdiv_C.next_cnt\[5\] net172 vssd1 vssd1
+ vccd1 vccd1 genblk1\[8\].osc.clkdiv_C.cnt\[5\] sky130_fd_sc_hd__dfrtp_4
XTAP_1366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_127_718 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11643_ _05540_ _05413_ genblk2\[8\].wave_shpr.div.acc\[24\] vssd1 vssd1 vccd1 vccd1
+ _05542_ sky130_fd_sc_hd__mux2_1
XFILLER_0_127_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_80_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11574_ _05386_ _05369_ vssd1 vssd1 vccd1 vccd1 _05491_ sky130_fd_sc_hd__or2b_1
XFILLER_0_25_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13313_ clknet_leaf_121_clk net242 net78 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10525_ _04655_ _04755_ _04756_ _04657_ net1108 vssd1 vssd1 vccd1 vccd1 _00513_ sky130_fd_sc_hd__a32o_1
XFILLER_0_80_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13244_ clknet_leaf_9_clk _00567_ net54 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.quo\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10456_ _04597_ _04706_ vssd1 vssd1 vccd1 vccd1 _04707_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10349__A1 _01757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11546__B1 _05444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13175_ clknet_leaf_129_clk _00500_ net67 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.acc\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07708__B _02403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10387_ _04651_ vssd1 vssd1 vccd1 vccd1 _04661_ sky130_fd_sc_hd__buf_2
XANTENNA__10415__A _04676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06612__B _01519_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11204__A2_N _01490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12126_ net858 _05876_ _05850_ _05882_ vssd1 vssd1 vccd1 vccd1 _00988_ sky130_fd_sc_hd__a22o_1
XANTENNA__07765__A2 _01309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06973__B1 _01311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12057_ _05819_ genblk1\[10\].osc.clkdiv_C.cnt\[11\] vssd1 vssd1 vccd1 vccd1 _05833_
+ sky130_fd_sc_hd__and2_1
X_11008_ _05094_ _04989_ vssd1 vssd1 vccd1 vccd1 _05095_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10521__A1 _04651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10150__A _04455_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_87_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12959_ clknet_leaf_136_clk _00288_ net42 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.b1\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_142_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06480_ net29 _01407_ vssd1 vssd1 vccd1 vccd1 _01408_ sky130_fd_sc_hd__nor2_1
XTAP_2590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08150_ genblk1\[3\].osc.clkdiv_C.cnt\[3\] _01234_ _02854_ _02855_ _02856_ vssd1
+ vssd1 vccd1 vccd1 _02857_ sky130_fd_sc_hd__o221a_1
XFILLER_0_16_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09089__C _01197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07101_ genblk1\[8\].osc.clkdiv_C.cnt\[11\] _01904_ _01907_ vssd1 vssd1 vccd1 vccd1
+ genblk1\[8\].osc.clkdiv_C.next_cnt\[11\] sky130_fd_sc_hd__o21a_1
X_08081_ _02752_ _02753_ _02755_ _02786_ _02787_ vssd1 vssd1 vccd1 vccd1 _02788_ sky130_fd_sc_hd__o221a_1
XFILLER_0_113_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06256__A2 _01210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07032_ _01851_ vssd1 vssd1 vccd1 vccd1 genblk1\[7\].osc.clkdiv_C.next_cnt\[16\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_70_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_11_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_3_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_101_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_113_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07618__B _02064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_197 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08983_ sig_norm.quo\[8\] _01098_ _03667_ vssd1 vssd1 vccd1 vccd1 _03668_ sky130_fd_sc_hd__a21bo_1
X_07934_ genblk2\[8\].wave_shpr.div.fin_quo\[4\] _02640_ vssd1 vssd1 vccd1 vccd1 _02641_
+ sky130_fd_sc_hd__nor2_1
X_07865_ _02216_ _02552_ genblk2\[0\].wave_shpr.div.fin_quo\[0\] vssd1 vssd1 vccd1
+ vccd1 _02572_ sky130_fd_sc_hd__and3_1
XANTENNA__06796__A2_N _01666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09604_ genblk2\[1\].wave_shpr.div.acc\[10\] _04104_ _04095_ vssd1 vssd1 vccd1 vccd1
+ _04105_ sky130_fd_sc_hd__mux2_1
X_06816_ genblk1\[5\].osc.clkdiv_C.cnt\[12\] _01355_ vssd1 vssd1 vccd1 vccd1 _01688_
+ sky130_fd_sc_hd__or2_1
X_07796_ _02496_ _02497_ vssd1 vssd1 vccd1 vccd1 _02503_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwire30 _02635_ vssd1 vssd1 vccd1 vccd1 net30 sky130_fd_sc_hd__clkbuf_2
X_06747_ genblk1\[4\].osc.clkdiv_C.cnt\[7\] genblk1\[4\].osc.clkdiv_C.cnt\[6\] _01616_
+ genblk1\[4\].osc.clkdiv_C.cnt\[8\] vssd1 vssd1 vccd1 vccd1 _01629_ sky130_fd_sc_hd__a31o_1
X_09535_ _03719_ vssd1 vssd1 vccd1 vccd1 _04058_ sky130_fd_sc_hd__buf_4
XANTENNA__12265__A1 _01240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10995__A _05023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09466_ net1247 _01327_ _03822_ vssd1 vssd1 vccd1 vccd1 _04021_ sky130_fd_sc_hd__mux2_1
XFILLER_0_149_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06678_ genblk1\[4\].osc.clkdiv_C.cnt\[1\] vssd1 vssd1 vccd1 vccd1 _01568_ sky130_fd_sc_hd__inv_2
XANTENNA__06684__S _01188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08417_ _03085_ _03123_ vssd1 vssd1 vccd1 vccd1 _03124_ sky130_fd_sc_hd__xnor2_1
X_09397_ genblk2\[1\].wave_shpr.div.acc\[10\] genblk2\[1\].wave_shpr.div.b1\[10\]
+ vssd1 vssd1 vccd1 vccd1 _03961_ sky130_fd_sc_hd__or2b_1
XFILLER_0_108_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_863 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08184__B _02885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08348_ _03054_ vssd1 vssd1 vccd1 vccd1 _03055_ sky130_fd_sc_hd__inv_2
XFILLER_0_117_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08279_ genblk2\[9\].wave_shpr.div.fin_quo\[4\] _02303_ _02264_ _02223_ vssd1 vssd1
+ vccd1 vccd1 _02986_ sky130_fd_sc_hd__a31o_1
XFILLER_0_21_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10310_ genblk2\[4\].wave_shpr.div.acc\[25\] genblk2\[4\].wave_shpr.div.acc\[24\]
+ genblk2\[4\].wave_shpr.div.acc\[26\] _04621_ vssd1 vssd1 vccd1 vccd1 _04622_ sky130_fd_sc_hd__or4b_4
XFILLER_0_62_899 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07995__A2 _01484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11290_ net988 _05279_ _05283_ _05291_ vssd1 vssd1 vccd1 vccd1 _00743_ sky130_fd_sc_hd__a22o_1
X_10241_ genblk2\[3\].wave_shpr.div.i\[1\] genblk2\[3\].wave_shpr.div.i\[0\] vssd1
+ vssd1 vccd1 vccd1 _04557_ sky130_fd_sc_hd__or2_1
X_10172_ _04419_ vssd1 vssd1 vccd1 vccd1 _04507_ sky130_fd_sc_hd__buf_4
Xfanout150 net171 vssd1 vssd1 vccd1 vccd1 net150 sky130_fd_sc_hd__clkbuf_4
Xfanout161 net162 vssd1 vssd1 vccd1 vccd1 net161 sky130_fd_sc_hd__buf_2
Xfanout172 net173 vssd1 vssd1 vccd1 vccd1 net172 sky130_fd_sc_hd__clkbuf_4
Xfanout183 net185 vssd1 vssd1 vccd1 vccd1 net183 sky130_fd_sc_hd__clkbuf_4
Xfanout194 net195 vssd1 vssd1 vccd1 vccd1 net194 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08172__A2 _01498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06183__A1 _01099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12813_ clknet_leaf_58_clk _00146_ net192 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.quo\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10806__A2 _04858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_97_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12744_ clknet_leaf_49_clk genblk1\[11\].osc.clkdiv_C.next_cnt\[3\] net108 vssd1
+ vssd1 vccd1 vccd1 genblk1\[11\].osc.clkdiv_C.cnt\[3\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__07132__B1 _01349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12008__A1 _01483_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12675_ clknet_leaf_90_clk genblk1\[7\].osc.clkdiv_C.next_cnt\[6\] net141 vssd1 vssd1
+ vccd1 vccd1 genblk1\[7\].osc.clkdiv_C.cnt\[6\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_53_800 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_127_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11626_ net1114 _05507_ _05445_ _05530_ vssd1 vssd1 vccd1 vccd1 _00840_ sky130_fd_sc_hd__a22o_1
XFILLER_0_108_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11557_ _05378_ _05373_ vssd1 vssd1 vccd1 vccd1 _05478_ sky130_fd_sc_hd__or2b_1
XFILLER_0_108_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_69_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10508_ net472 _04744_ _04745_ vssd1 vssd1 vccd1 vccd1 _04746_ sky130_fd_sc_hd__a21o_1
Xhold609 genblk2\[1\].wave_shpr.div.acc\[8\] vssd1 vssd1 vccd1 vccd1 net827 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11488_ _03726_ _05439_ _03736_ vssd1 vssd1 vccd1 vccd1 _00793_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_100_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09188__A1 _03714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_0_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10439_ _04580_ _04590_ vssd1 vssd1 vccd1 vccd1 _04694_ sky130_fd_sc_hd__xor2_1
X_13227_ clknet_leaf_127_clk _00550_ net67 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10145__A _04451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_903 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_914 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13158_ clknet_leaf_121_clk _00483_ net78 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.quo\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_925 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12109_ net1035 _05844_ _05850_ _05869_ vssd1 vssd1 vccd1 vccd1 _00984_ sky130_fd_sc_hd__a22o_1
XTAP_958 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13089_ clknet_leaf_137_clk _00416_ net40 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.acc\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_969 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07454__A _02147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11298__A2 _05279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08163__A2 _01498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07650_ genblk2\[11\].wave_shpr.div.fin_quo\[6\] _02349_ _02351_ _02356_ vssd1 vssd1
+ vccd1 vccd1 _02357_ sky130_fd_sc_hd__and4_1
X_06601_ genblk1\[3\].osc.clkdiv_C.cnt\[12\] _01507_ _01508_ genblk1\[3\].osc.clkdiv_C.cnt\[11\]
+ vssd1 vssd1 vccd1 vccd1 _01509_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__07910__A2 _01564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07581_ _01186_ _01437_ _01226_ _01171_ genblk1\[9\].osc.clkdiv_C.cnt\[0\] vssd1
+ vssd1 vccd1 vccd1 _02288_ sky130_fd_sc_hd__o311a_1
X_09320_ _03835_ vssd1 vssd1 vccd1 vccd1 _03903_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_87_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06532_ _01452_ _01454_ _01455_ vssd1 vssd1 vccd1 vccd1 genblk1\[2\].osc.clkdiv_C.next_cnt\[2\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_88_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_146_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_118_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09251_ genblk2\[0\].wave_shpr.div.quo\[18\] _03845_ _03847_ net410 _03854_ vssd1
+ vssd1 vccd1 vccd1 _00141_ sky130_fd_sc_hd__a221o_1
X_06463_ genblk1\[1\].osc.clkdiv_C.cnt\[10\] _01394_ _01396_ _01374_ vssd1 vssd1 vccd1
+ vccd1 genblk1\[1\].osc.clkdiv_C.next_cnt\[10\] sky130_fd_sc_hd__o211a_1
XFILLER_0_7_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08202_ _02906_ _02907_ _02908_ _02416_ vssd1 vssd1 vccd1 vccd1 _02909_ sky130_fd_sc_hd__a211o_1
XFILLER_0_118_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_885 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_8_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09182_ net1273 _01214_ _03722_ vssd1 vssd1 vccd1 vccd1 _03818_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06394_ genblk1\[1\].osc.clkdiv_C.cnt\[15\] _01210_ _01337_ genblk1\[1\].osc.clkdiv_C.cnt\[12\]
+ vssd1 vssd1 vccd1 vccd1 _01338_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_43_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_7_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_145_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08133_ genblk2\[4\].wave_shpr.div.fin_quo\[2\] _02839_ vssd1 vssd1 vccd1 vccd1 _02840_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_55_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11222__A2 _05246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_721 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout218_A net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08064_ genblk1\[5\].osc.clkdiv_C.cnt\[3\] _01195_ _01254_ vssd1 vssd1 vccd1 vccd1
+ _02771_ sky130_fd_sc_hd__or3_1
XANTENNA__07629__A _01174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07015_ genblk1\[7\].osc.clkdiv_C.cnt\[10\] _01837_ genblk1\[7\].osc.clkdiv_C.cnt\[11\]
+ vssd1 vssd1 vccd1 vccd1 _01840_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06252__B _01188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07729__A2 net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_wire33_A _02348_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06401__A2 genblk1\[1\].osc.clkdiv_C.cnt\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08966_ sig_norm.quo\[5\] _03653_ _01155_ vssd1 vssd1 vccd1 vccd1 _03654_ sky130_fd_sc_hd__mux2_1
X_07917_ genblk1\[8\].osc.clkdiv_C.cnt\[5\] _01858_ _02621_ _02622_ _02623_ vssd1
+ vssd1 vccd1 vccd1 _02624_ sky130_fd_sc_hd__o221a_1
X_08897_ sig_norm.acc\[11\] sig_norm.acc\[12\] _03591_ _03594_ vssd1 vssd1 vccd1 vccd1
+ _03602_ sky130_fd_sc_hd__nor4_2
Xclkbuf_leaf_95_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_95_clk sky130_fd_sc_hd__clkbuf_16
X_07848_ _02509_ _02551_ _02554_ vssd1 vssd1 vccd1 vccd1 _02555_ sky130_fd_sc_hd__or3_1
XANTENNA__07901__A2 _01246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07779_ _01181_ genblk1\[0\].osc.clkdiv_C.cnt\[7\] _02485_ vssd1 vssd1 vccd1 vccd1
+ _02486_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_78_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39_627 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09518_ net460 _04043_ _04047_ genblk2\[1\].wave_shpr.div.quo\[7\] vssd1 vssd1 vccd1
+ vccd1 _00215_ sky130_fd_sc_hd__a22o_1
X_10790_ _04943_ _04944_ vssd1 vssd1 vccd1 vccd1 _04945_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09449_ _04012_ vssd1 vssd1 vccd1 vccd1 _00181_ sky130_fd_sc_hd__clkbuf_1
XPHY_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12460_ clknet_leaf_104_clk _00033_ net155 vssd1 vssd1 vccd1 vccd1 PWM.final_sample_in\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11749__B1 _05624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_136_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_46_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11411_ _05369_ _05385_ _05386_ vssd1 vssd1 vccd1 vccd1 _05387_ sky130_fd_sc_hd__a21o_1
XFILLER_0_152_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12391_ net785 _06039_ _06040_ _06065_ vssd1 vssd1 vccd1 vccd1 _01070_ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11342_ _05217_ _05273_ vssd1 vssd1 vccd1 vccd1 _05331_ sky130_fd_sc_hd__or2_1
XFILLER_0_132_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11273_ net1013 _05246_ _05250_ _05278_ vssd1 vssd1 vccd1 vccd1 _00739_ sky130_fd_sc_hd__a22o_1
X_10224_ _04416_ _04480_ _04543_ net524 vssd1 vssd1 vccd1 vccd1 _04546_ sky130_fd_sc_hd__a2bb2o_1
X_13012_ clknet_leaf_133_clk _00341_ net60 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.acc\[24\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__09754__A _01436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10155_ _04376_ _04387_ vssd1 vssd1 vccd1 vccd1 _04494_ sky130_fd_sc_hd__xor2_1
XFILLER_0_100_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold6 _00961_ vssd1 vssd1 vccd1 vccd1 net224 sky130_fd_sc_hd__dlygate4sd3_1
X_10086_ _04453_ vssd1 vssd1 vccd1 vccd1 _04455_ sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_86_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_86_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_57_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10988_ _03719_ genblk1\[6\].osc.clkdiv_C.cnt\[17\] vssd1 vssd1 vccd1 vccd1 _05080_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_146_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_84_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12727_ clknet_leaf_38_clk genblk1\[10\].osc.clkdiv_C.next_cnt\[4\] net113 vssd1
+ vssd1 vccd1 vccd1 genblk1\[10\].osc.clkdiv_C.cnt\[4\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_38_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_822 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10660__B1 _04857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12658_ clknet_leaf_27_clk genblk1\[6\].osc.clkdiv_C.next_cnt\[7\] net90 vssd1 vssd1
+ vccd1 vccd1 genblk1\[6\].osc.clkdiv_C.cnt\[7\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_154_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_115_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11609_ _05401_ _05517_ vssd1 vssd1 vccd1 vccd1 _05518_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_53_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12589_ clknet_leaf_14_clk genblk1\[2\].osc.clkdiv_C.next_cnt\[10\] net72 vssd1 vssd1
+ vccd1 vccd1 genblk1\[2\].osc.clkdiv_C.cnt\[10\] sky130_fd_sc_hd__dfrtp_2
Xclkbuf_leaf_10_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_10_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_111_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07959__A2 _01311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_105_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold406 _00639_ vssd1 vssd1 vccd1 vccd1 net624 sky130_fd_sc_hd__dlygate4sd3_1
Xhold417 _00389_ vssd1 vssd1 vccd1 vccd1 net635 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_20_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold428 genblk2\[9\].wave_shpr.div.acc\[22\] vssd1 vssd1 vccd1 vccd1 net646 sky130_fd_sc_hd__dlygate4sd3_1
Xhold439 genblk2\[3\].wave_shpr.div.acc\[18\] vssd1 vssd1 vccd1 vccd1 net657 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_110_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08820_ _03470_ _03472_ vssd1 vssd1 vccd1 vccd1 _03527_ sky130_fd_sc_hd__nor2_1
XFILLER_0_110_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06395__B2 genblk1\[1\].osc.clkdiv_C.cnt\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1106 genblk2\[10\].wave_shpr.div.quo\[5\] vssd1 vssd1 vccd1 vccd1 net1324 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1117 genblk2\[8\].wave_shpr.div.quo\[6\] vssd1 vssd1 vccd1 vccd1 net1335 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1128 genblk2\[3\].wave_shpr.div.quo\[5\] vssd1 vssd1 vccd1 vccd1 net1346 sky130_fd_sc_hd__dlygate4sd3_1
X_08751_ genblk2\[7\].wave_shpr.div.fin_quo\[0\] _02467_ vssd1 vssd1 vccd1 vccd1 _03458_
+ sky130_fd_sc_hd__nand2_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07615__C _01437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_77_clk clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_77_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_136_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07702_ _02406_ _02408_ vssd1 vssd1 vccd1 vccd1 _02409_ sky130_fd_sc_hd__nand2_1
X_08682_ genblk2\[2\].wave_shpr.div.fin_quo\[2\] _03113_ _03115_ _02224_ vssd1 vssd1
+ vccd1 vccd1 _03389_ sky130_fd_sc_hd__a31o_1
XFILLER_0_136_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07633_ genblk1\[11\].osc.clkdiv_C.cnt\[10\] _01262_ _01494_ _02128_ vssd1 vssd1
+ vccd1 vccd1 _02340_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA_fanout168_A net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07564_ _01930_ _01227_ _01732_ _02268_ _02270_ vssd1 vssd1 vccd1 vccd1 _02271_ sky130_fd_sc_hd__o221a_1
XANTENNA__07631__B _01179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09303_ net1049 _03870_ _03877_ _03890_ vssd1 vssd1 vccd1 vccd1 _00157_ sky130_fd_sc_hd__a22o_1
X_06515_ _01440_ vssd1 vssd1 vccd1 vccd1 _01441_ sky130_fd_sc_hd__buf_6
XFILLER_0_8_510 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07495_ _02216_ vssd1 vssd1 vccd1 vccd1 _02217_ sky130_fd_sc_hd__buf_2
XFILLER_0_119_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_660 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_61_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_822 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09839__A _04269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06446_ genblk1\[1\].osc.clkdiv_C.cnt\[5\] genblk1\[1\].osc.clkdiv_C.cnt\[4\] _01380_
+ vssd1 vssd1 vccd1 vccd1 _01385_ sky130_fd_sc_hd__and3_1
X_09234_ genblk2\[0\].wave_shpr.div.quo\[11\] _03841_ _03839_ net569 _03844_ vssd1
+ vssd1 vccd1 vccd1 _00134_ sky130_fd_sc_hd__a221o_1
XFILLER_0_91_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_63_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09165_ genblk2\[0\].wave_shpr.div.fin_quo\[4\] genblk2\[0\].wave_shpr.div.quo\[3\]
+ _00001_ vssd1 vssd1 vccd1 vccd1 _03809_ sky130_fd_sc_hd__mux2_1
XFILLER_0_17_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_90_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06377_ _01188_ _01191_ vssd1 vssd1 vccd1 vccd1 _01321_ sky130_fd_sc_hd__nand2b_4
XFILLER_0_133_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08116_ genblk1\[4\].osc.clkdiv_C.cnt\[1\] _01866_ genblk1\[4\].osc.clkdiv_C.cnt\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02823_ sky130_fd_sc_hd__o21a_1
XFILLER_0_44_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09096_ _03744_ _01490_ _03741_ vssd1 vssd1 vccd1 vccd1 _03745_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_32_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08047_ genblk1\[5\].osc.clkdiv_C.cnt\[12\] _01666_ _02753_ vssd1 vssd1 vccd1 vccd1
+ _02754_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold940 genblk2\[0\].wave_shpr.div.i\[3\] vssd1 vssd1 vccd1 vccd1 net1158 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold951 _02257_ vssd1 vssd1 vccd1 vccd1 net1169 sky130_fd_sc_hd__dlygate4sd3_1
Xhold962 genblk1\[6\].osc.clkdiv_C.cnt\[10\] vssd1 vssd1 vccd1 vccd1 net1180 sky130_fd_sc_hd__dlygate4sd3_1
Xhold973 genblk2\[8\].wave_shpr.div.b1\[17\] vssd1 vssd1 vccd1 vccd1 net1191 sky130_fd_sc_hd__dlygate4sd3_1
Xhold984 genblk2\[7\].wave_shpr.div.b1\[6\] vssd1 vssd1 vccd1 vccd1 net1202 sky130_fd_sc_hd__dlygate4sd3_1
Xhold995 genblk1\[2\].osc.clkdiv_C.cnt\[11\] vssd1 vssd1 vccd1 vccd1 net1213 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11903__B1 _03841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09998_ _04371_ _04392_ _04393_ vssd1 vssd1 vccd1 vccd1 _04394_ sky130_fd_sc_hd__a21o_1
X_08949_ _03638_ _03639_ sig_norm.quo\[2\] _01098_ vssd1 vssd1 vccd1 vccd1 _03640_
+ sky130_fd_sc_hd__a2bb2o_1
Xclkbuf_leaf_68_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_68_clk sky130_fd_sc_hd__clkbuf_16
X_11960_ genblk2\[10\].wave_shpr.div.acc\[18\] _05781_ vssd1 vssd1 vccd1 vccd1 _05782_
+ sky130_fd_sc_hd__or2_1
XANTENNA__08532__C1 _02364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07822__A net7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10911_ genblk2\[7\].wave_shpr.div.b1\[7\] _04444_ _04848_ vssd1 vssd1 vccd1 vccd1
+ _05040_ sky130_fd_sc_hd__mux2_1
XANTENNA__07886__B2 _02592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11891_ _05718_ _05715_ _05719_ vssd1 vssd1 vccd1 vccd1 _05720_ sky130_fd_sc_hd__o21ai_1
X_13630_ clknet_leaf_67_clk _00943_ net195 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.b1\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10842_ _04981_ genblk2\[6\].wave_shpr.div.acc\[2\] _04985_ vssd1 vssd1 vccd1 vccd1
+ _04986_ sky130_fd_sc_hd__o21a_1
XANTENNA__09088__B1 _01591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07638__A1 _01229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13561_ clknet_leaf_85_clk _00876_ net184 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.quo\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_632 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10773_ _04812_ _04764_ vssd1 vssd1 vccd1 vccd1 _04932_ sky130_fd_sc_hd__nor2_1
XFILLER_0_109_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12512_ clknet_leaf_84_clk _00074_ net202 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.i\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_82_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13492_ clknet_leaf_87_clk _00809_ net177 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.quo\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12443_ genblk2\[11\].wave_shpr.div.acc\[25\] _05980_ genblk2\[11\].wave_shpr.div.acc\[24\]
+ genblk2\[11\].wave_shpr.div.acc\[26\] vssd1 vssd1 vccd1 vccd1 _06103_ sky130_fd_sc_hd__or4b_1
XFILLER_0_35_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11198__A1 _05239_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12374_ net997 _06039_ _06040_ _06052_ vssd1 vssd1 vccd1 vccd1 _01066_ sky130_fd_sc_hd__a22o_1
XFILLER_0_151_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06604__C _01208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11325_ net805 _05311_ _05315_ _05318_ vssd1 vssd1 vccd1 vccd1 _00751_ sky130_fd_sc_hd__a22o_1
XANTENNA__06613__A2 _01256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_50_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_10_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11256_ _05260_ genblk1\[7\].osc.clkdiv_C.cnt\[13\] vssd1 vssd1 vccd1 vccd1 _05268_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_66_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09563__A1 _04045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10207_ genblk2\[3\].wave_shpr.div.acc\[16\] _04533_ _04507_ vssd1 vssd1 vccd1 vccd1
+ _04534_ sky130_fd_sc_hd__mux2_1
X_11187_ _05233_ vssd1 vssd1 vccd1 vccd1 _00698_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07574__B1 genblk1\[9\].osc.clkdiv_C.cnt\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10138_ _04480_ _04380_ genblk2\[3\].wave_shpr.div.b1\[0\] vssd1 vssd1 vccd1 vccd1
+ _04481_ sky130_fd_sc_hd__or3b_1
Xclkbuf_leaf_59_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_59_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__08118__A2 _01326_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10069_ net1205 _04444_ _04440_ vssd1 vssd1 vccd1 vccd1 _04445_ sky130_fd_sc_hd__mux2_1
XANTENNA__08828__A net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13759_ clknet_leaf_66_clk _01070_ net213 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.acc\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_06300_ _01261_ vssd1 vssd1 vccd1 vccd1 _01262_ sky130_fd_sc_hd__buf_4
XFILLER_0_127_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07280_ genblk1\[10\].osc.clkdiv_C.cnt\[10\] _02048_ genblk1\[10\].osc.clkdiv_C.cnt\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02051_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06231_ _01181_ _01192_ vssd1 vssd1 vccd1 vccd1 _01193_ sky130_fd_sc_hd__nand2_2
XFILLER_0_122_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06162_ net10 vssd1 vssd1 vccd1 vccd1 _01134_ sky130_fd_sc_hd__inv_2
XFILLER_0_53_482 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_131_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold203 genblk2\[7\].wave_shpr.div.quo\[7\] vssd1 vssd1 vccd1 vccd1 net421 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_142_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold214 genblk2\[10\].wave_shpr.div.quo\[9\] vssd1 vssd1 vccd1 vccd1 net432 sky130_fd_sc_hd__dlygate4sd3_1
Xhold225 genblk2\[11\].wave_shpr.div.quo\[12\] vssd1 vssd1 vccd1 vccd1 net443 sky130_fd_sc_hd__dlygate4sd3_1
Xhold236 genblk2\[0\].wave_shpr.div.quo\[23\] vssd1 vssd1 vccd1 vccd1 net454 sky130_fd_sc_hd__dlygate4sd3_1
Xhold247 _00461_ vssd1 vssd1 vccd1 vccd1 net465 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06518__A2_N _01442_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold258 genblk2\[0\].wave_shpr.div.quo\[22\] vssd1 vssd1 vccd1 vccd1 net476 sky130_fd_sc_hd__dlygate4sd3_1
X_09921_ net788 _04315_ _04322_ _04331_ vssd1 vssd1 vccd1 vccd1 _00334_ sky130_fd_sc_hd__a22o_1
Xhold269 genblk2\[7\].wave_shpr.div.quo\[22\] vssd1 vssd1 vccd1 vccd1 net487 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08357__A2 _02521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09852_ _04277_ _04278_ net782 _04248_ vssd1 vssd1 vccd1 vccd1 _00318_ sky130_fd_sc_hd__a2bb2o_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07565__B1 _01799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08803_ _03204_ _03205_ _03216_ vssd1 vssd1 vccd1 vccd1 _03510_ sky130_fd_sc_hd__o21ba_1
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09783_ _03732_ net1152 _04241_ vssd1 vssd1 vccd1 vccd1 _00286_ sky130_fd_sc_hd__o21a_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06995_ genblk1\[7\].osc.clkdiv_C.cnt\[3\] _01825_ vssd1 vssd1 vccd1 vccd1 _01828_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__08109__A2 _01323_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08734_ _03202_ _03440_ _03405_ _03406_ vssd1 vssd1 vccd1 vccd1 _03441_ sky130_fd_sc_hd__o211ai_2
XANTENNA__07642__A net33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08665_ _02932_ _02839_ genblk2\[4\].wave_shpr.div.fin_quo\[2\] vssd1 vssd1 vccd1
+ vccd1 _03372_ sky130_fd_sc_hd__a21oi_1
XANTENNA__10479__S _04704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07616_ _02318_ _02319_ _02320_ _02321_ _02322_ vssd1 vssd1 vccd1 vccd1 _02323_ sky130_fd_sc_hd__o311a_1
XFILLER_0_49_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08596_ _02798_ _03299_ _03301_ vssd1 vssd1 vccd1 vccd1 _03303_ sky130_fd_sc_hd__a21oi_1
X_07547_ PWM.final_sample_in\[5\] net1168 PWM.start vssd1 vssd1 vccd1 vccd1 _02257_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_48_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07478_ _02204_ vssd1 vssd1 vccd1 vccd1 _00023_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_64_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09217_ _03838_ vssd1 vssd1 vccd1 vccd1 _03839_ sky130_fd_sc_hd__clkbuf_4
X_06429_ _01372_ vssd1 vssd1 vccd1 vccd1 _01373_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_106_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06705__B _01196_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09148_ _03747_ _03794_ _03795_ vssd1 vssd1 vccd1 vccd1 _03796_ sky130_fd_sc_hd__a21o_1
XFILLER_0_115_860 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10927__A1 _01365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09079_ _03708_ _01210_ vssd1 vssd1 vccd1 vccd1 _03733_ sky130_fd_sc_hd__nand2_8
XFILLER_0_32_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_20_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11110_ genblk2\[7\].wave_shpr.div.acc\[11\] genblk2\[7\].wave_shpr.div.b1\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05170_ sky130_fd_sc_hd__or2b_1
X_12090_ _05854_ _05753_ vssd1 vssd1 vccd1 vccd1 _05855_ sky130_fd_sc_hd__xnor2_1
Xhold770 genblk2\[7\].wave_shpr.div.acc\[6\] vssd1 vssd1 vccd1 vccd1 net988 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold781 genblk2\[9\].wave_shpr.div.acc\[5\] vssd1 vssd1 vccd1 vccd1 net999 sky130_fd_sc_hd__dlygate4sd3_1
X_11041_ _05006_ _04971_ vssd1 vssd1 vccd1 vccd1 _05120_ sky130_fd_sc_hd__or2b_1
Xhold792 genblk2\[7\].wave_shpr.div.acc\[16\] vssd1 vssd1 vccd1 vccd1 net1010 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09751__B _01302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12992_ clknet_leaf_131_clk _00321_ net64 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.acc\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12301__B1 _06010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_hold929_A genblk2\[8\].wave_shpr.div.b1\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11943_ _05739_ _05763_ _05764_ vssd1 vssd1 vccd1 vccd1 _05765_ sky130_fd_sc_hd__a21o_1
X_11874_ genblk2\[9\].wave_shpr.div.acc\[19\] _05608_ _05707_ vssd1 vssd1 vccd1 vccd1
+ _05708_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_67_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13613_ clknet_leaf_94_clk _00926_ net159 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.fin_quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10825_ genblk2\[6\].wave_shpr.div.acc\[14\] genblk2\[6\].wave_shpr.div.b1\[14\]
+ vssd1 vssd1 vccd1 vccd1 _04969_ sky130_fd_sc_hd__or2b_1
XANTENNA__11802__A _03693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13544_ clknet_leaf_101_clk _00859_ net164 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.fin_quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10756_ _04804_ _04768_ vssd1 vssd1 vccd1 vccd1 _04919_ sky130_fd_sc_hd__or2b_1
XFILLER_0_82_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_54_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11521__B genblk1\[8\].osc.clkdiv_C.cnt\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13475_ clknet_leaf_71_clk _00792_ net216 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.b1\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10687_ _04869_ genblk1\[5\].osc.clkdiv_C.cnt\[9\] vssd1 vssd1 vccd1 vccd1 _04871_
+ sky130_fd_sc_hd__and2_1
XANTENNA__11013__S _05023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12426_ _05978_ net20 vssd1 vssd1 vccd1 vccd1 _06092_ sky130_fd_sc_hd__nor2_1
XANTENNA__08036__A1 genblk2\[6\].wave_shpr.div.fin_quo\[7\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_112_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10918__A1 net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12357_ _03942_ vssd1 vssd1 vccd1 vccd1 _06039_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_121_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11308_ _05201_ _05171_ vssd1 vssd1 vccd1 vccd1 _05305_ sky130_fd_sc_hd__or2b_1
X_12288_ genblk2\[1\].wave_shpr.div.b1\[12\] _06005_ _05994_ vssd1 vssd1 vccd1 vccd1
+ _06006_ sky130_fd_sc_hd__mux2_1
XANTENNA__08339__A2 _02467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11239_ _05074_ genblk1\[7\].osc.clkdiv_C.cnt\[5\] vssd1 vssd1 vccd1 vccd1 _05259_
+ sky130_fd_sc_hd__and2_1
XANTENNA__11894__A2 _03696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06780_ genblk1\[4\].osc.clkdiv_C.cnt\[16\] _01652_ vssd1 vssd1 vccd1 vccd1 _01654_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_26_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08450_ _03155_ _03156_ genblk2\[8\].wave_shpr.div.fin_quo\[4\] _02521_ vssd1 vssd1
+ vccd1 vccd1 _03157_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_147_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07401_ genblk2\[0\].wave_shpr.div.start vssd1 vssd1 vccd1 vccd1 _02147_ sky130_fd_sc_hd__buf_8
XFILLER_0_148_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08381_ genblk1\[2\].osc.clkdiv_C.cnt\[1\] _01209_ _02336_ genblk1\[2\].osc.clkdiv_C.cnt\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03088_ sky130_fd_sc_hd__a22o_1
XFILLER_0_9_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07332_ genblk1\[11\].osc.clkdiv_C.cnt\[1\] genblk1\[11\].osc.clkdiv_C.cnt\[0\] vssd1
+ vssd1 vccd1 vccd1 _02095_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06806__A _01336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07263_ genblk1\[10\].osc.clkdiv_C.cnt\[4\] _02034_ genblk1\[10\].osc.clkdiv_C.cnt\[5\]
+ vssd1 vssd1 vccd1 vccd1 _02040_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_155_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09002_ net1172 net1176 _01154_ vssd1 vssd1 vccd1 vccd1 _03681_ sky130_fd_sc_hd__mux2_1
X_06214_ freq_div.state\[2\] vssd1 vssd1 vccd1 vccd1 _01176_ sky130_fd_sc_hd__buf_4
XANTENNA__09224__B1 _03840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07194_ genblk1\[9\].osc.clkdiv_C.cnt\[13\] genblk1\[9\].osc.clkdiv_C.cnt\[12\] _01978_
+ vssd1 vssd1 vccd1 vccd1 _01981_ sky130_fd_sc_hd__and3_1
XANTENNA__10909__A1 _04432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09775__A1 _02336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06145_ _01114_ _01116_ vssd1 vssd1 vccd1 vccd1 _01117_ sky130_fd_sc_hd__or2_1
XFILLER_0_77_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout200_A net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09904_ net953 _04315_ _04289_ _04318_ vssd1 vssd1 vccd1 vccd1 _00330_ sky130_fd_sc_hd__a22o_1
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09835_ _02147_ vssd1 vssd1 vccd1 vccd1 _04268_ sky130_fd_sc_hd__buf_4
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09766_ _01302_ _03727_ vssd1 vssd1 vccd1 vccd1 _04233_ sky130_fd_sc_hd__nor2_4
X_06978_ genblk1\[7\].osc.clkdiv_C.cnt\[17\] vssd1 vssd1 vccd1 vccd1 _01814_ sky130_fd_sc_hd__inv_2
XANTENNA__09063__S _03722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08717_ _03386_ _03392_ vssd1 vssd1 vccd1 vccd1 _03424_ sky130_fd_sc_hd__nand2_1
XANTENNA__11098__B1 _05057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09697_ _04171_ genblk2\[2\].wave_shpr.div.acc\[2\] _04176_ vssd1 vssd1 vccd1 vccd1
+ _04177_ sky130_fd_sc_hd__o21a_1
XTAP_2216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08648_ _03280_ _03292_ _03354_ vssd1 vssd1 vccd1 vccd1 _03355_ sky130_fd_sc_hd__a21oi_1
XTAP_1515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_49_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08579_ _03285_ _02404_ vssd1 vssd1 vccd1 vccd1 _03286_ sky130_fd_sc_hd__nor2_1
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10610_ genblk2\[6\].wave_shpr.div.b1\[0\] _01189_ _04637_ vssd1 vssd1 vccd1 vccd1
+ _04830_ sky130_fd_sc_hd__mux2_1
XFILLER_0_119_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11590_ net908 _05447_ _05484_ _05503_ vssd1 vssd1 vccd1 vccd1 _00831_ sky130_fd_sc_hd__a22o_1
XFILLER_0_119_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10073__A1 _04242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10541_ genblk2\[5\].wave_shpr.div.acc\[11\] genblk2\[5\].wave_shpr.div.b1\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04769_ sky130_fd_sc_hd__or2b_1
XFILLER_0_106_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_791 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13260_ clknet_leaf_0_clk _00583_ net38 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.acc\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10472_ _04606_ _04570_ vssd1 vssd1 vccd1 vccd1 _04719_ sky130_fd_sc_hd__or2b_1
XFILLER_0_121_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12211_ genblk2\[11\].wave_shpr.div.b1\[4\] genblk2\[11\].wave_shpr.div.acc\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05949_ sky130_fd_sc_hd__and2b_1
XFILLER_0_32_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13191_ clknet_leaf_122_clk net735 net78 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.i\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_121_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold879_A genblk2\[5\].wave_shpr.div.b1\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12142_ genblk2\[10\].wave_shpr.div.acc\[16\] _05894_ _05865_ vssd1 vssd1 vccd1 vccd1
+ _05895_ sky130_fd_sc_hd__mux2_1
XFILLER_0_102_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07792__A3 _01344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09518__B2 genblk2\[1\].wave_shpr.div.quo\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12073_ genblk2\[10\].wave_shpr.div.b1\[0\] _05787_ genblk2\[10\].wave_shpr.div.acc\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05842_ sky130_fd_sc_hd__a21oi_1
X_11024_ _04998_ _04975_ vssd1 vssd1 vccd1 vccd1 _05107_ sky130_fd_sc_hd__or2b_1
XANTENNA__11089__B1 _05055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12975_ clknet_leaf_124_clk _00304_ net71 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.quo\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11926_ genblk2\[10\].wave_shpr.div.b1\[1\] genblk2\[10\].wave_shpr.div.acc\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05748_ sky130_fd_sc_hd__and2b_1
XTAP_2750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11857_ _05602_ _05556_ vssd1 vssd1 vccd1 vccd1 _05695_ sky130_fd_sc_hd__or2b_1
XFILLER_0_129_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10808_ _04956_ vssd1 vssd1 vccd1 vccd1 _00596_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_82_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11788_ net306 _02203_ _03693_ net565 _05643_ vssd1 vssd1 vccd1 vccd1 _00889_ sky130_fd_sc_hd__a221o_1
XANTENNA__10064__A1 _01589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11261__B1 _05249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13527_ clknet_leaf_98_clk _00844_ net169 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.acc\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_421 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10739_ _04795_ _04905_ vssd1 vssd1 vccd1 vccd1 _04906_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_153_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11800__A2 _05623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13458_ clknet_leaf_99_clk _00775_ net165 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.fin_quo\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_35_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12409_ net897 _06072_ _06073_ _06079_ vssd1 vssd1 vccd1 vccd1 _01074_ sky130_fd_sc_hd__a22o_1
XFILLER_0_106_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13389_ clknet_leaf_78_clk _00708_ net205 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.b1\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07457__A _02189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06361__A _01223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07950_ _01556_ _01564_ genblk1\[7\].osc.clkdiv_C.cnt\[1\] vssd1 vssd1 vccd1 vccd1
+ _02657_ sky130_fd_sc_hd__a21o_1
X_06901_ _01748_ _01749_ _01752_ _01754_ vssd1 vssd1 vccd1 vccd1 _01755_ sky130_fd_sc_hd__or4_1
X_07881_ _02545_ _02518_ _02424_ _02541_ vssd1 vssd1 vccd1 vccd1 _02588_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_128_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09620_ _03998_ _03957_ vssd1 vssd1 vccd1 vccd1 _04117_ sky130_fd_sc_hd__or2b_1
XFILLER_0_37_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06832_ genblk1\[5\].osc.clkdiv_C.cnt\[3\] _01698_ vssd1 vssd1 vccd1 vccd1 _01701_
+ sky130_fd_sc_hd__nor2_1
XANTENNA__07904__B _01869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09551_ net340 _04042_ _04046_ net608 _04066_ vssd1 vssd1 vccd1 vccd1 _00229_ sky130_fd_sc_hd__a221o_1
X_06763_ genblk1\[4\].osc.clkdiv_C.cnt\[12\] _01637_ vssd1 vssd1 vccd1 vccd1 _01641_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_144_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08502_ _03198_ _03197_ vssd1 vssd1 vccd1 vccd1 _03209_ sky130_fd_sc_hd__and2b_1
X_09482_ genblk2\[2\].wave_shpr.div.b1\[8\] _01183_ _04024_ vssd1 vssd1 vccd1 vccd1
+ _04030_ sky130_fd_sc_hd__mux2_1
X_06694_ genblk1\[4\].osc.clkdiv_C.cnt\[11\] _01313_ _01561_ _01582_ _01583_ vssd1
+ vssd1 vccd1 vccd1 _01584_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_66_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_78_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08433_ _02310_ _03139_ _02314_ vssd1 vssd1 vccd1 vccd1 _03140_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout150_A net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08364_ _02846_ _03060_ _03064_ _03066_ _03070_ vssd1 vssd1 vccd1 vccd1 _03071_ sky130_fd_sc_hd__a32o_1
XFILLER_0_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_58_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_760 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10055__A1 _04436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07315_ genblk1\[11\].osc.clkdiv_C.cnt\[8\] _01211_ _02077_ genblk1\[11\].osc.clkdiv_C.cnt\[12\]
+ _02078_ vssd1 vssd1 vccd1 vccd1 _02079_ sky130_fd_sc_hd__o221a_1
X_08295_ _02998_ _03001_ vssd1 vssd1 vccd1 vccd1 _03002_ sky130_fd_sc_hd__nor2_1
XFILLER_0_34_728 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09847__A _04250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07246_ net1080 _02027_ vssd1 vssd1 vccd1 vccd1 genblk1\[10\].osc.clkdiv_C.next_cnt\[0\]
+ sky130_fd_sc_hd__nor2_1
XANTENNA__08751__A genblk2\[7\].wave_shpr.div.fin_quo\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_103_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_103_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07177_ genblk1\[9\].osc.clkdiv_C.cnt\[7\] _01967_ vssd1 vssd1 vccd1 vccd1 _01970_
+ sky130_fd_sc_hd__or2_1
XANTENNA__07759__B1 _02224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06128_ net13 net15 vssd1 vssd1 vccd1 vccd1 _01100_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07504__B_N net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09818_ _04250_ vssd1 vssd1 vccd1 vccd1 _04259_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_fanout63_A net85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09749_ genblk2\[2\].wave_shpr.div.fin_quo\[7\] net1197 _00009_ vssd1 vssd1 vccd1
+ vccd1 _04222_ sky130_fd_sc_hd__mux2_1
XTAP_2002 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2013 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2024 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10818__B1 _04858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12760_ clknet_leaf_93_clk _00001_ net146 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.done
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2035 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2046 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2057 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2068 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2079 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11711_ _05556_ _05601_ _05602_ vssd1 vssd1 vccd1 vccd1 _05603_ sky130_fd_sc_hd__a21oi_2
XTAP_1345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12691_ clknet_leaf_54_clk genblk1\[8\].osc.clkdiv_C.next_cnt\[4\] net174 vssd1 vssd1
+ vccd1 vccd1 genblk1\[8\].osc.clkdiv_C.cnt\[4\] sky130_fd_sc_hd__dfrtp_4
XTAP_1356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11642_ net946 _05448_ _05445_ _05541_ vssd1 vssd1 vccd1 vccd1 _00845_ sky130_fd_sc_hd__a22o_1
XFILLER_0_126_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_119_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11573_ net932 _05447_ _05484_ _05490_ vssd1 vssd1 vccd1 vccd1 _00827_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13312_ clknet_leaf_118_clk _00633_ net138 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10524_ genblk2\[4\].wave_shpr.div.i\[1\] genblk2\[4\].wave_shpr.div.i\[0\] vssd1
+ vssd1 vccd1 vccd1 _04756_ sky130_fd_sc_hd__nand2_1
XFILLER_0_135_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13243_ clknet_leaf_9_clk _00566_ net55 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.quo\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_150_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10455_ _04598_ _04574_ vssd1 vssd1 vccd1 vccd1 _04706_ sky130_fd_sc_hd__or2b_1
XFILLER_0_33_772 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13174_ clknet_leaf_129_clk _00499_ net65 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.acc\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10386_ net602 _04657_ _04655_ genblk2\[4\].wave_shpr.div.quo\[10\] _04660_ vssd1
+ vssd1 vccd1 vccd1 _00470_ sky130_fd_sc_hd__a221o_1
XFILLER_0_103_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12125_ genblk2\[10\].wave_shpr.div.acc\[12\] _05881_ _05865_ vssd1 vssd1 vccd1 vccd1
+ _05882_ sky130_fd_sc_hd__mux2_1
XANTENNA__09492__A _01411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12056_ net440 _05823_ _05825_ net518 _05832_ vssd1 vssd1 vccd1 vccd1 _00968_ sky130_fd_sc_hd__a221o_1
XFILLER_0_74_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11007_ _04990_ _04979_ vssd1 vssd1 vccd1 vccd1 _05094_ sky130_fd_sc_hd__or2b_1
XFILLER_0_74_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12958_ clknet_leaf_136_clk _00287_ net42 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.b1\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_90_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08478__B2 _02308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11909_ genblk2\[10\].wave_shpr.div.acc\[17\] genblk2\[10\].wave_shpr.div.b1\[17\]
+ vssd1 vssd1 vccd1 vccd1 _05731_ sky130_fd_sc_hd__or2b_1
XTAP_2580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12889_ clknet_leaf_30_clk _00220_ net96 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.quo\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12358__A _03941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11262__A _04676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12026__A2 _05813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_55_341 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09089__D _03738_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07100_ _01887_ _01906_ vssd1 vssd1 vccd1 vccd1 _01907_ sky130_fd_sc_hd__nor2_1
XFILLER_0_126_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_130_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08080_ _01200_ _01680_ _02748_ _02749_ vssd1 vssd1 vccd1 vccd1 _02787_ sky130_fd_sc_hd__o22a_1
XFILLER_0_126_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07031_ _01822_ _01849_ _01850_ vssd1 vssd1 vccd1 vccd1 _01851_ sky130_fd_sc_hd__and3b_1
XFILLER_0_130_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_113_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__13550__RESET_B net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08982_ _01097_ _03570_ _03666_ vssd1 vssd1 vccd1 vccd1 _03667_ sky130_fd_sc_hd__or3_1
X_07933_ genblk2\[8\].wave_shpr.div.fin_quo\[3\] _02639_ vssd1 vssd1 vccd1 vccd1 _02640_
+ sky130_fd_sc_hd__or2_1
XANTENNA_fanout198_A net218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07864_ _02517_ _02566_ _02570_ vssd1 vssd1 vccd1 vccd1 _02571_ sky130_fd_sc_hd__a21o_1
XANTENNA__10341__A _03701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09603_ _03989_ _04103_ vssd1 vssd1 vccd1 vccd1 _04104_ sky130_fd_sc_hd__xnor2_1
X_06815_ genblk1\[5\].osc.clkdiv_C.cnt\[12\] _01355_ vssd1 vssd1 vccd1 vccd1 _01687_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07795_ genblk1\[0\].osc.clkdiv_C.cnt\[9\] _01184_ vssd1 vssd1 vccd1 vccd1 _02502_
+ sky130_fd_sc_hd__nand2_1
Xwire20 _06088_ vssd1 vssd1 vccd1 vccd1 net20 sky130_fd_sc_hd__buf_1
Xwire31 _02508_ vssd1 vssd1 vccd1 vccd1 net31 sky130_fd_sc_hd__clkbuf_2
X_09534_ net511 _04052_ _04053_ net519 _04057_ vssd1 vssd1 vccd1 vccd1 _00221_ sky130_fd_sc_hd__a221o_1
X_06746_ _01627_ vssd1 vssd1 vccd1 vccd1 _01628_ sky130_fd_sc_hd__inv_2
XANTENNA__09666__B1 _04048_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10487__S _04704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09465_ _04020_ vssd1 vssd1 vccd1 vccd1 _00189_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06677_ genblk1\[4\].osc.clkdiv_C.cnt\[5\] _01565_ vssd1 vssd1 vccd1 vccd1 _01567_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_365 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08416_ _03114_ _03121_ _03122_ vssd1 vssd1 vccd1 vccd1 _03123_ sky130_fd_sc_hd__o21ai_1
X_09396_ genblk2\[1\].wave_shpr.div.acc\[11\] genblk2\[1\].wave_shpr.div.b1\[11\]
+ vssd1 vssd1 vccd1 vccd1 _03960_ sky130_fd_sc_hd__or2b_1
XFILLER_0_47_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11225__B1 _05250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08347_ _03030_ _03051_ _03052_ _03053_ vssd1 vssd1 vccd1 vccd1 _03054_ sky130_fd_sc_hd__o211a_1
XFILLER_0_47_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_117_763 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_61_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_116_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08278_ _02303_ _02264_ genblk2\[9\].wave_shpr.div.fin_quo\[4\] vssd1 vssd1 vccd1
+ vccd1 _02985_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_62_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_131_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07229_ _01229_ _01230_ vssd1 vssd1 vccd1 vccd1 _02011_ sky130_fd_sc_hd__nand2_4
XFILLER_0_15_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10240_ _04556_ vssd1 vssd1 vccd1 vccd1 _00428_ sky130_fd_sc_hd__clkbuf_1
X_10171_ _04394_ _04505_ vssd1 vssd1 vccd1 vccd1 _04506_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xfanout140 net145 vssd1 vssd1 vccd1 vccd1 net140 sky130_fd_sc_hd__clkbuf_4
Xfanout151 net152 vssd1 vssd1 vccd1 vccd1 net151 sky130_fd_sc_hd__clkbuf_4
Xfanout162 net163 vssd1 vssd1 vccd1 vccd1 net162 sky130_fd_sc_hd__clkbuf_2
Xfanout173 net174 vssd1 vssd1 vccd1 vccd1 net173 sky130_fd_sc_hd__clkbuf_4
Xfanout184 net185 vssd1 vssd1 vccd1 vccd1 net184 sky130_fd_sc_hd__buf_2
XANTENNA__10503__A2 _04715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_709 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout195 net198 vssd1 vssd1 vccd1 vccd1 net195 sky130_fd_sc_hd__clkbuf_2
X_12812_ clknet_leaf_58_clk net266 net192 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.quo\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_96_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_96_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_70_clk_A clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1120 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12743_ clknet_leaf_49_clk genblk1\[11\].osc.clkdiv_C.next_cnt\[2\] net108 vssd1
+ vssd1 vccd1 vccd1 genblk1\[11\].osc.clkdiv_C.cnt\[2\] sky130_fd_sc_hd__dfrtp_4
XTAP_1131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07132__B2 genblk1\[9\].osc.clkdiv_C.cnt\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_831 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12674_ clknet_leaf_90_clk genblk1\[7\].osc.clkdiv_C.next_cnt\[5\] net174 vssd1 vssd1
+ vccd1 vccd1 genblk1\[7\].osc.clkdiv_C.cnt\[5\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_154_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11625_ genblk2\[8\].wave_shpr.div.acc\[18\] _05529_ vssd1 vssd1 vccd1 vccd1 _05530_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__06891__B1 _01484_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_85_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11556_ _05449_ _05475_ _05477_ _05448_ net699 vssd1 vssd1 vccd1 vccd1 _00823_ sky130_fd_sc_hd__a32o_1
XFILLER_0_13_709 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06904__A _01576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_664 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10507_ _04619_ _04622_ vssd1 vssd1 vccd1 vccd1 _04745_ sky130_fd_sc_hd__and2b_1
XFILLER_0_107_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11487_ net713 vssd1 vssd1 vccd1 vccd1 _05439_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_720 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10990__A2 _05023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13226_ clknet_leaf_127_clk net254 net132 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_100_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10438_ net842 _04683_ _04690_ _04693_ vssd1 vssd1 vccd1 vccd1 _00489_ sky130_fd_sc_hd__a22o_1
XANTENNA__07199__A1 genblk1\[9\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08396__B1 _01209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_122_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_904 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13157_ clknet_leaf_121_clk _00482_ net78 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.quo\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_915 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10369_ _04654_ vssd1 vssd1 vccd1 vccd1 _04655_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_85_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_926 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12108_ genblk2\[10\].wave_shpr.div.acc\[8\] _05868_ _05865_ vssd1 vssd1 vccd1 vccd1
+ _05869_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_948 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13088_ clknet_leaf_137_clk _00415_ net40 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.acc\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_959 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08148__B1 _01513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_23_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12039_ _05812_ vssd1 vssd1 vccd1 vccd1 _05823_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_18_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_18_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_1_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_1_0_clk sky130_fd_sc_hd__clkbuf_8
X_06600_ _01241_ _01432_ vssd1 vssd1 vccd1 vccd1 _01508_ sky130_fd_sc_hd__nor2_2
X_07580_ _01432_ _01221_ genblk1\[9\].osc.clkdiv_C.cnt\[1\] vssd1 vssd1 vccd1 vccd1
+ _02287_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_38_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06531_ genblk1\[2\].osc.clkdiv_C.cnt\[1\] genblk1\[2\].osc.clkdiv_C.cnt\[0\] genblk1\[2\].osc.clkdiv_C.cnt\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01455_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_125_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09250_ _03853_ genblk1\[0\].osc.clkdiv_C.cnt\[9\] vssd1 vssd1 vccd1 vccd1 _03854_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_146_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06462_ genblk1\[1\].osc.clkdiv_C.cnt\[10\] _01394_ vssd1 vssd1 vccd1 vccd1 _01396_
+ sky130_fd_sc_hd__nand2_1
X_08201_ net17 _02552_ genblk2\[10\].wave_shpr.div.fin_quo\[6\] vssd1 vssd1 vccd1
+ vccd1 _02908_ sky130_fd_sc_hd__and3_1
XFILLER_0_90_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06882__B1 _01735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09181_ _03817_ vssd1 vssd1 vccd1 vccd1 _00108_ sky130_fd_sc_hd__clkbuf_1
X_06393_ _01336_ _01226_ vssd1 vssd1 vccd1 vccd1 _01337_ sky130_fd_sc_hd__nor2_4
XFILLER_0_29_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08132_ genblk2\[4\].wave_shpr.div.fin_quo\[0\] genblk2\[4\].wave_shpr.div.fin_quo\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02839_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_114_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08063_ genblk1\[5\].osc.clkdiv_C.cnt\[2\] _01238_ net35 vssd1 vssd1 vccd1 vccd1
+ _02770_ sky130_fd_sc_hd__or3_1
XFILLER_0_43_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07014_ genblk1\[7\].osc.clkdiv_C.cnt\[10\] _01837_ _01839_ vssd1 vssd1 vccd1 vccd1
+ genblk1\[7\].osc.clkdiv_C.next_cnt\[10\] sky130_fd_sc_hd__o21a_1
XFILLER_0_101_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_113_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_59_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08965_ _03650_ _03652_ vssd1 vssd1 vccd1 vccd1 _03653_ sky130_fd_sc_hd__xnor2_1
X_07916_ genblk1\[8\].osc.clkdiv_C.cnt\[4\] _01487_ vssd1 vssd1 vccd1 vccd1 _02623_
+ sky130_fd_sc_hd__or2_1
X_08896_ sig_norm.b1\[0\] _03578_ _03580_ vssd1 vssd1 vccd1 vccd1 _03601_ sky130_fd_sc_hd__nand3_1
X_07847_ _02217_ _02553_ genblk2\[0\].wave_shpr.div.fin_quo\[3\] vssd1 vssd1 vccd1
+ vccd1 _02554_ sky130_fd_sc_hd__and3_1
XFILLER_0_98_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07778_ _01181_ genblk1\[0\].osc.clkdiv_C.cnt\[7\] _01198_ vssd1 vssd1 vccd1 vccd1
+ _02485_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11446__A0 genblk2\[8\].wave_shpr.div.fin_quo\[2\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09517_ genblk2\[1\].wave_shpr.div.quo\[7\] _04043_ _04047_ net292 vssd1 vssd1 vccd1
+ vccd1 _00214_ sky130_fd_sc_hd__a22o_1
X_06729_ _01600_ _01613_ _01614_ vssd1 vssd1 vccd1 vccd1 _01615_ sky130_fd_sc_hd__and3_1
XANTENNA__13532__D _00023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11997__A1 _01556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09448_ genblk2\[1\].wave_shpr.div.fin_quo\[0\] _04011_ _00007_ vssd1 vssd1 vccd1
+ vccd1 _04012_ sky130_fd_sc_hd__mux2_1
XPHY_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09379_ _03942_ vssd1 vssd1 vccd1 vccd1 _03947_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_47_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11410_ genblk2\[8\].wave_shpr.div.b1\[6\] genblk2\[8\].wave_shpr.div.acc\[6\] vssd1
+ vssd1 vccd1 vccd1 _05386_ sky130_fd_sc_hd__and2b_1
X_12390_ genblk2\[11\].wave_shpr.div.acc\[10\] _06064_ _06055_ vssd1 vssd1 vccd1 vccd1
+ _06065_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_35_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_151_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11341_ net628 _05311_ _05315_ _05330_ vssd1 vssd1 vccd1 vccd1 _00755_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11272_ genblk2\[7\].wave_shpr.div.acc\[1\] _05277_ _05222_ vssd1 vssd1 vccd1 vccd1
+ _05278_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13011_ clknet_leaf_133_clk _00340_ net59 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.acc\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10223_ net524 _04518_ _04522_ _04545_ vssd1 vssd1 vccd1 vccd1 _00422_ sky130_fd_sc_hd__a22o_1
XANTENNA__09754__B _01925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10154_ net979 _04486_ _04490_ _04493_ vssd1 vssd1 vccd1 vccd1 _00405_ sky130_fd_sc_hd__a22o_1
XFILLER_0_100_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10085_ net794 _04452_ _04420_ _04454_ vssd1 vssd1 vccd1 vccd1 _00375_ sky130_fd_sc_hd__a22o_1
Xhold7 modein.delay_octave_down_in\[0\] vssd1 vssd1 vccd1 vccd1 net225 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11524__B genblk1\[8\].osc.clkdiv_C.cnt\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10987_ _05054_ vssd1 vssd1 vccd1 vccd1 _05079_ sky130_fd_sc_hd__inv_2
XANTENNA__11988__A1 _01946_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12726_ clknet_leaf_37_clk genblk1\[10\].osc.clkdiv_C.next_cnt\[3\] net113 vssd1
+ vssd1 vccd1 vccd1 genblk1\[10\].osc.clkdiv_C.cnt\[3\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_128_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12657_ clknet_leaf_27_clk genblk1\[6\].osc.clkdiv_C.next_cnt\[6\] net90 vssd1 vssd1
+ vccd1 vccd1 genblk1\[6\].osc.clkdiv_C.cnt\[6\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_154_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11608_ _05402_ _05361_ vssd1 vssd1 vccd1 vccd1 _05517_ sky130_fd_sc_hd__or2b_1
XFILLER_0_143_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08066__C1 genblk1\[5\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09802__B1 _04252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12588_ clknet_leaf_14_clk genblk1\[2\].osc.clkdiv_C.next_cnt\[9\] net72 vssd1 vssd1
+ vccd1 vccd1 genblk1\[2\].osc.clkdiv_C.cnt\[9\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_80_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07449__B _02153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11539_ _05464_ genblk1\[8\].osc.clkdiv_C.cnt\[13\] vssd1 vssd1 vccd1 vccd1 _05467_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_20_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold407 genblk2\[5\].wave_shpr.div.b1\[5\] vssd1 vssd1 vccd1 vccd1 net625 sky130_fd_sc_hd__dlygate4sd3_1
Xhold418 genblk2\[0\].wave_shpr.div.quo\[20\] vssd1 vssd1 vccd1 vccd1 net636 sky130_fd_sc_hd__dlygate4sd3_1
Xhold429 _00913_ vssd1 vssd1 vccd1 vccd1 net647 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_0_433 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13209_ clknet_leaf_25_clk _00532_ net86 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.b1\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_477 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06395__A2 _01210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08750_ _03455_ _03456_ vssd1 vssd1 vccd1 vccd1 _03457_ sky130_fd_sc_hd__or2_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1107 genblk2\[8\].wave_shpr.div.quo\[5\] vssd1 vssd1 vccd1 vccd1 net1325 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1118 genblk2\[5\].wave_shpr.div.quo\[1\] vssd1 vssd1 vccd1 vccd1 net1336 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1129 genblk2\[7\].wave_shpr.div.quo\[0\] vssd1 vssd1 vccd1 vccd1 net1347 sky130_fd_sc_hd__dlygate4sd3_1
X_07701_ genblk2\[10\].wave_shpr.div.fin_quo\[2\] _02407_ vssd1 vssd1 vccd1 vccd1
+ _02408_ sky130_fd_sc_hd__and2b_1
X_08681_ _03113_ _03115_ genblk2\[2\].wave_shpr.div.fin_quo\[2\] vssd1 vssd1 vccd1
+ vccd1 _03388_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_136_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08541__B1 _02308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07632_ genblk1\[11\].osc.clkdiv_C.cnt\[10\] _01262_ _02338_ vssd1 vssd1 vccd1 vccd1
+ _02339_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_136_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07563_ _01930_ _01556_ _01564_ _01801_ _01928_ vssd1 vssd1 vccd1 vccd1 _02270_ sky130_fd_sc_hd__a32o_1
XANTENNA__07631__C _01249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09302_ genblk2\[0\].wave_shpr.div.acc\[7\] _03888_ _03889_ vssd1 vssd1 vccd1 vccd1
+ _03890_ sky130_fd_sc_hd__mux2_1
XFILLER_0_152_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06514_ _01191_ vssd1 vssd1 vccd1 vccd1 _01440_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07494_ net17 vssd1 vssd1 vccd1 vccd1 _02216_ sky130_fd_sc_hd__buf_2
XANTENNA__10100__B1 _04454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_91_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_8_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_75_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09233_ _03725_ genblk1\[0\].osc.clkdiv_C.cnt\[2\] vssd1 vssd1 vccd1 vccd1 _03844_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_35_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06445_ _01384_ vssd1 vssd1 vccd1 vccd1 genblk1\[1\].osc.clkdiv_C.next_cnt\[4\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_29_683 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_146_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09164_ _03808_ vssd1 vssd1 vccd1 vccd1 _00100_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06376_ freq_div.state\[0\] _01178_ vssd1 vssd1 vccd1 vccd1 _01320_ sky130_fd_sc_hd__xnor2_4
XFILLER_0_127_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08115_ _01172_ _01180_ _01568_ vssd1 vssd1 vccd1 vccd1 _02822_ sky130_fd_sc_hd__a21oi_1
XANTENNA__06607__B1 _01514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_133_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08072__A2 _01309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09095_ _01211_ _01556_ _03743_ vssd1 vssd1 vccd1 vccd1 _03744_ sky130_fd_sc_hd__mux2_1
XFILLER_0_142_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_761 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09855__A _04214_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08046_ genblk1\[5\].osc.clkdiv_C.cnt\[13\] _01674_ _01666_ genblk1\[5\].osc.clkdiv_C.cnt\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02753_ sky130_fd_sc_hd__o22a_1
XFILLER_0_31_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold930 genblk2\[3\].wave_shpr.div.i\[3\] vssd1 vssd1 vccd1 vccd1 net1148 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold941 genblk1\[2\].osc.clkdiv_C.cnt\[10\] vssd1 vssd1 vccd1 vccd1 net1159 sky130_fd_sc_hd__dlygate4sd3_1
Xhold952 sig_norm.quo\[4\] vssd1 vssd1 vccd1 vccd1 net1170 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold963 genblk2\[7\].wave_shpr.div.i\[3\] vssd1 vssd1 vccd1 vccd1 net1181 sky130_fd_sc_hd__dlygate4sd3_1
Xhold974 genblk2\[4\].wave_shpr.div.b1\[11\] vssd1 vssd1 vccd1 vccd1 net1192 sky130_fd_sc_hd__dlygate4sd3_1
Xhold985 genblk2\[11\].wave_shpr.div.acc\[20\] vssd1 vssd1 vccd1 vccd1 net1203 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11903__A1 _03839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold996 genblk2\[8\].wave_shpr.div.b1\[3\] vssd1 vssd1 vccd1 vccd1 net1214 sky130_fd_sc_hd__dlygate4sd3_1
X_09997_ genblk2\[3\].wave_shpr.div.b1\[7\] genblk2\[3\].wave_shpr.div.acc\[7\] vssd1
+ vssd1 vccd1 vccd1 _04393_ sky130_fd_sc_hd__and2b_1
XANTENNA__07583__A1 genblk1\[9\].osc.clkdiv_C.cnt\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08948_ _01098_ _03559_ vssd1 vssd1 vccd1 vccd1 _03639_ sky130_fd_sc_hd__or2_1
X_08879_ _03575_ sig_norm.acc\[3\] _03584_ vssd1 vssd1 vccd1 vccd1 _03585_ sky130_fd_sc_hd__o21a_1
XANTENNA__08532__B1 net2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10910_ _05039_ vssd1 vssd1 vccd1 vccd1 _00615_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07822__B net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07886__A2 _02539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11890_ genblk2\[9\].wave_shpr.div.acc\[24\] _05646_ _05715_ vssd1 vssd1 vccd1 vccd1
+ _05719_ sky130_fd_sc_hd__or3b_1
X_10841_ _04982_ _04983_ _04984_ vssd1 vssd1 vccd1 vccd1 _04985_ sky130_fd_sc_hd__o21ai_1
X_13560_ clknet_leaf_84_clk net291 net184 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.quo\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10772_ net925 _04918_ _04922_ _04931_ vssd1 vssd1 vccd1 vccd1 _00585_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12511_ clknet_leaf_84_clk _00073_ net202 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.i\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_54_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10642__A1 _04645_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13491_ clknet_leaf_88_clk _00808_ net177 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.quo\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_81_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12442_ genblk2\[11\].wave_shpr.div.acc\[24\] _05980_ genblk2\[11\].wave_shpr.div.acc\[25\]
+ vssd1 vssd1 vccd1 vccd1 _06102_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_35_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_124_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12373_ genblk2\[11\].wave_shpr.div.acc\[6\] _06051_ _05982_ vssd1 vssd1 vccd1 vccd1
+ _06052_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10945__A2 _05052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11324_ genblk2\[7\].wave_shpr.div.acc\[13\] _05317_ _05300_ vssd1 vssd1 vccd1 vccd1
+ _05318_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11255_ genblk2\[7\].wave_shpr.div.quo\[21\] _05255_ _05256_ net527 _05267_ vssd1
+ vssd1 vccd1 vccd1 _00732_ sky130_fd_sc_hd__a221o_1
XFILLER_0_31_892 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10206_ _04532_ _04410_ vssd1 vssd1 vccd1 vccd1 _04533_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11519__B genblk1\[8\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11186_ genblk2\[8\].wave_shpr.div.b1\[5\] _01508_ _05042_ vssd1 vssd1 vccd1 vccd1
+ _05233_ sky130_fd_sc_hd__mux2_1
XANTENNA__07574__A1 _01336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10137_ _04417_ _04418_ vssd1 vssd1 vccd1 vccd1 _04480_ sky130_fd_sc_hd__nor2_2
X_10068_ _01325_ _01226_ vssd1 vssd1 vccd1 vccd1 _04444_ sky130_fd_sc_hd__nor2_2
XFILLER_0_82_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12130__S _05865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_85_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13758_ clknet_leaf_66_clk _01069_ net197 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.acc\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12083__B1 _05817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13394__RESET_B net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_57_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12709_ clknet_leaf_56_clk genblk1\[9\].osc.clkdiv_C.next_cnt\[4\] net181 vssd1 vssd1
+ vccd1 vccd1 genblk1\[9\].osc.clkdiv_C.cnt\[4\] sky130_fd_sc_hd__dfrtp_4
X_13689_ clknet_leaf_57_clk _00004_ net184 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.busy
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_759 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06230_ _01175_ _01191_ vssd1 vssd1 vccd1 vccd1 _01192_ sky130_fd_sc_hd__nand2_4
XFILLER_0_127_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_26_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06161_ _01130_ _01132_ vssd1 vssd1 vccd1 vccd1 _01133_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold204 _00719_ vssd1 vssd1 vccd1 vccd1 net422 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold215 _00958_ vssd1 vssd1 vccd1 vccd1 net433 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07801__A2 _01577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold226 _01045_ vssd1 vssd1 vccd1 vccd1 net444 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold237 _00147_ vssd1 vssd1 vccd1 vccd1 net455 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09920_ genblk2\[2\].wave_shpr.div.acc\[16\] _04330_ _04301_ vssd1 vssd1 vccd1 vccd1
+ _04331_ sky130_fd_sc_hd__mux2_1
Xhold248 genblk2\[0\].wave_shpr.div.quo\[18\] vssd1 vssd1 vccd1 vccd1 net466 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_22_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold259 genblk2\[6\].wave_shpr.div.quo\[9\] vssd1 vssd1 vccd1 vccd1 net477 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10149__B1 _04456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06811__B _01326_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09851_ genblk2\[2\].wave_shpr.div.b1\[0\] genblk2\[2\].wave_shpr.div.acc\[0\] _04214_
+ _04275_ vssd1 vssd1 vccd1 vccd1 _04278_ sky130_fd_sc_hd__a31o_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08802_ _03219_ _03222_ _03220_ _03221_ vssd1 vssd1 vccd1 vccd1 _03509_ sky130_fd_sc_hd__o211a_1
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11361__A2 _05248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06672__A2_N _01326_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09782_ _03702_ _01490_ vssd1 vssd1 vccd1 vccd1 _04241_ sky130_fd_sc_hd__nand2_4
X_06994_ genblk1\[7\].osc.clkdiv_C.cnt\[3\] _01825_ vssd1 vssd1 vccd1 vccd1 _01827_
+ sky130_fd_sc_hd__and2_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08733_ _03175_ _03201_ _03200_ vssd1 vssd1 vccd1 vccd1 _03440_ sky130_fd_sc_hd__o21a_1
XANTENNA_fanout180_A net185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08664_ _02798_ _03370_ vssd1 vssd1 vccd1 vccd1 _03371_ sky130_fd_sc_hd__nand2_1
XFILLER_0_139_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_07615_ genblk1\[11\].osc.clkdiv_C.cnt\[2\] _01186_ _01437_ _01225_ vssd1 vssd1 vccd1
+ vccd1 _02322_ sky130_fd_sc_hd__or4_1
XTAP_1719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08595_ _02798_ _03299_ _03301_ vssd1 vssd1 vccd1 vccd1 _03302_ sky130_fd_sc_hd__and3_1
XFILLER_0_76_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07546_ _02256_ vssd1 vssd1 vccd1 vccd1 _00034_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09490__A1 _04034_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07477_ _02201_ _02153_ genblk2\[9\].wave_shpr.div.busy vssd1 vssd1 vccd1 vccd1 _02204_
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_63_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11180__A _03708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_146_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09216_ _03837_ vssd1 vssd1 vccd1 vccd1 _03838_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_17_642 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06428_ genblk1\[1\].osc.clkdiv_C.cnt\[0\] _01304_ _01319_ _01331_ _01371_ vssd1
+ vssd1 vccd1 vccd1 _01372_ sky130_fd_sc_hd__a2111oi_2
XFILLER_0_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_44_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09147_ genblk2\[0\].wave_shpr.div.b1\[16\] genblk2\[0\].wave_shpr.div.acc\[16\]
+ vssd1 vssd1 vccd1 vccd1 _03795_ sky130_fd_sc_hd__and2b_1
XFILLER_0_32_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08045__A2 _01675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06359_ _01179_ _01222_ _01302_ vssd1 vssd1 vccd1 vccd1 _01303_ sky130_fd_sc_hd__or3_1
XFILLER_0_32_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_115_872 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_20_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09078_ _03702_ vssd1 vssd1 vccd1 vccd1 _03732_ sky130_fd_sc_hd__buf_8
XFILLER_0_102_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08029_ genblk2\[6\].wave_shpr.div.fin_quo\[2\] _02735_ vssd1 vssd1 vccd1 vccd1 _02736_
+ sky130_fd_sc_hd__or2_1
XANTENNA__07817__B net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold760 genblk2\[8\].wave_shpr.div.acc\[8\] vssd1 vssd1 vccd1 vccd1 net978 sky130_fd_sc_hd__dlygate4sd3_1
Xhold771 genblk2\[10\].wave_shpr.div.acc\[2\] vssd1 vssd1 vccd1 vccd1 net989 sky130_fd_sc_hd__dlygate4sd3_1
Xhold782 genblk2\[3\].wave_shpr.div.acc\[23\] vssd1 vssd1 vccd1 vccd1 net1000 sky130_fd_sc_hd__dlygate4sd3_1
X_11040_ _05051_ vssd1 vssd1 vccd1 vccd1 _05119_ sky130_fd_sc_hd__clkbuf_4
Xhold793 _00753_ vssd1 vssd1 vccd1 vccd1 net1011 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11888__B1 _03696_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12991_ clknet_leaf_130_clk _00320_ net65 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.acc\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08505__B1 _02224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11942_ genblk2\[10\].wave_shpr.div.b1\[9\] genblk2\[10\].wave_shpr.div.acc\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05764_ sky130_fd_sc_hd__and2b_1
XFILLER_0_99_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_98_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11873_ genblk2\[9\].wave_shpr.div.acc\[19\] _05704_ vssd1 vssd1 vccd1 vccd1 _05707_
+ sky130_fd_sc_hd__or2_1
X_13612_ clknet_leaf_94_clk _00925_ net159 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.fin_quo\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10824_ genblk2\[6\].wave_shpr.div.acc\[15\] genblk2\[6\].wave_shpr.div.b1\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04968_ sky130_fd_sc_hd__or2b_1
XANTENNA__12065__B1 _05815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10615__A1 _01684_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13543_ clknet_leaf_101_clk _00858_ net164 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.fin_quo\[5\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_54_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_512 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10755_ _02183_ vssd1 vssd1 vccd1 vccd1 _04918_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_55_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_94_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06295__A1 _01188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10091__A2 _04452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13474_ clknet_leaf_71_clk _00791_ net215 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.b1\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_10686_ net235 _04861_ _04862_ net378 _04870_ vssd1 vssd1 vccd1 vccd1 _00560_ sky130_fd_sc_hd__a221o_1
XFILLER_0_82_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12425_ net641 _06072_ _06073_ _06091_ vssd1 vssd1 vccd1 vccd1 _01078_ sky130_fd_sc_hd__a22o_1
XFILLER_0_63_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_125_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08036__A2 _02539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_140_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12356_ net1020 _06009_ _06010_ _06038_ vssd1 vssd1 vccd1 vccd1 _01062_ sky130_fd_sc_hd__a22o_1
X_11307_ net797 _05279_ _05283_ _05304_ vssd1 vssd1 vccd1 vccd1 _00747_ sky130_fd_sc_hd__a22o_1
XFILLER_0_121_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12125__S _05865_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10434__A _04654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12287_ _01337_ vssd1 vssd1 vccd1 vccd1 _06005_ sky130_fd_sc_hd__inv_2
X_11238_ net640 _05255_ _05256_ net670 _05258_ vssd1 vssd1 vccd1 vccd1 _00724_ sky130_fd_sc_hd__a221o_1
X_11169_ genblk2\[7\].wave_shpr.div.fin_quo\[3\] genblk2\[7\].wave_shpr.div.quo\[2\]
+ _00019_ vssd1 vssd1 vccd1 vccd1 _05226_ sky130_fd_sc_hd__mux2_1
XFILLER_0_117_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06359__A _01179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07400_ net1220 _02145_ vssd1 vssd1 vccd1 vccd1 genblk1\[11\].osc.clkdiv_C.next_cnt\[17\]
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_9_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08380_ genblk1\[2\].osc.clkdiv_C.cnt\[1\] _01209_ _02425_ genblk1\[2\].osc.clkdiv_C.cnt\[0\]
+ vssd1 vssd1 vccd1 vccd1 _03087_ sky130_fd_sc_hd__o211a_1
XFILLER_0_92_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07331_ genblk1\[11\].osc.clkdiv_C.cnt\[1\] genblk1\[11\].osc.clkdiv_C.cnt\[0\] vssd1
+ vssd1 vccd1 vccd1 _02094_ sky130_fd_sc_hd__or2_1
XFILLER_0_128_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08275__A2 _02361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_73_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06806__B _01564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07262_ genblk1\[10\].osc.clkdiv_C.cnt\[5\] genblk1\[10\].osc.clkdiv_C.cnt\[4\] _02034_
+ vssd1 vssd1 vccd1 vccd1 _02039_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_834 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09001_ _03680_ vssd1 vssd1 vccd1 vccd1 _00065_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06213_ freq_div.state\[1\] vssd1 vssd1 vccd1 vccd1 _01175_ sky130_fd_sc_hd__buf_4
X_07193_ net1296 _01978_ _01980_ vssd1 vssd1 vccd1 vccd1 genblk1\[9\].osc.clkdiv_C.next_cnt\[12\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_131_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_133 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06144_ _01113_ _01115_ vssd1 vssd1 vccd1 vccd1 _01116_ sky130_fd_sc_hd__nand2_1
XANTENNA__07918__A _01489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10344__A _01678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09903_ genblk2\[2\].wave_shpr.div.acc\[12\] _04317_ _04301_ vssd1 vssd1 vccd1 vccd1
+ _04318_ sky130_fd_sc_hd__mux2_1
Xwire5 _02589_ vssd1 vssd1 vccd1 vccd1 net1354 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09834_ genblk2\[2\].wave_shpr.div.quo\[20\] _04257_ _04259_ net322 _04267_ vssd1
+ vssd1 vccd1 vccd1 _00311_ sky130_fd_sc_hd__a221o_1
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09765_ _04232_ vssd1 vssd1 vccd1 vccd1 _00277_ sky130_fd_sc_hd__clkbuf_1
X_06977_ genblk1\[7\].osc.clkdiv_C.cnt\[16\] vssd1 vssd1 vccd1 vccd1 _01813_ sky130_fd_sc_hd__inv_2
X_08716_ _03387_ _03391_ vssd1 vssd1 vccd1 vccd1 _03423_ sky130_fd_sc_hd__or2b_1
XANTENNA__11098__A1 _05055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09696_ _04174_ _04175_ _04172_ vssd1 vssd1 vccd1 vccd1 _04176_ sky130_fd_sc_hd__o21ai_1
XTAP_2206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06269__A _01229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08647_ _03289_ _03290_ _02419_ _03284_ vssd1 vssd1 vccd1 vccd1 _03354_ sky130_fd_sc_hd__o211a_1
XFILLER_0_68_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08578_ genblk2\[10\].wave_shpr.div.fin_quo\[0\] vssd1 vssd1 vccd1 vccd1 _03285_
+ sky130_fd_sc_hd__inv_2
XTAP_1549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07529_ _01099_ _02245_ _02246_ vssd1 vssd1 vccd1 vccd1 _02247_ sky130_fd_sc_hd__and3_1
XFILLER_0_9_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10540_ genblk2\[5\].wave_shpr.div.acc\[12\] genblk2\[5\].wave_shpr.div.b1\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04768_ sky130_fd_sc_hd__or2b_1
XFILLER_0_119_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_134_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10471_ net778 _04715_ _04690_ _04718_ vssd1 vssd1 vccd1 vccd1 _00497_ sky130_fd_sc_hd__a22o_1
X_12210_ _05939_ _05946_ _05947_ vssd1 vssd1 vccd1 vccd1 _05948_ sky130_fd_sc_hd__a21o_1
XFILLER_0_121_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13190_ clknet_leaf_118_clk _00513_ net138 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.i\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_12141_ _05893_ _05777_ vssd1 vssd1 vccd1 vccd1 _05894_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_60_795 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_102_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09518__A2 _04043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12072_ genblk2\[10\].wave_shpr.div.acc\[0\] _00002_ _05840_ net247 _05841_ vssd1
+ vssd1 vccd1 vccd1 _00975_ sky130_fd_sc_hd__o221a_1
Xhold590 genblk2\[7\].wave_shpr.div.acc\[13\] vssd1 vssd1 vccd1 vccd1 net808 sky130_fd_sc_hd__dlygate4sd3_1
X_11023_ net867 _05086_ _05093_ _05106_ vssd1 vssd1 vccd1 vccd1 _00661_ sky130_fd_sc_hd__a22o_1
XANTENNA__10533__B1 _03855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12974_ clknet_leaf_124_clk net554 net71 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.quo\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11925_ genblk2\[10\].wave_shpr.div.acc\[0\] genblk2\[10\].wave_shpr.div.b1\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05747_ sky130_fd_sc_hd__or2b_1
XTAP_2740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12038__B1 _05816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06517__A2_N _01439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11856_ net912 _05684_ _05685_ _05694_ vssd1 vssd1 vccd1 vccd1 _00906_ sky130_fd_sc_hd__a22o_1
XTAP_2784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_704 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_68_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_74_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_670 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10807_ _04856_ _02183_ genblk2\[5\].wave_shpr.div.i\[0\] vssd1 vssd1 vccd1 vccd1
+ _04956_ sky130_fd_sc_hd__mux2_1
X_11787_ _05631_ genblk1\[9\].osc.clkdiv_C.cnt\[15\] vssd1 vssd1 vccd1 vccd1 _05643_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_94_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10738_ _04796_ _04772_ vssd1 vssd1 vccd1 vccd1 _04905_ sky130_fd_sc_hd__or2b_1
X_13526_ clknet_leaf_98_clk _00843_ net169 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.acc\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_293 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_125_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_36_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13457_ clknet_leaf_99_clk _00774_ net165 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.fin_quo\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_10669_ genblk2\[5\].wave_shpr.div.quo\[10\] _04858_ _04855_ net310 _04860_ vssd1
+ vssd1 vccd1 vccd1 _00553_ sky130_fd_sc_hd__a221o_1
XANTENNA__11549__C1 _05472_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08841__B _03544_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12408_ genblk2\[11\].wave_shpr.div.acc\[14\] _06078_ _06055_ vssd1 vssd1 vccd1 vccd1
+ _06079_ sky130_fd_sc_hd__mux2_1
X_13388_ clknet_leaf_78_clk _00707_ net208 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.b1\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_23_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12339_ net434 _03942_ _03941_ net438 _06027_ vssd1 vssd1 vccd1 vccd1 _01056_ sky130_fd_sc_hd__a221o_1
XANTENNA__06361__B _01226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_121_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06900_ _01753_ genblk1\[6\].osc.clkdiv_C.cnt\[0\] _01363_ genblk1\[6\].osc.clkdiv_C.cnt\[15\]
+ genblk1\[6\].osc.clkdiv_C.cnt\[17\] vssd1 vssd1 vccd1 vccd1 _01754_ sky130_fd_sc_hd__a221o_1
X_07880_ _02424_ _02471_ _02519_ vssd1 vssd1 vccd1 vccd1 _02587_ sky130_fd_sc_hd__o21a_1
X_06831_ genblk1\[5\].osc.clkdiv_C.cnt\[3\] _01698_ vssd1 vssd1 vccd1 vccd1 _01700_
+ sky130_fd_sc_hd__and2_1
X_09550_ _04055_ genblk1\[1\].osc.clkdiv_C.cnt\[13\] vssd1 vssd1 vccd1 vccd1 _04066_
+ sky130_fd_sc_hd__and2_1
X_06762_ genblk1\[4\].osc.clkdiv_C.cnt\[12\] _01637_ vssd1 vssd1 vccd1 vccd1 _01640_
+ sky130_fd_sc_hd__or2_1
X_08501_ net24 _03207_ vssd1 vssd1 vccd1 vccd1 _03208_ sky130_fd_sc_hd__or2b_1
X_09481_ _04029_ vssd1 vssd1 vccd1 vccd1 _00196_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_144_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06693_ genblk1\[4\].osc.clkdiv_C.cnt\[11\] _01313_ _01340_ genblk1\[4\].osc.clkdiv_C.cnt\[8\]
+ vssd1 vssd1 vccd1 vccd1 _01583_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_53_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08432_ _03137_ _03138_ genblk2\[9\].wave_shpr.div.fin_quo\[3\] _02308_ vssd1 vssd1
+ vccd1 vccd1 _03139_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12029__B1 _05817_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08363_ _02939_ _03069_ _02943_ vssd1 vssd1 vccd1 vccd1 _03070_ sky130_fd_sc_hd__o21a_1
XFILLER_0_19_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_901 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout143_A net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07314_ genblk1\[11\].osc.clkdiv_C.cnt\[12\] _02077_ genblk1\[11\].osc.clkdiv_C.cnt\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02078_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_34_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_731 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08294_ _02998_ _02999_ _03000_ vssd1 vssd1 vccd1 vccd1 _03001_ sky130_fd_sc_hd__nor3_1
XFILLER_0_46_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12638__RESET_B net109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07245_ _02026_ vssd1 vssd1 vccd1 vccd1 _02027_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_280 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08751__B _02467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07176_ genblk1\[9\].osc.clkdiv_C.cnt\[7\] _01967_ vssd1 vssd1 vccd1 vccd1 _01969_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06127_ _01098_ vssd1 vssd1 vccd1 vccd1 _01099_ sky130_fd_sc_hd__buf_2
XFILLER_0_2_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_100_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11307__A2 _05279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09074__S _03722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09817_ net553 _04257_ _04251_ genblk2\[2\].wave_shpr.div.quo\[11\] _04258_ vssd1
+ vssd1 vccd1 vccd1 _00303_ sky130_fd_sc_hd__a221o_1
X_09748_ _04221_ vssd1 vssd1 vccd1 vccd1 _00271_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_69_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout56_A net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2003 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10818__A1 _04855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2014 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2025 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09679_ genblk2\[2\].wave_shpr.div.acc\[14\] genblk2\[2\].wave_shpr.div.b1\[14\]
+ vssd1 vssd1 vccd1 vccd1 _04159_ sky130_fd_sc_hd__or2b_1
XTAP_2036 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2047 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2058 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11710_ genblk2\[9\].wave_shpr.div.b1\[15\] genblk2\[9\].wave_shpr.div.acc\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05602_ sky130_fd_sc_hd__and2b_1
XTAP_1324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2069 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12690_ clknet_leaf_53_clk genblk1\[8\].osc.clkdiv_C.next_cnt\[3\] net174 vssd1 vssd1
+ vccd1 vccd1 genblk1\[8\].osc.clkdiv_C.cnt\[3\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_hold522_A genblk2\[10\].wave_shpr.div.quo\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_139_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11641_ genblk2\[8\].wave_shpr.div.acc\[23\] _05412_ _05540_ vssd1 vssd1 vccd1 vccd1
+ _05541_ sky130_fd_sc_hd__a21o_1
XTAP_1379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11572_ genblk2\[8\].wave_shpr.div.acc\[5\] _05489_ _05417_ vssd1 vssd1 vccd1 vccd1
+ _05490_ sky130_fd_sc_hd__mux2_1
XFILLER_0_37_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13311_ clknet_leaf_118_clk net721 net137 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_91_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10523_ genblk2\[4\].wave_shpr.div.i\[1\] genblk2\[4\].wave_shpr.div.i\[0\] vssd1
+ vssd1 vccd1 vccd1 _04755_ sky130_fd_sc_hd__or2_1
XFILLER_0_150_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13242_ clknet_leaf_9_clk net246 net55 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.quo\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10454_ net891 _04683_ _04690_ _04705_ vssd1 vssd1 vccd1 vccd1 _00493_ sky130_fd_sc_hd__a22o_1
XANTENNA__06462__A genblk1\[1\].osc.clkdiv_C.cnt\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11546__A2 _05441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13173_ clknet_leaf_128_clk _00498_ net66 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.acc\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10385_ _04477_ genblk1\[4\].osc.clkdiv_C.cnt\[2\] vssd1 vssd1 vccd1 vccd1 _04660_
+ sky130_fd_sc_hd__and2_1
X_12124_ _05769_ _05880_ vssd1 vssd1 vccd1 vccd1 _05881_ sky130_fd_sc_hd__xnor2_1
XANTENNA__06973__A2 _01363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12055_ _05819_ genblk1\[10\].osc.clkdiv_C.cnt\[10\] vssd1 vssd1 vccd1 vccd1 _05832_
+ sky130_fd_sc_hd__and2_1
X_11006_ _05054_ vssd1 vssd1 vccd1 vccd1 _05093_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12957_ clknet_leaf_114_clk _00286_ net132 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.b1\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11482__A1 _02656_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11908_ net273 _05729_ _05730_ vssd1 vssd1 vccd1 vccd1 _00922_ sky130_fd_sc_hd__a21oi_1
XTAP_2570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_59_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12888_ clknet_leaf_30_clk _00219_ net96 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.quo\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07150__A2 _01799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09013__A _02171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11839_ _05594_ _05560_ vssd1 vssd1 vccd1 vccd1 _05681_ sky130_fd_sc_hd__or2b_1
XFILLER_0_145_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_117_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_353 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13509_ clknet_leaf_80_clk _00826_ net205 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.acc\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07030_ genblk1\[7\].osc.clkdiv_C.cnt\[16\] _01847_ vssd1 vssd1 vccd1 vccd1 _01850_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__07468__A _02147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_2_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08402__A2 _01411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08981_ _03525_ _03568_ _03569_ vssd1 vssd1 vccd1 vccd1 _03666_ sky130_fd_sc_hd__and3_1
X_07932_ genblk2\[8\].wave_shpr.div.fin_quo\[0\] genblk2\[8\].wave_shpr.div.fin_quo\[1\]
+ genblk2\[8\].wave_shpr.div.fin_quo\[2\] vssd1 vssd1 vccd1 vccd1 _02639_ sky130_fd_sc_hd__or3_1
X_07863_ _02469_ _02569_ _02529_ vssd1 vssd1 vccd1 vccd1 _02570_ sky130_fd_sc_hd__o21a_1
XANTENNA__07913__A1 genblk1\[8\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09602_ _03990_ _03961_ vssd1 vssd1 vccd1 vccd1 _04103_ sky130_fd_sc_hd__or2b_1
X_06814_ genblk1\[5\].osc.clkdiv_C.cnt\[6\] _01242_ _01682_ _01683_ _01685_ vssd1
+ vssd1 vccd1 vccd1 _01686_ sky130_fd_sc_hd__a221o_1
X_07794_ _02478_ _02492_ _02495_ _02500_ vssd1 vssd1 vccd1 vccd1 _02501_ sky130_fd_sc_hd__or4b_1
XANTENNA__09622__S _04095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07931__A net30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09533_ _04055_ genblk1\[1\].osc.clkdiv_C.cnt\[5\] vssd1 vssd1 vccd1 vccd1 _04057_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06745_ genblk1\[4\].osc.clkdiv_C.cnt\[8\] genblk1\[4\].osc.clkdiv_C.cnt\[7\] _01620_
+ vssd1 vssd1 vccd1 vccd1 _01627_ sky130_fd_sc_hd__and3_1
Xwire32 _02302_ vssd1 vssd1 vccd1 vccd1 net32 sky130_fd_sc_hd__clkbuf_2
XANTENNA__09666__A1 _04045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09464_ genblk2\[2\].wave_shpr.div.b1\[0\] net35 _03822_ vssd1 vssd1 vccd1 vccd1
+ _04020_ sky130_fd_sc_hd__mux2_1
XANTENNA__11473__A1 _04230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06676_ genblk1\[4\].osc.clkdiv_C.cnt\[5\] _01565_ vssd1 vssd1 vccd1 vccd1 _01566_
+ sky130_fd_sc_hd__and2_1
X_08415_ net8 _02744_ _02365_ vssd1 vssd1 vccd1 vccd1 _03122_ sky130_fd_sc_hd__and3_2
XFILLER_0_65_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09395_ genblk2\[1\].wave_shpr.div.acc\[12\] genblk2\[1\].wave_shpr.div.b1\[12\]
+ vssd1 vssd1 vccd1 vccd1 _03959_ sky130_fd_sc_hd__or2b_1
XFILLER_0_80_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_148_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08346_ _02993_ _02994_ _02995_ vssd1 vssd1 vccd1 vccd1 _03053_ sky130_fd_sc_hd__a21o_1
XFILLER_0_80_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08277_ _02977_ _02983_ vssd1 vssd1 vccd1 vccd1 _02984_ sky130_fd_sc_hd__and2b_1
XFILLER_0_117_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_15_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10984__B1 _05054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07228_ genblk1\[10\].osc.clkdiv_C.cnt\[7\] _01235_ _01227_ genblk1\[10\].osc.clkdiv_C.cnt\[9\]
+ vssd1 vssd1 vccd1 vccd1 _02010_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_132_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_120_907 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07159_ _01957_ vssd1 vssd1 vccd1 vccd1 genblk1\[9\].osc.clkdiv_C.next_cnt\[1\] sky130_fd_sc_hd__clkbuf_1
XANTENNA__07062__D1 genblk1\[8\].osc.clkdiv_C.cnt\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10170_ _04395_ _04370_ vssd1 vssd1 vccd1 vccd1 _04505_ sky130_fd_sc_hd__or2b_1
Xfanout130 net131 vssd1 vssd1 vccd1 vccd1 net130 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10532__A _03690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout141 net145 vssd1 vssd1 vccd1 vccd1 net141 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xfanout152 net158 vssd1 vssd1 vccd1 vccd1 net152 sky130_fd_sc_hd__clkbuf_4
Xfanout163 net171 vssd1 vssd1 vccd1 vccd1 net163 sky130_fd_sc_hd__clkbuf_2
Xfanout174 net218 vssd1 vssd1 vccd1 vccd1 net174 sky130_fd_sc_hd__buf_2
Xfanout185 net218 vssd1 vssd1 vccd1 vccd1 net185 sky130_fd_sc_hd__clkbuf_2
XANTENNA__13260__RESET_B net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06707__A2 _01304_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout196 net198 vssd1 vssd1 vccd1 vccd1 net196 sky130_fd_sc_hd__clkbuf_4
X_12811_ clknet_leaf_59_clk _00144_ net192 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.quo\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1110 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11464__A1 net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07668__B1 _02013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_1121 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12742_ clknet_leaf_50_clk genblk1\[11\].osc.clkdiv_C.next_cnt\[1\] net108 vssd1
+ vssd1 vccd1 vccd1 genblk1\[11\].osc.clkdiv_C.cnt\[1\] sky130_fd_sc_hd__dfrtp_4
XTAP_1132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12673_ clknet_leaf_90_clk genblk1\[7\].osc.clkdiv_C.next_cnt\[4\] net173 vssd1 vssd1
+ vccd1 vccd1 genblk1\[7\].osc.clkdiv_C.cnt\[4\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_38_843 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11624_ _05409_ _05416_ vssd1 vssd1 vccd1 vccd1 _05529_ sky130_fd_sc_hd__nand2b_1
XFILLER_0_92_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11555_ _05417_ _05476_ vssd1 vssd1 vccd1 vccd1 _05477_ sky130_fd_sc_hd__nand2_1
XANTENNA__08391__B _01302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06904__B _01757_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10506_ genblk2\[4\].wave_shpr.div.acc\[20\] _04740_ vssd1 vssd1 vccd1 vccd1 _04744_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_52_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_378 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11486_ _03831_ net390 _03717_ vssd1 vssd1 vccd1 vccd1 _00792_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_80_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_553 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13225_ clknet_leaf_114_clk _00548_ net133 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10437_ genblk2\[4\].wave_shpr.div.acc\[3\] _04692_ _04623_ vssd1 vssd1 vccd1 vccd1
+ _04693_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13156_ clknet_leaf_121_clk net666 net78 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.quo\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_905 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10368_ _04653_ vssd1 vssd1 vccd1 vccd1 _04654_ sky130_fd_sc_hd__clkbuf_4
XTAP_916 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12107_ _05761_ _05867_ vssd1 vssd1 vccd1 vccd1 _05868_ sky130_fd_sc_hd__xnor2_1
XTAP_927 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_938 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13087_ clknet_leaf_136_clk _00414_ net42 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.acc\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_949 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10299_ _04568_ _04609_ _04610_ vssd1 vssd1 vccd1 vccd1 _04611_ sky130_fd_sc_hd__a21o_1
X_12038_ net223 _05818_ _05816_ net398 _05822_ vssd1 vssd1 vccd1 vccd1 _00960_ sky130_fd_sc_hd__a221o_1
XFILLER_0_18_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06530_ genblk1\[2\].osc.clkdiv_C.cnt\[2\] genblk1\[2\].osc.clkdiv_C.cnt\[1\] genblk1\[2\].osc.clkdiv_C.cnt\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01454_ sky130_fd_sc_hd__and3_1
XANTENNA__07470__B _02153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_629 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12912__RESET_B net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08320__B2 _02362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_75_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06461_ _01373_ _01394_ _01395_ vssd1 vssd1 vccd1 vccd1 genblk1\[1\].osc.clkdiv_C.next_cnt\[9\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_146_837 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08200_ _02405_ _02403_ _02410_ _02524_ vssd1 vssd1 vccd1 vccd1 _02907_ sky130_fd_sc_hd__o31a_1
XFILLER_0_145_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_118_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09180_ net1249 _01356_ _03722_ vssd1 vssd1 vccd1 vccd1 _03817_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_90_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06392_ _01179_ vssd1 vssd1 vccd1 vccd1 _01336_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_50_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08131_ _02221_ _02837_ vssd1 vssd1 vccd1 vccd1 _02838_ sky130_fd_sc_hd__nor2_2
XFILLER_0_50_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_114_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10617__A _03701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08062_ _02766_ _02768_ vssd1 vssd1 vccd1 vccd1 _02769_ sky130_fd_sc_hd__nand2_1
XANTENNA__07831__B1 _02224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07013_ genblk1\[7\].osc.clkdiv_C.cnt\[10\] _01837_ _01822_ vssd1 vssd1 vccd1 vccd1
+ _01839_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_732 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_789 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_fanout106_A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07595__C1 genblk1\[9\].osc.clkdiv_C.cnt\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08964_ _03651_ _03646_ _03506_ vssd1 vssd1 vccd1 vccd1 _03652_ sky130_fd_sc_hd__a21oi_1
X_07915_ genblk1\[8\].osc.clkdiv_C.cnt\[3\] _01866_ _01487_ genblk1\[8\].osc.clkdiv_C.cnt\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02622_ sky130_fd_sc_hd__a22o_1
X_08895_ net629 _03596_ vssd1 vssd1 vccd1 vccd1 _03600_ sky130_fd_sc_hd__or2_1
X_07846_ _02552_ vssd1 vssd1 vccd1 vccd1 _02553_ sky130_fd_sc_hd__clkbuf_2
XANTENNA__07898__B1 _01576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07777_ genblk1\[0\].osc.clkdiv_C.cnt\[4\] _01258_ vssd1 vssd1 vccd1 vccd1 _02484_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_67_905 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09516_ net292 _04043_ _04047_ net771 vssd1 vssd1 vccd1 vccd1 _00213_ sky130_fd_sc_hd__a22o_1
X_06728_ genblk1\[4\].osc.clkdiv_C.cnt\[4\] _01609_ vssd1 vssd1 vccd1 vccd1 _01614_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_78_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09447_ _04010_ vssd1 vssd1 vccd1 vccd1 _04011_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_66_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06659_ _01522_ _01551_ vssd1 vssd1 vccd1 vccd1 _01552_ sky130_fd_sc_hd__nor2_1
XPHY_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_149_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09378_ genblk2\[11\].wave_shpr.div.i\[1\] genblk2\[11\].wave_shpr.div.i\[0\] vssd1
+ vssd1 vccd1 vccd1 _03946_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_19_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11749__A2 _05623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08329_ genblk2\[7\].wave_shpr.div.fin_quo\[4\] vssd1 vssd1 vccd1 vccd1 _03036_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_323 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08075__B1 _01726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11340_ genblk2\[7\].wave_shpr.div.acc\[17\] _05329_ _05300_ vssd1 vssd1 vccd1 vccd1
+ _05330_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11271_ _05184_ _05276_ vssd1 vssd1 vccd1 vccd1 _05277_ sky130_fd_sc_hd__nor2_1
X_13010_ clknet_leaf_133_clk _00339_ net59 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.acc\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10222_ _04543_ _04544_ vssd1 vssd1 vccd1 vccd1 _04545_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10153_ genblk2\[3\].wave_shpr.div.acc\[3\] _04492_ _04420_ vssd1 vssd1 vccd1 vccd1
+ _04493_ sky130_fd_sc_hd__mux2_1
X_10084_ _04453_ vssd1 vssd1 vccd1 vccd1 _04454_ sky130_fd_sc_hd__buf_4
Xhold8 genblk2\[9\].wave_shpr.div.quo\[22\] vssd1 vssd1 vccd1 vccd1 net226 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10488__A2 _04715_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07571__A genblk1\[9\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06187__A _01157_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10986_ net283 _05051_ _05054_ net668 _05078_ vssd1 vssd1 vccd1 vccd1 _00652_ sky130_fd_sc_hd__a221o_1
X_13774_ clknet_leaf_73_clk _01085_ net213 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.acc\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12725_ clknet_leaf_37_clk genblk1\[10\].osc.clkdiv_C.next_cnt\[2\] net113 vssd1
+ vssd1 vccd1 vccd1 genblk1\[10\].osc.clkdiv_C.cnt\[2\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_155_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10660__A2 _04853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12656_ clknet_leaf_27_clk genblk1\[6\].osc.clkdiv_C.next_cnt\[5\] net90 vssd1 vssd1
+ vccd1 vccd1 genblk1\[6\].osc.clkdiv_C.cnt\[5\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_154_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_707 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_846 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_509 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08066__B1 _01171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11607_ net846 _05507_ _05484_ _05516_ vssd1 vssd1 vccd1 vccd1 _00835_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12587_ clknet_leaf_14_clk genblk1\[2\].osc.clkdiv_C.next_cnt\[8\] net72 vssd1 vssd1
+ vccd1 vccd1 genblk1\[2\].osc.clkdiv_C.cnt\[8\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_154_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11538_ net575 _05454_ _05458_ net660 _05466_ vssd1 vssd1 vccd1 vccd1 _00816_ sky130_fd_sc_hd__a221o_1
XFILLER_0_41_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xhold408 genblk2\[4\].wave_shpr.div.quo\[20\] vssd1 vssd1 vccd1 vccd1 net626 sky130_fd_sc_hd__dlygate4sd3_1
Xhold419 genblk2\[4\].wave_shpr.div.quo\[13\] vssd1 vssd1 vccd1 vccd1 net637 sky130_fd_sc_hd__dlygate4sd3_1
X_11469_ _05431_ vssd1 vssd1 vccd1 vccd1 _00782_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09566__B1 _04047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13208_ clknet_leaf_8_clk _00531_ net88 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.b1\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_110_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_489 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13139_ clknet_leaf_115_clk net750 net133 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1108 genblk2\[5\].wave_shpr.div.quo\[3\] vssd1 vssd1 vccd1 vccd1 net1326 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1119 genblk2\[8\].wave_shpr.div.quo\[2\] vssd1 vssd1 vccd1 vccd1 net1337 sky130_fd_sc_hd__dlygate4sd3_1
X_07700_ genblk2\[10\].wave_shpr.div.fin_quo\[0\] genblk2\[10\].wave_shpr.div.fin_quo\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02407_ sky130_fd_sc_hd__nor2_1
X_08680_ _03307_ _03330_ _03328_ vssd1 vssd1 vccd1 vccd1 _03387_ sky130_fd_sc_hd__a21oi_1
XANTENNA__08541__A1 genblk2\[8\].wave_shpr.div.fin_quo\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_136_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08541__B2 genblk2\[8\].wave_shpr.div.fin_quo\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_07631_ _02128_ _01179_ _01249_ vssd1 vssd1 vccd1 vccd1 _02338_ sky130_fd_sc_hd__or3_1
XFILLER_0_45_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07562_ genblk1\[9\].osc.clkdiv_C.cnt\[11\] _01799_ _01731_ _02268_ vssd1 vssd1 vccd1
+ vccd1 _02269_ sky130_fd_sc_hd__a2bb2o_1
X_09301_ _03803_ vssd1 vssd1 vccd1 vccd1 _03889_ sky130_fd_sc_hd__buf_4
XFILLER_0_75_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06513_ _01213_ vssd1 vssd1 vccd1 vccd1 _01439_ sky130_fd_sc_hd__buf_4
XFILLER_0_152_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07493_ modein.delay_in\[0\] vssd1 vssd1 vccd1 vccd1 _02215_ sky130_fd_sc_hd__inv_2
XFILLER_0_76_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_779 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09232_ net569 _03841_ _03839_ net598 _03843_ vssd1 vssd1 vccd1 vccd1 _00133_ sky130_fd_sc_hd__a221o_1
XFILLER_0_145_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06444_ _01374_ _01382_ _01383_ vssd1 vssd1 vccd1 vccd1 _01384_ sky130_fd_sc_hd__and3_1
XFILLER_0_152_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_645 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10545__B_N genblk2\[5\].wave_shpr.div.b1\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_8_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_29_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09163_ genblk2\[0\].wave_shpr.div.fin_quo\[3\] net1314 _00001_ vssd1 vssd1 vccd1
+ vccd1 _03808_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06375_ _01306_ _01315_ _01316_ _01318_ vssd1 vssd1 vccd1 vccd1 _01319_ sky130_fd_sc_hd__or4b_1
X_08114_ _02811_ _02820_ vssd1 vssd1 vccd1 vccd1 _02821_ sky130_fd_sc_hd__nand2_1
X_09094_ _01367_ _03739_ vssd1 vssd1 vccd1 vccd1 _03743_ sky130_fd_sc_hd__or2_1
XFILLER_0_43_175 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08072__A3 _01180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_337 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08045_ genblk1\[5\].osc.clkdiv_C.cnt\[13\] _01675_ _02748_ _02751_ vssd1 vssd1 vccd1
+ vccd1 _02752_ sky130_fd_sc_hd__a211o_1
Xhold920 genblk2\[6\].wave_shpr.div.acc\[20\] vssd1 vssd1 vccd1 vccd1 net1138 sky130_fd_sc_hd__dlygate4sd3_1
Xhold931 genblk2\[9\].wave_shpr.div.i\[2\] vssd1 vssd1 vccd1 vccd1 net1149 sky130_fd_sc_hd__dlygate4sd3_1
Xhold942 genblk2\[4\].wave_shpr.div.i\[3\] vssd1 vssd1 vccd1 vccd1 net1160 sky130_fd_sc_hd__dlygate4sd3_1
Xhold953 genblk2\[10\].wave_shpr.div.b1\[2\] vssd1 vssd1 vccd1 vccd1 net1171 sky130_fd_sc_hd__dlygate4sd3_1
Xhold964 genblk1\[8\].osc.clkdiv_C.cnt\[13\] vssd1 vssd1 vccd1 vccd1 net1182 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold975 genblk1\[3\].osc.clkdiv_C.cnt\[12\] vssd1 vssd1 vccd1 vccd1 net1193 sky130_fd_sc_hd__dlygate4sd3_1
Xhold986 genblk2\[11\].wave_shpr.div.b1\[10\] vssd1 vssd1 vccd1 vccd1 net1204 sky130_fd_sc_hd__dlygate4sd3_1
Xhold997 genblk2\[7\].wave_shpr.div.fin_quo\[7\] vssd1 vssd1 vccd1 vccd1 net1215 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10082__A _04451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09996_ _04372_ _04390_ _04391_ vssd1 vssd1 vccd1 vccd1 _04392_ sky130_fd_sc_hd__a21o_1
XFILLER_0_110_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07583__A2 _01234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08947_ _03557_ _03558_ _03546_ _03551_ vssd1 vssd1 vccd1 vccd1 _03638_ sky130_fd_sc_hd__o211a_1
XANTENNA_clkbuf_leaf_84_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11906__A _03690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08878_ _03576_ sig_norm.acc\[2\] _03583_ vssd1 vssd1 vccd1 vccd1 _03584_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07829_ _02530_ _02535_ vssd1 vssd1 vccd1 vccd1 _02536_ sky130_fd_sc_hd__nor2_1
X_10840_ genblk2\[6\].wave_shpr.div.b1\[1\] genblk2\[6\].wave_shpr.div.acc\[1\] vssd1
+ vssd1 vccd1 vccd1 _04984_ sky130_fd_sc_hd__or2b_1
XFILLER_0_67_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_99_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10771_ genblk2\[5\].wave_shpr.div.acc\[15\] _04930_ _04907_ vssd1 vssd1 vccd1 vccd1
+ _04931_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_66_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_82_705 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12510_ clknet_leaf_84_clk net1040 net202 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.i\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_136_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13490_ clknet_leaf_88_clk _00807_ net177 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.quo\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12441_ net1078 _03947_ _03944_ _06101_ vssd1 vssd1 vccd1 vccd1 _01084_ sky130_fd_sc_hd__a22o_1
XANTENNA_clkbuf_leaf_22_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_35_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12372_ _05952_ _06050_ vssd1 vssd1 vccd1 vccd1 _06051_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_23_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_849 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11323_ _05206_ _05316_ vssd1 vssd1 vccd1 vccd1 _05317_ sky130_fd_sc_hd__xnor2_1
Xclkbuf_4_0_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_0_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_105_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11254_ _05260_ genblk1\[7\].osc.clkdiv_C.cnt\[12\] vssd1 vssd1 vccd1 vccd1 _05267_
+ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_37_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06470__A genblk1\[1\].osc.clkdiv_C.cnt\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07559__C1 genblk1\[9\].osc.clkdiv_C.cnt\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_120_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10205_ _04411_ _04362_ vssd1 vssd1 vccd1 vccd1 _04532_ sky130_fd_sc_hd__nor2_1
XFILLER_0_120_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11185_ _03727_ _01432_ net593 _03687_ vssd1 vssd1 vccd1 vccd1 _00697_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__07574__A2 _01437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10136_ _03819_ net436 _00010_ genblk2\[3\].wave_shpr.div.acc\[0\] _04479_ vssd1
+ vssd1 vccd1 vccd1 _00401_ sky130_fd_sc_hd__o221a_1
XFILLER_0_100_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10067_ _04443_ vssd1 vssd1 vccd1 vccd1 _00368_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__11535__B genblk1\[8\].osc.clkdiv_C.cnt\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_309 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_58_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13757_ clknet_leaf_70_clk _01068_ net213 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.acc\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_136_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_136_clk
+ sky130_fd_sc_hd__clkbuf_16
X_10969_ net582 _05062_ _05064_ net595 _05069_ vssd1 vssd1 vccd1 vccd1 _00644_ sky130_fd_sc_hd__a221o_1
XANTENNA__10094__B1 _04456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12708_ clknet_leaf_56_clk genblk1\[9\].osc.clkdiv_C.next_cnt\[3\] net181 vssd1 vssd1
+ vccd1 vccd1 genblk1\[9\].osc.clkdiv_C.cnt\[3\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_73_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13688_ clknet_leaf_63_clk _01001_ net190 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.acc\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12639_ clknet_leaf_16_clk genblk1\[5\].osc.clkdiv_C.next_cnt\[6\] net73 vssd1 vssd1
+ vccd1 vccd1 genblk1\[5\].osc.clkdiv_C.cnt\[6\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_109_870 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_110_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_127_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06160_ _01117_ _01131_ vssd1 vssd1 vccd1 vccd1 _01132_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_5_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_130_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold205 genblk2\[5\].wave_shpr.div.quo\[8\] vssd1 vssd1 vccd1 vccd1 net423 sky130_fd_sc_hd__dlygate4sd3_1
Xhold216 genblk2\[11\].wave_shpr.div.quo\[23\] vssd1 vssd1 vccd1 vccd1 net434 sky130_fd_sc_hd__dlygate4sd3_1
Xhold227 genblk2\[8\].wave_shpr.div.quo\[24\] vssd1 vssd1 vccd1 vccd1 net445 sky130_fd_sc_hd__dlygate4sd3_1
Xhold238 genblk2\[8\].wave_shpr.div.acc\[22\] vssd1 vssd1 vccd1 vccd1 net456 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07476__A _02203_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold249 genblk2\[11\].wave_shpr.div.quo\[10\] vssd1 vssd1 vccd1 vccd1 net467 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_22_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09850_ genblk2\[2\].wave_shpr.div.b1\[0\] _04214_ genblk2\[2\].wave_shpr.div.acc\[0\]
+ vssd1 vssd1 vccd1 vccd1 _04277_ sky130_fd_sc_hd__a21oi_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_798 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07565__A2 _01328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08801_ _03451_ _03506_ _03507_ vssd1 vssd1 vccd1 vccd1 _03508_ sky130_fd_sc_hd__o21bai_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09781_ _04240_ vssd1 vssd1 vccd1 vccd1 _00285_ sky130_fd_sc_hd__clkbuf_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06993_ _01823_ _01825_ _01826_ vssd1 vssd1 vccd1 vccd1 genblk1\[7\].osc.clkdiv_C.next_cnt\[2\]
+ sky130_fd_sc_hd__nor3_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08732_ _03431_ _03438_ vssd1 vssd1 vccd1 vccd1 _03439_ sky130_fd_sc_hd__xnor2_1
X_08663_ genblk2\[5\].wave_shpr.div.fin_quo\[3\] _02521_ _02791_ _03369_ vssd1 vssd1
+ vccd1 vccd1 _03370_ sky130_fd_sc_hd__a211o_1
XANTENNA__07722__C1 _01172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07614_ _01171_ _01192_ _01208_ genblk1\[11\].osc.clkdiv_C.cnt\[3\] vssd1 vssd1 vccd1
+ vccd1 _02321_ sky130_fd_sc_hd__a31o_1
X_08594_ net10 _02364_ _03300_ vssd1 vssd1 vccd1 vccd1 _03301_ sky130_fd_sc_hd__and3_1
XTAP_1709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09630__S _04095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07545_ PWM.final_sample_in\[4\] net1150 PWM.start vssd1 vssd1 vccd1 vccd1 _02256_
+ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_127_clk clknet_4_2_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_127_clk
+ sky130_fd_sc_hd__clkbuf_16
XANTENNA__10085__B1 _04420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07476_ _02203_ vssd1 vssd1 vccd1 vccd1 _00022_ sky130_fd_sc_hd__inv_2
XFILLER_0_36_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_656 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_17_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11180__B genblk2\[8\].wave_shpr.div.b1\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06427_ _01335_ _01353_ _01357_ _01370_ vssd1 vssd1 vccd1 vccd1 _01371_ sky130_fd_sc_hd__or4b_1
X_09215_ _02152_ genblk2\[0\].wave_shpr.div.busy _02149_ vssd1 vssd1 vccd1 vccd1 _03837_
+ sky130_fd_sc_hd__and3_1
XFILLER_0_17_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09146_ _03748_ _03792_ _03793_ vssd1 vssd1 vccd1 vccd1 _03794_ sky130_fd_sc_hd__a21o_1
XANTENNA__09866__A _04250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09501__B1_N _03717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06358_ _01301_ vssd1 vssd1 vccd1 vccd1 _01302_ sky130_fd_sc_hd__buf_6
XFILLER_0_16_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09077_ _03731_ vssd1 vssd1 vccd1 vccd1 _00090_ sky130_fd_sc_hd__clkbuf_1
X_06289_ _01246_ _01250_ vssd1 vssd1 vccd1 vccd1 _01251_ sky130_fd_sc_hd__nand2_1
XFILLER_0_130_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_32_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08028_ genblk2\[6\].wave_shpr.div.fin_quo\[0\] genblk2\[6\].wave_shpr.div.fin_quo\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02735_ sky130_fd_sc_hd__or2_1
XFILLER_0_102_545 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold750 genblk2\[2\].wave_shpr.div.acc\[22\] vssd1 vssd1 vccd1 vccd1 net968 sky130_fd_sc_hd__dlygate4sd3_1
Xhold761 genblk2\[3\].wave_shpr.div.acc\[4\] vssd1 vssd1 vccd1 vccd1 net979 sky130_fd_sc_hd__dlygate4sd3_1
Xhold772 genblk2\[1\].wave_shpr.div.acc\[2\] vssd1 vssd1 vccd1 vccd1 net990 sky130_fd_sc_hd__dlygate4sd3_1
Xhold783 genblk2\[6\].wave_shpr.div.acc\[21\] vssd1 vssd1 vccd1 vccd1 net1001 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold794 genblk2\[5\].wave_shpr.div.acc\[23\] vssd1 vssd1 vccd1 vccd1 net1012 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11888__A1 _03694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout86_A net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09950__B1 _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09979_ genblk2\[3\].wave_shpr.div.acc\[4\] genblk2\[3\].wave_shpr.div.b1\[4\] vssd1
+ vssd1 vccd1 vccd1 _04375_ sky130_fd_sc_hd__or2b_1
X_12990_ clknet_leaf_131_clk _00319_ net65 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.acc\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07308__A2 _01513_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12301__A2 _06009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11941_ _05740_ _05761_ _05762_ vssd1 vssd1 vccd1 vccd1 _05763_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11872_ net1023 _05684_ _05685_ _05706_ vssd1 vssd1 vccd1 vccd1 _00910_ sky130_fd_sc_hd__a22o_1
X_13611_ clknet_leaf_93_clk _00924_ net159 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.fin_quo\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_39_234 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10823_ genblk2\[6\].wave_shpr.div.b1\[16\] genblk2\[6\].wave_shpr.div.acc\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04967_ sky130_fd_sc_hd__xor2_1
Xclkbuf_leaf_118_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_118_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_95_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_109_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_55_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13542_ clknet_leaf_101_clk _00857_ net165 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.fin_quo\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10754_ net1014 _04886_ _04890_ _04917_ vssd1 vssd1 vccd1 vccd1 _00581_ sky130_fd_sc_hd__a22o_1
XANTENNA__06465__A genblk1\[1\].osc.clkdiv_C.cnt\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_109_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_70_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10685_ _04869_ genblk1\[5\].osc.clkdiv_C.cnt\[8\] vssd1 vssd1 vccd1 vccd1 _04870_
+ sky130_fd_sc_hd__and2_1
X_13473_ clknet_leaf_74_clk _00790_ net215 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.b1\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06184__B _01095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12424_ _06089_ _06090_ vssd1 vssd1 vccd1 vccd1 _06091_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_124_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08441__B1 _02361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12355_ genblk2\[11\].wave_shpr.div.acc\[2\] _06037_ _05982_ vssd1 vssd1 vccd1 vccd1
+ _06038_ sky130_fd_sc_hd__mux2_1
X_11306_ genblk2\[7\].wave_shpr.div.acc\[9\] _05303_ _05300_ vssd1 vssd1 vccd1 vccd1
+ _05304_ sky130_fd_sc_hd__mux2_1
X_12286_ _03726_ _01312_ _06004_ vssd1 vssd1 vccd1 vccd1 _01026_ sky130_fd_sc_hd__a21oi_1
X_11237_ _05074_ genblk1\[7\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 _05258_
+ sky130_fd_sc_hd__and2_1
X_11168_ _05225_ vssd1 vssd1 vccd1 vccd1 _00687_ sky130_fd_sc_hd__clkbuf_1
X_10119_ net451 _04461_ _04462_ genblk2\[3\].wave_shpr.div.quo\[17\] _04470_ vssd1
+ vssd1 vccd1 vccd1 _00393_ sky130_fd_sc_hd__a221o_1
X_11099_ _00016_ _05159_ net1177 vssd1 vssd1 vccd1 vccd1 _05161_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09016__A _02155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11500__B1 _05446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_77_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09450__S _00007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10596__S _00015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_109_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_109_clk
+ sky130_fd_sc_hd__clkbuf_16
X_07330_ _02093_ vssd1 vssd1 vccd1 vccd1 genblk1\[11\].osc.clkdiv_C.next_cnt\[0\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_45_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07261_ _02038_ vssd1 vssd1 vccd1 vccd1 genblk1\[10\].osc.clkdiv_C.next_cnt\[4\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_143_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09000_ net1102 net1126 _01154_ vssd1 vssd1 vccd1 vccd1 _03680_ sky130_fd_sc_hd__mux2_1
XFILLER_0_116_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06212_ _01173_ vssd1 vssd1 vccd1 vccd1 _01174_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_143_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_345 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07192_ _01953_ _01979_ vssd1 vssd1 vccd1 vccd1 _01980_ sky130_fd_sc_hd__nor2_1
XANTENNA__09224__A2 _03836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_115_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06143_ net14 _01112_ vssd1 vssd1 vccd1 vccd1 _01115_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_13_145 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07918__B genblk1\[8\].osc.clkdiv_C.cnt\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_41_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09902_ _04196_ _04316_ vssd1 vssd1 vccd1 vccd1 _04317_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_1_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_53 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09833_ _04069_ genblk1\[2\].osc.clkdiv_C.cnt\[11\] vssd1 vssd1 vccd1 vccd1 _04267_
+ sky130_fd_sc_hd__and2_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09764_ net1245 _01794_ _04039_ vssd1 vssd1 vccd1 vccd1 _04232_ sky130_fd_sc_hd__mux2_1
X_06976_ genblk1\[7\].osc.clkdiv_C.cnt\[12\] _01811_ vssd1 vssd1 vccd1 vccd1 _01812_
+ sky130_fd_sc_hd__xnor2_1
X_08715_ _03383_ _03395_ _03420_ _03421_ vssd1 vssd1 vccd1 vccd1 _03422_ sky130_fd_sc_hd__a211o_1
XANTENNA__12295__A1 _03687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09695_ genblk2\[2\].wave_shpr.div.acc\[0\] genblk2\[2\].wave_shpr.div.b1\[0\] vssd1
+ vssd1 vccd1 vccd1 _04175_ sky130_fd_sc_hd__and2b_1
XTAP_2207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08646_ _03140_ _03150_ vssd1 vssd1 vccd1 vccd1 _03353_ sky130_fd_sc_hd__xor2_1
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07171__B1 genblk1\[9\].osc.clkdiv_C.cnt\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07710__A2 _02362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08577_ _03141_ _03283_ _02901_ vssd1 vssd1 vccd1 vccd1 _03284_ sky130_fd_sc_hd__o21a_1
XANTENNA__12287__A _01337_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07528_ sig_norm.busy sig_norm.i\[0\] sig_norm.i\[1\] vssd1 vssd1 vccd1 vccd1 _02246_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07459_ _02190_ genblk2\[7\].wave_shpr.div.i\[1\] genblk2\[7\].wave_shpr.div.i\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02191_ sky130_fd_sc_hd__or3b_1
X_10470_ genblk2\[4\].wave_shpr.div.acc\[11\] _04717_ _04704_ vssd1 vssd1 vccd1 vccd1
+ _04718_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09129_ genblk2\[0\].wave_shpr.div.b1\[7\] genblk2\[0\].wave_shpr.div.acc\[7\] vssd1
+ vssd1 vccd1 vccd1 _03777_ sky130_fd_sc_hd__and2b_1
X_12140_ _05778_ _05732_ vssd1 vssd1 vccd1 vccd1 _05893_ sky130_fd_sc_hd__nor2_1
XFILLER_0_20_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_103_854 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_130_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12071_ _03719_ genblk1\[10\].osc.clkdiv_C.cnt\[17\] vssd1 vssd1 vccd1 vccd1 _05841_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_4_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold580 _00747_ vssd1 vssd1 vccd1 vccd1 net798 sky130_fd_sc_hd__dlygate4sd3_1
Xhold591 genblk2\[7\].wave_shpr.div.acc\[15\] vssd1 vssd1 vccd1 vccd1 net809 sky130_fd_sc_hd__dlygate4sd3_1
X_11022_ genblk2\[6\].wave_shpr.div.acc\[7\] _05104_ _05105_ vssd1 vssd1 vccd1 vccd1
+ _05106_ sky130_fd_sc_hd__mux2_1
XANTENNA_hold934_A genblk2\[3\].wave_shpr.div.b1\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11089__A2 _05057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12286__A1 _03726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12973_ clknet_leaf_124_clk net442 net71 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.quo\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11924_ genblk2\[10\].wave_shpr.div.acc\[1\] genblk2\[10\].wave_shpr.div.b1\[1\]
+ vssd1 vssd1 vccd1 vccd1 _05746_ sky130_fd_sc_hd__xnor2_1
XTAP_2730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11855_ genblk2\[9\].wave_shpr.div.acc\[14\] _05693_ _05673_ vssd1 vssd1 vccd1 vccd1
+ _05694_ sky130_fd_sc_hd__mux2_1
XFILLER_0_129_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08394__B _01411_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_716 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10806_ net392 _04858_ _04855_ _04955_ vssd1 vssd1 vccd1 vccd1 _00595_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11786_ genblk2\[9\].wave_shpr.div.quo\[23\] _02203_ _03693_ net226 _05642_ vssd1
+ vssd1 vccd1 vccd1 _00888_ sky130_fd_sc_hd__a221o_1
XFILLER_0_144_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13525_ clknet_leaf_98_clk _00842_ net169 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.acc\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10737_ net927 _04886_ _04890_ _04904_ vssd1 vssd1 vccd1 vccd1 _00577_ sky130_fd_sc_hd__a22o_1
XANTENNA__11261__A2 _05245_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_83_888 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13456_ clknet_leaf_100_clk _00773_ net164 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.fin_quo\[4\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_36_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10668_ _04672_ genblk1\[5\].osc.clkdiv_C.cnt\[1\] vssd1 vssd1 vccd1 vccd1 _04860_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_113_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_253 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_140_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12407_ _05968_ _06077_ vssd1 vssd1 vccd1 vccd1 _06078_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07738__B _02013_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07217__B2 _01342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10599_ _04824_ vssd1 vssd1 vccd1 vccd1 _00519_ sky130_fd_sc_hd__clkbuf_1
X_13387_ clknet_leaf_83_clk _00706_ net200 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.b1\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_112_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_774 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12338_ _03833_ _02081_ vssd1 vssd1 vccd1 vccd1 _06027_ sky130_fd_sc_hd__nor2_1
XFILLER_0_121_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12269_ _05995_ vssd1 vssd1 vccd1 vccd1 _01018_ sky130_fd_sc_hd__clkbuf_1
X_06830_ _01693_ _01698_ _01699_ vssd1 vssd1 vccd1 vccd1 genblk1\[5\].osc.clkdiv_C.next_cnt\[2\]
+ sky130_fd_sc_hd__nor3_1
X_06761_ _01639_ vssd1 vssd1 vccd1 vccd1 genblk1\[4\].osc.clkdiv_C.next_cnt\[11\]
+ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12277__A1 _02001_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08500_ _02520_ _02587_ _03206_ vssd1 vssd1 vccd1 vccd1 _03207_ sky130_fd_sc_hd__o21ai_1
X_09480_ genblk2\[2\].wave_shpr.div.b1\[7\] _04028_ _04024_ vssd1 vssd1 vccd1 vccd1
+ _04029_ sky130_fd_sc_hd__mux2_1
X_06692_ _01562_ _01573_ _01579_ _01581_ vssd1 vssd1 vccd1 vccd1 _01582_ sky130_fd_sc_hd__or4b_1
XANTENNA__09180__S _03722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08431_ genblk2\[9\].wave_shpr.div.fin_quo\[2\] net32 _02262_ _02222_ vssd1 vssd1
+ vccd1 vccd1 _03138_ sky130_fd_sc_hd__a31o_1
XFILLER_0_59_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12029__B2 genblk2\[10\].wave_shpr.div.quo\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06900__B1 _01363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_19_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08362_ genblk2\[3\].wave_shpr.div.fin_quo\[5\] _02539_ _03068_ _02592_ vssd1 vssd1
+ vccd1 vccd1 _03069_ sky130_fd_sc_hd__a22o_1
XFILLER_0_58_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11788__B1 _03693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07313_ _01308_ _01439_ vssd1 vssd1 vccd1 vccd1 _02077_ sky130_fd_sc_hd__nand2_2
X_08293_ _02921_ _02997_ _02992_ _02996_ vssd1 vssd1 vccd1 vccd1 _03000_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_73_354 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_fanout136_A net171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_743 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07244_ _01990_ _01991_ _02009_ _02010_ _02025_ vssd1 vssd1 vccd1 vccd1 _02026_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_27_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07929__A _02221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_730 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07175_ _01953_ _01967_ _01968_ vssd1 vssd1 vccd1 vccd1 genblk1\[9\].osc.clkdiv_C.next_cnt\[6\]
+ sky130_fd_sc_hd__nor3_1
X_06126_ _01097_ vssd1 vssd1 vccd1 vccd1 _01098_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_14_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_41_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08708__B2 _02468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10802__B _04880_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09816_ _04058_ _01410_ vssd1 vssd1 vccd1 vccd1 _04258_ sky130_fd_sc_hd__nor2_1
X_09747_ genblk2\[2\].wave_shpr.div.fin_quo\[6\] genblk2\[2\].wave_shpr.div.quo\[5\]
+ _00009_ vssd1 vssd1 vccd1 vccd1 _04221_ sky130_fd_sc_hd__mux2_1
XANTENNA__12268__A1 _01589_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06959_ genblk1\[7\].osc.clkdiv_C.cnt\[0\] net34 genblk1\[7\].osc.clkdiv_C.cnt\[10\]
+ vssd1 vssd1 vccd1 vccd1 _01795_ sky130_fd_sc_hd__and3b_1
XTAP_2004 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2015 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09678_ genblk2\[2\].wave_shpr.div.acc\[15\] genblk2\[2\].wave_shpr.div.b1\[15\]
+ vssd1 vssd1 vccd1 vccd1 _04158_ sky130_fd_sc_hd__or2b_1
XTAP_2026 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2037 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout49_A net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2048 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2059 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08629_ _02734_ _02735_ genblk2\[6\].wave_shpr.div.fin_quo\[2\] vssd1 vssd1 vccd1
+ vccd1 _03336_ sky130_fd_sc_hd__a21oi_1
XTAP_1325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11640_ _05413_ _05416_ vssd1 vssd1 vccd1 vccd1 _05540_ sky130_fd_sc_hd__and2b_1
XFILLER_0_37_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11571_ _05488_ _05383_ vssd1 vssd1 vccd1 vccd1 _05489_ sky130_fd_sc_hd__xnor2_1
X_13310_ clknet_leaf_118_clk net272 net137 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.quo\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10522_ _04754_ vssd1 vssd1 vccd1 vccd1 _00512_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_24_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_847 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_713 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10453_ net1340 _04703_ _04704_ vssd1 vssd1 vccd1 vccd1 _04705_ sky130_fd_sc_hd__mux2_1
X_13241_ clknet_leaf_10_clk _00564_ net55 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.quo\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_122_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13172_ clknet_leaf_128_clk _00497_ net66 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.acc\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10384_ net672 _04657_ _04655_ genblk2\[4\].wave_shpr.div.quo\[9\] _04659_ vssd1
+ vssd1 vccd1 vccd1 _00469_ sky130_fd_sc_hd__a221o_1
XFILLER_0_32_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12123_ _05770_ _05736_ vssd1 vssd1 vccd1 vccd1 _05880_ sky130_fd_sc_hd__or2b_1
X_12054_ net518 _05823_ _05825_ net547 _05831_ vssd1 vssd1 vccd1 vccd1 _00967_ sky130_fd_sc_hd__a221o_1
X_11005_ net986 _05086_ _05056_ _05092_ vssd1 vssd1 vccd1 vccd1 _00657_ sky130_fd_sc_hd__a22o_1
XANTENNA__06186__A1 _01155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_88_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_87_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_99_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12956_ clknet_leaf_136_clk _00285_ net42 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.b1\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07135__B1 _01925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11543__B genblk1\[8\].osc.clkdiv_C.cnt\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11907_ net273 _05729_ _03855_ vssd1 vssd1 vccd1 vccd1 _05730_ sky130_fd_sc_hd__o21ai_1
XTAP_2560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12887_ clknet_leaf_30_clk _00218_ net96 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.quo\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_74_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11838_ net807 _05652_ _05653_ _05680_ vssd1 vssd1 vccd1 vccd1 _00902_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_126_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11769_ _05631_ genblk1\[9\].osc.clkdiv_C.cnt\[6\] vssd1 vssd1 vccd1 vccd1 _05634_
+ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_40_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_40_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_28_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13508_ clknet_leaf_79_clk _00825_ net205 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.acc\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_15_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_573 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13439_ clknet_leaf_94_clk _00758_ net162 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.acc\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_141_746 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_70_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08980_ _01157_ _03664_ _03665_ vssd1 vssd1 vccd1 vccd1 _00059_ sky130_fd_sc_hd__o21ai_1
X_07931_ net30 vssd1 vssd1 vccd1 vccd1 _02638_ sky130_fd_sc_hd__buf_2
XFILLER_0_48_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07862_ _02525_ _02567_ _02568_ _02361_ genblk2\[1\].wave_shpr.div.fin_quo\[2\] vssd1
+ vssd1 vccd1 vccd1 _02569_ sky130_fd_sc_hd__a32o_1
X_09601_ net813 _04076_ _04080_ _04102_ vssd1 vssd1 vccd1 vccd1 _00243_ sky130_fd_sc_hd__a22o_1
XANTENNA__07913__A2 _01309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06813_ genblk1\[5\].osc.clkdiv_C.cnt\[0\] _01684_ vssd1 vssd1 vccd1 vccd1 _01685_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_155_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07793_ _02496_ _02497_ _02498_ _02499_ vssd1 vssd1 vccd1 vccd1 _02500_ sky130_fd_sc_hd__and4_1
X_09532_ net519 _04052_ _04053_ net537 _04056_ vssd1 vssd1 vccd1 vccd1 _00220_ sky130_fd_sc_hd__a221o_1
X_06744_ _01626_ vssd1 vssd1 vccd1 vccd1 genblk1\[4\].osc.clkdiv_C.next_cnt\[7\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_97 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07126__B1 _01855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xwire33 _02348_ vssd1 vssd1 vccd1 vccd1 net33 sky130_fd_sc_hd__buf_2
XFILLER_0_148_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08746__C genblk2\[6\].wave_shpr.div.fin_quo\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_94_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09463_ _04019_ vssd1 vssd1 vccd1 vccd1 _00188_ sky130_fd_sc_hd__clkbuf_1
X_06675_ _01187_ _01564_ vssd1 vssd1 vccd1 vccd1 _01565_ sky130_fd_sc_hd__nand2_4
X_08414_ genblk2\[2\].wave_shpr.div.fin_quo\[7\] _02468_ _03120_ _02592_ vssd1 vssd1
+ vccd1 vccd1 _03121_ sky130_fd_sc_hd__a22o_1
X_09394_ genblk2\[1\].wave_shpr.div.acc\[13\] genblk2\[1\].wave_shpr.div.b1\[13\]
+ vssd1 vssd1 vccd1 vccd1 _03958_ sky130_fd_sc_hd__or2b_1
XFILLER_0_93_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_710 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_19_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08345_ _02993_ _02994_ _02995_ vssd1 vssd1 vccd1 vccd1 _03052_ sky130_fd_sc_hd__nand3_1
XANTENNA__11225__A2 _05246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_31_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_31_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_73_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08276_ _02416_ _02982_ _02419_ vssd1 vssd1 vccd1 vccd1 _02983_ sky130_fd_sc_hd__o21ai_2
XANTENNA__07659__A net3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07227_ genblk1\[10\].osc.clkdiv_C.cnt\[5\] _01992_ _02008_ vssd1 vssd1 vccd1 vccd1
+ _02009_ sky130_fd_sc_hd__o21a_1
XFILLER_0_131_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06282__B _01242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_116_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_131_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07158_ _01954_ _01955_ _01956_ vssd1 vssd1 vccd1 vccd1 _01957_ sky130_fd_sc_hd__and3_1
XFILLER_0_120_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_267 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_30_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06109_ _01089_ vssd1 vssd1 vccd1 vccd1 smpl_rt_clkdiv.clkDiv_inst.next_hzX sky130_fd_sc_hd__clkbuf_1
XANTENNA__07062__C1 _01490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_610 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07089_ net1185 _01897_ _01899_ vssd1 vssd1 vccd1 vccd1 genblk1\[8\].osc.clkdiv_C.next_cnt\[7\]
+ sky130_fd_sc_hd__a21oi_1
Xfanout120 net122 vssd1 vssd1 vccd1 vccd1 net120 sky130_fd_sc_hd__buf_2
XFILLER_0_100_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout131 net136 vssd1 vssd1 vccd1 vccd1 net131 sky130_fd_sc_hd__clkbuf_2
Xclkbuf_leaf_98_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_98_clk sky130_fd_sc_hd__clkbuf_16
Xfanout142 net145 vssd1 vssd1 vccd1 vccd1 net142 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08157__A2 _01361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout153 net155 vssd1 vssd1 vccd1 vccd1 net153 sky130_fd_sc_hd__clkbuf_4
Xfanout164 net165 vssd1 vssd1 vccd1 vccd1 net164 sky130_fd_sc_hd__clkbuf_4
Xfanout175 net176 vssd1 vssd1 vccd1 vccd1 net175 sky130_fd_sc_hd__clkbuf_4
Xfanout186 net188 vssd1 vssd1 vccd1 vccd1 net186 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08562__C1 genblk2\[7\].wave_shpr.div.fin_quo\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout197 net198 vssd1 vssd1 vccd1 vccd1 net197 sky130_fd_sc_hd__buf_2
X_12810_ clknet_leaf_59_clk net299 net187 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.quo\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_96_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1100 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_906 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12741_ clknet_leaf_49_clk genblk1\[11\].osc.clkdiv_C.next_cnt\[0\] net108 vssd1
+ vssd1 vccd1 vccd1 genblk1\[11\].osc.clkdiv_C.cnt\[0\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__08865__B1 _02248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1111 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1122 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12672_ clknet_leaf_90_clk genblk1\[7\].osc.clkdiv_C.next_cnt\[3\] net173 vssd1 vssd1
+ vccd1 vccd1 genblk1\[7\].osc.clkdiv_C.cnt\[3\] sky130_fd_sc_hd__dfrtp_2
XTAP_1166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_38_855 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11623_ net1222 _05507_ _05445_ _05528_ vssd1 vssd1 vccd1 vccd1 _00839_ sky130_fd_sc_hd__a22o_1
XFILLER_0_53_814 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_22_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_22_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_52_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11554_ _05374_ _05375_ vssd1 vssd1 vccd1 vccd1 _05476_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_25_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06473__A genblk1\[1\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10505_ net472 _04715_ _04722_ _04743_ vssd1 vssd1 vccd1 vccd1 _00506_ sky130_fd_sc_hd__a22o_1
XFILLER_0_122_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11485_ _03831_ net374 _03728_ vssd1 vssd1 vccd1 vccd1 _00791_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_100_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12177__B1 _05818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13224_ clknet_leaf_114_clk _00547_ net132 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.quo\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09784__A _01490_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10436_ _04588_ _04691_ vssd1 vssd1 vccd1 vccd1 _04692_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_61_891 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_20_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08396__A2 _01349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13155_ clknet_leaf_121_clk net627 net80 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.quo\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10367_ _02152_ genblk2\[4\].wave_shpr.div.busy _02175_ vssd1 vssd1 vccd1 vccd1 _04653_
+ sky130_fd_sc_hd__and3_1
XTAP_906 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_917 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12106_ _05762_ _05740_ vssd1 vssd1 vccd1 vccd1 _05867_ sky130_fd_sc_hd__or2b_1
XTAP_928 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13086_ clknet_leaf_136_clk net943 net42 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.acc\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10298_ genblk2\[4\].wave_shpr.div.b1\[14\] genblk2\[4\].wave_shpr.div.acc\[14\]
+ vssd1 vssd1 vccd1 vccd1 _04610_ sky130_fd_sc_hd__and2b_1
XTAP_939 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_89_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_89_clk sky130_fd_sc_hd__clkbuf_16
X_12037_ _05819_ genblk1\[10\].osc.clkdiv_C.cnt\[2\] vssd1 vssd1 vccd1 vccd1 _05822_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_109_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13388__RESET_B net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__13317__RESET_B net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09024__A _02203_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12939_ clknet_leaf_110_clk _00268_ net136 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.fin_quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10663__B1 _04857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06460_ genblk1\[1\].osc.clkdiv_C.cnt\[9\] _01392_ vssd1 vssd1 vccd1 vccd1 _01395_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_146_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_87_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_91_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_146_849 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06391_ genblk1\[1\].osc.clkdiv_C.cnt\[10\] _01334_ vssd1 vssd1 vccd1 vccd1 _01335_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_145_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_13_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_13_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_141_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_56_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08130_ _02819_ _02836_ genblk1\[4\].osc.clkdiv_C.cnt\[16\] genblk1\[4\].osc.clkdiv_C.cnt\[17\]
+ vssd1 vssd1 vccd1 vccd1 _02837_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_83_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09281__B1 _03840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_154_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08061_ genblk1\[5\].osc.clkdiv_C.cnt\[4\] net36 _02767_ vssd1 vssd1 vccd1 vccd1
+ _02768_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_113_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07012_ _01823_ _01837_ _01838_ vssd1 vssd1 vccd1 vccd1 genblk1\[7\].osc.clkdiv_C.next_cnt\[9\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_24_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09033__B1 _03702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_51_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07595__B1 genblk1\[9\].osc.clkdiv_C.cnt\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08963_ _03559_ _03563_ _03564_ vssd1 vssd1 vccd1 vccd1 _03651_ sky130_fd_sc_hd__a21o_1
XFILLER_0_11_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07914_ genblk1\[8\].osc.clkdiv_C.cnt\[3\] _01866_ _02619_ _01489_ _02620_ vssd1
+ vssd1 vccd1 vccd1 _02621_ sky130_fd_sc_hd__o221a_1
X_08894_ net629 _02260_ _03599_ vssd1 vssd1 vccd1 vccd1 _00039_ sky130_fd_sc_hd__a21o_1
X_07845_ net18 vssd1 vssd1 vccd1 vccd1 _02552_ sky130_fd_sc_hd__buf_2
XFILLER_0_75_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07898__B2 genblk1\[8\].osc.clkdiv_C.cnt\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07776_ _01229_ _01359_ vssd1 vssd1 vccd1 vccd1 _02483_ sky130_fd_sc_hd__nand2_1
X_09515_ genblk2\[1\].wave_shpr.div.quo\[5\] _04043_ _04047_ net414 vssd1 vssd1 vccd1
+ vccd1 _00212_ sky130_fd_sc_hd__a22o_1
XFILLER_0_39_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06727_ genblk1\[4\].osc.clkdiv_C.cnt\[4\] _01609_ vssd1 vssd1 vccd1 vccd1 _01613_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_79_788 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06277__B _01188_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10654__B1 _04821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_66_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_82 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09446_ genblk2\[1\].wave_shpr.div.acc\[25\] genblk2\[1\].wave_shpr.div.acc\[26\]
+ _04009_ vssd1 vssd1 vccd1 vccd1 _04010_ sky130_fd_sc_hd__or3_2
XPHY_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06658_ genblk1\[3\].osc.clkdiv_C.cnt\[15\] genblk1\[3\].osc.clkdiv_C.cnt\[14\] _01547_
+ vssd1 vssd1 vccd1 vccd1 _01551_ sky130_fd_sc_hd__and3_1
XPHY_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06873__A2 _01726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09377_ genblk2\[11\].wave_shpr.div.i\[1\] genblk2\[11\].wave_shpr.div.i\[0\] vssd1
+ vssd1 vccd1 vccd1 _03945_ sky130_fd_sc_hd__or2_1
XFILLER_0_81_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06589_ _01191_ _01233_ vssd1 vssd1 vccd1 vccd1 _01497_ sky130_fd_sc_hd__or2_1
XFILLER_0_93_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_90_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08328_ _02688_ vssd1 vssd1 vccd1 vccd1 _03035_ sky130_fd_sc_hd__inv_2
XFILLER_0_74_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06293__A _01196_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_61_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_7_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_62_666 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_104_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08259_ _02848_ _02894_ vssd1 vssd1 vccd1 vccd1 _02966_ sky130_fd_sc_hd__xor2_2
XFILLER_0_104_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_392 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11270_ genblk2\[7\].wave_shpr.div.b1\[0\] _05182_ _05183_ vssd1 vssd1 vccd1 vccd1
+ _05276_ sky130_fd_sc_hd__and3_1
X_10221_ genblk2\[3\].wave_shpr.div.acc\[20\] _04541_ vssd1 vssd1 vccd1 vccd1 _04544_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_120_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10152_ _04385_ _04491_ vssd1 vssd1 vccd1 vccd1 _04492_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_100_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10083_ _02170_ genblk2\[3\].wave_shpr.div.busy _02167_ vssd1 vssd1 vccd1 vccd1 _04453_
+ sky130_fd_sc_hd__and3_1
Xhold9 _00888_ vssd1 vssd1 vccd1 vccd1 net227 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13773_ clknet_leaf_74_clk _01084_ net213 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.acc\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_10985_ _05074_ genblk1\[6\].osc.clkdiv_C.cnt\[16\] vssd1 vssd1 vccd1 vccd1 _05078_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_29_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12724_ clknet_leaf_37_clk genblk1\[10\].osc.clkdiv_C.next_cnt\[1\] net113 vssd1
+ vssd1 vccd1 vccd1 genblk1\[10\].osc.clkdiv_C.cnt\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_155_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_641 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_84_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_38_652 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12655_ clknet_leaf_27_clk genblk1\[6\].osc.clkdiv_C.next_cnt\[4\] net90 vssd1 vssd1
+ vccd1 vccd1 genblk1\[6\].osc.clkdiv_C.cnt\[4\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__10718__A _04856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__08066__A1 _01179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11606_ genblk2\[8\].wave_shpr.div.acc\[13\] _05515_ _05493_ vssd1 vssd1 vccd1 vccd1
+ _05516_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12586_ clknet_leaf_14_clk genblk1\[2\].osc.clkdiv_C.next_cnt\[7\] net74 vssd1 vssd1
+ vccd1 vccd1 genblk1\[2\].osc.clkdiv_C.cnt\[7\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_26_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09802__A2 _04248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_135_370 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11537_ _05464_ genblk1\[8\].osc.clkdiv_C.cnt\[12\] vssd1 vssd1 vccd1 vccd1 _05466_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_151_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold409 _00480_ vssd1 vssd1 vccd1 vccd1 net627 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_123_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11468_ net1208 _01811_ _05237_ vssd1 vssd1 vccd1 vccd1 _05431_ sky130_fd_sc_hd__mux2_1
XFILLER_0_110_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13207_ clknet_leaf_25_clk _00530_ net86 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.b1\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10419_ _04654_ vssd1 vssd1 vccd1 vccd1 _04679_ sky130_fd_sc_hd__inv_2
XFILLER_0_21_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11399_ genblk2\[8\].wave_shpr.div.acc\[0\] genblk2\[8\].wave_shpr.div.b1\[0\] vssd1
+ vssd1 vccd1 vccd1 _05375_ sky130_fd_sc_hd__and2b_1
XFILLER_0_110_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_21 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13138_ clknet_leaf_115_clk net733 net135 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.quo\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13069_ clknet_leaf_24_clk net546 net93 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.quo\[21\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1109 genblk2\[2\].wave_shpr.div.quo\[3\] vssd1 vssd1 vccd1 vccd1 net1327 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_leaf_2_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_2_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__08541__A2 _02526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07630_ genblk1\[11\].osc.clkdiv_C.cnt\[8\] _02336_ net34 vssd1 vssd1 vccd1 vccd1
+ _02337_ sky130_fd_sc_hd__and3_1
XFILLER_0_136_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06378__A net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07561_ genblk1\[9\].osc.clkdiv_C.cnt\[10\] vssd1 vssd1 vccd1 vccd1 _02268_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09300_ _03776_ _03887_ vssd1 vssd1 vccd1 vccd1 _03888_ sky130_fd_sc_hd__xnor2_1
X_06512_ genblk1\[2\].osc.clkdiv_C.cnt\[6\] _01437_ vssd1 vssd1 vccd1 vccd1 _01438_
+ sky130_fd_sc_hd__xor2_1
X_07492_ _02214_ vssd1 vssd1 vccd1 vccd1 _00005_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__10100__A2 _04457_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09231_ _03725_ genblk1\[0\].osc.clkdiv_C.cnt\[1\] vssd1 vssd1 vccd1 vccd1 _03843_
+ sky130_fd_sc_hd__and2_1
X_06443_ genblk1\[1\].osc.clkdiv_C.cnt\[4\] _01380_ vssd1 vssd1 vccd1 vccd1 _01383_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_146_657 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06825__B genblk1\[5\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09162_ _03807_ vssd1 vssd1 vccd1 vccd1 _00099_ sky130_fd_sc_hd__clkbuf_1
X_06374_ _01307_ _01311_ _01312_ genblk1\[1\].osc.clkdiv_C.cnt\[11\] _01317_ vssd1
+ vssd1 vccd1 vccd1 _01318_ sky130_fd_sc_hd__o221a_1
XFILLER_0_145_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08113_ genblk1\[4\].osc.clkdiv_C.cnt\[9\] _01323_ _01592_ genblk1\[4\].osc.clkdiv_C.cnt\[8\]
+ vssd1 vssd1 vccd1 vccd1 _02820_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_32_817 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09093_ _01367_ _03739_ _03741_ _01342_ _03742_ vssd1 vssd1 vccd1 vccd1 _00095_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_688 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout216_A net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_187 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08044_ _01181_ _01680_ _02749_ _02750_ vssd1 vssd1 vccd1 vccd1 _02751_ sky130_fd_sc_hd__o211ai_1
Xhold910 PWM.final_in\[7\] vssd1 vssd1 vccd1 vccd1 net1128 sky130_fd_sc_hd__dlygate4sd3_1
Xhold921 genblk2\[0\].wave_shpr.div.acc\[2\] vssd1 vssd1 vccd1 vccd1 net1139 sky130_fd_sc_hd__dlygate4sd3_1
Xhold932 PWM.final_in\[4\] vssd1 vssd1 vccd1 vccd1 net1150 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold943 sig_norm.b1\[0\] vssd1 vssd1 vccd1 vccd1 net1161 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10363__A _03833_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold954 PWM.final_in\[3\] vssd1 vssd1 vccd1 vccd1 net1172 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07656__B _02362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold965 genblk1\[10\].osc.clkdiv_C.cnt\[8\] vssd1 vssd1 vccd1 vccd1 net1183 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07568__B1 _01246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_101_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold976 genblk1\[9\].osc.clkdiv_C.cnt\[17\] vssd1 vssd1 vccd1 vccd1 net1194 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_101_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold987 genblk2\[4\].wave_shpr.div.b1\[12\] vssd1 vssd1 vccd1 vccd1 net1205 sky130_fd_sc_hd__dlygate4sd3_1
Xhold998 _05230_ vssd1 vssd1 vccd1 vccd1 net1216 sky130_fd_sc_hd__dlygate4sd3_1
X_09995_ genblk2\[3\].wave_shpr.div.b1\[6\] genblk2\[3\].wave_shpr.div.acc\[6\] vssd1
+ vssd1 vccd1 vccd1 _04391_ sky130_fd_sc_hd__and2b_1
X_08946_ _03637_ vssd1 vssd1 vccd1 vccd1 _00053_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__12313__B1 _03944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07672__A _01308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08877_ _03577_ _03581_ _03582_ vssd1 vssd1 vccd1 vccd1 _03583_ sky130_fd_sc_hd__a21oi_1
XANTENNA__11194__A _03707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_99_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07828_ _02533_ _02534_ _02518_ vssd1 vssd1 vccd1 vccd1 _02535_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_98_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06288__A _01248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07740__B1 _01356_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07759_ genblk2\[1\].wave_shpr.div.fin_quo\[5\] _02461_ _02464_ _02224_ vssd1 vssd1
+ vccd1 vccd1 _02466_ sky130_fd_sc_hd__a31o_1
XFILLER_0_79_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12092__A2 _05844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10770_ _04809_ _04929_ vssd1 vssd1 vccd1 vccd1 _04930_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_55_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09429_ _03960_ _03991_ _03992_ vssd1 vssd1 vccd1 vccd1 _03993_ sky130_fd_sc_hd__a21o_1
XFILLER_0_109_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_717 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_109_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12440_ _06099_ _05980_ genblk2\[11\].wave_shpr.div.acc\[24\] vssd1 vssd1 vccd1 vccd1
+ _06101_ sky130_fd_sc_hd__mux2_1
X_12371_ _05953_ _05936_ vssd1 vssd1 vccd1 vccd1 _06050_ sky130_fd_sc_hd__or2b_1
XFILLER_0_151_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11322_ _05207_ _05168_ vssd1 vssd1 vccd1 vccd1 _05316_ sky130_fd_sc_hd__or2b_1
XFILLER_0_105_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_132_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11253_ genblk2\[7\].wave_shpr.div.quo\[20\] _05255_ _05256_ net231 _05266_ vssd1
+ vssd1 vccd1 vccd1 _00731_ sky130_fd_sc_hd__a221o_1
XANTENNA__07559__B1 _01361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06470__B genblk1\[1\].osc.clkdiv_C.cnt\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10204_ net1016 _04518_ _04522_ _04531_ vssd1 vssd1 vccd1 vccd1 _00417_ sky130_fd_sc_hd__a22o_1
X_11184_ _05232_ vssd1 vssd1 vccd1 vccd1 _00696_ sky130_fd_sc_hd__clkbuf_1
X_10135_ genblk2\[3\].wave_shpr.div.acc_next\[0\] _04455_ vssd1 vssd1 vccd1 vccd1
+ _04479_ sky130_fd_sc_hd__or2b_1
XANTENNA__07574__A3 _01226_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12304__B1 _06010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07582__A genblk1\[9\].osc.clkdiv_C.cnt\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10066_ net1192 _04229_ _04440_ vssd1 vssd1 vccd1 vccd1 _04443_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13756_ clknet_leaf_69_clk _01067_ net212 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.acc\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12083__A2 _05844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10968_ _05059_ genblk1\[6\].osc.clkdiv_C.cnt\[8\] vssd1 vssd1 vccd1 vccd1 _05069_
+ sky130_fd_sc_hd__and2_1
XANTENNA__10094__A1 net401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06298__B1 _01240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12707_ clknet_leaf_56_clk genblk1\[9\].osc.clkdiv_C.next_cnt\[2\] net181 vssd1 vssd1
+ vccd1 vccd1 genblk1\[9\].osc.clkdiv_C.cnt\[2\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_155_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13687_ clknet_leaf_63_clk _01000_ net191 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.acc\[25\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_38_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10899_ _03687_ _05033_ _04233_ vssd1 vssd1 vccd1 vccd1 _00610_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_128_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_622 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_116_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12638_ clknet_leaf_19_clk genblk1\[5\].osc.clkdiv_C.next_cnt\[5\] net109 vssd1 vssd1
+ vccd1 vccd1 genblk1\[5\].osc.clkdiv_C.cnt\[5\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_155_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_26_655 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09787__A1 _01365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12569_ clknet_leaf_27_clk genblk1\[1\].osc.clkdiv_C.next_cnt\[8\] net90 vssd1 vssd1
+ vccd1 vccd1 genblk1\[1\].osc.clkdiv_C.cnt\[8\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_14_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_80_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09448__S _00007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold206 genblk2\[11\].wave_shpr.div.b1\[15\] vssd1 vssd1 vccd1 vccd1 net424 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_80_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_885 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold217 _01057_ vssd1 vssd1 vccd1 vccd1 net435 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_513 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold228 genblk2\[10\].wave_shpr.div.quo\[24\] vssd1 vssd1 vccd1 vccd1 net446 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11279__A _05249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold239 genblk2\[2\].wave_shpr.div.quo\[13\] vssd1 vssd1 vccd1 vccd1 net457 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_111_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_0_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_40_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08800_ _03450_ _03449_ _03427_ _03422_ vssd1 vssd1 vccd1 vccd1 _03507_ sky130_fd_sc_hd__o211a_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06222__B1 _01183_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08762__A2 _02539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09780_ net1285 _01858_ _04238_ vssd1 vssd1 vccd1 vccd1 _04240_ sky130_fd_sc_hd__mux2_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06992_ net1252 net1058 genblk1\[7\].osc.clkdiv_C.cnt\[2\] vssd1 vssd1 vccd1 vccd1
+ _01826_ sky130_fd_sc_hd__a21oi_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07492__A _02214_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08731_ _03433_ _03437_ vssd1 vssd1 vccd1 vccd1 _03438_ sky130_fd_sc_hd__xnor2_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08662_ genblk2\[5\].wave_shpr.div.fin_quo\[2\] _03367_ _03368_ vssd1 vssd1 vccd1
+ vccd1 _03369_ sky130_fd_sc_hd__o21a_1
XANTENNA__07722__B1 _01591_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07613_ genblk1\[11\].osc.clkdiv_C.cnt\[1\] _01186_ _01354_ _01321_ genblk1\[11\].osc.clkdiv_C.cnt\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02320_ sky130_fd_sc_hd__o311a_1
X_08593_ genblk2\[4\].wave_shpr.div.fin_quo\[0\] _02526_ _02361_ genblk2\[4\].wave_shpr.div.fin_quo\[1\]
+ _02838_ vssd1 vssd1 vccd1 vccd1 _03300_ sky130_fd_sc_hd__a221o_1
XFILLER_0_89_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout166_A net170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07544_ _02255_ vssd1 vssd1 vccd1 vccd1 _00033_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10085__A1 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10085__B2 _04454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07475_ _02155_ _02202_ vssd1 vssd1 vccd1 vccd1 _02203_ sky130_fd_sc_hd__nor2_4
XFILLER_0_45_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09214_ _03835_ vssd1 vssd1 vccd1 vccd1 _03836_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_119_668 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06426_ _01197_ _01364_ _01368_ genblk1\[1\].osc.clkdiv_C.cnt\[7\] _01369_ vssd1
+ vssd1 vccd1 vccd1 _01370_ sky130_fd_sc_hd__o221a_1
XFILLER_0_8_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09227__B1 _03840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_91_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09778__A1 _01487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09145_ genblk2\[0\].wave_shpr.div.b1\[15\] genblk2\[0\].wave_shpr.div.acc\[15\]
+ vssd1 vssd1 vccd1 vccd1 _03793_ sky130_fd_sc_hd__and2b_1
XFILLER_0_16_154 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06357_ freq_div.state\[2\] freq_div.state\[0\] vssd1 vssd1 vccd1 vccd1 _01301_ sky130_fd_sc_hd__and2b_1
XANTENNA__07667__A _01308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09076_ net1291 _01483_ _03722_ vssd1 vssd1 vccd1 vccd1 _03731_ sky130_fd_sc_hd__mux2_1
X_06288_ _01248_ _01249_ vssd1 vssd1 vccd1 vccd1 _01250_ sky130_fd_sc_hd__nor2_2
XANTENNA__08450__B2 _02521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08027_ _02733_ vssd1 vssd1 vccd1 vccd1 _02734_ sky130_fd_sc_hd__buf_2
XFILLER_0_130_844 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold740 genblk2\[11\].wave_shpr.div.acc\[5\] vssd1 vssd1 vccd1 vccd1 net958 sky130_fd_sc_hd__dlygate4sd3_1
Xhold751 genblk2\[10\].wave_shpr.div.acc\[3\] vssd1 vssd1 vccd1 vccd1 net969 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_557 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold762 genblk2\[8\].wave_shpr.div.acc\[4\] vssd1 vssd1 vccd1 vccd1 net980 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold773 genblk2\[8\].wave_shpr.div.acc\[17\] vssd1 vssd1 vccd1 vccd1 net991 sky130_fd_sc_hd__dlygate4sd3_1
Xhold784 genblk2\[2\].wave_shpr.div.acc\[14\] vssd1 vssd1 vccd1 vccd1 net1002 sky130_fd_sc_hd__dlygate4sd3_1
Xhold795 genblk2\[7\].wave_shpr.div.acc\[2\] vssd1 vssd1 vccd1 vccd1 net1013 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13073__RESET_B net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06425__A1_N genblk1\[1\].osc.clkdiv_C.cnt\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09978_ genblk2\[3\].wave_shpr.div.b1\[4\] genblk2\[3\].wave_shpr.div.acc\[4\] vssd1
+ vssd1 vccd1 vccd1 _04374_ sky130_fd_sc_hd__or2b_1
XANTENNA_fanout79_A net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08929_ sig_norm.acc\[10\] _03622_ vssd1 vssd1 vccd1 vccd1 _03625_ sky130_fd_sc_hd__and2b_1
X_11940_ genblk2\[10\].wave_shpr.div.b1\[8\] genblk2\[10\].wave_shpr.div.acc\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05762_ sky130_fd_sc_hd__and2b_1
XFILLER_0_99_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11871_ _05704_ _05705_ vssd1 vssd1 vccd1 vccd1 _05706_ sky130_fd_sc_hd__nand2_1
XFILLER_0_67_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13610_ clknet_leaf_93_clk _00923_ net159 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.fin_quo\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_39_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10822_ genblk2\[6\].wave_shpr.div.acc\[17\] genblk2\[6\].wave_shpr.div.b1\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04966_ sky130_fd_sc_hd__or2b_1
XFILLER_0_67_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_79_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_39_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13541_ clknet_leaf_101_clk _00856_ net165 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.fin_quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11273__B1 _05250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10753_ genblk2\[5\].wave_shpr.div.acc\[11\] _04916_ _04907_ vssd1 vssd1 vccd1 vccd1
+ _04917_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06465__B genblk1\[1\].osc.clkdiv_C.cnt\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_137_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_82_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09218__B1 _03804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13472_ clknet_leaf_74_clk _00789_ net212 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.b1\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10684_ _04268_ vssd1 vssd1 vccd1 vccd1 _04869_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_137_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06184__C _01096_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12423_ _05976_ net20 genblk2\[11\].wave_shpr.div.acc\[18\] vssd1 vssd1 vccd1 vccd1
+ _06090_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_124_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_35_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08441__A1 _02525_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12354_ _05944_ _06036_ vssd1 vssd1 vccd1 vccd1 _06037_ sky130_fd_sc_hd__xnor2_1
XANTENNA__07244__A2 _01991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11305_ _05198_ _05302_ vssd1 vssd1 vccd1 vccd1 _05303_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_132_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10207__S _04507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12285_ _03702_ net1121 vssd1 vssd1 vccd1 vccd1 _06004_ sky130_fd_sc_hd__nor2_1
X_11236_ genblk2\[7\].wave_shpr.div.quo\[12\] _05255_ _05256_ net370 _05257_ vssd1
+ vssd1 vccd1 vccd1 _00723_ sky130_fd_sc_hd__a221o_1
XFILLER_0_120_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_120_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold7_A modein.delay_octave_down_in\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11167_ genblk2\[7\].wave_shpr.div.fin_quo\[2\] net1311 _00019_ vssd1 vssd1 vccd1
+ vccd1 _05225_ sky130_fd_sc_hd__mux2_1
X_10118_ _04465_ genblk1\[3\].osc.clkdiv_C.cnt\[9\] vssd1 vssd1 vccd1 vccd1 _04470_
+ sky130_fd_sc_hd__and2_1
XANTENNA__08201__A net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11098_ _05055_ _05158_ _05160_ _05057_ net739 vssd1 vssd1 vccd1 vccd1 _00682_ sky130_fd_sc_hd__a32o_1
XFILLER_0_89_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10049_ _04433_ vssd1 vssd1 vccd1 vccd1 _00360_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_117_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06359__C _01302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_58_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09032__A _03701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13739_ clknet_leaf_46_clk _01050_ net119 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.quo\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_27_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09209__B1 _03736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07260_ _02028_ _02036_ _02037_ vssd1 vssd1 vccd1 vccd1 _02038_ sky130_fd_sc_hd__and3_1
XFILLER_0_38_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06211_ freq_div.state\[0\] vssd1 vssd1 vccd1 vccd1 _01173_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__06691__B1 _01498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07191_ genblk1\[9\].osc.clkdiv_C.cnt\[12\] _01978_ vssd1 vssd1 vccd1 vccd1 _01979_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_6_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10906__A _01805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_357 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_83_clk_A clknet_4_14_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_14_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06142_ net2 vssd1 vssd1 vccd1 vccd1 _01114_ sky130_fd_sc_hd__inv_2
XANTENNA__09178__S _03722_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_14_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06391__A genblk1\[1\].osc.clkdiv_C.cnt\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08432__B2 _02308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_1_541 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09901_ _04197_ _04161_ vssd1 vssd1 vccd1 vccd1 _04316_ sky130_fd_sc_hd__or2b_1
XFILLER_0_1_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_65 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_98_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08196__B1 _02222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09832_ net322 _04257_ _04259_ net339 _04266_ vssd1 vssd1 vccd1 vccd1 _00310_ sky130_fd_sc_hd__a221o_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10641__A _03707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09763_ _04231_ vssd1 vssd1 vccd1 vccd1 _00276_ sky130_fd_sc_hd__clkbuf_1
X_06975_ _01365_ _01355_ vssd1 vssd1 vccd1 vccd1 _01811_ sky130_fd_sc_hd__nor2_4
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_21_clk_A clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08714_ _03408_ _03419_ _03418_ vssd1 vssd1 vccd1 vccd1 _03421_ sky130_fd_sc_hd__a21oi_2
X_09694_ _04172_ _04173_ vssd1 vssd1 vccd1 vccd1 _04174_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08645_ _03349_ _03350_ _03340_ vssd1 vssd1 vccd1 vccd1 _03352_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07171__A1 genblk1\[9\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11472__A _03707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08576_ _02525_ _03281_ _03282_ _02361_ genblk2\[11\].wave_shpr.div.fin_quo\[2\]
+ vssd1 vssd1 vccd1 vccd1 _03283_ sky130_fd_sc_hd__a32o_1
XANTENNA_clkbuf_leaf_36_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07527_ sig_norm.i\[1\] _02243_ vssd1 vssd1 vccd1 vccd1 _02245_ sky130_fd_sc_hd__nand2_1
XFILLER_0_147_741 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_92_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07458_ genblk2\[7\].wave_shpr.div.i\[2\] genblk2\[7\].wave_shpr.div.i\[3\] genblk2\[7\].wave_shpr.div.i\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02190_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_17_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_119_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_45_761 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06682__B1 _01340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06409_ _01338_ _01339_ _01346_ _01352_ vssd1 vssd1 vccd1 vccd1 _01353_ sky130_fd_sc_hd__or4b_1
XFILLER_0_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07389_ _02081_ _02136_ vssd1 vssd1 vccd1 vccd1 _02139_ sky130_fd_sc_hd__nor2_1
XFILLER_0_150_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09128_ _03757_ _03774_ _03775_ vssd1 vssd1 vccd1 vccd1 _03776_ sky130_fd_sc_hd__a21o_1
XFILLER_0_121_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09059_ _01229_ genblk2\[0\].wave_shpr.div.b1\[8\] _03719_ vssd1 vssd1 vccd1 vccd1
+ _03720_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12070_ _05815_ vssd1 vssd1 vccd1 vccd1 _05840_ sky130_fd_sc_hd__inv_2
Xhold570 genblk2\[2\].wave_shpr.div.acc\[17\] vssd1 vssd1 vccd1 vccd1 net788 sky130_fd_sc_hd__dlygate4sd3_1
Xhold581 genblk2\[9\].wave_shpr.div.acc\[14\] vssd1 vssd1 vccd1 vccd1 net799 sky130_fd_sc_hd__dlygate4sd3_1
Xhold592 PWM.counter\[5\] vssd1 vssd1 vccd1 vccd1 net810 sky130_fd_sc_hd__dlygate4sd3_1
X_11021_ _05022_ vssd1 vssd1 vccd1 vccd1 _05105_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_109_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12972_ clknet_leaf_125_clk _00301_ net71 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.quo\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_11923_ genblk2\[10\].wave_shpr.div.acc\[2\] genblk2\[10\].wave_shpr.div.b1\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05745_ sky130_fd_sc_hd__or2b_1
XTAP_2720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11854_ _05599_ _05692_ vssd1 vssd1 vccd1 vccd1 _05693_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_129_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12038__A2 _05818_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10805_ genblk2\[5\].wave_shpr.div.acc\[25\] _04953_ vssd1 vssd1 vccd1 vccd1 _04955_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_138_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_28_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11785_ _05631_ genblk1\[9\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 _05642_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_103_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13524_ clknet_leaf_98_clk _00841_ net169 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.acc\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_137_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10736_ genblk2\[5\].wave_shpr.div.acc\[7\] _04903_ _04821_ vssd1 vssd1 vccd1 vccd1
+ _04904_ sky130_fd_sc_hd__mux2_1
XFILLER_0_138_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13455_ clknet_leaf_99_clk _00772_ net168 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.fin_quo\[3\]
+ sky130_fd_sc_hd__dfrtp_2
X_10667_ net310 _04858_ _04855_ net423 _04859_ vssd1 vssd1 vccd1 vccd1 _00552_ sky130_fd_sc_hd__a221o_1
XFILLER_0_125_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12406_ _05969_ _05928_ vssd1 vssd1 vccd1 vccd1 _06077_ sky130_fd_sc_hd__or2b_1
XFILLER_0_152_265 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_742 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07217__A2 _01996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_140_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08414__B2 _02592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13386_ clknet_leaf_86_clk _00705_ net183 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.b1\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10598_ genblk2\[5\].wave_shpr.div.fin_quo\[2\] net1336 _00015_ vssd1 vssd1 vccd1
+ vccd1 _04824_ sky130_fd_sc_hd__mux2_1
XANTENNA__06425__B1 _01340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12337_ net438 _03942_ _03941_ net504 _06026_ vssd1 vssd1 vccd1 vccd1 _01055_ sky130_fd_sc_hd__a221o_1
XFILLER_0_133_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12268_ net1235 _01589_ _05994_ vssd1 vssd1 vccd1 vccd1 _05995_ sky130_fd_sc_hd__mux2_1
X_11219_ genblk2\[7\].wave_shpr.div.quo\[2\] _05246_ _05250_ net563 vssd1 vssd1 vccd1
+ vccd1 _00713_ sky130_fd_sc_hd__a22o_1
XFILLER_0_120_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12199_ genblk2\[11\].wave_shpr.div.acc\[5\] genblk2\[11\].wave_shpr.div.b1\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05937_ sky130_fd_sc_hd__or2b_1
X_06760_ _01599_ _01636_ _01638_ vssd1 vssd1 vccd1 vccd1 _01639_ sky130_fd_sc_hd__and3_1
XFILLER_0_78_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06691_ genblk1\[4\].osc.clkdiv_C.cnt\[0\] _01210_ _01498_ genblk1\[4\].osc.clkdiv_C.cnt\[14\]
+ _01580_ vssd1 vssd1 vccd1 vccd1 _01581_ sky130_fd_sc_hd__o221a_1
XANTENNA__08350__B1 _02527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08430_ _02303_ _02262_ genblk2\[9\].wave_shpr.div.fin_quo\[2\] vssd1 vssd1 vccd1
+ vccd1 _03137_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_144_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12029__A2 _05813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_801 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08361_ genblk2\[3\].wave_shpr.div.fin_quo\[4\] _03067_ vssd1 vssd1 vccd1 vccd1 _03068_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_59_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07312_ genblk1\[11\].osc.clkdiv_C.cnt\[14\] _01210_ _01578_ genblk1\[11\].osc.clkdiv_C.cnt\[16\]
+ _02075_ vssd1 vssd1 vccd1 vccd1 _02076_ sky130_fd_sc_hd__o221a_1
XANTENNA__13765__RESET_B net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08292_ _02945_ _02967_ vssd1 vssd1 vccd1 vccd1 _02999_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_143_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07243_ genblk1\[10\].osc.clkdiv_C.cnt\[7\] _01235_ _02020_ _02022_ _02024_ vssd1
+ vssd1 vccd1 vccd1 _02025_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_144_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07929__B net30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_143_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07174_ genblk1\[9\].osc.clkdiv_C.cnt\[6\] _01965_ vssd1 vssd1 vccd1 vccd1 _01968_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06125_ _01094_ _01095_ _01096_ vssd1 vssd1 vccd1 vccd1 _01097_ sky130_fd_sc_hd__nor3_2
XFILLER_0_131_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_2_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_100_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_78_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10371__A _04654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09815_ _04247_ vssd1 vssd1 vccd1 vccd1 _04257_ sky130_fd_sc_hd__clkbuf_4
X_09746_ _04220_ vssd1 vssd1 vccd1 vccd1 _00270_ sky130_fd_sc_hd__clkbuf_1
X_06958_ _01228_ _01220_ _01233_ vssd1 vssd1 vccd1 vccd1 _01794_ sky130_fd_sc_hd__a21oi_4
XANTENNA__07680__A _01181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2005 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09677_ genblk2\[2\].wave_shpr.div.acc\[16\] genblk2\[2\].wave_shpr.div.b1\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04157_ sky130_fd_sc_hd__or2b_1
XTAP_2016 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06889_ genblk1\[6\].osc.clkdiv_C.cnt\[12\] _01519_ _01742_ genblk1\[6\].osc.clkdiv_C.cnt\[10\]
+ vssd1 vssd1 vccd1 vccd1 _01743_ sky130_fd_sc_hd__a2bb2o_1
XTAP_2027 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12298__A _03941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2038 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08628_ _03275_ _03276_ _03295_ vssd1 vssd1 vccd1 vccd1 _03335_ sky130_fd_sc_hd__nand3_2
XTAP_2049 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06296__A _01238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11228__B1 _05248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08559_ _03264_ _03265_ vssd1 vssd1 vccd1 vccd1 _03266_ sky130_fd_sc_hd__nor2_1
XTAP_1359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11570_ _05384_ _05370_ vssd1 vssd1 vccd1 vccd1 _05488_ sky130_fd_sc_hd__or2b_1
XFILLER_0_92_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_52_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10521_ _04654_ _04651_ genblk2\[4\].wave_shpr.div.i\[0\] vssd1 vssd1 vccd1 vccd1
+ _04754_ sky130_fd_sc_hd__mux2_1
XFILLER_0_135_766 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_107_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13240_ clknet_leaf_11_clk net234 net57 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.quo\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_150_725 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10452_ _04622_ vssd1 vssd1 vccd1 vccd1 _04704_ sky130_fd_sc_hd__buf_4
XFILLER_0_33_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13171_ clknet_leaf_126_clk _00496_ net66 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.acc\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10383_ _04058_ _01568_ vssd1 vssd1 vccd1 vccd1 _04659_ sky130_fd_sc_hd__nor2_1
X_12122_ net957 _05876_ _05850_ _05879_ vssd1 vssd1 vccd1 vccd1 _00987_ sky130_fd_sc_hd__a22o_1
X_12053_ _05819_ genblk1\[10\].osc.clkdiv_C.cnt\[9\] vssd1 vssd1 vccd1 vccd1 _05831_
+ sky130_fd_sc_hd__and2_1
X_11004_ genblk2\[6\].wave_shpr.div.acc\[3\] _05091_ _05023_ vssd1 vssd1 vccd1 vccd1
+ _05092_ sky130_fd_sc_hd__mux2_1
X_12955_ clknet_leaf_136_clk _00284_ net62 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.b1\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_59_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07135__A1 genblk1\[9\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07135__B2 genblk1\[9\].osc.clkdiv_C.cnt\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11906_ _03690_ _05728_ _05729_ vssd1 vssd1 vccd1 vccd1 _00921_ sky130_fd_sc_hd__nor3_1
XTAP_2550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12886_ clknet_leaf_30_clk _00217_ net98 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.quo\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11219__B1 _05250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11837_ genblk2\[9\].wave_shpr.div.acc\[10\] _05679_ _05673_ vssd1 vssd1 vccd1 vccd1
+ _05680_ sky130_fd_sc_hd__mux2_1
XTAP_2594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1871 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1882 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1893 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11768_ net485 _05628_ _05629_ net541 _05633_ vssd1 vssd1 vccd1 vccd1 _00879_ sky130_fd_sc_hd__a221o_1
XFILLER_0_138_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10719_ _04787_ _04779_ vssd1 vssd1 vccd1 vccd1 _04891_ sky130_fd_sc_hd__or2b_1
X_13507_ clknet_leaf_80_clk _00824_ net205 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.acc\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11699_ _05562_ _05589_ _05590_ vssd1 vssd1 vccd1 vccd1 _05591_ sky130_fd_sc_hd__a21o_1
XFILLER_0_125_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13438_ clknet_leaf_95_clk _00757_ net159 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.acc\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_153_585 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_758 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_51_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_113_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_786 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_140_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13369_ clknet_leaf_116_clk _00688_ net140 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.fin_quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09456__S _00007_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_11_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07930_ genblk2\[8\].wave_shpr.div.fin_quo\[5\] vssd1 vssd1 vccd1 vccd1 _02637_ sky130_fd_sc_hd__inv_2
XANTENNA__07484__B _02153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07861_ genblk2\[1\].wave_shpr.div.fin_quo\[0\] _02458_ _02459_ genblk2\[1\].wave_shpr.div.fin_quo\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02568_ sky130_fd_sc_hd__a31o_1
X_09600_ genblk2\[1\].wave_shpr.div.acc\[9\] _04101_ _04095_ vssd1 vssd1 vccd1 vccd1
+ _04102_ sky130_fd_sc_hd__mux2_1
XANTENNA__08571__B1 _02316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06812_ _01189_ _01678_ vssd1 vssd1 vccd1 vccd1 _01684_ sky130_fd_sc_hd__nor2_2
XANTENNA__07913__A3 _01855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07792_ _01246_ _01439_ _01344_ _01169_ vssd1 vssd1 vccd1 vccd1 _02499_ sky130_fd_sc_hd__a31o_1
X_09531_ _04055_ genblk1\[1\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 _04056_
+ sky130_fd_sc_hd__and2_1
X_06743_ _01599_ _01624_ _01625_ vssd1 vssd1 vccd1 vccd1 _01626_ sky130_fd_sc_hd__and3_1
XANTENNA__07126__A1 genblk1\[9\].osc.clkdiv_C.cnt\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07126__B2 genblk1\[9\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09462_ genblk2\[1\].wave_shpr.div.fin_quo\[7\] genblk2\[1\].wave_shpr.div.quo\[6\]
+ _00007_ vssd1 vssd1 vccd1 vccd1 _04019_ sky130_fd_sc_hd__mux2_1
X_06674_ _01563_ vssd1 vssd1 vccd1 vccd1 _01564_ sky130_fd_sc_hd__buf_6
XFILLER_0_66_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_78_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08413_ genblk2\[2\].wave_shpr.div.fin_quo\[6\] _03119_ vssd1 vssd1 vccd1 vccd1 _03120_
+ sky130_fd_sc_hd__xnor2_1
X_09393_ genblk2\[1\].wave_shpr.div.acc\[14\] genblk2\[1\].wave_shpr.div.b1\[14\]
+ vssd1 vssd1 vccd1 vccd1 _03957_ sky130_fd_sc_hd__or2b_1
XFILLER_0_93_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08344_ _03048_ _03049_ _03050_ vssd1 vssd1 vccd1 vccd1 _03051_ sky130_fd_sc_hd__and3_2
XFILLER_0_74_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_117_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_675 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_744 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07659__B _02364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08275_ genblk2\[10\].wave_shpr.div.fin_quo\[5\] _02361_ _02980_ _02981_ vssd1 vssd1
+ vccd1 vccd1 _02982_ sky130_fd_sc_hd__a22o_1
XANTENNA__10366__A _04651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__10984__A2 _05051_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07226_ genblk1\[10\].osc.clkdiv_C.cnt\[5\] _01992_ _02007_ vssd1 vssd1 vccd1 vccd1
+ _02008_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_104_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07157_ genblk1\[9\].osc.clkdiv_C.cnt\[1\] genblk1\[9\].osc.clkdiv_C.cnt\[0\] vssd1
+ vssd1 vccd1 vccd1 _01956_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06108_ net1179 net395 _01088_ vssd1 vssd1 vccd1 vccd1 _01089_ sky130_fd_sc_hd__and3_1
XFILLER_0_131_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07088_ genblk1\[8\].osc.clkdiv_C.cnt\[7\] _01897_ _01886_ vssd1 vssd1 vccd1 vccd1
+ _01899_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_100_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout110 net111 vssd1 vssd1 vccd1 vccd1 net110 sky130_fd_sc_hd__clkbuf_4
Xfanout121 net122 vssd1 vssd1 vccd1 vccd1 net121 sky130_fd_sc_hd__clkbuf_4
Xfanout132 net133 vssd1 vssd1 vccd1 vccd1 net132 sky130_fd_sc_hd__clkbuf_4
Xfanout143 net145 vssd1 vssd1 vccd1 vccd1 net143 sky130_fd_sc_hd__clkbuf_4
Xfanout154 net155 vssd1 vssd1 vccd1 vccd1 net154 sky130_fd_sc_hd__buf_2
Xfanout165 net170 vssd1 vssd1 vccd1 vccd1 net165 sky130_fd_sc_hd__clkbuf_4
Xfanout176 net218 vssd1 vssd1 vccd1 vccd1 net176 sky130_fd_sc_hd__clkbuf_2
Xfanout187 net188 vssd1 vssd1 vccd1 vccd1 net187 sky130_fd_sc_hd__clkbuf_4
Xfanout198 net218 vssd1 vssd1 vccd1 vccd1 net198 sky130_fd_sc_hd__buf_2
XFILLER_0_97_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09729_ genblk2\[2\].wave_shpr.div.acc\[18\] _04208_ vssd1 vssd1 vccd1 vccd1 _04209_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_97_712 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_97_756 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12740_ clknet_leaf_48_clk genblk1\[10\].osc.clkdiv_C.next_cnt\[17\] net119 vssd1
+ vssd1 vccd1 vccd1 genblk1\[10\].osc.clkdiv_C.cnt\[17\] sky130_fd_sc_hd__dfrtp_1
XTAP_1101 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07668__A2 _02374_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1112 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1123 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12671_ clknet_leaf_89_clk genblk1\[7\].osc.clkdiv_C.next_cnt\[2\] net173 vssd1 vssd1
+ vccd1 vccd1 genblk1\[7\].osc.clkdiv_C.cnt\[2\] sky130_fd_sc_hd__dfrtp_4
XTAP_1156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11622_ genblk2\[8\].wave_shpr.div.acc\[17\] _05527_ _05416_ vssd1 vssd1 vccd1 vccd1
+ _05528_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09814__B1 _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11553_ genblk2\[8\].wave_shpr.div.acc\[1\] _05416_ vssd1 vssd1 vccd1 vccd1 _05475_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_123_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10504_ genblk2\[4\].wave_shpr.div.acc\[20\] _04740_ vssd1 vssd1 vccd1 vccd1 _04743_
+ sky130_fd_sc_hd__xnor2_1
X_11484_ _03727_ _01490_ _03687_ net478 vssd1 vssd1 vccd1 vccd1 _00790_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__12177__A1 _05816_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_561 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13223_ clknet_leaf_114_clk _00546_ net132 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10435_ _04589_ _04581_ vssd1 vssd1 vccd1 vccd1 _04691_ sky130_fd_sc_hd__or2b_1
XFILLER_0_150_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07053__B1 _01870_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13154_ clknet_leaf_121_clk _00479_ net77 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.quo\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10366_ _04651_ vssd1 vssd1 vccd1 vccd1 _04652_ sky130_fd_sc_hd__buf_2
X_12105_ net954 _05844_ _05850_ _05866_ vssd1 vssd1 vccd1 vccd1 _00983_ sky130_fd_sc_hd__a22o_1
XTAP_907 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06800__B1 _01666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13085_ clknet_leaf_135_clk _00412_ net62 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.acc\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_929 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10297_ _04569_ _04607_ _04608_ vssd1 vssd1 vccd1 vccd1 _04609_ sky130_fd_sc_hd__a21o_1
X_12036_ net398 _05818_ _05816_ net432 _05821_ vssd1 vssd1 vccd1 vccd1 _00959_ sky130_fd_sc_hd__a221o_1
XANTENNA__08553__B1 _02261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_907 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12938_ clknet_leaf_111_clk _00267_ net136 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.fin_quo\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10663__A1 net308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12869_ clknet_leaf_134_clk _00200_ net60 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.b1\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_133_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_205 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_28_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_653 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06390_ _01333_ vssd1 vssd1 vccd1 vccd1 _01334_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__09805__B1 _04252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09040__A _03707_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_826 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08060_ genblk1\[5\].osc.clkdiv_C.cnt\[5\] _01238_ vssd1 vssd1 vccd1 vccd1 _02767_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_43_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07011_ genblk1\[7\].osc.clkdiv_C.cnt\[9\] _01835_ vssd1 vssd1 vccd1 vccd1 _01838_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07495__A _02216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08962_ _03507_ _03451_ vssd1 vssd1 vccd1 vccd1 _03650_ sky130_fd_sc_hd__nor2_1
XANTENNA__08103__B _01574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07913_ genblk1\[8\].osc.clkdiv_C.cnt\[0\] _01309_ _01855_ genblk1\[8\].osc.clkdiv_C.cnt\[1\]
+ genblk1\[8\].osc.clkdiv_C.cnt\[2\] vssd1 vssd1 vccd1 vccd1 _02620_ sky130_fd_sc_hd__a311o_1
X_08893_ _01099_ _03574_ _03598_ vssd1 vssd1 vccd1 vccd1 _03599_ sky130_fd_sc_hd__and3_1
XANTENNA_fanout196_A net198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07844_ genblk2\[0\].wave_shpr.div.fin_quo\[2\] _02549_ _02550_ vssd1 vssd1 vccd1
+ vccd1 _02551_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_98_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09215__A _02152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07775_ genblk1\[0\].osc.clkdiv_C.cnt\[2\] _01227_ _02479_ _02480_ _02481_ vssd1
+ vssd1 vccd1 vccd1 _02482_ sky130_fd_sc_hd__o221a_1
X_09514_ net414 _04043_ _04047_ net701 vssd1 vssd1 vccd1 vccd1 _00211_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_79_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06726_ _01612_ vssd1 vssd1 vccd1 vccd1 genblk1\[4\].osc.clkdiv_C.next_cnt\[3\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_149_644 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09445_ genblk2\[1\].wave_shpr.div.acc\[24\] _04008_ vssd1 vssd1 vccd1 vccd1 _04009_
+ sky130_fd_sc_hd__or2_2
XFILLER_0_148_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10654__B2 _04855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06657_ net1195 _01547_ _01550_ vssd1 vssd1 vccd1 vccd1 genblk1\[3\].osc.clkdiv_C.next_cnt\[14\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_91_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_19_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09376_ _03940_ vssd1 vssd1 vccd1 vccd1 _03944_ sky130_fd_sc_hd__clkbuf_4
X_06588_ _01437_ _01225_ vssd1 vssd1 vccd1 vccd1 _01496_ sky130_fd_sc_hd__or2_4
XFILLER_0_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__12296__B1_N _03735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_686 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08327_ genblk2\[8\].wave_shpr.div.fin_quo\[5\] _02467_ _03033_ _02636_ vssd1 vssd1
+ vccd1 vccd1 _03034_ sky130_fd_sc_hd__a211o_1
XANTENNA__10096__A _04451_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08075__A2 _01678_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09272__B2 _03836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08258_ _02958_ _02963_ _02964_ vssd1 vssd1 vccd1 vccd1 _02965_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_62_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07209_ _01556_ _01564_ vssd1 vssd1 vccd1 vccd1 _01991_ sky130_fd_sc_hd__nand2_8
X_08189_ _02849_ _02894_ _02895_ vssd1 vssd1 vccd1 vccd1 _02896_ sky130_fd_sc_hd__o21a_1
XFILLER_0_15_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10220_ genblk2\[3\].wave_shpr.div.acc\[20\] _04541_ vssd1 vssd1 vccd1 vccd1 _04543_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_42_391 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07035__B1 _01248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_30_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10151_ _04386_ _04377_ vssd1 vssd1 vccd1 vccd1 _04491_ sky130_fd_sc_hd__or2b_1
XFILLER_0_30_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10082_ _04451_ vssd1 vssd1 vccd1 vccd1 _04452_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_89_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07571__C _01355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_69_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_97_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13772_ clknet_leaf_73_clk _01083_ net215 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.acc\[24\]
+ sky130_fd_sc_hd__dfrtp_2
X_10984_ genblk2\[6\].wave_shpr.div.quo\[24\] _05051_ _05054_ net385 _05077_ vssd1
+ vssd1 vccd1 vccd1 _00651_ sky130_fd_sc_hd__a221o_1
XFILLER_0_139_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10645__A1 _01365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12723_ clknet_leaf_37_clk genblk1\[10\].osc.clkdiv_C.next_cnt\[0\] net113 vssd1
+ vssd1 vccd1 vccd1 genblk1\[10\].osc.clkdiv_C.cnt\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_84_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_128_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_128_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12654_ clknet_leaf_27_clk genblk1\[6\].osc.clkdiv_C.next_cnt\[3\] net90 vssd1 vssd1
+ vccd1 vccd1 genblk1\[6\].osc.clkdiv_C.cnt\[3\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_84_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11605_ _05399_ _05514_ vssd1 vssd1 vccd1 vccd1 _05515_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_155_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07299__B _01235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12585_ clknet_leaf_124_clk genblk1\[2\].osc.clkdiv_C.next_cnt\[6\] net76 vssd1 vssd1
+ vccd1 vccd1 genblk1\[2\].osc.clkdiv_C.cnt\[6\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_111_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09795__A _02152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11536_ net660 _05454_ _05458_ net677 _05465_ vssd1 vssd1 vccd1 vccd1 _00815_ sky130_fd_sc_hd__a221o_1
XFILLER_0_135_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11740__A1_N _01099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_34_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11467_ _05430_ vssd1 vssd1 vccd1 vccd1 _00781_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_111_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13206_ clknet_leaf_25_clk _00529_ net88 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.b1\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10418_ net643 _04651_ _04654_ genblk2\[4\].wave_shpr.div.quo\[24\] _04678_ vssd1
+ vssd1 vccd1 vccd1 _00484_ sky130_fd_sc_hd__a221o_1
XFILLER_0_110_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09566__A2 _04043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11398_ genblk2\[8\].wave_shpr.div.acc\[1\] genblk2\[8\].wave_shpr.div.b1\[1\] vssd1
+ vssd1 vccd1 vccd1 _05374_ sky130_fd_sc_hd__xor2_1
X_13137_ clknet_leaf_115_clk _00462_ net135 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.quo\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_33 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10349_ net1266 _01757_ _04637_ vssd1 vssd1 vccd1 vccd1 _04642_ sky130_fd_sc_hd__mux2_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13068_ clknet_leaf_24_clk net297 net93 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.quo\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11565__A _05444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12019_ _05814_ vssd1 vssd1 vccd1 vccd1 _05815_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__10333__B1 _01262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09035__A _02171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07560_ genblk1\[9\].osc.clkdiv_C.cnt\[13\] _01245_ _01328_ genblk1\[9\].osc.clkdiv_C.cnt\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02267_ sky130_fd_sc_hd__o22a_1
X_06511_ _01332_ vssd1 vssd1 vccd1 vccd1 _01437_ sky130_fd_sc_hd__buf_4
XFILLER_0_88_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07491_ _02211_ _02152_ genblk2\[11\].wave_shpr.div.busy vssd1 vssd1 vccd1 vccd1
+ _02214_ sky130_fd_sc_hd__and3b_1
XFILLER_0_76_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06304__A2 _01235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09230_ genblk2\[0\].wave_shpr.div.quo\[9\] _03841_ _03839_ net277 _03842_ vssd1
+ vssd1 vccd1 vccd1 _00132_ sky130_fd_sc_hd__a221o_1
X_06442_ genblk1\[1\].osc.clkdiv_C.cnt\[4\] _01380_ vssd1 vssd1 vccd1 vccd1 _01382_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_119_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_29_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_669 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09161_ genblk2\[0\].wave_shpr.div.fin_quo\[2\] net1322 _00001_ vssd1 vssd1 vccd1
+ vccd1 _03807_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06373_ genblk1\[1\].osc.clkdiv_C.cnt\[2\] _01240_ vssd1 vssd1 vccd1 vccd1 _01317_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_127_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_16_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_44_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08112_ _02804_ _02806_ _02808_ _02817_ _02818_ vssd1 vssd1 vccd1 vccd1 _02819_ sky130_fd_sc_hd__o221a_1
X_09092_ _01367_ _03740_ vssd1 vssd1 vccd1 vccd1 _03742_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_678 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08043_ genblk1\[5\].osc.clkdiv_C.cnt\[14\] _01360_ vssd1 vssd1 vccd1 vccd1 _02750_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_fanout111_A net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold900 genblk2\[10\].wave_shpr.div.acc\[1\] vssd1 vssd1 vccd1 vccd1 net1118 sky130_fd_sc_hd__dlygate4sd3_1
Xhold911 genblk2\[4\].wave_shpr.div.acc\[1\] vssd1 vssd1 vccd1 vccd1 net1129 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_840 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold922 genblk2\[7\].wave_shpr.div.b1\[1\] vssd1 vssd1 vccd1 vccd1 net1140 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_728 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout209_A net210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12010__B1 _03733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold933 _03682_ vssd1 vssd1 vccd1 vccd1 net1151 sky130_fd_sc_hd__dlygate4sd3_1
Xhold944 genblk1\[8\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 net1162 sky130_fd_sc_hd__dlygate4sd3_1
Xhold955 genblk2\[10\].wave_shpr.div.b1\[6\] vssd1 vssd1 vccd1 vccd1 net1173 sky130_fd_sc_hd__dlygate4sd3_1
Xhold966 genblk2\[0\].wave_shpr.div.b1\[10\] vssd1 vssd1 vccd1 vccd1 net1184 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07568__B2 genblk1\[9\].osc.clkdiv_C.cnt\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold977 genblk1\[3\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 net1195 sky130_fd_sc_hd__dlygate4sd3_1
X_09994_ _04373_ _04388_ _04389_ vssd1 vssd1 vccd1 vccd1 _04390_ sky130_fd_sc_hd__a21o_1
Xhold988 genblk2\[4\].wave_shpr.div.b1\[8\] vssd1 vssd1 vccd1 vccd1 net1206 sky130_fd_sc_hd__dlygate4sd3_1
Xhold999 genblk2\[11\].wave_shpr.div.b1\[9\] vssd1 vssd1 vccd1 vccd1 net1217 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06240__A1 _01201_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08945_ sig_norm.quo\[2\] _03636_ _00024_ vssd1 vssd1 vccd1 vccd1 _03637_ sky130_fd_sc_hd__mux2_1
X_08876_ sig_norm.b1\[2\] sig_norm.acc\[2\] vssd1 vssd1 vccd1 vccd1 _03582_ sky130_fd_sc_hd__xor2_1
X_07827_ genblk2\[0\].wave_shpr.div.fin_quo\[4\] _02309_ _02509_ vssd1 vssd1 vccd1
+ vccd1 _02534_ sky130_fd_sc_hd__a21o_1
XANTENNA__06288__B _01249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07740__A1 genblk1\[1\].osc.clkdiv_C.cnt\[9\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__13208__RESET_B net88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07740__B2 genblk1\[1\].osc.clkdiv_C.cnt\[8\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07758_ _02461_ _02464_ genblk2\[1\].wave_shpr.div.fin_quo\[5\] vssd1 vssd1 vccd1
+ vccd1 _02465_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_66_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_726 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06709_ _01558_ _01560_ _01584_ _01598_ vssd1 vssd1 vccd1 vccd1 _01599_ sky130_fd_sc_hd__or4_4
XANTENNA__09493__A1 _04036_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07689_ genblk1\[10\].osc.clkdiv_C.cnt\[10\] _02005_ _02394_ _02395_ vssd1 vssd1
+ vccd1 vccd1 _02396_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_66_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09428_ genblk2\[1\].wave_shpr.div.b1\[11\] genblk2\[1\].wave_shpr.div.acc\[11\]
+ vssd1 vssd1 vccd1 vccd1 _03992_ sky130_fd_sc_hd__and2b_1
XFILLER_0_125_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09359_ net933 _03903_ _03910_ _03932_ vssd1 vssd1 vccd1 vccd1 _00171_ sky130_fd_sc_hd__a22o_1
XFILLER_0_137_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_118_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_35_667 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12370_ net841 _06039_ _06040_ _06049_ vssd1 vssd1 vccd1 vccd1 _01065_ sky130_fd_sc_hd__a22o_1
XFILLER_0_105_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11321_ _05249_ vssd1 vssd1 vccd1 vccd1 _05315_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_90_795 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11252_ _05260_ genblk1\[7\].osc.clkdiv_C.cnt\[11\] vssd1 vssd1 vccd1 vccd1 _05266_
+ sky130_fd_sc_hd__and2_1
XANTENNA__07559__A1 _01200_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10203_ genblk2\[3\].wave_shpr.div.acc\[15\] _04530_ _04507_ vssd1 vssd1 vccd1 vccd1
+ _04531_ sky130_fd_sc_hd__mux2_1
X_11183_ net1214 _04242_ _05042_ vssd1 vssd1 vccd1 vccd1 _05232_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10134_ genblk2\[3\].wave_shpr.div.acc_next\[0\] _04451_ _04455_ net561 _04478_ vssd1
+ vssd1 vccd1 vccd1 _00400_ sky130_fd_sc_hd__a221o_1
X_10065_ _04442_ vssd1 vssd1 vccd1 vccd1 _00367_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_106_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09484__A1 _01302_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10967_ net595 _05062_ _05064_ net594 _05068_ vssd1 vssd1 vccd1 vccd1 _00643_ sky130_fd_sc_hd__a221o_1
X_13755_ clknet_leaf_68_clk _01066_ net212 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.acc\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06298__A1 genblk1\[0\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10094__A2 _04452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_73_707 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12706_ clknet_leaf_86_clk genblk1\[9\].osc.clkdiv_C.next_cnt\[1\] net183 vssd1 vssd1
+ vccd1 vccd1 genblk1\[9\].osc.clkdiv_C.cnt\[1\] sky130_fd_sc_hd__dfrtp_4
X_13686_ clknet_leaf_63_clk _00999_ net191 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.acc\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10898_ net1140 vssd1 vssd1 vccd1 vccd1 _05033_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12637_ clknet_leaf_16_clk genblk1\[5\].osc.clkdiv_C.next_cnt\[4\] net73 vssd1 vssd1
+ vccd1 vccd1 genblk1\[5\].osc.clkdiv_C.cnt\[4\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_143_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_26_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_517 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_667 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12568_ clknet_leaf_27_clk genblk1\[1\].osc.clkdiv_C.next_cnt\[7\] net90 vssd1 vssd1
+ vccd1 vccd1 genblk1\[1\].osc.clkdiv_C.cnt\[7\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_135_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11519_ _05450_ genblk1\[8\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 _05456_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_124_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_151_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12499_ clknet_leaf_103_clk _00061_ net156 vssd1 vssd1 vccd1 vccd1 sig_norm.quo\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_123_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold207 genblk2\[1\].wave_shpr.div.b1\[16\] vssd1 vssd1 vccd1 vccd1 net425 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold218 genblk1\[3\].osc.clkdiv_C.cnt\[17\] vssd1 vssd1 vccd1 vccd1 net436 sky130_fd_sc_hd__buf_1
XFILLER_0_124_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold229 _00973_ vssd1 vssd1 vccd1 vccd1 net447 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_1_734 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09464__S _03822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06222__A1 _01172_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06991_ genblk1\[7\].osc.clkdiv_C.cnt\[2\] genblk1\[7\].osc.clkdiv_C.cnt\[1\] genblk1\[7\].osc.clkdiv_C.cnt\[0\]
+ vssd1 vssd1 vccd1 vccd1 _01825_ sky130_fd_sc_hd__and3_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08730_ _03114_ _03436_ _03122_ vssd1 vssd1 vccd1 vccd1 _03437_ sky130_fd_sc_hd__o21a_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06389__A _01179_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08661_ _03176_ _02789_ _03177_ _02525_ vssd1 vssd1 vccd1 vccd1 _03368_ sky130_fd_sc_hd__o31a_1
X_07612_ _01186_ _01354_ genblk1\[11\].osc.clkdiv_C.cnt\[1\] vssd1 vssd1 vccd1 vccd1
+ _02319_ sky130_fd_sc_hd__o21a_1
X_08592_ genblk2\[5\].wave_shpr.div.fin_quo\[0\] _02527_ _02521_ genblk2\[5\].wave_shpr.div.fin_quo\[1\]
+ _02791_ vssd1 vssd1 vccd1 vccd1 _03299_ sky130_fd_sc_hd__a221o_1
XFILLER_0_49_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07543_ PWM.final_sample_in\[3\] net1172 PWM.start vssd1 vssd1 vccd1 vccd1 _02255_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_49_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09475__A1 _01248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12074__A3 _05787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10085__A2 _04452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07474_ genblk2\[9\].wave_shpr.div.busy _02201_ vssd1 vssd1 vccd1 vccd1 _02202_ sky130_fd_sc_hd__and2_2
X_09213_ _02151_ vssd1 vssd1 vccd1 vccd1 _03835_ sky130_fd_sc_hd__buf_2
X_06425_ genblk1\[1\].osc.clkdiv_C.cnt\[7\] _01368_ _01340_ genblk1\[1\].osc.clkdiv_C.cnt\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01369_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_146_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_134_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09144_ _03749_ _03790_ _03791_ vssd1 vssd1 vccd1 vccd1 _03792_ sky130_fd_sc_hd__a21o_1
X_06356_ genblk1\[0\].osc.clkdiv_C.cnt\[17\] _01298_ _01300_ _01270_ vssd1 vssd1 vccd1
+ vccd1 genblk1\[0\].osc.clkdiv_C.next_cnt\[17\] sky130_fd_sc_hd__o211a_1
XFILLER_0_32_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_16_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09075_ _03730_ vssd1 vssd1 vccd1 vccd1 _00089_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06287_ _01173_ _01188_ vssd1 vssd1 vccd1 vccd1 _01249_ sky130_fd_sc_hd__nor2_4
XFILLER_0_114_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_102_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_114_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08026_ _02712_ _02731_ _02732_ vssd1 vssd1 vccd1 vccd1 _02733_ sky130_fd_sc_hd__o21a_4
XFILLER_0_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold730 genblk2\[3\].wave_shpr.div.acc\[17\] vssd1 vssd1 vccd1 vccd1 net948 sky130_fd_sc_hd__dlygate4sd3_1
Xhold741 genblk2\[10\].wave_shpr.div.b1\[16\] vssd1 vssd1 vccd1 vccd1 net959 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold752 genblk2\[4\].wave_shpr.div.acc\[5\] vssd1 vssd1 vccd1 vccd1 net970 sky130_fd_sc_hd__dlygate4sd3_1
Xhold763 genblk2\[5\].wave_shpr.div.acc\[13\] vssd1 vssd1 vccd1 vccd1 net981 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_569 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold774 genblk2\[7\].wave_shpr.div.acc\[3\] vssd1 vssd1 vccd1 vccd1 net992 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_130_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold785 genblk2\[6\].wave_shpr.div.acc\[10\] vssd1 vssd1 vccd1 vccd1 net1003 sky130_fd_sc_hd__dlygate4sd3_1
Xhold796 genblk2\[5\].wave_shpr.div.acc\[12\] vssd1 vssd1 vccd1 vccd1 net1014 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07683__A _01174_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09950__A2 _04253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09977_ genblk2\[3\].wave_shpr.div.acc\[5\] genblk2\[3\].wave_shpr.div.b1\[5\] vssd1
+ vssd1 vccd1 vccd1 _04373_ sky130_fd_sc_hd__or2b_1
XANTENNA__06407__A2_N _01349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08928_ net663 _02260_ _03624_ vssd1 vssd1 vccd1 vccd1 _00048_ sky130_fd_sc_hd__a21o_1
XFILLER_0_99_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_99_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08859_ _03427_ _03505_ _03500_ _03504_ vssd1 vssd1 vccd1 vccd1 _03566_ sky130_fd_sc_hd__a211oi_1
X_11870_ _05607_ _05646_ genblk2\[9\].wave_shpr.div.acc\[18\] vssd1 vssd1 vccd1 vccd1
+ _05705_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_86_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10821_ net856 _04965_ vssd1 vssd1 vccd1 vccd1 _00600_ sky130_fd_sc_hd__nor2_1
XFILLER_0_79_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09466__A1 _01327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10752_ _04801_ _04915_ vssd1 vssd1 vccd1 vccd1 _04916_ sky130_fd_sc_hd__xnor2_1
X_13540_ clknet_leaf_101_clk _00855_ net164 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.fin_quo\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_39_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_55_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13471_ clknet_leaf_75_clk _00788_ net204 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.b1\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10683_ net378 _04861_ _04862_ net551 _04868_ vssd1 vssd1 vccd1 vccd1 _00559_ sky130_fd_sc_hd__a221o_1
XANTENNA__09218__A1 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09218__B2 _03839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12422_ _05977_ net20 vssd1 vssd1 vccd1 vccd1 _06089_ sky130_fd_sc_hd__or2_1
XFILLER_0_152_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07858__A _02216_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_63_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_853 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12353_ genblk2\[11\].wave_shpr.div.b1\[2\] genblk2\[11\].wave_shpr.div.acc\[2\]
+ vssd1 vssd1 vccd1 vccd1 _06036_ sky130_fd_sc_hd__xor2_1
X_11304_ _05199_ _05172_ vssd1 vssd1 vccd1 vccd1 _05302_ sky130_fd_sc_hd__or2b_1
XFILLER_0_133_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12284_ _06003_ vssd1 vssd1 vccd1 vccd1 _01025_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_132_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11235_ _05074_ genblk1\[7\].osc.clkdiv_C.cnt\[3\] vssd1 vssd1 vccd1 vccd1 _05257_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_30_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09284__S _03804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09941__A2 _04253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11166_ _05224_ vssd1 vssd1 vccd1 vccd1 _00686_ sky130_fd_sc_hd__clkbuf_1
X_10117_ genblk2\[3\].wave_shpr.div.quo\[17\] _04461_ _04462_ net376 _04469_ vssd1
+ vssd1 vccd1 vccd1 _00392_ sky130_fd_sc_hd__a221o_1
X_11097_ _05159_ vssd1 vssd1 vccd1 vccd1 _05160_ sky130_fd_sc_hd__inv_2
X_10048_ genblk2\[4\].wave_shpr.div.b1\[3\] _01223_ _04238_ vssd1 vssd1 vccd1 vccd1
+ _04433_ sky130_fd_sc_hd__mux2_1
Xhold90 genblk2\[5\].wave_shpr.div.quo\[7\] vssd1 vssd1 vccd1 vccd1 net308 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_89_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11843__A _02203_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_821 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11999_ _03687_ net420 _03705_ vssd1 vssd1 vccd1 vccd1 _00939_ sky130_fd_sc_hd__a21bo_1
X_13738_ clknet_leaf_46_clk net352 net119 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.quo\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_128_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09209__A1 _03714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13669_ clknet_leaf_41_clk _00982_ net125 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.acc\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_06210_ _01171_ vssd1 vssd1 vccd1 vccd1 _01172_ sky130_fd_sc_hd__clkbuf_8
X_07190_ _01953_ _01977_ _01978_ vssd1 vssd1 vccd1 vccd1 genblk1\[9\].osc.clkdiv_C.next_cnt\[11\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_14_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_143_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06141_ net14 _01112_ vssd1 vssd1 vccd1 vccd1 _01113_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_412 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_13_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06391__B _01334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_856 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_112_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09900_ _04247_ vssd1 vssd1 vccd1 vccd1 _04315_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08599__A net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09194__S _03822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_1_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09831_ _04069_ genblk1\[2\].osc.clkdiv_C.cnt\[10\] vssd1 vssd1 vccd1 vccd1 _04266_
+ sky130_fd_sc_hd__and2_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09762_ net1290 _04230_ _04039_ vssd1 vssd1 vccd1 vccd1 _04231_ sky130_fd_sc_hd__mux2_1
X_06974_ genblk1\[7\].osc.clkdiv_C.cnt\[14\] _01675_ vssd1 vssd1 vccd1 vccd1 _01810_
+ sky130_fd_sc_hd__xor2_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08713_ _03408_ _03418_ _03419_ vssd1 vssd1 vccd1 vccd1 _03420_ sky130_fd_sc_hd__and3_2
X_09693_ genblk2\[2\].wave_shpr.div.acc\[1\] genblk2\[2\].wave_shpr.div.b1\[1\] vssd1
+ vssd1 vccd1 vccd1 _04173_ sky130_fd_sc_hd__or2b_1
XFILLER_0_20_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08644_ _03340_ _03349_ _03350_ vssd1 vssd1 vccd1 vccd1 _03351_ sky130_fd_sc_hd__nand3_1
XFILLER_0_96_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_95_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_95_117 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08575_ genblk2\[11\].wave_shpr.div.fin_quo\[0\] genblk2\[11\].wave_shpr.div.fin_quo\[1\]
+ _02349_ _02351_ vssd1 vssd1 vccd1 vccd1 _03282_ sky130_fd_sc_hd__nand4_1
XTAP_1519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10369__A _04654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09448__A1 _04011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_76_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07526_ sig_norm.busy net939 _01099_ _02244_ vssd1 vssd1 vccd1 vccd1 _00026_ sky130_fd_sc_hd__o211a_1
XFILLER_0_64_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_729 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08120__A1 _01224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_147_753 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07457_ _02189_ vssd1 vssd1 vccd1 vccd1 _00017_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_8_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_119_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_797 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06408_ genblk1\[1\].osc.clkdiv_C.cnt\[3\] _01323_ _01347_ _01348_ _01351_ vssd1
+ vssd1 vccd1 vccd1 _01352_ sky130_fd_sc_hd__o221a_1
XFILLER_0_146_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_17_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_45_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07388_ _02081_ _02136_ vssd1 vssd1 vccd1 vccd1 _02138_ sky130_fd_sc_hd__nand2_1
XFILLER_0_106_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06582__A _01489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09127_ genblk2\[0\].wave_shpr.div.b1\[6\] genblk2\[0\].wave_shpr.div.acc\[6\] vssd1
+ vssd1 vccd1 vccd1 _03775_ sky130_fd_sc_hd__and2b_1
X_06339_ genblk1\[0\].osc.clkdiv_C.cnt\[11\] genblk1\[0\].osc.clkdiv_C.cnt\[10\] _01286_
+ vssd1 vssd1 vccd1 vccd1 _01290_ sky130_fd_sc_hd__and3_1
XFILLER_0_44_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09058_ _02170_ vssd1 vssd1 vccd1 vccd1 _03719_ sky130_fd_sc_hd__buf_6
X_08009_ _02713_ _02714_ _02715_ vssd1 vssd1 vccd1 vccd1 _02716_ sky130_fd_sc_hd__o21ba_1
Xhold560 genblk2\[4\].wave_shpr.div.acc\[12\] vssd1 vssd1 vccd1 vccd1 net778 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10518__B1 _04655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold571 genblk2\[9\].wave_shpr.div.i\[3\] vssd1 vssd1 vccd1 vccd1 net789 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout91_A net127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold582 genblk2\[5\].wave_shpr.div.b1\[14\] vssd1 vssd1 vccd1 vccd1 net800 sky130_fd_sc_hd__dlygate4sd3_1
X_11020_ _04995_ _05103_ vssd1 vssd1 vccd1 vccd1 _05104_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09384__B1 _03947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold593 _01165_ vssd1 vssd1 vccd1 vccd1 net811 sky130_fd_sc_hd__dlygate4sd3_1
X_12971_ clknet_leaf_125_clk net301 net71 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.quo\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_99_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11922_ genblk2\[10\].wave_shpr.div.acc\[3\] genblk2\[10\].wave_shpr.div.b1\[3\]
+ vssd1 vssd1 vccd1 vccd1 _05744_ sky130_fd_sc_hd__or2b_1
XTAP_2710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_99_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_86_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11853_ _05600_ _05557_ vssd1 vssd1 vccd1 vccd1 _05692_ sky130_fd_sc_hd__or2b_1
XTAP_2765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06476__B genblk1\[1\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10804_ net1041 _04858_ _04855_ _04954_ vssd1 vssd1 vccd1 vccd1 _00594_ sky130_fd_sc_hd__a22o_1
XFILLER_0_95_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11784_ net226 _02203_ _03693_ net416 _05641_ vssd1 vssd1 vccd1 vccd1 _00887_ sky130_fd_sc_hd__a221o_1
X_13523_ clknet_leaf_98_clk _00840_ net169 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.acc\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_10735_ _04793_ _04902_ vssd1 vssd1 vccd1 vccd1 _04903_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_103_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_94_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13454_ clknet_leaf_99_clk _00771_ net164 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.fin_quo\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_10666_ _04672_ genblk1\[5\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 _04859_
+ sky130_fd_sc_hd__and2_1
XANTENNA__06492__A _01229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12405_ net993 _06072_ _06073_ _06076_ vssd1 vssd1 vccd1 vccd1 _01073_ sky130_fd_sc_hd__a22o_1
X_13385_ clknet_leaf_83_clk _00704_ net200 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.b1\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10597_ _04823_ vssd1 vssd1 vccd1 vccd1 _00518_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08414__A2 _02468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_277 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12336_ _03689_ genblk1\[11\].osc.clkdiv_C.cnt\[13\] vssd1 vssd1 vccd1 vccd1 _06026_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_23_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12267_ _03707_ vssd1 vssd1 vccd1 vccd1 _05994_ sky130_fd_sc_hd__buf_4
XFILLER_0_10_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11218_ net563 _05246_ _05250_ net822 vssd1 vssd1 vccd1 vccd1 _00712_ sky130_fd_sc_hd__a22o_1
X_12198_ genblk2\[11\].wave_shpr.div.acc\[6\] genblk2\[11\].wave_shpr.div.b1\[6\]
+ vssd1 vssd1 vccd1 vccd1 _05936_ sky130_fd_sc_hd__or2b_1
XANTENNA__11182__B1 _04241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11149_ genblk2\[7\].wave_shpr.div.b1\[14\] genblk2\[7\].wave_shpr.div.acc\[14\]
+ vssd1 vssd1 vccd1 vccd1 _05209_ sky130_fd_sc_hd__and2b_1
XFILLER_0_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11485__A1 _03831_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06690_ genblk1\[4\].osc.clkdiv_C.cnt\[0\] _01209_ _01578_ genblk1\[4\].osc.clkdiv_C.cnt\[16\]
+ vssd1 vssd1 vccd1 vccd1 _01580_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__06667__A _01556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08360_ _02885_ _02886_ vssd1 vssd1 vccd1 vccd1 _03067_ sky130_fd_sc_hd__or2b_1
XFILLER_0_19_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07311_ genblk1\[11\].osc.clkdiv_C.cnt\[8\] _01211_ _01262_ genblk1\[11\].osc.clkdiv_C.cnt\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02075_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__11788__A2 _02203_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08291_ _02992_ _02996_ _02921_ _02997_ vssd1 vssd1 vccd1 vccd1 _02998_ sky130_fd_sc_hd__o211a_1
XFILLER_0_144_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_46_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10996__B1 _05057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07242_ genblk1\[10\].osc.clkdiv_C.cnt\[0\] _01321_ _01183_ _02023_ vssd1 vssd1 vccd1
+ vccd1 _02024_ sky130_fd_sc_hd__o22a_1
XFILLER_0_15_902 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_6_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07173_ genblk1\[9\].osc.clkdiv_C.cnt\[6\] _01965_ vssd1 vssd1 vccd1 vccd1 _01967_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_131_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08405__A2 _01578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08106__B _01574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06124_ genblk2\[1\].wave_shpr.div.done genblk2\[0\].wave_shpr.div.done genblk2\[3\].wave_shpr.div.done
+ genblk2\[2\].wave_shpr.div.done vssd1 vssd1 vccd1 vccd1 _01096_ sky130_fd_sc_hd__or4_2
XFILLER_0_131_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_631 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06967__A2 _01574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10652__A _02170_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_100_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09366__B1 _03839_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_651 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_10_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09814_ genblk2\[2\].wave_shpr.div.quo\[11\] _04253_ _04251_ net441 _04256_ vssd1
+ vssd1 vccd1 vccd1 _00302_ sky130_fd_sc_hd__a221o_1
X_09745_ genblk2\[2\].wave_shpr.div.fin_quo\[5\] genblk2\[2\].wave_shpr.div.quo\[4\]
+ _00009_ vssd1 vssd1 vccd1 vccd1 _04220_ sky130_fd_sc_hd__mux2_1
XFILLER_0_94_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06957_ genblk1\[7\].osc.clkdiv_C.cnt\[2\] _01227_ _01732_ genblk1\[7\].osc.clkdiv_C.cnt\[3\]
+ _01792_ vssd1 vssd1 vccd1 vccd1 _01793_ sky130_fd_sc_hd__a221oi_1
XFILLER_0_69_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2006 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09676_ genblk2\[2\].wave_shpr.div.acc\[17\] _04041_ vssd1 vssd1 vccd1 vccd1 _04156_
+ sky130_fd_sc_hd__or2_1
X_06888_ _01658_ _01675_ vssd1 vssd1 vccd1 vccd1 _01742_ sky130_fd_sc_hd__nand2_2
XFILLER_0_96_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2017 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2028 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2039 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08627_ _03293_ _03294_ vssd1 vssd1 vccd1 vccd1 _03334_ sky130_fd_sc_hd__or2b_1
XTAP_1305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10099__A _04269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_448 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08558_ genblk2\[8\].wave_shpr.div.fin_quo\[0\] genblk2\[8\].wave_shpr.div.fin_quo\[1\]
+ _02638_ _02223_ vssd1 vssd1 vccd1 vccd1 _03265_ sky130_fd_sc_hd__a31o_1
XFILLER_0_77_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07509_ _02228_ PWM.final_sample_in\[6\] vssd1 vssd1 vccd1 vccd1 _02229_ sky130_fd_sc_hd__and2_1
X_08489_ _03182_ _03186_ _03195_ vssd1 vssd1 vccd1 vccd1 _03196_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_135_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_91_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10520_ net763 _04657_ _04655_ _04753_ vssd1 vssd1 vccd1 vccd1 _00511_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_745 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_784 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10451_ _04595_ _04702_ vssd1 vssd1 vccd1 vccd1 _04703_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09054__C1 _03717_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_737 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_32_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13170_ clknet_leaf_126_clk _00495_ net68 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.acc\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06407__B2 _01342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10382_ genblk2\[4\].wave_shpr.div.quo\[9\] _04657_ _04655_ net251 _04658_ vssd1
+ vssd1 vccd1 vccd1 _00468_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12121_ genblk2\[10\].wave_shpr.div.acc\[11\] _05878_ _05865_ vssd1 vssd1 vccd1 vccd1
+ _05879_ sky130_fd_sc_hd__mux2_1
XANTENNA__07080__A1 genblk1\[8\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12052_ genblk2\[10\].wave_shpr.div.quo\[17\] _05823_ _05825_ net353 _05830_ vssd1
+ vssd1 vccd1 vccd1 _00966_ sky130_fd_sc_hd__a221o_1
Xhold390 genblk2\[1\].wave_shpr.div.quo\[21\] vssd1 vssd1 vccd1 vccd1 net608 sky130_fd_sc_hd__dlygate4sd3_1
X_11003_ _04987_ _05090_ vssd1 vssd1 vccd1 vccd1 _05091_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10911__A0 genblk2\[7\].wave_shpr.div.b1\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06591__B1 _01498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_82_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12954_ clknet_leaf_136_clk _00283_ net62 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.b1\[10\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1090 genblk2\[6\].wave_shpr.div.b1\[8\] vssd1 vssd1 vccd1 vccd1 net1308 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07135__A2 _01311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11905_ genblk2\[0\].wave_shpr.div.i\[3\] _02150_ _05726_ vssd1 vssd1 vccd1 vccd1
+ _05729_ sky130_fd_sc_hd__and3_1
XTAP_2540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12885_ clknet_leaf_30_clk _00216_ net97 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.quo\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_114_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11836_ _05591_ _05678_ vssd1 vssd1 vccd1 vccd1 _05679_ sky130_fd_sc_hd__xnor2_1
XTAP_2595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_97_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1872 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_138_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1883 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1894 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11767_ _05631_ genblk1\[9\].osc.clkdiv_C.cnt\[5\] vssd1 vssd1 vccd1 vccd1 _05633_
+ sky130_fd_sc_hd__and2_1
X_13506_ clknet_leaf_98_clk _00823_ net167 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.acc\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10718_ _04856_ vssd1 vssd1 vccd1 vccd1 _04890_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__07843__B1 _02527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11698_ genblk2\[9\].wave_shpr.div.b1\[9\] genblk2\[9\].wave_shpr.div.acc\[9\] vssd1
+ vssd1 vccd1 vccd1 _05590_ sky130_fd_sc_hd__and2b_1
XFILLER_0_126_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07111__A genblk1\[8\].osc.clkdiv_C.cnt\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_778 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13437_ clknet_leaf_95_clk _00756_ net161 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.acc\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_20_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10649_ _02171_ genblk2\[6\].wave_shpr.div.b1\[17\] vssd1 vssd1 vccd1 vccd1 _04852_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_113_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_153_597 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09737__S _00009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_23_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13368_ clknet_leaf_116_clk _00687_ net139 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.fin_quo\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_12319_ net342 _06014_ _06015_ net443 _06017_ vssd1 vssd1 vccd1 vccd1 _01046_ sky130_fd_sc_hd__a221o_1
X_13299_ clknet_leaf_84_clk _00620_ net202 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.b1\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_clkbuf_leaf_35_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09038__A _02336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07860_ genblk2\[1\].wave_shpr.div.fin_quo\[0\] genblk2\[1\].wave_shpr.div.fin_quo\[1\]
+ _02458_ _02459_ vssd1 vssd1 vccd1 vccd1 _02567_ sky130_fd_sc_hd__nand4_1
X_06811_ genblk1\[5\].osc.clkdiv_C.cnt\[8\] _01326_ vssd1 vssd1 vccd1 vccd1 _01683_
+ sky130_fd_sc_hd__or2_1
X_07791_ genblk1\[0\].osc.clkdiv_C.cnt\[11\] _01263_ vssd1 vssd1 vccd1 vccd1 _02498_
+ sky130_fd_sc_hd__nand2_1
X_06742_ genblk1\[4\].osc.clkdiv_C.cnt\[7\] _01620_ vssd1 vssd1 vccd1 vccd1 _01625_
+ sky130_fd_sc_hd__or2_1
XANTENNA__11458__A1 _02064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09530_ _03707_ vssd1 vssd1 vccd1 vccd1 _04055_ sky130_fd_sc_hd__clkbuf_2
XANTENNA__07126__A2 _01925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09461_ _04018_ vssd1 vssd1 vccd1 vccd1 _00187_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__06828__C genblk1\[5\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire35 _01239_ vssd1 vssd1 vccd1 vccd1 net35 sky130_fd_sc_hd__buf_2
X_06673_ _01175_ _01194_ vssd1 vssd1 vccd1 vccd1 _01563_ sky130_fd_sc_hd__or2b_1
X_08412_ _03118_ genblk2\[2\].wave_shpr.div.fin_quo\[5\] net25 vssd1 vssd1 vccd1 vccd1
+ _03119_ sky130_fd_sc_hd__or3b_1
XFILLER_0_148_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09392_ genblk2\[1\].wave_shpr.div.acc\[15\] genblk2\[1\].wave_shpr.div.b1\[15\]
+ vssd1 vssd1 vccd1 vccd1 _03956_ sky130_fd_sc_hd__or2b_1
XFILLER_0_65_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08343_ _03013_ _03029_ vssd1 vssd1 vccd1 vccd1 _03050_ sky130_fd_sc_hd__xor2_1
XFILLER_0_129_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout141_A net145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_108_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_80_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08274_ _02979_ _02404_ _02978_ _02525_ vssd1 vssd1 vccd1 vccd1 _02981_ sky130_fd_sc_hd__o31a_1
XANTENNA__07659__C _02365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_55_890 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07225_ _01994_ _02000_ _02004_ _02006_ vssd1 vssd1 vccd1 vccd1 _02007_ sky130_fd_sc_hd__or4_1
XFILLER_0_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_116_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_497 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07156_ genblk1\[9\].osc.clkdiv_C.cnt\[1\] genblk1\[9\].osc.clkdiv_C.cnt\[0\] vssd1
+ vssd1 vccd1 vccd1 _01955_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06107_ smpl_rt_clkdiv.clkDiv_inst.cnt\[5\] smpl_rt_clkdiv.clkDiv_inst.cnt\[4\] _01087_
+ vssd1 vssd1 vccd1 vccd1 _01088_ sky130_fd_sc_hd__and3_1
XANTENNA__07062__A1 genblk1\[8\].osc.clkdiv_C.cnt\[6\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_30_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07087_ _01887_ _01897_ _01898_ vssd1 vssd1 vccd1 vccd1 genblk1\[8\].osc.clkdiv_C.next_cnt\[6\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_2_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_100_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xfanout100 net101 vssd1 vssd1 vccd1 vccd1 net100 sky130_fd_sc_hd__clkbuf_2
Xfanout111 net112 vssd1 vssd1 vccd1 vccd1 net111 sky130_fd_sc_hd__clkbuf_2
Xfanout122 net126 vssd1 vssd1 vccd1 vccd1 net122 sky130_fd_sc_hd__buf_2
Xfanout133 net135 vssd1 vssd1 vccd1 vccd1 net133 sky130_fd_sc_hd__clkbuf_4
Xfanout144 net145 vssd1 vssd1 vccd1 vccd1 net144 sky130_fd_sc_hd__buf_2
Xfanout155 net157 vssd1 vssd1 vccd1 vccd1 net155 sky130_fd_sc_hd__clkbuf_4
Xfanout166 net170 vssd1 vssd1 vccd1 vccd1 net166 sky130_fd_sc_hd__clkbuf_4
Xfanout177 net180 vssd1 vssd1 vccd1 vccd1 net177 sky130_fd_sc_hd__clkbuf_4
Xfanout188 net198 vssd1 vssd1 vccd1 vccd1 net188 sky130_fd_sc_hd__buf_2
Xfanout199 net210 vssd1 vssd1 vccd1 vccd1 net199 sky130_fd_sc_hd__clkbuf_4
X_07989_ _02692_ _02693_ _02694_ _02695_ vssd1 vssd1 vccd1 vccd1 _02696_ sky130_fd_sc_hd__a211o_1
X_09728_ _04156_ _04206_ _04207_ vssd1 vssd1 vccd1 vccd1 _04208_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout54_A net58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_97_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09511__B1 _04047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09659_ _04009_ genblk2\[1\].wave_shpr.div.acc\[25\] genblk2\[1\].wave_shpr.div.acc\[26\]
+ vssd1 vssd1 vccd1 vccd1 _04145_ sky130_fd_sc_hd__or3b_1
XTAP_1102 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1113 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12670_ clknet_leaf_90_clk genblk1\[7\].osc.clkdiv_C.next_cnt\[1\] net173 vssd1 vssd1
+ vccd1 vccd1 genblk1\[7\].osc.clkdiv_C.cnt\[1\] sky130_fd_sc_hd__dfrtp_4
XTAP_1157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11621_ _05407_ _05526_ vssd1 vssd1 vccd1 vccd1 _05527_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08617__A2 _02362_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_64_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07825__B1 _02223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11552_ _05473_ _05474_ net1116 _05442_ vssd1 vssd1 vccd1 vccd1 _00822_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__08027__A _02733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_18_570 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10503_ net694 _04715_ _04722_ _04742_ vssd1 vssd1 vccd1 vccd1 _00505_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11483_ _05438_ vssd1 vssd1 vccd1 vccd1 _00789_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_107_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13222_ clknet_leaf_114_clk net880 net132 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.quo\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10434_ _04654_ vssd1 vssd1 vccd1 vccd1 _04690_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__07866__A net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10365_ _02177_ vssd1 vssd1 vccd1 vccd1 _04651_ sky130_fd_sc_hd__clkbuf_4
X_13153_ clknet_leaf_121_clk net256 net77 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.quo\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07053__B2 genblk1\[8\].osc.clkdiv_C.cnt\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_131_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12104_ genblk2\[10\].wave_shpr.div.acc\[7\] _05864_ _05865_ vssd1 vssd1 vccd1 vccd1
+ _05866_ sky130_fd_sc_hd__mux2_1
XTAP_908 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_130_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13084_ clknet_leaf_135_clk _00411_ net62 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.acc\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_919 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10296_ genblk2\[4\].wave_shpr.div.b1\[13\] genblk2\[4\].wave_shpr.div.acc\[13\]
+ vssd1 vssd1 vccd1 vccd1 _04608_ sky130_fd_sc_hd__and2b_1
XFILLER_0_20_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_20_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_109_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12035_ _05819_ genblk1\[10\].osc.clkdiv_C.cnt\[1\] vssd1 vssd1 vccd1 vccd1 _05821_
+ sky130_fd_sc_hd__and2_1
XANTENNA__08002__B1 _01666_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08553__A1 genblk2\[6\].wave_shpr.div.fin_quo\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__07817__A_N net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12937_ clknet_leaf_111_clk _00266_ net130 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.fin_quo\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_125_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10663__A2 _04853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_87_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12868_ clknet_leaf_134_clk _00199_ net60 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.b1\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11819_ _05583_ _05665_ vssd1 vssd1 vccd1 vccd1 _05666_ sky130_fd_sc_hd__xnor2_1
XANTENNA__10467__A _04651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_7_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_83_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12799_ clknet_leaf_59_clk net278 net192 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.quo\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_665 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_126_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_28_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_43_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11997__S _05802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09018__C1 _03690_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07010_ genblk1\[7\].osc.clkdiv_C.cnt\[9\] _01835_ vssd1 vssd1 vccd1 vccd1 _01837_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_113_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07776__A _01229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_52_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08241__B1 _02527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_59_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08961_ _03649_ vssd1 vssd1 vccd1 vccd1 _00056_ sky130_fd_sc_hd__clkbuf_1
X_07912_ _01233_ _02617_ _02618_ vssd1 vssd1 vccd1 vccd1 _02619_ sky130_fd_sc_hd__o21ba_1
X_08892_ sig_norm.acc\[0\] _03597_ vssd1 vssd1 vccd1 vccd1 _03598_ sky130_fd_sc_hd__xnor2_1
X_07843_ genblk2\[0\].wave_shpr.div.fin_quo\[2\] _02549_ _02527_ vssd1 vssd1 vccd1
+ vccd1 _02550_ sky130_fd_sc_hd__o21ai_1
X_07774_ genblk1\[0\].osc.clkdiv_C.cnt\[3\] _01215_ vssd1 vssd1 vccd1 vccd1 _02481_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_78_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09513_ net701 _04043_ _04047_ net755 vssd1 vssd1 vccd1 vccd1 _00210_ sky130_fd_sc_hd__a22o_1
X_06725_ _01600_ _01610_ _01611_ vssd1 vssd1 vccd1 vccd1 _01612_ sky130_fd_sc_hd__and3_1
XFILLER_0_149_634 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11761__A _03693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09444_ genblk2\[1\].wave_shpr.div.acc\[23\] genblk2\[1\].wave_shpr.div.acc\[22\]
+ genblk2\[1\].wave_shpr.div.acc\[21\] _04007_ vssd1 vssd1 vccd1 vccd1 _04008_ sky130_fd_sc_hd__or4_1
XANTENNA__10654__A2 _04853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06656_ _01523_ _01549_ vssd1 vssd1 vccd1 vccd1 _01550_ sky130_fd_sc_hd__nor2_1
XPHY_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_148_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_109_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_93_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06587_ genblk1\[3\].osc.clkdiv_C.cnt\[7\] _01494_ vssd1 vssd1 vccd1 vccd1 _01495_
+ sky130_fd_sc_hd__xnor2_1
X_09375_ _03943_ vssd1 vssd1 vccd1 vccd1 _00176_ sky130_fd_sc_hd__clkbuf_1
X_08326_ _03031_ _03032_ vssd1 vssd1 vccd1 vccd1 _03033_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_117_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_698 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_7_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08257_ _02946_ _02957_ _02951_ vssd1 vssd1 vccd1 vccd1 _02964_ sky130_fd_sc_hd__or3_1
XFILLER_0_105_715 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07208_ genblk1\[10\].osc.clkdiv_C.cnt\[9\] vssd1 vssd1 vccd1 vccd1 _01990_ sky130_fd_sc_hd__inv_2
X_08188_ _02799_ _02847_ vssd1 vssd1 vccd1 vccd1 _02895_ sky130_fd_sc_hd__or2_1
XFILLER_0_104_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11367__B1 _05248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07139_ genblk1\[9\].osc.clkdiv_C.cnt\[14\] _01246_ _01196_ _01937_ _01938_ vssd1
+ vssd1 vccd1 vccd1 _01939_ sky130_fd_sc_hd__o221a_1
XFILLER_0_132_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10150_ _04455_ vssd1 vssd1 vccd1 vccd1 _04490_ sky130_fd_sc_hd__clkbuf_4
X_10081_ _02169_ vssd1 vssd1 vccd1 vccd1 _04451_ sky130_fd_sc_hd__buf_4
XFILLER_0_100_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10342__A1 _01326_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12631__RESET_B net112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13771_ clknet_leaf_73_clk _01082_ net215 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.acc\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10983_ _05074_ genblk1\[6\].osc.clkdiv_C.cnt\[15\] vssd1 vssd1 vccd1 vccd1 _05077_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_97_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_139_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12722_ clknet_leaf_86_clk genblk1\[9\].osc.clkdiv_C.next_cnt\[17\] net183 vssd1
+ vssd1 vccd1 vccd1 genblk1\[9\].osc.clkdiv_C.cnt\[17\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_69_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_hold902_A genblk1\[5\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_69_289 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_85_738 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_38_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_790 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_139_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12653_ clknet_leaf_27_clk genblk1\[6\].osc.clkdiv_C.next_cnt\[2\] net89 vssd1 vssd1
+ vccd1 vccd1 genblk1\[6\].osc.clkdiv_C.cnt\[2\] sky130_fd_sc_hd__dfrtp_1
X_11604_ _05400_ _05362_ vssd1 vssd1 vccd1 vccd1 _05514_ sky130_fd_sc_hd__or2b_1
XFILLER_0_93_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12584_ clknet_leaf_124_clk genblk1\[2\].osc.clkdiv_C.next_cnt\[5\] net76 vssd1 vssd1
+ vccd1 vccd1 genblk1\[2\].osc.clkdiv_C.cnt\[5\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_93_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_142_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_209 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08471__B1 _02789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11535_ _05464_ genblk1\[8\].osc.clkdiv_C.cnt\[11\] vssd1 vssd1 vccd1 vccd1 _05465_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_111_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_108_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07596__A net32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_52_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_80_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_151_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_40_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11466_ net1268 _02433_ _05237_ vssd1 vssd1 vccd1 vccd1 _05430_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_33_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13205_ clknet_leaf_8_clk _00528_ net48 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.b1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_111_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10417_ _04672_ genblk1\[4\].osc.clkdiv_C.cnt\[16\] vssd1 vssd1 vccd1 vccd1 _04678_
+ sky130_fd_sc_hd__and2_1
X_11397_ genblk2\[8\].wave_shpr.div.acc\[2\] genblk2\[8\].wave_shpr.div.b1\[2\] vssd1
+ vssd1 vccd1 vccd1 _05373_ sky130_fd_sc_hd__or2b_1
XFILLER_0_96_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13136_ clknet_leaf_115_clk net465 net133 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.quo\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10348_ _04641_ vssd1 vssd1 vccd1 vccd1 _00451_ sky130_fd_sc_hd__clkbuf_1
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10279_ _04580_ _04590_ _04578_ vssd1 vssd1 vccd1 vccd1 _04591_ sky130_fd_sc_hd__o21ai_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13067_ clknet_leaf_22_clk _00394_ net93 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.quo\[19\]
+ sky130_fd_sc_hd__dfrtp_1
X_12018_ _02152_ genblk2\[10\].wave_shpr.div.busy _02206_ vssd1 vssd1 vccd1 vccd1
+ _05814_ sky130_fd_sc_hd__and3_1
XANTENNA__10333__A1 _03714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10333__B2 _03705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_88_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10896__S _04848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_139_clk clknet_4_0_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_139_clk
+ sky130_fd_sc_hd__clkbuf_16
X_06510_ _01349_ vssd1 vssd1 vccd1 vccd1 _01436_ sky130_fd_sc_hd__buf_4
XFILLER_0_48_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07490_ _02213_ vssd1 vssd1 vccd1 vccd1 _00004_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09051__A _03702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06441_ _01373_ _01380_ _01381_ vssd1 vssd1 vccd1 vccd1 genblk1\[1\].osc.clkdiv_C.next_cnt\[3\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_8_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_84_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_719 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09160_ _03806_ vssd1 vssd1 vccd1 vccd1 _00098_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06372_ genblk1\[1\].osc.clkdiv_C.cnt\[5\] _01305_ vssd1 vssd1 vccd1 vccd1 _01316_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_83_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08111_ genblk1\[4\].osc.clkdiv_C.cnt\[14\] _01361_ _02802_ _02803_ vssd1 vssd1 vccd1
+ vccd1 _02818_ sky130_fd_sc_hd__o31a_1
XFILLER_0_145_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09091_ _01201_ _03741_ vssd1 vssd1 vccd1 vccd1 _00094_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_114_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_127_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_154_681 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_4_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08042_ genblk1\[5\].osc.clkdiv_C.cnt\[14\] _01359_ vssd1 vssd1 vccd1 vccd1 _02749_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_71_487 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_114_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_101_60 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold901 genblk1\[10\].osc.clkdiv_C.cnt\[12\] vssd1 vssd1 vccd1 vccd1 net1119 sky130_fd_sc_hd__dlygate4sd3_1
Xhold912 genblk2\[6\].wave_shpr.div.i\[1\] vssd1 vssd1 vccd1 vccd1 net1130 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12010__A1 _03732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold923 sig_norm.acc\[11\] vssd1 vssd1 vccd1 vccd1 net1141 sky130_fd_sc_hd__dlygate4sd3_1
Xhold934 genblk2\[3\].wave_shpr.div.b1\[13\] vssd1 vssd1 vccd1 vccd1 net1152 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_852 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_141_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout104_A net107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold945 genblk2\[11\].wave_shpr.div.i\[3\] vssd1 vssd1 vccd1 vccd1 net1163 sky130_fd_sc_hd__dlygate4sd3_1
Xhold956 genblk2\[1\].wave_shpr.div.i\[3\] vssd1 vssd1 vccd1 vccd1 net1174 sky130_fd_sc_hd__dlygate4sd3_1
Xhold967 genblk1\[8\].osc.clkdiv_C.cnt\[7\] vssd1 vssd1 vccd1 vccd1 net1185 sky130_fd_sc_hd__dlygate4sd3_1
Xhold978 genblk1\[0\].osc.clkdiv_C.cnt\[16\] vssd1 vssd1 vccd1 vccd1 net1196 sky130_fd_sc_hd__dlygate4sd3_1
X_09993_ genblk2\[3\].wave_shpr.div.b1\[5\] genblk2\[3\].wave_shpr.div.acc\[5\] vssd1
+ vssd1 vccd1 vccd1 _04389_ sky130_fd_sc_hd__and2b_1
Xhold989 genblk1\[2\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 net1207 sky130_fd_sc_hd__dlygate4sd3_1
X_08944_ sig_norm.quo\[1\] _01098_ _03635_ vssd1 vssd1 vccd1 vccd1 _03636_ sky130_fd_sc_hd__a21o_1
XANTENNA__12313__A2 _03947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08875_ sig_norm.b1\[0\] _03578_ _03580_ vssd1 vssd1 vccd1 vccd1 _03581_ sky130_fd_sc_hd__a21o_1
XANTENNA__09190__A1 _03706_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07826_ _02531_ _02532_ vssd1 vssd1 vccd1 vccd1 _02533_ sky130_fd_sc_hd__nor2_1
XANTENNA__07740__A2 _01334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07757_ genblk2\[1\].wave_shpr.div.fin_quo\[4\] _02463_ vssd1 vssd1 vccd1 vccd1 _02464_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_79_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_149_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10088__B1 _04456_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_126_90 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06708_ _01585_ _01587_ _01590_ _01597_ vssd1 vssd1 vccd1 vccd1 _01598_ sky130_fd_sc_hd__or4b_1
X_07688_ genblk1\[10\].osc.clkdiv_C.cnt\[9\] _01215_ _02011_ genblk1\[10\].osc.clkdiv_C.cnt\[11\]
+ vssd1 vssd1 vccd1 vccd1 _02395_ sky130_fd_sc_hd__a22o_1
XFILLER_0_149_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09427_ _03961_ _03989_ _03990_ vssd1 vssd1 vccd1 vccd1 _03991_ sky130_fd_sc_hd__a21o_1
X_06639_ genblk1\[3\].osc.clkdiv_C.cnt\[7\] _01535_ genblk1\[3\].osc.clkdiv_C.cnt\[8\]
+ vssd1 vssd1 vccd1 vccd1 _01539_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_47_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09358_ genblk2\[0\].wave_shpr.div.acc\[21\] _03930_ _03931_ vssd1 vssd1 vccd1 vccd1
+ _03932_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_75_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_147 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_152_618 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_74_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08309_ genblk2\[11\].wave_shpr.div.fin_quo\[4\] _02361_ vssd1 vssd1 vccd1 vccd1
+ _03016_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_657 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08453__B1 _02526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09289_ genblk2\[0\].wave_shpr.div.acc\[4\] _03879_ _03804_ vssd1 vssd1 vccd1 vccd1
+ _03880_ sky130_fd_sc_hd__mux2_1
XFILLER_0_105_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11320_ net808 _05311_ _05283_ _05314_ vssd1 vssd1 vccd1 vccd1 _00750_ sky130_fd_sc_hd__a22o_1
XFILLER_0_34_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11251_ net231 _05255_ _05256_ net400 _05265_ vssd1 vssd1 vccd1 vccd1 _00730_ sky130_fd_sc_hd__a221o_1
XANTENNA__08205__B1 _02316_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07559__A2 genblk1\[9\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10202_ _04408_ _04529_ vssd1 vssd1 vccd1 vccd1 _04530_ sky130_fd_sc_hd__xnor2_1
X_11182_ _03732_ net389 _04241_ vssd1 vssd1 vccd1 vccd1 _00695_ sky130_fd_sc_hd__o21a_1
XANTENNA__07568__A1_N genblk1\[9\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
X_10133_ _04477_ genblk1\[3\].osc.clkdiv_C.cnt\[16\] vssd1 vssd1 vccd1 vccd1 _04478_
+ sky130_fd_sc_hd__and2_1
XANTENNA__12261__S _05802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12304__A2 _06009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10064_ net1232 _01589_ _04440_ vssd1 vssd1 vccd1 vccd1 _04442_ sky130_fd_sc_hd__mux2_1
XANTENNA__07582__C _01221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06519__B1 _01418_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09570__S _04011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07731__A2 _01360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13754_ clknet_leaf_68_clk _01065_ net212 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.acc\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10966_ _04676_ _01753_ vssd1 vssd1 vccd1 vccd1 _05068_ sky130_fd_sc_hd__nor2_1
X_12705_ clknet_leaf_86_clk genblk1\[9\].osc.clkdiv_C.next_cnt\[0\] net181 vssd1 vssd1
+ vccd1 vccd1 genblk1\[9\].osc.clkdiv_C.cnt\[0\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__13600__RESET_B net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06298__A2 _01256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13685_ clknet_leaf_63_clk _00998_ net191 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.acc\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_10897_ _05032_ vssd1 vssd1 vccd1 vccd1 _00609_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_128_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12636_ clknet_leaf_19_clk genblk1\[5\].osc.clkdiv_C.next_cnt\[3\] net109 vssd1 vssd1
+ vccd1 vccd1 genblk1\[5\].osc.clkdiv_C.cnt\[3\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_72_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_25_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_65_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_31_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_529 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12567_ clknet_leaf_27_clk genblk1\[1\].osc.clkdiv_C.next_cnt\[6\] net89 vssd1 vssd1
+ vccd1 vccd1 genblk1\[1\].osc.clkdiv_C.cnt\[6\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_108_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_136_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__10251__B1 _03855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11518_ net482 _05454_ _05449_ net506 _05455_ vssd1 vssd1 vccd1 vccd1 _00807_ sky130_fd_sc_hd__a221o_1
X_12498_ clknet_leaf_103_clk _00060_ net156 vssd1 vssd1 vccd1 vccd1 sig_norm.quo\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_41_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold208 genblk2\[1\].wave_shpr.div.quo\[18\] vssd1 vssd1 vccd1 vccd1 net426 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_151_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold219 _00401_ vssd1 vssd1 vccd1 vccd1 net437 sky130_fd_sc_hd__dlygate4sd3_1
X_11449_ _05421_ vssd1 vssd1 vccd1 vccd1 _00772_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09745__S _00009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11751__B1 _05624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13119_ clknet_leaf_2_clk _00444_ net51 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.b1\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__06222__A2 _01180_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06990_ _01823_ _01824_ vssd1 vssd1 vccd1 vccd1 genblk1\[7\].osc.clkdiv_C.next_cnt\[1\]
+ sky130_fd_sc_hd__nor2_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07970__A2 _01577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11503__B1 _05446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13759__RESET_B net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08660_ _02789_ _03177_ vssd1 vssd1 vccd1 vccd1 _03367_ sky130_fd_sc_hd__nor2_1
XANTENNA__07722__A2 _01262_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07611_ _01186_ _01437_ _01225_ genblk1\[11\].osc.clkdiv_C.cnt\[2\] vssd1 vssd1 vccd1
+ vccd1 _02318_ sky130_fd_sc_hd__o31a_1
X_08591_ _03246_ _03258_ _03296_ _03297_ vssd1 vssd1 vccd1 vccd1 _03298_ sky130_fd_sc_hd__a211o_2
X_07542_ _02254_ vssd1 vssd1 vccd1 vccd1 _00032_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07473_ genblk2\[9\].wave_shpr.div.i\[1\] _02200_ genblk2\[9\].wave_shpr.div.i\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02201_ sky130_fd_sc_hd__or3b_1
XFILLER_0_91_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09212_ _03834_ vssd1 vssd1 vccd1 vccd1 _00122_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06424_ _01365_ _01367_ vssd1 vssd1 vccd1 vccd1 _01368_ sky130_fd_sc_hd__nor2_2
XFILLER_0_29_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09227__A2 _03836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09143_ genblk2\[0\].wave_shpr.div.b1\[14\] genblk2\[0\].wave_shpr.div.acc\[14\]
+ vssd1 vssd1 vccd1 vccd1 _03791_ sky130_fd_sc_hd__and2b_1
X_06355_ genblk1\[0\].osc.clkdiv_C.cnt\[17\] _01298_ vssd1 vssd1 vccd1 vccd1 _01300_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_98_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_679 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_32_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09074_ genblk2\[0\].wave_shpr.div.b1\[13\] _01592_ _03722_ vssd1 vssd1 vccd1 vccd1
+ _03730_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06286_ _01247_ vssd1 vssd1 vccd1 vccd1 _01248_ sky130_fd_sc_hd__buf_4
X_08025_ genblk1\[6\].osc.clkdiv_C.cnt\[16\] genblk1\[6\].osc.clkdiv_C.cnt\[17\] vssd1
+ vssd1 vccd1 vccd1 _02732_ sky130_fd_sc_hd__nor2_1
Xhold720 genblk2\[9\].wave_shpr.div.acc\[6\] vssd1 vssd1 vccd1 vccd1 net938 sky130_fd_sc_hd__dlygate4sd3_1
Xhold731 genblk2\[11\].wave_shpr.div.acc\[13\] vssd1 vssd1 vccd1 vccd1 net949 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_61 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold742 genblk2\[11\].wave_shpr.div.acc\[26\] vssd1 vssd1 vccd1 vccd1 net960 sky130_fd_sc_hd__dlygate4sd3_1
Xhold753 genblk2\[4\].wave_shpr.div.acc\[7\] vssd1 vssd1 vccd1 vccd1 net971 sky130_fd_sc_hd__dlygate4sd3_1
Xhold764 genblk2\[5\].wave_shpr.div.acc\[20\] vssd1 vssd1 vccd1 vccd1 net982 sky130_fd_sc_hd__dlygate4sd3_1
Xhold775 genblk2\[11\].wave_shpr.div.acc\[14\] vssd1 vssd1 vccd1 vccd1 net993 sky130_fd_sc_hd__dlygate4sd3_1
Xhold786 genblk2\[0\].wave_shpr.div.acc\[11\] vssd1 vssd1 vccd1 vccd1 net1004 sky130_fd_sc_hd__dlygate4sd3_1
Xhold797 genblk2\[6\].wave_shpr.div.acc\[3\] vssd1 vssd1 vccd1 vccd1 net1015 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10390__A _04654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09976_ genblk2\[3\].wave_shpr.div.acc\[6\] genblk2\[3\].wave_shpr.div.b1\[6\] vssd1
+ vssd1 vccd1 vccd1 _04372_ sky130_fd_sc_hd__or2b_1
X_08927_ _01099_ _01156_ _03623_ vssd1 vssd1 vccd1 vccd1 _03624_ sky130_fd_sc_hd__and3_1
X_08858_ _03559_ _03563_ _03564_ vssd1 vssd1 vccd1 vccd1 _03565_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_99_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07809_ _02514_ _02515_ genblk2\[0\].wave_shpr.div.fin_quo\[6\] _02468_ vssd1 vssd1
+ vccd1 vccd1 _02516_ sky130_fd_sc_hd__a2bb2o_1
X_08789_ _03491_ _03495_ vssd1 vssd1 vccd1 vccd1 _03496_ sky130_fd_sc_hd__xnor2_1
X_10820_ net855 _02181_ _04962_ _03708_ vssd1 vssd1 vccd1 vccd1 _04965_ sky130_fd_sc_hd__a31o_1
XANTENNA__07204__A genblk1\[9\].osc.clkdiv_C.cnt\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10751_ _04802_ _04769_ vssd1 vssd1 vccd1 vccd1 _04915_ sky130_fd_sc_hd__or2b_1
XANTENNA__11273__A2 _05246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_39_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13470_ clknet_leaf_74_clk _00787_ net203 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.b1\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10682_ _04672_ genblk1\[5\].osc.clkdiv_C.cnt\[7\] vssd1 vssd1 vccd1 vccd1 _04868_
+ sky130_fd_sc_hd__and2_1
XANTENNA__09218__A2 _03836_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_47_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12421_ genblk2\[11\].wave_shpr.div.acc\[25\] genblk2\[11\].wave_shpr.div.acc\[24\]
+ genblk2\[11\].wave_shpr.div.acc\[26\] _05980_ vssd1 vssd1 vccd1 vccd1 _06088_ sky130_fd_sc_hd__nor4_1
XFILLER_0_118_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_50_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12352_ _03944_ _06033_ _06035_ _03947_ net1127 vssd1 vssd1 vccd1 vccd1 _01061_ sky130_fd_sc_hd__a32o_1
XANTENNA__08035__A _02221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_133_651 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11303_ net916 _05279_ _05283_ _05301_ vssd1 vssd1 vccd1 vccd1 _00746_ sky130_fd_sc_hd__a22o_1
X_12283_ genblk2\[1\].wave_shpr.div.b1\[10\] _01946_ _05994_ vssd1 vssd1 vccd1 vccd1
+ _06003_ sky130_fd_sc_hd__mux2_1
XANTENNA__08729__B2 _02468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09565__S _04011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11234_ _05249_ vssd1 vssd1 vccd1 vccd1 _05256_ sky130_fd_sc_hd__buf_2
XFILLER_0_31_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12930__D _00009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11165_ genblk2\[7\].wave_shpr.div.fin_quo\[1\] net1347 _00019_ vssd1 vssd1 vccd1
+ vccd1 _05224_ sky130_fd_sc_hd__mux2_1
XANTENNA__07952__A2 _01801_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10116_ _04465_ genblk1\[3\].osc.clkdiv_C.cnt\[8\] vssd1 vssd1 vccd1 vccd1 _04469_
+ sky130_fd_sc_hd__and2_1
X_11096_ genblk2\[6\].wave_shpr.div.i\[1\] genblk2\[6\].wave_shpr.div.i\[0\] genblk2\[6\].wave_shpr.div.i\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05159_ sky130_fd_sc_hd__and3_1
XFILLER_0_117_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10047_ _03727_ _04432_ net1075 _03687_ vssd1 vssd1 vccd1 vccd1 _00359_ sky130_fd_sc_hd__a2bb2o_1
Xhold80 genblk2\[0\].wave_shpr.div.quo\[19\] vssd1 vssd1 vccd1 vccd1 net298 sky130_fd_sc_hd__dlygate4sd3_1
Xhold91 _00551_ vssd1 vssd1 vccd1 vccd1 net309 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12020__A _05815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11998_ _05804_ vssd1 vssd1 vccd1 vccd1 _00938_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07114__A genblk1\[8\].osc.clkdiv_C.cnt\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13737_ clknet_leaf_47_clk _01048_ net119 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.quo\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10949_ _04869_ genblk1\[6\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 _05058_
+ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_70_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_70_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_27_900 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13668_ clknet_leaf_42_clk _00981_ net123 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.acc\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_144_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_39_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12619_ clknet_leaf_17_clk genblk1\[4\].osc.clkdiv_C.next_cnt\[4\] net83 vssd1 vssd1
+ vccd1 vccd1 genblk1\[4\].osc.clkdiv_C.cnt\[4\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__06691__A2 _01210_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13599_ clknet_leaf_77_clk _00914_ net208 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.acc\[23\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_14_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_06140_ _01103_ _01111_ vssd1 vssd1 vccd1 vccd1 _01112_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_108_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_54_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_41_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06979__B1 _01196_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_662 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_77_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07928__C1 genblk1\[8\].osc.clkdiv_C.cnt\[16\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08196__A2 net33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_111_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09830_ net339 _04257_ _04259_ net393 _04265_ vssd1 vssd1 vccd1 vccd1 _00309_ sky130_fd_sc_hd__a221o_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07943__A2 _01925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09761_ _01436_ _04229_ vssd1 vssd1 vccd1 vccd1 _04230_ sky130_fd_sc_hd__nand2_4
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06973_ genblk1\[7\].osc.clkdiv_C.cnt\[15\] _01363_ _01311_ genblk1\[7\].osc.clkdiv_C.cnt\[11\]
+ _01808_ vssd1 vssd1 vccd1 vccd1 _01809_ sky130_fd_sc_hd__a221o_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08712_ _03406_ _03407_ _03359_ _03381_ vssd1 vssd1 vccd1 vccd1 _03419_ sky130_fd_sc_hd__a211o_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09692_ genblk2\[2\].wave_shpr.div.b1\[1\] genblk2\[2\].wave_shpr.div.acc\[1\] vssd1
+ vssd1 vccd1 vccd1 _04172_ sky130_fd_sc_hd__or2b_1
X_08643_ _02604_ _03344_ _03348_ _02648_ vssd1 vssd1 vccd1 vccd1 _03350_ sky130_fd_sc_hd__a22o_1
XANTENNA_fanout171_A net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08574_ genblk2\[11\].wave_shpr.div.fin_quo\[0\] net33 _02350_ genblk2\[11\].wave_shpr.div.fin_quo\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03281_ sky130_fd_sc_hd__a31o_1
XFILLER_0_95_129 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07525_ _02243_ vssd1 vssd1 vccd1 vccd1 _02244_ sky130_fd_sc_hd__inv_2
XFILLER_0_88_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08656__B1 _02885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_76_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_61_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_61_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__08120__A2 _01249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_147_765 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_654 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07456_ _02186_ _02153_ genblk2\[6\].wave_shpr.div.busy vssd1 vssd1 vccd1 vccd1 _02189_
+ sky130_fd_sc_hd__and3b_1
XFILLER_0_29_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_676 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_45_741 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06407_ genblk1\[1\].osc.clkdiv_C.cnt\[16\] _01349_ _01350_ _01342_ vssd1 vssd1 vccd1
+ vccd1 _01351_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__06682__A2 _01439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10385__A _04477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07387_ _02137_ vssd1 vssd1 vccd1 vccd1 genblk1\[11\].osc.clkdiv_C.next_cnt\[13\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_09126_ _03758_ _03772_ _03773_ vssd1 vssd1 vccd1 vccd1 _03774_ sky130_fd_sc_hd__a21o_1
X_06338_ genblk1\[0\].osc.clkdiv_C.cnt\[10\] _01286_ genblk1\[0\].osc.clkdiv_C.cnt\[11\]
+ vssd1 vssd1 vccd1 vccd1 _01289_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12475__RESET_B net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06269_ _01229_ _01230_ vssd1 vssd1 vccd1 vccd1 _01231_ sky130_fd_sc_hd__nor2_4
XFILLER_0_103_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09057_ _03718_ vssd1 vssd1 vccd1 vccd1 _00083_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08008_ genblk1\[6\].osc.clkdiv_C.cnt\[3\] _01730_ _01758_ _01729_ vssd1 vssd1 vccd1
+ vccd1 _02715_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_103_879 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold550 genblk2\[8\].wave_shpr.div.b1\[7\] vssd1 vssd1 vccd1 vccd1 net768 sky130_fd_sc_hd__dlygate4sd3_1
Xhold561 genblk2\[3\].wave_shpr.div.quo\[3\] vssd1 vssd1 vccd1 vccd1 net779 sky130_fd_sc_hd__dlygate4sd3_1
Xhold572 genblk2\[3\].wave_shpr.div.acc\[10\] vssd1 vssd1 vccd1 vccd1 net790 sky130_fd_sc_hd__dlygate4sd3_1
Xhold583 genblk2\[7\].wave_shpr.div.i\[2\] vssd1 vssd1 vccd1 vccd1 net801 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09384__A1 _03944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold594 genblk2\[2\].wave_shpr.div.quo\[1\] vssd1 vssd1 vccd1 vccd1 net812 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11191__A1 _01556_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_fanout84_A net85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09959_ _04251_ _04355_ _04357_ _04253_ net711 vssd1 vssd1 vccd1 vccd1 _00346_ sky130_fd_sc_hd__a32o_1
X_12970_ clknet_leaf_113_clk net276 net128 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.quo\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_11921_ genblk2\[10\].wave_shpr.div.acc\[4\] genblk2\[10\].wave_shpr.div.b1\[4\]
+ vssd1 vssd1 vccd1 vccd1 _05743_ sky130_fd_sc_hd__and2b_1
XANTENNA__13263__RESET_B net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07860__C _02458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_99_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11852_ net799 _05684_ _05685_ _05691_ vssd1 vssd1 vccd1 vccd1 _00905_ sky130_fd_sc_hd__a22o_1
XTAP_2755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10803_ _04952_ _04949_ _04953_ vssd1 vssd1 vccd1 vccd1 _04954_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_67_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_68_866 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_877 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11783_ _05631_ genblk1\[9\].osc.clkdiv_C.cnt\[13\] vssd1 vssd1 vccd1 vccd1 _05641_
+ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_52_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_52_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_68_899 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08111__A2 _01361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13522_ clknet_leaf_79_clk _00839_ net206 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.acc\[18\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_138_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10734_ _04794_ _04773_ vssd1 vssd1 vccd1 vccd1 _04902_ sky130_fd_sc_hd__or2b_1
XFILLER_0_12_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07870__A1 _02221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13453_ clknet_leaf_99_clk _00770_ net168 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.fin_quo\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_24_903 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10665_ _02182_ vssd1 vssd1 vccd1 vccd1 _04858_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_35_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__06492__B _01182_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12404_ genblk2\[11\].wave_shpr.div.acc\[13\] _06075_ _06055_ vssd1 vssd1 vccd1 vccd1
+ _06076_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13384_ clknet_leaf_83_clk _00703_ net200 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.b1\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_10596_ genblk2\[5\].wave_shpr.div.fin_quo\[1\] genblk2\[5\].wave_shpr.div.quo\[0\]
+ _00015_ vssd1 vssd1 vccd1 vccd1 _04823_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12335_ genblk2\[11\].wave_shpr.div.quo\[21\] _06014_ _06015_ net239 _06025_ vssd1
+ vssd1 vccd1 vccd1 _01054_ sky130_fd_sc_hd__a221o_1
XFILLER_0_23_468 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_133_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12266_ _05993_ vssd1 vssd1 vccd1 vccd1 _01017_ sky130_fd_sc_hd__clkbuf_1
X_11217_ _05249_ vssd1 vssd1 vccd1 vccd1 _05250_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_120_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12197_ genblk2\[11\].wave_shpr.div.acc\[7\] genblk2\[11\].wave_shpr.div.b1\[7\]
+ vssd1 vssd1 vccd1 vccd1 _05935_ sky130_fd_sc_hd__or2b_1
XANTENNA__11182__A1 _03732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11148_ _05168_ _05206_ _05207_ vssd1 vssd1 vccd1 vccd1 _05208_ sky130_fd_sc_hd__a21o_1
X_11079_ genblk2\[6\].wave_shpr.div.acc\[22\] _05146_ vssd1 vssd1 vccd1 vccd1 _05148_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__07138__B1 genblk1\[9\].osc.clkdiv_C.cnt\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06667__B _01344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_721 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_43_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_43_clk sky130_fd_sc_hd__clkbuf_16
X_07310_ genblk1\[11\].osc.clkdiv_C.cnt\[10\] _02002_ vssd1 vssd1 vccd1 vccd1 _02074_
+ sky130_fd_sc_hd__xnor2_1
X_08290_ _02747_ _02919_ _02920_ vssd1 vssd1 vccd1 vccd1 _02997_ sky130_fd_sc_hd__a21o_1
XANTENNA__09850__A2 _04214_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10996__A1 _05055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_9_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_129_798 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07241_ genblk1\[10\].osc.clkdiv_C.cnt\[12\] vssd1 vssd1 vccd1 vccd1 _02023_ sky130_fd_sc_hd__inv_2
XFILLER_0_128_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_914 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_27_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_54_571 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07172_ _01953_ _01965_ _01966_ vssd1 vssd1 vccd1 vccd1 genblk1\[9\].osc.clkdiv_C.next_cnt\[5\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_82_891 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06123_ genblk2\[5\].wave_shpr.div.done genblk2\[4\].wave_shpr.div.done genblk2\[7\].wave_shpr.div.done
+ genblk2\[6\].wave_shpr.div.done vssd1 vssd1 vccd1 vccd1 _01095_ sky130_fd_sc_hd__or4_4
XFILLER_0_14_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_30_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_100_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_111_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__13774__RESET_B net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09813_ _04058_ _01414_ vssd1 vssd1 vccd1 vccd1 _04256_ sky130_fd_sc_hd__nor2_1
XANTENNA__10920__A1 _02433_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__11764__A _02155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09744_ _04219_ vssd1 vssd1 vccd1 vccd1 _00269_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07961__B _01360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06956_ genblk1\[7\].osc.clkdiv_C.cnt\[11\] _01311_ _01732_ genblk1\[7\].osc.clkdiv_C.cnt\[3\]
+ vssd1 vssd1 vccd1 vccd1 _01792_ sky130_fd_sc_hd__o22ai_1
X_09675_ net285 _04154_ _04155_ vssd1 vssd1 vccd1 vccd1 _00264_ sky130_fd_sc_hd__a21oi_1
X_06887_ genblk1\[6\].osc.clkdiv_C.cnt\[1\] _01738_ _01740_ vssd1 vssd1 vccd1 vccd1
+ _01741_ sky130_fd_sc_hd__a21bo_1
XTAP_2007 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2018 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2029 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08626_ _03331_ _03332_ _03298_ vssd1 vssd1 vccd1 vccd1 _03333_ sky130_fd_sc_hd__nand3b_2
XTAP_1306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_1317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08557_ genblk2\[8\].wave_shpr.div.fin_quo\[0\] _02638_ genblk2\[8\].wave_shpr.div.fin_quo\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03264_ sky130_fd_sc_hd__a21oi_1
Xclkbuf_leaf_34_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_34_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07508_ PWM.counter\[6\] vssd1 vssd1 vccd1 vccd1 _02228_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_696 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08488_ _03187_ _03194_ vssd1 vssd1 vccd1 vccd1 _03195_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_135_735 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07439_ _02147_ _02176_ vssd1 vssd1 vccd1 vccd1 _02177_ sky130_fd_sc_hd__nor2_1
XFILLER_0_107_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_134_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_18_796 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10450_ _04596_ _04575_ vssd1 vssd1 vccd1 vccd1 _04702_ sky130_fd_sc_hd__or2b_1
XFILLER_0_17_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09109_ genblk2\[0\].wave_shpr.div.acc\[6\] genblk2\[0\].wave_shpr.div.b1\[6\] vssd1
+ vssd1 vccd1 vccd1 _03757_ sky130_fd_sc_hd__or2b_1
XFILLER_0_150_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_21_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10381_ _04477_ genblk1\[4\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 _04658_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_103_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_32_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_60_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_103_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12120_ _05767_ _05877_ vssd1 vssd1 vccd1 vccd1 _05878_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_102_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12051_ _03833_ _02003_ vssd1 vssd1 vccd1 vccd1 _05830_ sky130_fd_sc_hd__nor2_1
XFILLER_0_2_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold380 genblk2\[0\].wave_shpr.div.quo\[9\] vssd1 vssd1 vccd1 vccd1 net598 sky130_fd_sc_hd__dlygate4sd3_1
Xhold391 genblk2\[6\].wave_shpr.div.quo\[22\] vssd1 vssd1 vccd1 vccd1 net609 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11002_ _04988_ _04980_ vssd1 vssd1 vccd1 vccd1 _05090_ sky130_fd_sc_hd__or2b_1
XANTENNA__10911__A1 _04444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12953_ clknet_leaf_136_clk _00282_ net62 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.b1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1080 genblk2\[3\].wave_shpr.div.b1\[8\] vssd1 vssd1 vccd1 vccd1 net1298 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1091 genblk2\[4\].wave_shpr.div.quo\[0\] vssd1 vssd1 vccd1 vccd1 net1309 sky130_fd_sc_hd__dlygate4sd3_1
X_11904_ _00000_ _05726_ net1158 vssd1 vssd1 vccd1 vccd1 _05728_ sky130_fd_sc_hd__a21oi_1
XTAP_2530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12884_ clknet_leaf_30_clk net461 net97 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.quo\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_87_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11219__A2 _05246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11835_ _05592_ _05561_ vssd1 vssd1 vccd1 vccd1 _05678_ sky130_fd_sc_hd__or2b_1
XTAP_1840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_25_clk clknet_4_4_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_25_clk sky130_fd_sc_hd__clkbuf_16
XTAP_2596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07599__A _02261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_95_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1873 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_324 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_95_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1884 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11766_ genblk2\[9\].wave_shpr.div.quo\[13\] _05628_ _05629_ net243 _05632_ vssd1
+ vssd1 vccd1 vccd1 _00878_ sky130_fd_sc_hd__a221o_1
XFILLER_0_28_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_83_655 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1895 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13505_ clknet_leaf_98_clk _00822_ net167 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.acc\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10717_ net961 _04886_ _04857_ _04889_ vssd1 vssd1 vccd1 vccd1 _00572_ sky130_fd_sc_hd__a22o_1
X_11697_ _05563_ _05587_ _05588_ vssd1 vssd1 vccd1 vccd1 _05589_ sky130_fd_sc_hd__a21o_1
X_13436_ clknet_leaf_95_clk _00755_ net159 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.acc\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07111__B genblk1\[8\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_919 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10648_ _03726_ _04851_ _03736_ vssd1 vssd1 vccd1 vccd1 _00541_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_70_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_113_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_125_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_140_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13367_ clknet_leaf_116_clk _00686_ net139 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.fin_quo\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_106_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10579_ _04767_ _04805_ _04806_ vssd1 vssd1 vccd1 vccd1 _04807_ sky130_fd_sc_hd__a21o_1
X_12318_ _05835_ genblk1\[11\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 _06017_
+ sky130_fd_sc_hd__and2_1
X_13298_ clknet_leaf_84_clk _00619_ net202 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.b1\[10\]
+ sky130_fd_sc_hd__dfrtp_1
X_12249_ genblk2\[11\].wave_shpr.div.fin_quo\[2\] net769 _00005_ vssd1 vssd1 vccd1
+ vccd1 _05985_ sky130_fd_sc_hd__mux2_1
XANTENNA__09038__B net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12352__B1 _03947_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10902__A1 _01923_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06810_ genblk1\[5\].osc.clkdiv_C.cnt\[8\] _01326_ vssd1 vssd1 vccd1 vccd1 _01682_
+ sky130_fd_sc_hd__nand2_1
X_07790_ genblk1\[0\].osc.clkdiv_C.cnt\[10\] _01996_ _01801_ vssd1 vssd1 vccd1 vccd1
+ _02497_ sky130_fd_sc_hd__or3_1
XFILLER_0_3_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06741_ genblk1\[4\].osc.clkdiv_C.cnt\[7\] _01620_ vssd1 vssd1 vccd1 vccd1 _01624_
+ sky130_fd_sc_hd__nand2_1
Xwire25 _03112_ vssd1 vssd1 vccd1 vccd1 net25 sky130_fd_sc_hd__clkbuf_2
X_09460_ genblk2\[1\].wave_shpr.div.fin_quo\[6\] genblk2\[1\].wave_shpr.div.quo\[5\]
+ _00007_ vssd1 vssd1 vccd1 vccd1 _04018_ sky130_fd_sc_hd__mux2_1
X_06672_ genblk1\[4\].osc.clkdiv_C.cnt\[3\] _01326_ _01498_ genblk1\[4\].osc.clkdiv_C.cnt\[14\]
+ vssd1 vssd1 vccd1 vccd1 _01562_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__08893__A _01099_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08411_ genblk2\[2\].wave_shpr.div.fin_quo\[4\] _03117_ vssd1 vssd1 vccd1 vccd1 _03118_
+ sky130_fd_sc_hd__or2_1
X_09391_ genblk2\[1\].wave_shpr.div.acc\[16\] genblk2\[1\].wave_shpr.div.b1\[16\]
+ vssd1 vssd1 vccd1 vccd1 _03955_ sky130_fd_sc_hd__and2b_1
Xclkbuf_leaf_16_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_16_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__10418__B1 _04654_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08342_ _03041_ _03042_ _03047_ vssd1 vssd1 vccd1 vccd1 _03049_ sky130_fd_sc_hd__a21o_1
XFILLER_0_19_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_80_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_86_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_129_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08273_ _02404_ _02978_ _02979_ vssd1 vssd1 vccd1 vccd1 _02980_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_74_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08117__B _01326_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07224_ genblk1\[10\].osc.clkdiv_C.cnt\[11\] _02005_ vssd1 vssd1 vccd1 vccd1 _02006_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_80_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07155_ _01952_ vssd1 vssd1 vccd1 vccd1 _01954_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_563 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06106_ smpl_rt_clkdiv.clkDiv_inst.cnt\[3\] _01086_ vssd1 vssd1 vccd1 vccd1 _01087_
+ sky130_fd_sc_hd__and2_1
XANTENNA__07062__A2 _01249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07086_ genblk1\[8\].osc.clkdiv_C.cnt\[6\] _01895_ vssd1 vssd1 vccd1 vccd1 _01898_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_112_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_2_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_1_181 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xfanout101 net107 vssd1 vssd1 vccd1 vccd1 net101 sky130_fd_sc_hd__clkbuf_2
XANTENNA__12343__B1 _03941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout112 net127 vssd1 vssd1 vccd1 vccd1 net112 sky130_fd_sc_hd__buf_2
Xfanout123 net125 vssd1 vssd1 vccd1 vccd1 net123 sky130_fd_sc_hd__clkbuf_4
Xfanout134 net135 vssd1 vssd1 vccd1 vccd1 net134 sky130_fd_sc_hd__clkbuf_4
Xfanout145 net171 vssd1 vssd1 vccd1 vccd1 net145 sky130_fd_sc_hd__clkbuf_4
Xfanout156 net157 vssd1 vssd1 vccd1 vccd1 net156 sky130_fd_sc_hd__clkbuf_4
Xfanout167 net170 vssd1 vssd1 vccd1 vccd1 net167 sky130_fd_sc_hd__clkbuf_4
XANTENNA__10602__S _00015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout178 net180 vssd1 vssd1 vccd1 vccd1 net178 sky130_fd_sc_hd__clkbuf_2
Xfanout189 net191 vssd1 vssd1 vccd1 vccd1 net189 sky130_fd_sc_hd__clkbuf_4
X_07988_ _02217_ _02553_ genblk2\[7\].wave_shpr.div.fin_quo\[7\] vssd1 vssd1 vccd1
+ vccd1 _02695_ sky130_fd_sc_hd__and3_1
XANTENNA__06588__A _01437_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09727_ genblk2\[2\].wave_shpr.div.acc\[17\] _04041_ vssd1 vssd1 vccd1 vccd1 _04207_
+ sky130_fd_sc_hd__and2_1
X_06939_ genblk1\[6\].osc.clkdiv_C.cnt\[12\] genblk1\[6\].osc.clkdiv_C.cnt\[11\] _01777_
+ vssd1 vssd1 vccd1 vccd1 _01781_ sky130_fd_sc_hd__and3_1
XFILLER_0_96_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10657__B1 _04857_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09511__B2 net764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09658_ net1228 _04048_ _04045_ _04144_ vssd1 vssd1 vccd1 vccd1 _00258_ sky130_fd_sc_hd__a22o_1
XTAP_1103 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1114 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout47_A net50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08609_ _03314_ _02789_ _03315_ vssd1 vssd1 vccd1 vccd1 _03316_ sky130_fd_sc_hd__o21a_1
XFILLER_0_139_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1125 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09589_ _03984_ _03964_ vssd1 vssd1 vccd1 vccd1 _04093_ sky130_fd_sc_hd__or2b_1
XTAP_1147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11620_ _05408_ _05358_ vssd1 vssd1 vccd1 vccd1 _05526_ sky130_fd_sc_hd__or2b_1
XFILLER_0_154_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12490__RESET_B net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_37_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09814__A2 _04253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_38_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11551_ genblk2\[8\].wave_shpr.div.b1\[0\] genblk2\[8\].wave_shpr.div.acc\[0\] _05417_
+ _05471_ vssd1 vssd1 vccd1 vccd1 _05474_ sky130_fd_sc_hd__a31o_1
XFILLER_0_9_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10502_ _04740_ _04741_ vssd1 vssd1 vccd1 vccd1 _04742_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11482_ genblk2\[9\].wave_shpr.div.b1\[12\] _02656_ _05433_ vssd1 vssd1 vccd1 vccd1
+ _05438_ sky130_fd_sc_hd__mux2_1
X_13221_ clknet_leaf_114_clk _00544_ net132 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.quo\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_850 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10433_ net1068 _04683_ _04656_ _04689_ vssd1 vssd1 vccd1 vccd1 _00488_ sky130_fd_sc_hd__a22o_1
XFILLER_0_21_703 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_33_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13152_ clknet_leaf_17_clk _00477_ net80 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.quo\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10364_ _04650_ vssd1 vssd1 vccd1 vccd1 _00458_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_21_747 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12103_ _05786_ vssd1 vssd1 vccd1 vccd1 _05865_ sky130_fd_sc_hd__buf_4
XFILLER_0_20_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_20_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_909 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13083_ clknet_leaf_135_clk _00410_ net61 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.acc\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_10295_ _04570_ _04605_ _04606_ vssd1 vssd1 vccd1 vccd1 _04607_ sky130_fd_sc_hd__a21o_1
X_12034_ net432 _05818_ _05816_ genblk2\[10\].wave_shpr.div.quo\[8\] _05820_ vssd1
+ vssd1 vccd1 vccd1 _00958_ sky130_fd_sc_hd__a221o_1
XFILLER_0_109_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08553__A2 genblk2\[6\].wave_shpr.div.fin_quo\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_125_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10648__B1 _03736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12936_ clknet_leaf_113_clk _00265_ net130 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.fin_quo\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_87_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12867_ clknet_leaf_134_clk _00198_ net60 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.b1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_2393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11818_ _05584_ _05565_ vssd1 vssd1 vccd1 vccd1 _05665_ sky130_fd_sc_hd__or2b_1
XFILLER_0_56_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09266__B1 _03838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12798_ clknet_leaf_57_clk _00131_ net183 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.quo\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09805__A2 _04248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11749_ net586 _05623_ _05624_ net700 vssd1 vssd1 vccd1 vccd1 _00869_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_50_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_56_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_55_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10820__B1 _03708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_114_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_198 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_119_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06961__A _01432_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_413 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13419_ clknet_leaf_91_clk _00738_ net147 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.acc\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07776__B _01359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_141_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11376__A1 _05248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_113_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_121_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08960_ sig_norm.quo\[5\] _03648_ _00024_ vssd1 vssd1 vccd1 vccd1 _03649_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_5_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_5_clk sky130_fd_sc_hd__clkbuf_16
X_07911_ _01228_ _01308_ _01440_ _01889_ _01879_ vssd1 vssd1 vccd1 vccd1 _02618_ sky130_fd_sc_hd__o41a_1
X_08891_ sig_norm.b1\[0\] _03596_ vssd1 vssd1 vccd1 vccd1 _03597_ sky130_fd_sc_hd__nand2_1
X_07842_ genblk2\[0\].wave_shpr.div.fin_quo\[0\] genblk2\[0\].wave_shpr.div.fin_quo\[1\]
+ _02510_ vssd1 vssd1 vccd1 vccd1 _02549_ sky130_fd_sc_hd__o21a_1
XANTENNA__11422__A_N genblk2\[8\].wave_shpr.div.b1\[12\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07773_ genblk1\[0\].osc.clkdiv_C.cnt\[2\] _01556_ _01564_ _01190_ genblk1\[0\].osc.clkdiv_C.cnt\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02480_ sky130_fd_sc_hd__a32o_1
XFILLER_0_79_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09512_ genblk2\[1\].wave_shpr.div.quo\[2\] _04043_ _04047_ net684 vssd1 vssd1 vccd1
+ vccd1 _00209_ sky130_fd_sc_hd__a22o_1
X_06724_ genblk1\[4\].osc.clkdiv_C.cnt\[3\] _01605_ vssd1 vssd1 vccd1 vccd1 _01611_
+ sky130_fd_sc_hd__or2_1
XANTENNA__12930__RESET_B net150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_79_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_149_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09443_ genblk2\[1\].wave_shpr.div.acc\[20\] genblk2\[1\].wave_shpr.div.acc\[19\]
+ _04006_ vssd1 vssd1 vccd1 vccd1 _04007_ sky130_fd_sc_hd__or3_1
X_06655_ genblk1\[3\].osc.clkdiv_C.cnt\[14\] _01547_ vssd1 vssd1 vccd1 vccd1 _01549_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_93_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09374_ _03941_ _03942_ genblk2\[11\].wave_shpr.div.i\[0\] vssd1 vssd1 vccd1 vccd1
+ _03943_ sky130_fd_sc_hd__mux2_1
X_06586_ _01342_ _01248_ vssd1 vssd1 vccd1 vccd1 _01494_ sky130_fd_sc_hd__nor2_4
XFILLER_0_47_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08325_ genblk2\[8\].wave_shpr.div.fin_quo\[4\] _02638_ _02640_ _02223_ vssd1 vssd1
+ vccd1 vccd1 _03032_ sky130_fd_sc_hd__a31o_1
XFILLER_0_90_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_129_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_145_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_34_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10811__B1 _04858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08256_ _02742_ _02962_ _02745_ vssd1 vssd1 vccd1 vccd1 _02963_ sky130_fd_sc_hd__o21a_1
XFILLER_0_144_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07207_ net1194 _01988_ vssd1 vssd1 vccd1 vccd1 genblk1\[9\].osc.clkdiv_C.next_cnt\[17\]
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__11489__A _02171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08187_ _02890_ _02891_ _02892_ _02893_ vssd1 vssd1 vccd1 vccd1 _02894_ sky130_fd_sc_hd__a31o_1
XANTENNA__10393__A _04477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_81_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_120_708 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_15_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07138_ genblk1\[9\].osc.clkdiv_C.cnt\[14\] _01246_ genblk1\[9\].osc.clkdiv_C.cnt\[17\]
+ vssd1 vssd1 vccd1 vccd1 _01938_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_112_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07069_ _01886_ vssd1 vssd1 vccd1 vccd1 _01887_ sky130_fd_sc_hd__clkbuf_4
X_10080_ _04450_ vssd1 vssd1 vccd1 vccd1 _00374_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_96_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13770_ clknet_leaf_71_clk _01081_ net215 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.acc\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_10982_ net385 _05051_ _05054_ net609 _05076_ vssd1 vssd1 vccd1 vccd1 _00650_ sky130_fd_sc_hd__a221o_1
XFILLER_0_97_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_706 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12721_ clknet_leaf_86_clk genblk1\[9\].osc.clkdiv_C.next_cnt\[16\] net183 vssd1
+ vssd1 vccd1 vccd1 genblk1\[9\].osc.clkdiv_C.cnt\[16\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_97_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_38_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_84_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12652_ clknet_leaf_27_clk genblk1\[6\].osc.clkdiv_C.next_cnt\[1\] net89 vssd1 vssd1
+ vccd1 vccd1 genblk1\[6\].osc.clkdiv_C.cnt\[1\] sky130_fd_sc_hd__dfrtp_4
XANTENNA_clkbuf_leaf_34_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_37_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08038__A net12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_806 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11603_ net833 _05507_ _05484_ _05513_ vssd1 vssd1 vccd1 vccd1 _00834_ sky130_fd_sc_hd__a22o_1
X_12583_ clknet_leaf_124_clk genblk1\[2\].osc.clkdiv_C.next_cnt\[4\] net72 vssd1 vssd1
+ vccd1 vccd1 genblk1\[2\].osc.clkdiv_C.cnt\[4\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_93_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11534_ _04268_ vssd1 vssd1 vccd1 vccd1 _05464_ sky130_fd_sc_hd__buf_2
XFILLER_0_20_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_658 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_151_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_80_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11465_ _05429_ vssd1 vssd1 vccd1 vccd1 _00780_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_49_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13204_ clknet_leaf_8_clk _00527_ net48 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.b1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_10416_ net714 _04651_ _04654_ net698 _04677_ vssd1 vssd1 vccd1 vccd1 _00483_ sky130_fd_sc_hd__a221o_1
XFILLER_0_33_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_0_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11396_ genblk2\[8\].wave_shpr.div.acc\[3\] genblk2\[8\].wave_shpr.div.b1\[3\] vssd1
+ vssd1 vccd1 vccd1 _05372_ sky130_fd_sc_hd__or2b_1
X_13135_ clknet_leaf_114_clk net419 net133 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.quo\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_0_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10347_ net1283 _01658_ _04637_ vssd1 vssd1 vccd1 vccd1 _04641_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12307__B1 _06010_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13066_ clknet_leaf_22_clk net452 net93 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.quo\[18\]
+ sky130_fd_sc_hd__dfrtp_1
X_10278_ _04581_ _04588_ _04589_ vssd1 vssd1 vccd1 vccd1 _04590_ sky130_fd_sc_hd__a21oi_1
X_12017_ _05812_ vssd1 vssd1 vccd1 vccd1 _05813_ sky130_fd_sc_hd__buf_4
XANTENNA_clkbuf_leaf_107_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xmax_cap1 _05138_ vssd1 vssd1 vccd1 vccd1 net1350 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_88_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_49_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11294__B1 _05283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12919_ clknet_leaf_39_clk _00250_ net115 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.acc\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06675__B _01564_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06440_ genblk1\[1\].osc.clkdiv_C.cnt\[3\] _01378_ vssd1 vssd1 vccd1 vccd1 _01381_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_0_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06371_ _01307_ _01311_ _01312_ genblk1\[1\].osc.clkdiv_C.cnt\[11\] _01314_ vssd1
+ vssd1 vccd1 vccd1 _01315_ sky130_fd_sc_hd__a221o_1
XFILLER_0_127_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_145_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_16_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08110_ genblk1\[4\].osc.clkdiv_C.cnt\[10\] _01313_ _02809_ _02810_ _02816_ vssd1
+ vssd1 vccd1 vccd1 _02817_ sky130_fd_sc_hd__o311a_1
XFILLER_0_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_44_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__13547__RESET_B net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_71_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_09090_ _03739_ _03740_ vssd1 vssd1 vccd1 vccd1 _03741_ sky130_fd_sc_hd__nor2b_1
XFILLER_0_142_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_32_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_733 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_08041_ genblk1\[5\].osc.clkdiv_C.cnt\[15\] _01576_ vssd1 vssd1 vccd1 vccd1 _02748_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_153_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_24_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold902 genblk1\[5\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 net1120 sky130_fd_sc_hd__dlygate4sd3_1
Xhold913 sig_norm.acc\[0\] vssd1 vssd1 vccd1 vccd1 net1131 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_114_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_12_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xhold924 PWM.final_sample_in\[7\] vssd1 vssd1 vccd1 vccd1 net1142 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_clkbuf_4_6_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold935 genblk2\[10\].wave_shpr.div.i\[3\] vssd1 vssd1 vccd1 vccd1 net1153 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_864 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold946 genblk2\[8\].wave_shpr.div.i\[3\] vssd1 vssd1 vccd1 vccd1 net1164 sky130_fd_sc_hd__dlygate4sd3_1
Xhold957 genblk2\[0\].wave_shpr.div.acc\[20\] vssd1 vssd1 vccd1 vccd1 net1175 sky130_fd_sc_hd__dlygate4sd3_1
Xhold968 genblk2\[4\].wave_shpr.div.b1\[9\] vssd1 vssd1 vccd1 vccd1 net1186 sky130_fd_sc_hd__dlygate4sd3_1
X_09992_ _04376_ _04387_ _04374_ vssd1 vssd1 vccd1 vccd1 _04388_ sky130_fd_sc_hd__o21ai_1
Xhold979 genblk2\[2\].wave_shpr.div.quo\[6\] vssd1 vssd1 vccd1 vccd1 net1197 sky130_fd_sc_hd__dlygate4sd3_1
X_08943_ _03545_ _03634_ _03546_ _01155_ vssd1 vssd1 vccd1 vccd1 _03635_ sky130_fd_sc_hd__o211a_1
XANTENNA__11756__B genblk1\[9\].osc.clkdiv_C.cnt\[1\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_4_15_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_15_0_clk sky130_fd_sc_hd__clkbuf_8
X_08874_ _03577_ _03579_ vssd1 vssd1 vccd1 vccd1 _03580_ sky130_fd_sc_hd__nand2_1
XFILLER_0_99_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07725__B1 _01313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07825_ genblk2\[0\].wave_shpr.div.fin_quo\[3\] _02510_ _02511_ _02223_ vssd1 vssd1
+ vccd1 vccd1 _02532_ sky130_fd_sc_hd__a31o_1
X_07756_ genblk2\[1\].wave_shpr.div.fin_quo\[2\] genblk2\[1\].wave_shpr.div.fin_quo\[3\]
+ _02462_ vssd1 vssd1 vccd1 vccd1 _02463_ sky130_fd_sc_hd__or3_1
XANTENNA__10088__B2 net794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06707_ genblk1\[4\].osc.clkdiv_C.cnt\[7\] _01304_ _01593_ _01594_ _01596_ vssd1
+ vssd1 vccd1 vccd1 _01597_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_79_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_67_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10388__A _04477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07687_ genblk1\[10\].osc.clkdiv_C.cnt\[11\] _02011_ _02005_ genblk1\[10\].osc.clkdiv_C.cnt\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02394_ sky130_fd_sc_hd__o22ai_2
X_09426_ genblk2\[1\].wave_shpr.div.b1\[10\] genblk2\[1\].wave_shpr.div.acc\[10\]
+ vssd1 vssd1 vccd1 vccd1 _03990_ sky130_fd_sc_hd__and2b_1
X_06638_ genblk1\[3\].osc.clkdiv_C.cnt\[8\] genblk1\[3\].osc.clkdiv_C.cnt\[7\] _01535_
+ vssd1 vssd1 vccd1 vccd1 _01538_ sky130_fd_sc_hd__and3_1
XFILLER_0_66_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09357_ genblk2\[0\].wave_shpr.div.acc\[21\] genblk2\[0\].wave_shpr.div.acc\[20\]
+ _03800_ net1352 vssd1 vssd1 vccd1 vccd1 _03931_ sky130_fd_sc_hd__or4_1
XFILLER_0_136_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_75_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06569_ net1167 _01476_ _01479_ vssd1 vssd1 vccd1 vccd1 genblk1\[2\].osc.clkdiv_C.next_cnt\[15\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_136_159 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07697__A _02403_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08308_ genblk2\[11\].wave_shpr.div.fin_quo\[3\] _02349_ _02351_ _02353_ _02222_
+ vssd1 vssd1 vccd1 vccd1 _03015_ sky130_fd_sc_hd__a41o_1
XFILLER_0_145_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09288_ _03878_ _03770_ vssd1 vssd1 vccd1 vccd1 _03879_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_117_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_145_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06464__B1 genblk1\[1\].osc.clkdiv_C.cnt\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08239_ _02646_ _02647_ vssd1 vssd1 vccd1 vccd1 _02946_ sky130_fd_sc_hd__or2_1
XFILLER_0_105_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11250_ _05260_ genblk1\[7\].osc.clkdiv_C.cnt\[10\] vssd1 vssd1 vccd1 vccd1 _05265_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_105_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10201_ _04409_ _04363_ vssd1 vssd1 vccd1 vccd1 _04529_ sky130_fd_sc_hd__or2b_1
X_11181_ _03819_ _01242_ _02064_ _05231_ vssd1 vssd1 vccd1 vccd1 _00694_ sky130_fd_sc_hd__o31a_1
XFILLER_0_31_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_101_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10132_ _04268_ vssd1 vssd1 vccd1 vccd1 _04477_ sky130_fd_sc_hd__buf_2
XFILLER_0_101_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10063_ _04441_ vssd1 vssd1 vccd1 vccd1 _00366_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10062__S _04440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07731__A3 net37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_98_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_85_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13753_ clknet_leaf_68_clk _01064_ net211 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.acc\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10965_ net594 _05062_ _05064_ net498 _05067_ vssd1 vssd1 vccd1 vccd1 _00642_ sky130_fd_sc_hd__a221o_1
X_12704_ clknet_leaf_89_clk genblk1\[8\].osc.clkdiv_C.next_cnt\[17\] net173 vssd1
+ vssd1 vccd1 vccd1 genblk1\[8\].osc.clkdiv_C.cnt\[17\] sky130_fd_sc_hd__dfrtp_1
X_13684_ clknet_leaf_63_clk _00997_ net191 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.acc\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_430 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10896_ genblk2\[7\].wave_shpr.div.b1\[0\] _01514_ _04848_ vssd1 vssd1 vccd1 vccd1
+ _05032_ sky130_fd_sc_hd__mux2_1
X_12635_ clknet_leaf_16_clk genblk1\[5\].osc.clkdiv_C.next_cnt\[2\] net74 vssd1 vssd1
+ vccd1 vccd1 genblk1\[5\].osc.clkdiv_C.cnt\[2\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_122_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_109_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12566_ clknet_leaf_28_clk genblk1\[1\].osc.clkdiv_C.next_cnt\[5\] net89 vssd1 vssd1
+ vccd1 vccd1 genblk1\[1\].osc.clkdiv_C.cnt\[5\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_31_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_25_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07400__A net1220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_41_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11517_ _05450_ genblk1\[8\].osc.clkdiv_C.cnt\[3\] vssd1 vssd1 vccd1 vccd1 _05455_
+ sky130_fd_sc_hd__and2_1
X_12497_ clknet_leaf_102_clk _00059_ net156 vssd1 vssd1 vccd1 vccd1 sig_norm.quo\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12018__A _02152_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_831 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold209 _00225_ vssd1 vssd1 vccd1 vccd1 net427 sky130_fd_sc_hd__dlygate4sd3_1
X_11448_ genblk2\[8\].wave_shpr.div.fin_quo\[3\] net1337 _00021_ vssd1 vssd1 vccd1
+ vccd1 _05421_ sky130_fd_sc_hd__mux2_1
XFILLER_0_151_685 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_150_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11379_ _03690_ _05355_ _05356_ vssd1 vssd1 vccd1 vccd1 _00767_ sky130_fd_sc_hd__nor3_1
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13118_ clknet_leaf_125_clk _00443_ net69 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.b1\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13049_ clknet_leaf_112_clk _00376_ net132 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.quo\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08380__B1 _02425_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_89_820 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07610_ genblk1\[11\].osc.clkdiv_C.cnt\[7\] _01211_ vssd1 vssd1 vccd1 vccd1 _02317_
+ sky130_fd_sc_hd__nand2_1
X_08590_ _03275_ _03276_ _03295_ vssd1 vssd1 vccd1 vccd1 _03297_ sky130_fd_sc_hd__a21oi_1
XANTENNA__09062__A _03701_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07541_ PWM.final_sample_in\[2\] net1102 PWM.start vssd1 vssd1 vccd1 vccd1 _02254_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_88_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_76_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_88_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07472_ genblk2\[9\].wave_shpr.div.i\[2\] genblk2\[9\].wave_shpr.div.i\[3\] genblk2\[9\].wave_shpr.div.i\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02200_ sky130_fd_sc_hd__nand3b_1
XANTENNA__08683__B2 _02468_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09211_ _03833_ net1302 vssd1 vssd1 vccd1 vccd1 _03834_ sky130_fd_sc_hd__and2_1
XFILLER_0_29_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_8_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06423_ _01366_ vssd1 vssd1 vccd1 vccd1 _01367_ sky130_fd_sc_hd__clkbuf_4
X_09142_ _03750_ _03788_ _03789_ vssd1 vssd1 vccd1 vccd1 _03790_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_44_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__08435__A1 net33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06354_ net1196 _01296_ _01299_ vssd1 vssd1 vccd1 vccd1 genblk1\[0\].osc.clkdiv_C.next_cnt\[16\]
+ sky130_fd_sc_hd__o21a_1
XANTENNA__07238__A2 _02011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_44_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_72_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06254__A1_N genblk1\[0\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08406__A net25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10703__B_N _04856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_127_682 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09073_ _03729_ vssd1 vssd1 vccd1 vccd1 _00088_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06285_ _01173_ _01191_ vssd1 vssd1 vccd1 vccd1 _01247_ sky130_fd_sc_hd__and2_1
XANTENNA_fanout214_A net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11990__A1 _04230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08024_ _02711_ _02724_ _02727_ _02730_ vssd1 vssd1 vccd1 vccd1 _02731_ sky130_fd_sc_hd__a31o_1
Xhold710 genblk2\[4\].wave_shpr.div.acc\[9\] vssd1 vssd1 vccd1 vccd1 net928 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_31_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold721 sig_norm.i\[0\] vssd1 vssd1 vccd1 vccd1 net939 sky130_fd_sc_hd__dlygate4sd3_1
Xhold732 genblk2\[8\].wave_shpr.div.acc\[7\] vssd1 vssd1 vccd1 vccd1 net950 sky130_fd_sc_hd__dlygate4sd3_1
Xhold743 genblk2\[5\].wave_shpr.div.acc\[3\] vssd1 vssd1 vccd1 vccd1 net961 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_97_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_13_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold754 _00492_ vssd1 vssd1 vccd1 vccd1 net972 sky130_fd_sc_hd__dlygate4sd3_1
Xhold765 genblk2\[1\].wave_shpr.div.acc\[19\] vssd1 vssd1 vccd1 vccd1 net983 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold776 _01073_ vssd1 vssd1 vccd1 vccd1 net994 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11742__A1 _02248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold787 genblk2\[8\].wave_shpr.div.b1\[13\] vssd1 vssd1 vccd1 vccd1 net1005 sky130_fd_sc_hd__dlygate4sd3_1
X_09975_ genblk2\[3\].wave_shpr.div.acc\[7\] genblk2\[3\].wave_shpr.div.b1\[7\] vssd1
+ vssd1 vccd1 vccd1 _04371_ sky130_fd_sc_hd__or2b_1
Xhold798 genblk2\[3\].wave_shpr.div.acc\[16\] vssd1 vssd1 vccd1 vccd1 net1016 sky130_fd_sc_hd__dlygate4sd3_1
X_08926_ sig_norm.acc\[9\] _03589_ _03622_ vssd1 vssd1 vccd1 vccd1 _03623_ sky130_fd_sc_hd__a21o_1
X_08857_ _03562_ _03557_ _03560_ _03561_ vssd1 vssd1 vccd1 vccd1 _03564_ sky130_fd_sc_hd__o211a_1
XFILLER_0_99_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07808_ genblk2\[0\].wave_shpr.div.fin_quo\[5\] _02510_ _02513_ _02224_ vssd1 vssd1
+ vccd1 vccd1 _02515_ sky130_fd_sc_hd__a31o_1
XANTENNA__10610__S _04637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08788_ _03114_ _03494_ _03122_ vssd1 vssd1 vccd1 vccd1 _03495_ sky130_fd_sc_hd__o21a_1
X_07739_ genblk1\[1\].osc.clkdiv_C.cnt\[9\] _01334_ _01312_ genblk1\[1\].osc.clkdiv_C.cnt\[10\]
+ vssd1 vssd1 vccd1 vccd1 _02446_ sky130_fd_sc_hd__a22o_1
XFILLER_0_79_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08123__B1 _01565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10750_ net1061 _04886_ _04890_ _04914_ vssd1 vssd1 vccd1 vccd1 _00580_ sky130_fd_sc_hd__a22o_1
XFILLER_0_94_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09409_ _03970_ _03971_ _03972_ vssd1 vssd1 vccd1 vccd1 _03973_ sky130_fd_sc_hd__a21o_1
X_10681_ genblk2\[5\].wave_shpr.div.quo\[15\] _04861_ _04862_ net249 _04867_ vssd1
+ vssd1 vccd1 vccd1 _00558_ sky130_fd_sc_hd__a221o_1
XFILLER_0_137_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12420_ net576 _06072_ _06073_ _06087_ vssd1 vssd1 vccd1 vccd1 _01077_ sky130_fd_sc_hd__a22o_1
XFILLER_0_118_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07220__A _01365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12351_ _05982_ _06034_ vssd1 vssd1 vccd1 vccd1 _06035_ sky130_fd_sc_hd__nand2_1
XFILLER_0_133_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_23_628 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10057__S _04238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_63_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08035__B _02733_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11302_ genblk2\[7\].wave_shpr.div.acc\[8\] _05299_ _05300_ vssd1 vssd1 vccd1 vccd1
+ _05301_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12282_ _06002_ vssd1 vssd1 vccd1 vccd1 _01024_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_105_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11233_ _05245_ vssd1 vssd1 vccd1 vccd1 _05255_ sky130_fd_sc_hd__buf_2
X_11164_ _05223_ vssd1 vssd1 vccd1 vccd1 _00685_ sky130_fd_sc_hd__clkbuf_1
X_10115_ net376 _04461_ _04462_ net514 _04468_ vssd1 vssd1 vccd1 vccd1 _00391_ sky130_fd_sc_hd__a221o_1
X_11095_ genblk2\[6\].wave_shpr.div.i\[1\] genblk2\[6\].wave_shpr.div.i\[0\] genblk2\[6\].wave_shpr.div.i\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05158_ sky130_fd_sc_hd__a21o_1
X_10046_ _01325_ _01996_ vssd1 vssd1 vccd1 vccd1 _04432_ sky130_fd_sc_hd__nor2_2
XFILLER_0_117_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold70 genblk2\[11\].wave_shpr.div.i\[4\] vssd1 vssd1 vccd1 vccd1 net288 sky130_fd_sc_hd__dlygate4sd3_1
Xhold81 _00143_ vssd1 vssd1 vccd1 vccd1 net299 sky130_fd_sc_hd__dlygate4sd3_1
Xhold92 genblk2\[5\].wave_shpr.div.quo\[9\] vssd1 vssd1 vccd1 vccd1 net310 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_58_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_85_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11997_ net1275 _01556_ _05802_ vssd1 vssd1 vccd1 vccd1 _05804_ sky130_fd_sc_hd__mux2_1
XFILLER_0_133_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10948_ _05051_ vssd1 vssd1 vccd1 vccd1 _05057_ sky130_fd_sc_hd__clkbuf_4
X_13736_ clknet_leaf_47_clk net343 net119 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.quo\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_85_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09610__A _04042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_912 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_42_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13667_ clknet_leaf_42_clk _00980_ net124 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.acc\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_10879_ _05022_ vssd1 vssd1 vccd1 vccd1 _05023_ sky130_fd_sc_hd__buf_4
XFILLER_0_85_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_144_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_26_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12618_ clknet_leaf_17_clk genblk1\[4\].osc.clkdiv_C.next_cnt\[3\] net80 vssd1 vssd1
+ vccd1 vccd1 genblk1\[4\].osc.clkdiv_C.cnt\[3\] sky130_fd_sc_hd__dfrtp_4
X_13598_ clknet_leaf_76_clk net647 net208 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.acc\[22\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_775 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_693 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12549_ clknet_leaf_60_clk genblk1\[0\].osc.clkdiv_C.next_cnt\[6\] net186 vssd1 vssd1
+ vccd1 vccd1 genblk1\[0\].osc.clkdiv_C.cnt\[6\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_13_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_108_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_1 _01487_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_111_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08196__A3 _02350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09760_ _01325_ _01423_ vssd1 vssd1 vccd1 vccd1 _04229_ sky130_fd_sc_hd__nor2_4
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06972_ genblk1\[7\].osc.clkdiv_C.cnt\[13\] _01214_ vssd1 vssd1 vccd1 vccd1 _01808_
+ sky130_fd_sc_hd__xnor2_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08711_ _03410_ _03417_ vssd1 vssd1 vccd1 vccd1 _03418_ sky130_fd_sc_hd__xor2_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11488__B1 _03736_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09691_ genblk2\[2\].wave_shpr.div.b1\[2\] vssd1 vssd1 vccd1 vccd1 _04171_ sky130_fd_sc_hd__inv_2
X_08642_ _02604_ _02648_ _03344_ _03348_ vssd1 vssd1 vccd1 vccd1 _03349_ sky130_fd_sc_hd__nand4_1
XFILLER_0_89_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08573_ _02310_ _03279_ _02314_ vssd1 vssd1 vccd1 vccd1 _03280_ sky130_fd_sc_hd__o21a_1
XFILLER_0_107_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_89_694 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_107_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07524_ _01152_ sig_norm.i\[0\] sig_norm.busy vssd1 vssd1 vccd1 vccd1 _02243_ sky130_fd_sc_hd__and3b_1
XFILLER_0_49_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_901 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09520__A _03855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_8_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07455_ _02188_ vssd1 vssd1 vccd1 vccd1 _00016_ sky130_fd_sc_hd__inv_2
XANTENNA__11660__B1 _03855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10666__A _04672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_147_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06406_ _01201_ genblk1\[1\].osc.clkdiv_C.cnt\[13\] genblk1\[1\].osc.clkdiv_C.cnt\[8\]
+ vssd1 vssd1 vccd1 vccd1 _01350_ sky130_fd_sc_hd__o21a_1
XFILLER_0_8_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_134_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07386_ _02091_ _02135_ _02136_ vssd1 vssd1 vccd1 vccd1 _02137_ sky130_fd_sc_hd__and3_1
XFILLER_0_146_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07040__A _01489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_60_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09125_ genblk2\[0\].wave_shpr.div.b1\[5\] genblk2\[0\].wave_shpr.div.acc\[5\] vssd1
+ vssd1 vccd1 vccd1 _03773_ sky130_fd_sc_hd__and2b_1
X_06337_ genblk1\[0\].osc.clkdiv_C.cnt\[10\] _01286_ _01288_ _01270_ vssd1 vssd1 vccd1
+ vccd1 genblk1\[0\].osc.clkdiv_C.next_cnt\[10\] sky130_fd_sc_hd__o211a_1
XFILLER_0_127_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__09081__A1 _03704_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_663 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09056_ net1289 _01201_ _03708_ vssd1 vssd1 vccd1 vccd1 _03718_ sky130_fd_sc_hd__mux2_1
X_06268_ _01220_ vssd1 vssd1 vccd1 vccd1 _01230_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_115_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__11497__A _05444_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08007_ _01729_ _01758_ _01735_ genblk1\[6\].osc.clkdiv_C.cnt\[1\] vssd1 vssd1 vccd1
+ vccd1 _02714_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_103_858 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_114_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold540 genblk2\[7\].wave_shpr.div.b1\[16\] vssd1 vssd1 vccd1 vccd1 net758 sky130_fd_sc_hd__dlygate4sd3_1
X_06199_ PWM.counter\[5\] PWM.counter\[4\] _01161_ vssd1 vssd1 vccd1 vccd1 _01164_
+ sky130_fd_sc_hd__and3_1
Xhold551 genblk2\[11\].wave_shpr.div.quo\[1\] vssd1 vssd1 vccd1 vccd1 net769 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10518__A2 _04657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07919__B1 _01858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_677 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold562 _00379_ vssd1 vssd1 vccd1 vccd1 net780 sky130_fd_sc_hd__dlygate4sd3_1
Xhold573 genblk2\[3\].wave_shpr.div.acc\[11\] vssd1 vssd1 vccd1 vccd1 net791 sky130_fd_sc_hd__dlygate4sd3_1
Xhold584 genblk2\[8\].wave_shpr.div.acc\[16\] vssd1 vssd1 vccd1 vccd1 net802 sky130_fd_sc_hd__dlygate4sd3_1
Xhold595 genblk2\[1\].wave_shpr.div.acc\[10\] vssd1 vssd1 vccd1 vccd1 net813 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08592__B1 _02521_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09958_ _04356_ vssd1 vssd1 vccd1 vccd1 _04357_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout77_A net84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08909_ _03587_ net26 vssd1 vssd1 vccd1 vccd1 _03611_ sky130_fd_sc_hd__or2_1
X_09889_ _04190_ _04306_ vssd1 vssd1 vccd1 vccd1 _04307_ sky130_fd_sc_hd__xnor2_1
X_11920_ genblk2\[10\].wave_shpr.div.acc\[5\] genblk2\[10\].wave_shpr.div.b1\[5\]
+ vssd1 vssd1 vccd1 vccd1 _05742_ sky130_fd_sc_hd__and2b_1
XFILLER_0_99_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__07860__D _02459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11851_ genblk2\[9\].wave_shpr.div.acc\[13\] _05690_ _05673_ vssd1 vssd1 vccd1 vccd1
+ _05691_ sky130_fd_sc_hd__mux2_1
XTAP_2734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10802_ genblk2\[5\].wave_shpr.div.acc\[24\] _04880_ _04949_ vssd1 vssd1 vccd1 vccd1
+ _04953_ sky130_fd_sc_hd__or3b_1
XTAP_2778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11782_ net416 _05628_ _05629_ net533 _05640_ vssd1 vssd1 vccd1 vccd1 _00886_ sky130_fd_sc_hd__a221o_1
XTAP_2789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09844__B1 _04250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_137_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10733_ net1037 _04886_ _04890_ _04901_ vssd1 vssd1 vccd1 vccd1 _00576_ sky130_fd_sc_hd__a22o_1
X_13521_ clknet_leaf_79_clk _00838_ net206 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.acc\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_755 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_83_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_48_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_12_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13452_ clknet_leaf_99_clk _00769_ net166 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.fin_quo\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_10664_ genblk2\[5\].wave_shpr.div.quo\[8\] _04853_ _04857_ net308 vssd1 vssd1 vccd1
+ vccd1 _00551_ sky130_fd_sc_hd__a22o_1
XFILLER_0_82_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_4_14_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12403_ _05966_ _06074_ vssd1 vssd1 vccd1 vccd1 _06075_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_915 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_141_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_51_712 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09072__A1 _01340_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_809 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13383_ clknet_leaf_83_clk _00702_ net200 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.b1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10595_ _04822_ vssd1 vssd1 vccd1 vccd1 _00517_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__07885__A _02526_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07083__B1 genblk1\[8\].osc.clkdiv_C.cnt\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12334_ _03689_ genblk1\[11\].osc.clkdiv_C.cnt\[12\] vssd1 vssd1 vccd1 vccd1 _06025_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_50_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_121_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12265_ net1295 _01240_ _05802_ vssd1 vssd1 vccd1 vccd1 _05993_ sky130_fd_sc_hd__mux2_1
XANTENNA__10509__A2 _04657_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11216_ _05247_ vssd1 vssd1 vccd1 vccd1 _05249_ sky130_fd_sc_hd__clkbuf_4
X_12196_ genblk2\[11\].wave_shpr.div.acc\[8\] genblk2\[11\].wave_shpr.div.b1\[8\]
+ vssd1 vssd1 vccd1 vccd1 _05934_ sky130_fd_sc_hd__or2b_1
X_11147_ genblk2\[7\].wave_shpr.div.b1\[13\] genblk2\[7\].wave_shpr.div.acc\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05207_ sky130_fd_sc_hd__and2b_1
XFILLER_0_37_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11078_ net1031 _05119_ _05126_ _05147_ vssd1 vssd1 vccd1 vccd1 _00675_ sky130_fd_sc_hd__a22o_1
XANTENNA__07138__A1 genblk1\[9\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10029_ genblk2\[3\].wave_shpr.div.fin_quo\[1\] genblk2\[3\].wave_shpr.div.quo\[0\]
+ _04422_ vssd1 vssd1 vccd1 vccd1 _04424_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_801 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_53_23 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_845 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_86_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13719_ clknet_leaf_36_clk _01030_ net105 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.b1\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11185__A1_N _03727_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_128_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07240_ genblk1\[10\].osc.clkdiv_C.cnt\[3\] _02013_ _02021_ vssd1 vssd1 vccd1 vccd1
+ _02022_ sky130_fd_sc_hd__a21oi_1
XANTENNA__07861__A2 _02458_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_6_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_27_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_113 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_143_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_6_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07171_ genblk1\[9\].osc.clkdiv_C.cnt\[4\] _01960_ genblk1\[9\].osc.clkdiv_C.cnt\[5\]
+ vssd1 vssd1 vccd1 vccd1 _01966_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_27_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_54_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07304__A2_N _02064_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_143_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06122_ genblk2\[9\].wave_shpr.div.done genblk2\[8\].wave_shpr.div.done genblk2\[11\].wave_shpr.div.done
+ genblk2\[10\].wave_shpr.div.done vssd1 vssd1 vccd1 vccd1 _01094_ sky130_fd_sc_hd__or4_2
XFILLER_0_14_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09366__A2 _03841_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09812_ net441 _04253_ _04251_ net574 _04255_ vssd1 vssd1 vccd1 vccd1 _00301_ sky130_fd_sc_hd__a221o_1
X_09743_ genblk2\[2\].wave_shpr.div.fin_quo\[4\] net1327 _00009_ vssd1 vssd1 vccd1
+ vccd1 _04219_ sky130_fd_sc_hd__mux2_1
X_06955_ net1063 _01790_ vssd1 vssd1 vccd1 vccd1 genblk1\[6\].osc.clkdiv_C.next_cnt\[17\]
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_94_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__10160__S _04420_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09674_ net285 _04154_ _03819_ vssd1 vssd1 vccd1 vccd1 _04155_ sky130_fd_sc_hd__o21ai_1
X_06886_ genblk1\[6\].osc.clkdiv_C.cnt\[1\] _01738_ _01739_ genblk1\[6\].osc.clkdiv_C.cnt\[8\]
+ vssd1 vssd1 vccd1 vccd1 _01740_ sky130_fd_sc_hd__o22a_1
XTAP_2008 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08625_ _03296_ _03297_ _03246_ _03258_ vssd1 vssd1 vccd1 vccd1 _03332_ sky130_fd_sc_hd__o211ai_2
XTAP_2019 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08556_ _02742_ _03261_ _03262_ _02745_ vssd1 vssd1 vccd1 vccd1 _03263_ sky130_fd_sc_hd__o31a_1
XTAP_1329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_76_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07507_ PWM.counter\[7\] vssd1 vssd1 vccd1 vccd1 _02227_ sky130_fd_sc_hd__inv_2
XANTENNA__09250__A _03853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_92_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12087__S _05787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08487_ _02939_ _03193_ _02943_ vssd1 vssd1 vccd1 vccd1 _03194_ sky130_fd_sc_hd__o21a_1
XFILLER_0_65_837 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07438_ genblk2\[4\].wave_shpr.div.busy _02175_ vssd1 vssd1 vccd1 vccd1 _02176_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_753 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_119_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_134_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07852__A2 _02309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_9_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_17_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_123_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07369_ _02123_ vssd1 vssd1 vccd1 vccd1 _02124_ sky130_fd_sc_hd__inv_2
XANTENNA__09054__A1 _03714_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_32_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_122_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09108_ genblk2\[0\].wave_shpr.div.acc\[7\] genblk2\[0\].wave_shpr.div.b1\[7\] vssd1
+ vssd1 vccd1 vccd1 _03756_ sky130_fd_sc_hd__or2b_1
XANTENNA__07604__A2 _02309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10380_ _04651_ vssd1 vssd1 vccd1 vccd1 _04657_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__12625__RESET_B net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_103_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09039_ _02147_ vssd1 vssd1 vccd1 vccd1 _03707_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_32_288 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12050_ net353 _05823_ _05825_ net357 _05829_ vssd1 vssd1 vccd1 vccd1 _00965_ sky130_fd_sc_hd__a221o_1
Xhold370 genblk2\[1\].wave_shpr.div.acc_next\[0\] vssd1 vssd1 vccd1 vccd1 net588 sky130_fd_sc_hd__dlygate4sd3_1
Xhold381 genblk2\[0\].wave_shpr.div.quo\[11\] vssd1 vssd1 vccd1 vccd1 net599 sky130_fd_sc_hd__dlygate4sd3_1
X_11001_ net1015 _05086_ _05056_ _05089_ vssd1 vssd1 vccd1 vccd1 _00656_ sky130_fd_sc_hd__a22o_1
Xhold392 genblk2\[1\].wave_shpr.div.quo\[10\] vssd1 vssd1 vccd1 vccd1 net610 sky130_fd_sc_hd__dlygate4sd3_1
X_12952_ clknet_leaf_125_clk _00281_ net61 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.b1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1070 genblk2\[7\].wave_shpr.div.b1\[2\] vssd1 vssd1 vccd1 vccd1 net1288 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1081 genblk2\[1\].wave_shpr.div.b1\[13\] vssd1 vssd1 vccd1 vccd1 net1299 sky130_fd_sc_hd__dlygate4sd3_1
Xhold1092 genblk2\[11\].wave_shpr.div.quo\[0\] vssd1 vssd1 vccd1 vccd1 net1310 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_87_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06879__B1 _01732_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11903_ _03839_ _05725_ _05727_ _03841_ net775 vssd1 vssd1 vccd1 vccd1 _00920_ sky130_fd_sc_hd__a32o_1
XTAP_2520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12883_ clknet_leaf_55_clk net293 net176 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.quo\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_2542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11834_ net884 _05652_ _05653_ _05677_ vssd1 vssd1 vccd1 vccd1 _00901_ sky130_fd_sc_hd__a22o_1
XTAP_2575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09817__B1 _04251_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11765_ _05631_ genblk1\[9\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 _05632_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_95_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1874 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1885 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1896 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10716_ genblk2\[5\].wave_shpr.div.acc\[2\] _04888_ _04821_ vssd1 vssd1 vccd1 vccd1
+ _04889_ sky130_fd_sc_hd__mux2_1
X_13504_ clknet_leaf_81_clk _00821_ net199 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.acc\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_138_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_138_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11696_ genblk2\[9\].wave_shpr.div.b1\[8\] genblk2\[9\].wave_shpr.div.acc\[8\] vssd1
+ vssd1 vccd1 vccd1 _05588_ sky130_fd_sc_hd__and2b_1
XFILLER_0_24_701 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_689 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10647_ net1096 vssd1 vssd1 vccd1 vccd1 _04851_ sky130_fd_sc_hd__inv_2
X_13435_ clknet_leaf_95_clk _00754_ net161 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.acc\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_130_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09045__A1 _01991_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13366_ clknet_leaf_91_clk _00685_ net143 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.fin_quo\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_10578_ genblk2\[5\].wave_shpr.div.b1\[13\] genblk2\[5\].wave_shpr.div.acc\[13\]
+ vssd1 vssd1 vccd1 vccd1 _04806_ sky130_fd_sc_hd__and2b_1
XFILLER_0_106_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12317_ net443 _06014_ _06015_ genblk2\[11\].wave_shpr.div.quo\[11\] _06016_ vssd1
+ vssd1 vccd1 vccd1 _01045_ sky130_fd_sc_hd__a221o_1
XFILLER_0_133_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13297_ clknet_leaf_86_clk _00618_ net179 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.b1\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_12248_ _05984_ vssd1 vssd1 vccd1 vccd1 _01008_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__12352__A1 _03944_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12179_ genblk2\[10\].wave_shpr.div.i\[1\] genblk2\[10\].wave_shpr.div.i\[0\] genblk2\[10\].wave_shpr.div.i\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05920_ sky130_fd_sc_hd__and3_1
XFILLER_0_48_89 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08308__B1 _02222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06740_ _01623_ vssd1 vssd1 vccd1 vccd1 genblk1\[4\].osc.clkdiv_C.next_cnt\[6\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_155_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06671_ genblk1\[4\].osc.clkdiv_C.cnt\[2\] _01559_ vssd1 vssd1 vccd1 vccd1 _01561_
+ sky130_fd_sc_hd__nor2_1
X_08410_ genblk2\[2\].wave_shpr.div.fin_quo\[3\] _03116_ vssd1 vssd1 vccd1 vccd1 _03117_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_149_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09390_ genblk2\[1\].wave_shpr.div.acc\[17\] genblk2\[1\].wave_shpr.div.b1\[17\]
+ vssd1 vssd1 vccd1 vccd1 _03954_ sky130_fd_sc_hd__or2b_1
XFILLER_0_58_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_47_815 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09070__A _03702_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08341_ _03041_ _03042_ _03047_ vssd1 vssd1 vccd1 vccd1 _03048_ sky130_fd_sc_hd__nand3_1
XFILLER_0_86_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_73_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08272_ genblk2\[10\].wave_shpr.div.fin_quo\[4\] vssd1 vssd1 vccd1 vccd1 _02979_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_80_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_104_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_129_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_144_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07223_ _01174_ _01230_ _01196_ vssd1 vssd1 vccd1 vccd1 _02005_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_105_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_14_211 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_144_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_fanout127_A net16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07154_ net1136 _01953_ vssd1 vssd1 vccd1 vccd1 genblk1\[9\].osc.clkdiv_C.next_cnt\[0\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_131_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_70_884 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_73_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_06105_ smpl_rt_clkdiv.clkDiv_inst.cnt\[1\] smpl_rt_clkdiv.clkDiv_inst.cnt\[0\] smpl_rt_clkdiv.clkDiv_inst.cnt\[2\]
+ vssd1 vssd1 vccd1 vccd1 _01086_ sky130_fd_sc_hd__and3_1
XFILLER_0_30_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07085_ genblk1\[8\].osc.clkdiv_C.cnt\[6\] _01895_ vssd1 vssd1 vccd1 vccd1 _01897_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_120_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12343__A1 genblk2\[11\].wave_shpr.div.acc_next\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout102 net104 vssd1 vssd1 vccd1 vccd1 net102 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_193 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08547__B1 _02309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout113 net114 vssd1 vssd1 vccd1 vccd1 net113 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_100_669 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11775__A _04676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout124 net125 vssd1 vssd1 vccd1 vccd1 net124 sky130_fd_sc_hd__clkbuf_4
XANTENNA__08011__A2 _01367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout135 net136 vssd1 vssd1 vccd1 vccd1 net135 sky130_fd_sc_hd__buf_2
Xfanout146 net150 vssd1 vssd1 vccd1 vccd1 net146 sky130_fd_sc_hd__clkbuf_4
Xfanout157 net158 vssd1 vssd1 vccd1 vccd1 net157 sky130_fd_sc_hd__clkbuf_2
Xfanout168 net170 vssd1 vssd1 vccd1 vccd1 net168 sky130_fd_sc_hd__clkbuf_4
X_07987_ _02225_ _02681_ vssd1 vssd1 vccd1 vccd1 _02694_ sky130_fd_sc_hd__and2_1
Xfanout179 net180 vssd1 vssd1 vccd1 vccd1 net179 sky130_fd_sc_hd__clkbuf_4
X_09726_ _04157_ _04204_ _04205_ vssd1 vssd1 vccd1 vccd1 _04206_ sky130_fd_sc_hd__a21o_1
X_06938_ genblk1\[6\].osc.clkdiv_C.cnt\[11\] _01777_ _01780_ vssd1 vssd1 vccd1 vccd1
+ genblk1\[6\].osc.clkdiv_C.next_cnt\[11\] sky130_fd_sc_hd__o21a_1
XANTENNA__09511__A2 _04043_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09657_ _04009_ _04129_ _04143_ vssd1 vssd1 vccd1 vccd1 _04144_ sky130_fd_sc_hd__o21ai_1
X_06869_ _01694_ _01723_ _01724_ vssd1 vssd1 vccd1 vccd1 _01725_ sky130_fd_sc_hd__and3_1
XFILLER_0_96_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1104 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08608_ genblk2\[5\].wave_shpr.div.fin_quo\[1\] vssd1 vssd1 vccd1 vccd1 _03315_ sky130_fd_sc_hd__inv_2
XTAP_1115 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1126 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09588_ net995 _04076_ _04080_ _04092_ vssd1 vssd1 vccd1 vccd1 _00240_ sky130_fd_sc_hd__a22o_1
XTAP_1137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_155_809 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08539_ _03235_ _03245_ vssd1 vssd1 vccd1 vccd1 _03246_ sky130_fd_sc_hd__or2b_1
XFILLER_0_49_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_100 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_148_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11550_ genblk2\[8\].wave_shpr.div.b1\[0\] _05417_ genblk2\[8\].wave_shpr.div.acc\[0\]
+ vssd1 vssd1 vccd1 vccd1 _05473_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_147_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10501_ genblk2\[4\].wave_shpr.div.acc\[18\] _04738_ net591 vssd1 vssd1 vccd1 vccd1
+ _04741_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_52_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_626 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_108_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11481_ _05437_ vssd1 vssd1 vccd1 vccd1 _00788_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_80_648 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13220_ clknet_leaf_136_clk _00543_ net62 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.quo\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_107_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10432_ genblk2\[4\].wave_shpr.div.acc\[2\] _04688_ _04623_ vssd1 vssd1 vccd1 vccd1
+ _04689_ sky130_fd_sc_hd__mux2_1
XFILLER_0_104_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08786__B1 _02224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13151_ clknet_leaf_17_clk net532 net80 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.quo\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10363_ _03833_ net1223 vssd1 vssd1 vccd1 vccd1 _04650_ sky130_fd_sc_hd__and2_1
XANTENNA__08043__B _01360_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12102_ _05759_ _05863_ vssd1 vssd1 vccd1 vccd1 _05864_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_130_260 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13082_ clknet_leaf_126_clk _00409_ net61 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.acc\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_10294_ genblk2\[4\].wave_shpr.div.b1\[12\] genblk2\[4\].wave_shpr.div.acc\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04606_ sky130_fd_sc_hd__and2b_1
X_12033_ _05819_ genblk1\[10\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 _05820_
+ sky130_fd_sc_hd__and2_1
XANTENNA__08002__A2 _01675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_18_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_109_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10896__A1 _01514_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07210__B1 _01241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_8_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06498__B net36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10648__A1 _03726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12935_ clknet_leaf_30_clk _00264_ net102 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.i\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_125_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_87_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12866_ clknet_leaf_135_clk _00197_ net61 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.b1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08069__A2 _01592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11817_ net938 _05652_ _05653_ _05664_ vssd1 vssd1 vccd1 vccd1 _00897_ sky130_fd_sc_hd__a22o_1
XTAP_2394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12797_ clknet_leaf_57_clk net270 net183 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_141_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_28_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_56_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11748_ genblk2\[9\].wave_shpr.div.quo\[3\] _05623_ _05624_ net686 vssd1 vssd1 vccd1
+ vccd1 _00868_ sky130_fd_sc_hd__a22o_1
XFILLER_0_138_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_55_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_71_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06961__B _01221_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11679_ genblk2\[9\].wave_shpr.div.acc\[2\] genblk2\[9\].wave_shpr.div.b1\[2\] vssd1
+ vssd1 vccd1 vccd1 _05571_ sky130_fd_sc_hd__or2b_1
XFILLER_0_114_717 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_52_840 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13418_ clknet_leaf_119_clk _00737_ net141 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.acc\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_3_425 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_469 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13349_ clknet_leaf_4_clk _00670_ net45 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.acc\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__09764__S _04039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_770 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11595__A _05441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07910_ _01230_ _01564_ _01889_ _01238_ vssd1 vssd1 vccd1 vccd1 _02617_ sky130_fd_sc_hd__a211oi_1
X_08890_ _03595_ vssd1 vssd1 vccd1 vccd1 _03596_ sky130_fd_sc_hd__buf_2
XFILLER_0_75_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07841_ _02530_ _02535_ vssd1 vssd1 vccd1 vccd1 _02548_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_75_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07772_ genblk1\[0\].osc.clkdiv_C.cnt\[1\] _01190_ net34 genblk1\[0\].osc.clkdiv_C.cnt\[0\]
+ _02336_ vssd1 vssd1 vccd1 vccd1 _02479_ sky130_fd_sc_hd__o2111a_1
X_09511_ net684 _04043_ _04047_ net764 vssd1 vssd1 vccd1 vccd1 _00208_ sky130_fd_sc_hd__a22o_1
XANTENNA__10639__A1 _04225_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06723_ _01609_ vssd1 vssd1 vccd1 vccd1 _01610_ sky130_fd_sc_hd__inv_2
XFILLER_0_78_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10939__A _05054_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09442_ genblk2\[1\].wave_shpr.div.acc\[18\] _04005_ vssd1 vssd1 vccd1 vccd1 _04006_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_78_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_4_2_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06654_ genblk1\[3\].osc.clkdiv_C.cnt\[13\] _01545_ _01548_ vssd1 vssd1 vccd1 vccd1
+ genblk1\[3\].osc.clkdiv_C.next_cnt\[13\] sky130_fd_sc_hd__o21a_1
XFILLER_0_66_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_47_601 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_75_910 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_93_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07313__A _01308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09373_ _02213_ vssd1 vssd1 vccd1 vccd1 _03942_ sky130_fd_sc_hd__buf_4
X_06585_ _01490_ genblk1\[3\].osc.clkdiv_C.cnt\[13\] _01363_ genblk1\[3\].osc.clkdiv_C.cnt\[15\]
+ vssd1 vssd1 vccd1 vccd1 _01493_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_47_645 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_86_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08324_ _02638_ _02640_ genblk2\[8\].wave_shpr.div.fin_quo\[4\] vssd1 vssd1 vccd1
+ vccd1 _03031_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_129_393 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_853 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08255_ _02960_ _02961_ genblk2\[6\].wave_shpr.div.fin_quo\[6\] _02539_ vssd1 vssd1
+ vccd1 vccd1 _02962_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_46_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10811__A1 _04855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_74_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12365__S _05982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10674__A _04672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07206_ _01989_ vssd1 vssd1 vccd1 vccd1 genblk1\[9\].osc.clkdiv_C.next_cnt\[16\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_104_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12013__B1 _03735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08186_ net9 _02744_ _02365_ vssd1 vssd1 vccd1 vccd1 _02893_ sky130_fd_sc_hd__nand3_1
XFILLER_0_6_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_873 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_70_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07137_ genblk1\[9\].osc.clkdiv_C.cnt\[16\] _01936_ vssd1 vssd1 vccd1 vccd1 _01937_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_113_772 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06243__A1 genblk1\[0\].osc.clkdiv_C.cnt\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07068_ _01862_ _01885_ vssd1 vssd1 vccd1 vccd1 _01886_ sky130_fd_sc_hd__nor2_2
XFILLER_0_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10613__S _04637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06599__A _01441_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09709_ genblk2\[2\].wave_shpr.div.b1\[8\] genblk2\[2\].wave_shpr.div.acc\[8\] vssd1
+ vssd1 vccd1 vccd1 _04189_ sky130_fd_sc_hd__and2b_1
XFILLER_0_97_512 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10981_ _05074_ genblk1\[6\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 _05076_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_69_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_12720_ clknet_leaf_86_clk genblk1\[9\].osc.clkdiv_C.next_cnt\[15\] net183 vssd1
+ vssd1 vccd1 vccd1 genblk1\[9\].osc.clkdiv_C.cnt\[15\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_139_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12651_ clknet_leaf_28_clk genblk1\[6\].osc.clkdiv_C.next_cnt\[0\] net89 vssd1 vssd1
+ vccd1 vccd1 genblk1\[6\].osc.clkdiv_C.cnt\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_155_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_740 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_65_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11602_ genblk2\[8\].wave_shpr.div.acc\[12\] _05512_ _05493_ vssd1 vssd1 vccd1 vccd1
+ _05513_ sky130_fd_sc_hd__mux2_1
XFILLER_0_108_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12582_ clknet_leaf_14_clk genblk1\[2\].osc.clkdiv_C.next_cnt\[3\] net74 vssd1 vssd1
+ vccd1 vccd1 genblk1\[2\].osc.clkdiv_C.cnt\[3\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_93_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_108_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_37_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11533_ genblk2\[8\].wave_shpr.div.quo\[19\] _05454_ _05458_ net617 _05463_ vssd1
+ vssd1 vccd1 vccd1 _00814_ sky130_fd_sc_hd__a221o_1
XFILLER_0_135_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_37_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_123_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12004__A0 genblk2\[11\].wave_shpr.div.b1\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11464_ net1230 net34 _05237_ vssd1 vssd1 vccd1 vccd1 _05429_ sky130_fd_sc_hd__mux2_1
XFILLER_0_150_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13203_ clknet_leaf_8_clk _00526_ net48 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.b1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_10415_ _04676_ _01650_ vssd1 vssd1 vccd1 vccd1 _04677_ sky130_fd_sc_hd__nor2_1
XFILLER_0_151_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_33_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08223__A2 _02308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11395_ genblk2\[8\].wave_shpr.div.acc\[4\] genblk2\[8\].wave_shpr.div.b1\[4\] vssd1
+ vssd1 vccd1 vccd1 _05371_ sky130_fd_sc_hd__or2b_1
XFILLER_0_110_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13134_ clknet_leaf_115_clk _00459_ net133 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.quo\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10346_ _04640_ vssd1 vssd1 vccd1 vccd1 _00450_ sky130_fd_sc_hd__clkbuf_1
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12307__A1 net355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13065_ clknet_leaf_22_clk net377 net95 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.quo\[17\]
+ sky130_fd_sc_hd__dfrtp_1
X_10277_ genblk2\[4\].wave_shpr.div.b1\[3\] genblk2\[4\].wave_shpr.div.acc\[3\] vssd1
+ vssd1 vccd1 vccd1 _04589_ sky130_fd_sc_hd__and2b_1
XFILLER_0_29_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12016_ _02208_ vssd1 vssd1 vccd1 vccd1 _05812_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_136_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_45_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap2 _04335_ vssd1 vssd1 vccd1 vccd1 net1351 sky130_fd_sc_hd__buf_1
XANTENNA__09487__A1 _04032_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_88_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12918_ clknet_leaf_39_clk _00249_ net115 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.acc\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_88_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_29_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_2180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12849_ clknet_leaf_58_clk _00180_ net194 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.i\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_131_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_145_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_61_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06370_ genblk1\[1\].osc.clkdiv_C.cnt\[4\] _01313_ vssd1 vssd1 vccd1 vccd1 _01314_
+ sky130_fd_sc_hd__xnor2_1
XTAP_1490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_44_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_71_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_28_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_126_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_127_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_126_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08040_ _02697_ _02698_ _02746_ vssd1 vssd1 vccd1 vccd1 _02747_ sky130_fd_sc_hd__nand3_1
XFILLER_0_127_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_24_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_40_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold903 genblk2\[1\].wave_shpr.div.b1\[11\] vssd1 vssd1 vccd1 vccd1 net1121 sky130_fd_sc_hd__dlygate4sd3_1
Xhold914 PWM.final_in\[6\] vssd1 vssd1 vccd1 vccd1 net1132 sky130_fd_sc_hd__dlygate4sd3_1
Xhold925 genblk1\[10\].osc.clkdiv_C.cnt\[15\] vssd1 vssd1 vccd1 vccd1 net1143 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold936 genblk2\[5\].wave_shpr.div.i\[2\] vssd1 vssd1 vccd1 vccd1 net1154 sky130_fd_sc_hd__dlygate4sd3_1
Xhold947 genblk2\[6\].wave_shpr.div.acc\[2\] vssd1 vssd1 vccd1 vccd1 net1165 sky130_fd_sc_hd__dlygate4sd3_1
Xhold958 sig_norm.quo\[2\] vssd1 vssd1 vccd1 vccd1 net1176 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__13516__RESET_B net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09991_ _04377_ _04385_ _04386_ vssd1 vssd1 vccd1 vccd1 _04387_ sky130_fd_sc_hd__a21oi_1
Xhold969 genblk2\[9\].wave_shpr.div.b1\[6\] vssd1 vssd1 vccd1 vccd1 net1187 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_110_731 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08942_ _03551_ _03633_ vssd1 vssd1 vccd1 vccd1 _03634_ sky130_fd_sc_hd__and2_1
X_08873_ sig_norm.acc\[1\] sig_norm.b1\[1\] vssd1 vssd1 vccd1 vccd1 _03579_ sky130_fd_sc_hd__or2b_1
XFILLER_0_36_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07824_ _02510_ _02511_ genblk2\[0\].wave_shpr.div.fin_quo\[3\] vssd1 vssd1 vccd1
+ vccd1 _02531_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_79_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07755_ genblk2\[1\].wave_shpr.div.fin_quo\[0\] genblk2\[1\].wave_shpr.div.fin_quo\[1\]
+ vssd1 vssd1 vccd1 vccd1 _02462_ sky130_fd_sc_hd__or2_1
XANTENNA__10088__A2 _04452_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06706_ genblk1\[4\].osc.clkdiv_C.cnt\[13\] _01595_ vssd1 vssd1 vccd1 vccd1 _01596_
+ sky130_fd_sc_hd__xnor2_1
X_07686_ _02023_ _02386_ _02388_ _02389_ _02392_ vssd1 vssd1 vccd1 vccd1 _02393_ sky130_fd_sc_hd__o221a_1
XANTENNA__08139__A net10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_67_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09425_ _03962_ _03987_ _03988_ vssd1 vssd1 vccd1 vccd1 _03989_ sky130_fd_sc_hd__a21o_1
X_06637_ net1095 _01535_ _01537_ vssd1 vssd1 vccd1 vccd1 genblk1\[3\].osc.clkdiv_C.next_cnt\[7\]
+ sky130_fd_sc_hd__a21oi_1
XFILLER_0_19_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_109_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_820 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09356_ genblk2\[0\].wave_shpr.div.acc\[20\] _03800_ net1352 vssd1 vssd1 vccd1 vccd1
+ _03930_ sky130_fd_sc_hd__or3_1
X_06568_ _01451_ _01478_ vssd1 vssd1 vccd1 vccd1 _01479_ sky130_fd_sc_hd__nor2_1
XFILLER_0_75_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_81_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08307_ _02349_ _02351_ _02353_ genblk2\[11\].wave_shpr.div.fin_quo\[3\] vssd1 vssd1
+ vccd1 vccd1 _03014_ sky130_fd_sc_hd__a31oi_1
XANTENNA__12095__S _05787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09287_ _03771_ _03759_ vssd1 vssd1 vccd1 vccd1 _03878_ sky130_fd_sc_hd__or2b_1
XANTENNA__10608__S _00015_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06499_ genblk1\[2\].osc.clkdiv_C.cnt\[13\] genblk1\[2\].osc.clkdiv_C.cnt\[0\] net35
+ vssd1 vssd1 vccd1 vccd1 _01425_ sky130_fd_sc_hd__nor3_1
XFILLER_0_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_823 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08238_ _02798_ _02931_ _02936_ _02938_ _02944_ vssd1 vssd1 vccd1 vccd1 _02945_ sky130_fd_sc_hd__a32o_1
XFILLER_0_62_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06464__A1 genblk1\[1\].osc.clkdiv_C.cnt\[10\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07661__B1 _01235_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_34_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_105_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08169_ genblk1\[3\].osc.clkdiv_C.cnt\[8\] _01423_ _02870_ _02871_ _02875_ vssd1
+ vssd1 vccd1 vccd1 _02876_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_133_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10200_ net930 _04518_ _04522_ _04528_ vssd1 vssd1 vccd1 vccd1 _00416_ sky130_fd_sc_hd__a22o_1
X_11180_ _03708_ genblk2\[8\].wave_shpr.div.b1\[1\] vssd1 vssd1 vccd1 vccd1 _05231_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_30_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10131_ genblk2\[3\].wave_shpr.div.quo\[24\] _04451_ _04455_ net490 _04476_ vssd1
+ vssd1 vccd1 vccd1 _00399_ sky130_fd_sc_hd__a221o_1
X_10062_ net1186 _01240_ _04440_ vssd1 vssd1 vccd1 vccd1 _04441_ sky130_fd_sc_hd__mux2_1
XANTENNA_hold838_A genblk2\[5\].wave_shpr.div.quo\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09469__A1 _01231_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_106_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12892__RESET_B net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_98_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_15_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13752_ clknet_leaf_68_clk _01063_ net211 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.acc\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10964_ _05059_ genblk1\[6\].osc.clkdiv_C.cnt\[6\] vssd1 vssd1 vccd1 vccd1 _05067_
+ sky130_fd_sc_hd__and2_1
XANTENNA__06495__C _01327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12703_ clknet_leaf_89_clk genblk1\[8\].osc.clkdiv_C.next_cnt\[16\] net173 vssd1
+ vssd1 vccd1 vccd1 genblk1\[8\].osc.clkdiv_C.cnt\[16\] sky130_fd_sc_hd__dfrtp_4
X_13683_ clknet_leaf_63_clk _00996_ net190 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.acc\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_10895_ _05031_ vssd1 vssd1 vccd1 vccd1 _00608_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_38_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_127_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09579__S _04011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12634_ clknet_leaf_16_clk genblk1\[5\].osc.clkdiv_C.next_cnt\[1\] net74 vssd1 vssd1
+ vccd1 vccd1 genblk1\[5\].osc.clkdiv_C.cnt\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_31_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_38_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12565_ clknet_leaf_28_clk genblk1\[1\].osc.clkdiv_C.next_cnt\[4\] net89 vssd1 vssd1
+ vccd1 vccd1 genblk1\[1\].osc.clkdiv_C.cnt\[4\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_109_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_81_765 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11516_ _05441_ vssd1 vssd1 vccd1 vccd1 _05454_ sky130_fd_sc_hd__buf_2
XFILLER_0_13_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_53_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12496_ clknet_leaf_102_clk _00058_ net158 vssd1 vssd1 vccd1 vccd1 sig_norm.quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_80_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_150_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_80_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_34_692 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11447_ _05420_ vssd1 vssd1 vccd1 vccd1 _00771_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_151_697 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11200__A1 _01565_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_0_225 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09944__A2 _04253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11378_ genblk2\[7\].wave_shpr.div.i\[3\] _02192_ _05353_ vssd1 vssd1 vccd1 vccd1
+ _05356_ sky130_fd_sc_hd__and3_1
XFILLER_0_21_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11751__A2 _05623_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10329_ _04632_ vssd1 vssd1 vccd1 vccd1 _00441_ sky130_fd_sc_hd__clkbuf_1
X_13117_ clknet_leaf_13_clk _00442_ net52 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.b1\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13048_ clknet_leaf_135_clk _00375_ net62 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.quo\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_832 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_88_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07540_ _02253_ vssd1 vssd1 vccd1 vccd1 _00031_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_clkbuf_leaf_80_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11179__B1_N _03705_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_49_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07471_ _02199_ vssd1 vssd1 vccd1 vccd1 _00021_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11812__S _05613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09210_ _02170_ vssd1 vssd1 vccd1 vccd1 _03833_ sky130_fd_sc_hd__clkbuf_8
X_06422_ _01233_ _01249_ vssd1 vssd1 vccd1 vccd1 _01366_ sky130_fd_sc_hd__nor2_1
XANTENNA__07798__A genblk1\[0\].osc.clkdiv_C.cnt\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_57_762 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_17_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09141_ genblk2\[0\].wave_shpr.div.b1\[13\] genblk2\[0\].wave_shpr.div.acc\[13\]
+ vssd1 vssd1 vccd1 vccd1 _03789_ sky130_fd_sc_hd__and2b_1
XANTENNA_clkbuf_leaf_95_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06353_ _01268_ _01298_ vssd1 vssd1 vccd1 vccd1 _01299_ sky130_fd_sc_hd__nor2_1
XANTENNA__13768__RESET_B net217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08435__A2 _02350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_115_823 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09072_ genblk2\[0\].wave_shpr.div.b1\[12\] _01340_ _03722_ vssd1 vssd1 vccd1 vccd1
+ _03729_ sky130_fd_sc_hd__mux2_1
XANTENNA__07310__B _02002_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06284_ _01245_ vssd1 vssd1 vccd1 vccd1 _01246_ sky130_fd_sc_hd__buf_4
XFILLER_0_4_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_21_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08023_ _01229_ _01749_ _02729_ vssd1 vssd1 vccd1 vccd1 _02730_ sky130_fd_sc_hd__a21o_1
XFILLER_0_115_878 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold700 genblk2\[2\].wave_shpr.div.acc\[3\] vssd1 vssd1 vccd1 vccd1 net918 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_141_152 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold711 genblk2\[10\].wave_shpr.div.acc\[7\] vssd1 vssd1 vccd1 vccd1 net929 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_fanout207_A net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold722 _00026_ vssd1 vssd1 vccd1 vccd1 net940 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold733 genblk2\[10\].wave_shpr.div.acc\[10\] vssd1 vssd1 vccd1 vccd1 net951 sky130_fd_sc_hd__dlygate4sd3_1
Xhold744 genblk2\[2\].wave_shpr.div.acc\[26\] vssd1 vssd1 vccd1 vccd1 net962 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__11767__B genblk1\[9\].osc.clkdiv_C.cnt\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold755 genblk2\[1\].wave_shpr.div.acc\[17\] vssd1 vssd1 vccd1 vccd1 net973 sky130_fd_sc_hd__dlygate4sd3_1
Xhold766 genblk2\[9\].wave_shpr.div.acc\[7\] vssd1 vssd1 vccd1 vccd1 net984 sky130_fd_sc_hd__dlygate4sd3_1
Xhold777 genblk2\[1\].wave_shpr.div.acc\[7\] vssd1 vssd1 vccd1 vccd1 net995 sky130_fd_sc_hd__dlygate4sd3_1
Xhold788 genblk2\[9\].wave_shpr.div.acc\[3\] vssd1 vssd1 vccd1 vccd1 net1006 sky130_fd_sc_hd__dlygate4sd3_1
X_09974_ genblk2\[3\].wave_shpr.div.acc\[8\] genblk2\[3\].wave_shpr.div.b1\[8\] vssd1
+ vssd1 vccd1 vccd1 _04370_ sky130_fd_sc_hd__or2b_1
Xhold799 genblk2\[3\].wave_shpr.div.acc\[13\] vssd1 vssd1 vccd1 vccd1 net1017 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10950__B1 _05055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_792 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_33_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08925_ _03590_ _03602_ vssd1 vssd1 vccd1 vccd1 _03622_ sky130_fd_sc_hd__nor2_1
X_08856_ _03560_ _03561_ _03562_ _03557_ vssd1 vssd1 vccd1 vccd1 _03563_ sky130_fd_sc_hd__a211o_1
XANTENNA__10702__B1 _04856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09253__A _03855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07807_ _02510_ _02513_ genblk2\[0\].wave_shpr.div.fin_quo\[5\] vssd1 vssd1 vccd1
+ vccd1 _02514_ sky130_fd_sc_hd__a21oi_1
X_08787_ _03492_ _03493_ genblk2\[2\].wave_shpr.div.fin_quo\[2\] _02468_ vssd1 vssd1
+ vccd1 vccd1 _03494_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__10399__A _04477_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_79_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_48_clk_A clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07738_ _02444_ _02013_ vssd1 vssd1 vccd1 vccd1 _02445_ sky130_fd_sc_hd__nor2_1
X_07669_ _01188_ _01440_ genblk1\[10\].osc.clkdiv_C.cnt\[3\] vssd1 vssd1 vccd1 vccd1
+ _02376_ sky130_fd_sc_hd__and3_1
XFILLER_0_149_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__11722__S _00023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09408_ genblk2\[1\].wave_shpr.div.b1\[1\] genblk2\[1\].wave_shpr.div.acc\[1\] vssd1
+ vssd1 vccd1 vccd1 _03972_ sky130_fd_sc_hd__and2b_1
X_10680_ _04676_ _01670_ vssd1 vssd1 vccd1 vccd1 _04867_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_63_710 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_137_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09339_ _03917_ _03794_ vssd1 vssd1 vccd1 vccd1 _03918_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_leaf_106_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_51_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07220__B _01189_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12350_ _05941_ _05942_ vssd1 vssd1 vccd1 vccd1 _06034_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_50_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_105_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_16_681 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11301_ _05221_ vssd1 vssd1 vccd1 vccd1 _05300_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_22_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_106_889 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12281_ genblk2\[1\].wave_shpr.div.b1\[9\] _02013_ _05994_ vssd1 vssd1 vccd1 vccd1
+ _06002_ sky130_fd_sc_hd__mux2_1
XFILLER_0_132_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11232_ net370 _05251_ _05248_ net736 _05254_ vssd1 vssd1 vccd1 vccd1 _00722_ sky130_fd_sc_hd__a221o_1
XFILLER_0_132_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_31_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10073__S _04440_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11163_ genblk2\[7\].wave_shpr.div.fin_quo\[0\] _05222_ _00019_ vssd1 vssd1 vccd1
+ vccd1 _05223_ sky130_fd_sc_hd__mux2_1
XANTENNA__10941__B1 _05056_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10114_ _04465_ genblk1\[3\].osc.clkdiv_C.cnt\[7\] vssd1 vssd1 vccd1 vccd1 _04468_
+ sky130_fd_sc_hd__and2_1
X_11094_ _05055_ _05156_ _05157_ _05057_ net1130 vssd1 vssd1 vccd1 vccd1 _00681_ sky130_fd_sc_hd__a32o_1
X_10045_ _03714_ _04431_ _03717_ vssd1 vssd1 vccd1 vccd1 _00358_ sky130_fd_sc_hd__o21ai_1
XANTENNA_clkbuf_4_10_0_clk_A clknet_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold60 _00132_ vssd1 vssd1 vccd1 vccd1 net278 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold71 genblk2\[10\].wave_shpr.div.i\[4\] vssd1 vssd1 vccd1 vccd1 net289 sky130_fd_sc_hd__dlygate4sd3_1
Xhold82 genblk2\[2\].wave_shpr.div.quo\[8\] vssd1 vssd1 vccd1 vccd1 net300 sky130_fd_sc_hd__clkdlybuf4s25_1
XANTENNA__08362__B2 _02592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold93 _00553_ vssd1 vssd1 vccd1 vccd1 net311 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_86_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_98_684 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11996_ _05803_ vssd1 vssd1 vccd1 vccd1 _00937_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_97_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13735_ clknet_leaf_46_clk _01046_ net119 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.quo\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_133_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10947_ net515 _05052_ _05056_ net523 vssd1 vssd1 vccd1 vccd1 _00635_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13666_ clknet_leaf_41_clk net869 net123 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.acc\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10878_ genblk2\[6\].wave_shpr.div.acc\[25\] genblk2\[6\].wave_shpr.div.acc\[24\]
+ genblk2\[6\].wave_shpr.div.acc\[26\] _05021_ vssd1 vssd1 vccd1 vccd1 _05022_ sky130_fd_sc_hd__or4_2
XFILLER_0_38_261 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_807 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12617_ clknet_leaf_18_clk genblk1\[4\].osc.clkdiv_C.next_cnt\[2\] net80 vssd1 vssd1
+ vccd1 vccd1 genblk1\[4\].osc.clkdiv_C.cnt\[2\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_109_661 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_155_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_4_14_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_14_0_clk sky130_fd_sc_hd__clkbuf_8
X_13597_ clknet_leaf_77_clk _00912_ net208 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.acc\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_108_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07625__B1 _01576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_54_787 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12548_ clknet_leaf_61_clk genblk1\[0\].osc.clkdiv_C.next_cnt\[5\] net186 vssd1 vssd1
+ vccd1 vccd1 genblk1\[0\].osc.clkdiv_C.cnt\[5\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__06979__A2 _01363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12479_ clknet_leaf_108_clk _00041_ net152 vssd1 vssd1 vccd1 vccd1 sig_norm.acc\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_41_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_2 _01507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_124_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_10_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09772__S _04039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06971_ genblk1\[7\].osc.clkdiv_C.cnt\[6\] _01802_ _01805_ genblk1\[7\].osc.clkdiv_C.cnt\[5\]
+ _01806_ vssd1 vssd1 vccd1 vccd1 _01807_ sky130_fd_sc_hd__o221a_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08710_ _03412_ _03416_ vssd1 vssd1 vccd1 vccd1 _03417_ sky130_fd_sc_hd__xnor2_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10711__S _04821_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11488__A1 _03726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09690_ genblk2\[2\].wave_shpr.div.acc\[3\] genblk2\[2\].wave_shpr.div.b1\[3\] vssd1
+ vssd1 vccd1 vccd1 _04170_ sky130_fd_sc_hd__or2b_1
XFILLER_0_83_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08641_ _03345_ _03346_ _03347_ _02694_ vssd1 vssd1 vccd1 vccd1 _03348_ sky130_fd_sc_hd__a211o_1
X_08572_ _03277_ _03278_ genblk2\[9\].wave_shpr.div.fin_quo\[2\] _02362_ vssd1 vssd1
+ vccd1 vccd1 _03279_ sky130_fd_sc_hd__a2bb2o_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07523_ _02227_ net286 _02242_ vssd1 vssd1 vccd1 vccd1 PWM.next_pwm_out sky130_fd_sc_hd__a21o_1
XFILLER_0_76_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA_fanout157_A net158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07454_ _02147_ _02187_ vssd1 vssd1 vccd1 vccd1 _02188_ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_18_913 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_64_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_119_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__10666__B genblk1\[5\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06405_ _01172_ vssd1 vssd1 vccd1 vccd1 _01349_ sky130_fd_sc_hd__buf_4
XFILLER_0_91_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07385_ genblk1\[11\].osc.clkdiv_C.cnt\[13\] _02132_ vssd1 vssd1 vccd1 vccd1 _02136_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_146_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_17_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_8_177 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09124_ _03759_ _03770_ _03771_ vssd1 vssd1 vccd1 vccd1 _03772_ sky130_fd_sc_hd__a21o_1
XANTENNA__07040__B _01344_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06336_ genblk1\[0\].osc.clkdiv_C.cnt\[10\] _01286_ vssd1 vssd1 vccd1 vccd1 _01288_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_127_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_60_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_5_851 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_72_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09055_ _03704_ net394 _03715_ vssd1 vssd1 vccd1 vccd1 _00082_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_4_350 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06267_ _01228_ vssd1 vssd1 vccd1 vccd1 _01229_ sky130_fd_sc_hd__buf_6
XANTENNA__12373__S _05982_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_142_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_60_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10682__A _04672_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_130_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_115_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08006_ genblk1\[6\].osc.clkdiv_C.cnt\[1\] _01735_ _01738_ genblk1\[6\].osc.clkdiv_C.cnt\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02713_ sky130_fd_sc_hd__o211a_1
Xhold530 genblk2\[10\].wave_shpr.div.i\[2\] vssd1 vssd1 vccd1 vccd1 net748 sky130_fd_sc_hd__dlygate4sd3_1
X_06198_ _01163_ _01161_ vssd1 vssd1 vccd1 vccd1 PWM.next_counter\[4\] sky130_fd_sc_hd__xnor2_1
XFILLER_0_13_673 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold541 genblk2\[10\].wave_shpr.div.b1\[14\] vssd1 vssd1 vccd1 vccd1 net759 sky130_fd_sc_hd__dlygate4sd3_1
Xhold552 genblk2\[5\].wave_shpr.div.quo\[6\] vssd1 vssd1 vccd1 vccd1 net770 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07919__A1 genblk1\[8\].osc.clkdiv_C.cnt\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold563 genblk2\[4\].wave_shpr.div.quo\[5\] vssd1 vssd1 vccd1 vccd1 net781 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07919__B2 genblk1\[8\].osc.clkdiv_C.cnt\[5\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold574 genblk2\[6\].wave_shpr.div.quo\[0\] vssd1 vssd1 vccd1 vccd1 net792 sky130_fd_sc_hd__clkbuf_2
Xhold585 genblk2\[1\].wave_shpr.div.acc\[23\] vssd1 vssd1 vccd1 vccd1 net803 sky130_fd_sc_hd__dlygate4sd3_1
Xhold596 genblk2\[3\].wave_shpr.div.quo\[5\] vssd1 vssd1 vccd1 vccd1 net814 sky130_fd_sc_hd__dlygate4sd3_1
X_09957_ genblk2\[2\].wave_shpr.div.i\[1\] genblk2\[2\].wave_shpr.div.i\[0\] genblk2\[2\].wave_shpr.div.i\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04356_ sky130_fd_sc_hd__and3_1
X_08908_ _03610_ vssd1 vssd1 vccd1 vccd1 _00042_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10621__S _04834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_890 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09888_ _04191_ _04164_ vssd1 vssd1 vccd1 vccd1 _04306_ sky130_fd_sc_hd__or2b_1
X_08839_ _03540_ _03545_ vssd1 vssd1 vccd1 vccd1 _03546_ sky130_fd_sc_hd__nand2_1
XTAP_2702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_802 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11850_ _05597_ _05689_ vssd1 vssd1 vccd1 vccd1 _05690_ sky130_fd_sc_hd__xnor2_1
XTAP_2735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10801_ genblk2\[5\].wave_shpr.div.acc\[24\] vssd1 vssd1 vccd1 vccd1 _04952_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_172 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_2779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11781_ _05631_ genblk1\[9\].osc.clkdiv_C.cnt\[12\] vssd1 vssd1 vccd1 vccd1 _05640_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_137_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13520_ clknet_leaf_79_clk _00837_ net206 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.acc\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10732_ genblk2\[5\].wave_shpr.div.acc\[6\] _04900_ _04821_ vssd1 vssd1 vccd1 vccd1
+ _04901_ sky130_fd_sc_hd__mux2_1
XFILLER_0_82_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13451_ clknet_leaf_119_clk _00768_ net143 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.i\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_35_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10663_ net308 _04853_ _04857_ net770 vssd1 vssd1 vccd1 vccd1 _00550_ sky130_fd_sc_hd__a22o_1
XFILLER_0_125_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_36_754 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_35_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12402_ _05967_ _05929_ vssd1 vssd1 vccd1 vccd1 _06074_ sky130_fd_sc_hd__or2b_1
X_10594_ genblk2\[5\].wave_shpr.div.fin_quo\[0\] _04821_ _00015_ vssd1 vssd1 vccd1
+ vccd1 _04822_ sky130_fd_sc_hd__mux2_1
X_13382_ clknet_leaf_83_clk _00701_ net200 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.b1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07083__A1 genblk1\[8\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12333_ net239 _06014_ _06015_ net483 _06024_ vssd1 vssd1 vccd1 vccd1 _01053_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_105_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12264_ _05992_ vssd1 vssd1 vccd1 vccd1 _01016_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08032__B1 _02261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11215_ net822 _05246_ _05222_ _05248_ vssd1 vssd1 vccd1 vccd1 _00711_ sky130_fd_sc_hd__a22o_1
X_12195_ genblk2\[11\].wave_shpr.div.acc\[9\] genblk2\[11\].wave_shpr.div.b1\[9\]
+ vssd1 vssd1 vccd1 vccd1 _05933_ sky130_fd_sc_hd__or2b_1
XFILLER_0_102_881 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09592__S _04095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11146_ _05169_ _05204_ _05205_ vssd1 vssd1 vccd1 vccd1 _05206_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11077_ genblk2\[6\].wave_shpr.div.acc\[21\] _05145_ _05146_ vssd1 vssd1 vccd1 vccd1
+ _05147_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_37_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07138__A2 _01246_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10028_ _04423_ vssd1 vssd1 vccd1 vccd1 _00349_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__06346__B1 genblk1\[0\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_813 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_53_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_57 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08099__B1 _02805_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_86_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11979_ _05794_ vssd1 vssd1 vccd1 vccd1 _00929_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_805 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06964__B _01799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_85_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13718_ clknet_leaf_36_clk _01029_ net105 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.b1\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_117_918 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13649_ clknet_leaf_38_clk _00962_ net126 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.quo\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_54_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07861__A3 _02459_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_860 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_125 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07170_ genblk1\[9\].osc.clkdiv_C.cnt\[5\] genblk1\[9\].osc.clkdiv_C.cnt\[4\] _01960_
+ vssd1 vssd1 vccd1 vccd1 _01965_ sky130_fd_sc_hd__and3_1
X_06121_ smpl_rt_clkdiv.clkDiv_inst.next_hzX _01093_ vssd1 vssd1 vccd1 vccd1 smpl_rt_clkdiv.clkDiv_inst.next_cnt\[7\]
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_5_169 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_41_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_152_781 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_120_clk clknet_4_3_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_120_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_41_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_111_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_78_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09396__B_N genblk2\[1\].wave_shpr.div.b1\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09811_ _04069_ genblk1\[2\].osc.clkdiv_C.cnt\[1\] vssd1 vssd1 vccd1 vccd1 _04255_
+ sky130_fd_sc_hd__and2_1
XANTENNA__06585__B1 _01363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09742_ _04218_ vssd1 vssd1 vccd1 vccd1 _00268_ sky130_fd_sc_hd__clkbuf_1
X_06954_ _01791_ vssd1 vssd1 vccd1 vccd1 genblk1\[6\].osc.clkdiv_C.next_cnt\[16\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_94_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__09523__B1 _04045_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09673_ _03690_ _04153_ _04154_ vssd1 vssd1 vccd1 vccd1 _00263_ sky130_fd_sc_hd__nor3_1
X_06885_ _01349_ _01209_ _01439_ vssd1 vssd1 vccd1 vccd1 _01739_ sky130_fd_sc_hd__and3_2
XFILLER_0_118_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_2009 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08624_ _03307_ _03330_ vssd1 vssd1 vccd1 vccd1 _03331_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_96_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08555_ _02217_ _02553_ genblk2\[6\].wave_shpr.div.fin_quo\[2\] vssd1 vssd1 vccd1
+ vccd1 _03262_ sky130_fd_sc_hd__and3_1
XANTENNA__11272__S _05222_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06874__B _01578_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_77_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_147_520 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07506_ _02218_ _02221_ _02224_ _02226_ vssd1 vssd1 vccd1 vccd1 FSM.next_mode\[1\]
+ sky130_fd_sc_hd__a31oi_1
X_08486_ genblk2\[3\].wave_shpr.div.fin_quo\[4\] _02467_ _03192_ _02592_ vssd1 vssd1
+ vccd1 vccd1 _03193_ sky130_fd_sc_hd__a22o_1
XFILLER_0_64_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_164 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07051__A _01336_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07437_ genblk2\[4\].wave_shpr.div.i\[1\] _02174_ genblk2\[4\].wave_shpr.div.i\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02175_ sky130_fd_sc_hd__or3b_1
XFILLER_0_64_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_17_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_80_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_18_776 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_91_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07368_ genblk1\[11\].osc.clkdiv_C.cnt\[9\] _02119_ vssd1 vssd1 vccd1 vccd1 _02123_
+ sky130_fd_sc_hd__and2_1
XANTENNA__07065__A1 genblk1\[8\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09107_ genblk2\[0\].wave_shpr.div.acc\[8\] genblk2\[0\].wave_shpr.div.b1\[8\] vssd1
+ vssd1 vccd1 vccd1 _03755_ sky130_fd_sc_hd__or2b_1
X_06319_ _01269_ _01276_ _01277_ vssd1 vssd1 vccd1 vccd1 genblk1\[0\].osc.clkdiv_C.next_cnt\[3\]
+ sky130_fd_sc_hd__nor3_1
Xclkbuf_leaf_111_clk clknet_4_8_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_111_clk
+ sky130_fd_sc_hd__clkbuf_16
X_07299_ genblk1\[11\].osc.clkdiv_C.cnt\[9\] _01235_ vssd1 vssd1 vccd1 vccd1 _02063_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_115_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_143_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_33_768 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09038_ _02336_ net34 vssd1 vssd1 vccd1 vccd1 _03706_ sky130_fd_sc_hd__nand2_2
XFILLER_0_60_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold360 genblk2\[0\].wave_shpr.div.acc_next\[0\] vssd1 vssd1 vccd1 vccd1 net578 sky130_fd_sc_hd__dlygate4sd3_1
Xhold371 _00232_ vssd1 vssd1 vccd1 vccd1 net589 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08565__A1 _02261_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold382 genblk2\[0\].wave_shpr.div.quo\[4\] vssd1 vssd1 vccd1 vccd1 net600 sky130_fd_sc_hd__dlygate4sd3_1
X_11000_ genblk2\[6\].wave_shpr.div.acc\[2\] _05088_ _05023_ vssd1 vssd1 vccd1 vccd1
+ _05089_ sky130_fd_sc_hd__mux2_1
Xhold393 genblk2\[8\].wave_shpr.div.quo\[15\] vssd1 vssd1 vccd1 vccd1 net611 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12113__A2 _05844_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09514__B1 _04047_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12951_ clknet_leaf_125_clk _00280_ net71 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.b1\[7\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1060 genblk2\[11\].wave_shpr.div.b1\[17\] vssd1 vssd1 vccd1 vccd1 net1278 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_99_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold1071 genblk2\[0\].wave_shpr.div.b1\[7\] vssd1 vssd1 vccd1 vccd1 net1289 sky130_fd_sc_hd__dlygate4sd3_1
X_11902_ _05726_ vssd1 vssd1 vccd1 vccd1 _05727_ sky130_fd_sc_hd__inv_2
XTAP_2510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1082 sig_norm.quo\[7\] vssd1 vssd1 vccd1 vccd1 net1300 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_59_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold1093 genblk2\[7\].wave_shpr.div.quo\[1\] vssd1 vssd1 vccd1 vccd1 net1311 sky130_fd_sc_hd__dlygate4sd3_1
X_12882_ clknet_leaf_91_clk _00213_ net146 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_hold918_A genblk1\[9\].osc.clkdiv_C.cnt\[0\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11833_ genblk2\[9\].wave_shpr.div.acc\[9\] _05676_ _05673_ vssd1 vssd1 vccd1 vccd1
+ _05677_ sky130_fd_sc_hd__mux2_1
XTAP_2565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_1831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_114_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11764_ _02155_ vssd1 vssd1 vccd1 vccd1 _05631_ sky130_fd_sc_hd__clkbuf_2
XTAP_1875 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_82_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13503_ clknet_leaf_87_clk _00820_ net180 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.acc_next\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1886 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10715_ _04784_ _04887_ vssd1 vssd1 vccd1 vccd1 _04888_ sky130_fd_sc_hd__xnor2_1
XTAP_1897 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_153_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11695_ _05564_ _05585_ _05586_ vssd1 vssd1 vccd1 vccd1 _05587_ sky130_fd_sc_hd__a21o_1
XFILLER_0_125_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09587__S _04011_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07896__A net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13434_ clknet_leaf_81_clk net1011 net199 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.acc\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_713 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10646_ _04850_ vssd1 vssd1 vccd1 vccd1 _00540_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_82_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_141_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_23_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_102_clk clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_102_clk
+ sky130_fd_sc_hd__clkbuf_16
XFILLER_0_24_757 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_3_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13365_ clknet_leaf_12_clk _00684_ net53 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.i\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_10577_ _04768_ _04803_ _04804_ vssd1 vssd1 vccd1 vccd1 _04805_ sky130_fd_sc_hd__a21o_1
XFILLER_0_106_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12316_ _05835_ genblk1\[11\].osc.clkdiv_C.cnt\[3\] vssd1 vssd1 vccd1 vccd1 _06016_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_23_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13296_ clknet_leaf_87_clk _00617_ net179 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.b1\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_139_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12247_ genblk2\[11\].wave_shpr.div.fin_quo\[1\] net1310 _00005_ vssd1 vssd1 vccd1
+ vccd1 _05984_ sky130_fd_sc_hd__mux2_1
XFILLER_0_121_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_48_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12178_ genblk2\[10\].wave_shpr.div.i\[1\] genblk2\[10\].wave_shpr.div.i\[0\] genblk2\[10\].wave_shpr.div.i\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05919_ sky130_fd_sc_hd__a21o_1
XANTENNA__11560__B1 _05446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06959__B net34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11129_ _05180_ _05187_ _05188_ vssd1 vssd1 vccd1 vccd1 _05189_ sky130_fd_sc_hd__a21oi_1
XANTENNA__12042__A _05815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_3_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_14 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_64_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07136__A genblk1\[9\].osc.clkdiv_C.cnt\[15\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_155_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06670_ genblk1\[4\].osc.clkdiv_C.cnt\[2\] _01559_ _01557_ genblk1\[4\].osc.clkdiv_C.cnt\[6\]
+ vssd1 vssd1 vccd1 vccd1 _01560_ sky130_fd_sc_hd__a22o_1
XANTENNA__11791__B_N _03693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xwire27 _01692_ vssd1 vssd1 vccd1 vccd1 net27 sky130_fd_sc_hd__buf_1
XANTENNA__06975__A _01365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_59_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08340_ _03045_ _03046_ _02745_ vssd1 vssd1 vccd1 vccd1 _03047_ sky130_fd_sc_hd__o21a_1
XANTENNA__10418__A2 _04651_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09070__B _01996_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_59_687 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_19_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08271_ _02409_ vssd1 vssd1 vccd1 vccd1 _02978_ sky130_fd_sc_hd__inv_2
XFILLER_0_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_104_51 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11820__S _05613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_117_748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07222_ genblk1\[10\].osc.clkdiv_C.cnt\[1\] _02001_ _02002_ _02003_ vssd1 vssd1 vccd1
+ vccd1 _02004_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_13_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_55_882 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_61_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_15_724 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_116_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_116_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_14_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07153_ _01952_ vssd1 vssd1 vccd1 vccd1 _01953_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_144_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_125_781 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_124_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_42_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07084_ _01887_ _01895_ _01896_ vssd1 vssd1 vccd1 vccd1 genblk1\[8\].osc.clkdiv_C.next_cnt\[5\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_120_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_30_749 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08156__A2_N _01361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_1_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_112_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_100_637 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08547__A1 genblk2\[6\].wave_shpr.div.fin_quo\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
Xfanout103 net104 vssd1 vssd1 vccd1 vccd1 net103 sky130_fd_sc_hd__clkbuf_2
XANTENNA__08547__B2 genblk2\[6\].wave_shpr.div.fin_quo\[1\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XANTENNA__12343__A2 _03942_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_659 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09526__A _04042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xfanout114 net126 vssd1 vssd1 vccd1 vccd1 net114 sky130_fd_sc_hd__clkbuf_4
Xfanout125 net126 vssd1 vssd1 vccd1 vccd1 net125 sky130_fd_sc_hd__buf_2
Xfanout136 net171 vssd1 vssd1 vccd1 vccd1 net136 sky130_fd_sc_hd__clkbuf_4
Xfanout147 net171 vssd1 vssd1 vccd1 vccd1 net147 sky130_fd_sc_hd__buf_2
Xfanout158 net171 vssd1 vssd1 vccd1 vccd1 net158 sky130_fd_sc_hd__clkbuf_2
X_07986_ _02691_ _02682_ _02690_ _02527_ vssd1 vssd1 vccd1 vccd1 _02693_ sky130_fd_sc_hd__o31a_1
Xfanout169 net170 vssd1 vssd1 vccd1 vccd1 net169 sky130_fd_sc_hd__clkbuf_4
XANTENNA__07770__A2 _01240_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09725_ genblk2\[2\].wave_shpr.div.b1\[16\] genblk2\[2\].wave_shpr.div.acc\[16\]
+ vssd1 vssd1 vccd1 vccd1 _04205_ sky130_fd_sc_hd__and2b_1
X_06937_ net28 _01779_ vssd1 vssd1 vccd1 vccd1 _01780_ sky130_fd_sc_hd__nor2_1
XANTENNA__11303__B1 _05283_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_97_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09656_ genblk2\[1\].wave_shpr.div.acc\[24\] _04008_ vssd1 vssd1 vccd1 vccd1 _04143_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__10657__A2 _04853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06868_ genblk1\[5\].osc.clkdiv_C.cnt\[16\] _01721_ vssd1 vssd1 vccd1 vccd1 _01724_
+ sky130_fd_sc_hd__nand2_1
XANTENNA__06885__A _01349_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_96_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09261__A _03853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08607_ genblk2\[5\].wave_shpr.div.fin_quo\[0\] vssd1 vssd1 vccd1 vccd1 _03314_ sky130_fd_sc_hd__inv_2
XTAP_1105 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_96_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1116 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09587_ genblk2\[1\].wave_shpr.div.acc\[6\] _04091_ _04011_ vssd1 vssd1 vccd1 vccd1
+ _04092_ sky130_fd_sc_hd__mux2_1
XTAP_1127 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06799_ genblk1\[5\].osc.clkdiv_C.cnt\[14\] _01210_ _01304_ genblk1\[5\].osc.clkdiv_C.cnt\[1\]
+ _01670_ vssd1 vssd1 vccd1 vccd1 _01671_ sky130_fd_sc_hd__a221o_1
XTAP_1138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08538_ _03243_ _03244_ vssd1 vssd1 vccd1 vccd1 _03245_ sky130_fd_sc_hd__and2_1
XFILLER_0_154_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_64_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08469_ genblk2\[5\].wave_shpr.div.fin_quo\[2\] vssd1 vssd1 vccd1 vccd1 _03176_ sky130_fd_sc_hd__inv_2
XANTENNA__11730__S _00023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10500_ _04618_ _04738_ vssd1 vssd1 vccd1 vccd1 _04740_ sky130_fd_sc_hd__or2_1
XFILLER_0_64_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_107_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11480_ genblk2\[9\].wave_shpr.div.b1\[11\] _01732_ _05433_ vssd1 vssd1 vccd1 vccd1
+ _05437_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_830 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07038__A1 _01436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10431_ _04586_ _04687_ vssd1 vssd1 vccd1 vccd1 _04688_ sky130_fd_sc_hd__xnor2_1
XANTENNA__08235__B1 _02467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_123_729 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_122_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__12127__A _05815_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_33_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_13150_ clknet_leaf_121_clk net681 net80 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.quo\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10362_ _03726_ _04649_ _03736_ vssd1 vssd1 vccd1 vccd1 _00457_ sky130_fd_sc_hd__o21ai_1
X_12101_ _05760_ _05741_ vssd1 vssd1 vccd1 vccd1 _05863_ sky130_fd_sc_hd__or2b_1
XANTENNA__11790__B1 _03693_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_130_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13081_ clknet_leaf_126_clk _00408_ net63 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.acc\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10293_ _04571_ _04603_ _04604_ vssd1 vssd1 vccd1 vccd1 _04605_ sky130_fd_sc_hd__a21o_1
XFILLER_0_130_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_12032_ _02155_ vssd1 vssd1 vccd1 vccd1 _05819_ sky130_fd_sc_hd__clkbuf_2
Xhold190 genblk2\[4\].wave_shpr.div.quo\[7\] vssd1 vssd1 vccd1 vccd1 net408 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07210__A1 _01359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07303__A2_N _01256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12934_ clknet_leaf_30_clk _00263_ net102 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.i\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_125_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12865_ clknet_leaf_135_clk _00196_ net61 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.b1\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_11816_ genblk2\[9\].wave_shpr.div.acc\[5\] _05663_ _05613_ vssd1 vssd1 vccd1 vccd1
+ _05664_ sky130_fd_sc_hd__mux2_1
XTAP_2384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_max_cap34_A _01794_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12796_ clknet_leaf_92_clk _00129_ net149 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_145_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_141_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11747_ genblk2\[9\].wave_shpr.div.quo\[2\] _05623_ _05624_ net649 vssd1 vssd1 vccd1
+ vccd1 _00867_ sky130_fd_sc_hd__a22o_1
XTAP_1694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12270__A1 _04229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_139_895 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_4_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11678_ genblk2\[9\].wave_shpr.div.acc\[3\] genblk2\[9\].wave_shpr.div.b1\[3\] vssd1
+ vssd1 vccd1 vccd1 _05570_ sky130_fd_sc_hd__or2b_1
X_13417_ clknet_leaf_119_clk _00736_ net141 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.acc_next\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_10629_ _04841_ vssd1 vssd1 vccd1 vccd1 _00532_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_12_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_3_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_51_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13348_ clknet_leaf_5_clk _00669_ net45 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.acc\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_122_751 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_122_773 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13279_ clknet_leaf_11_clk _00600_ net56 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.i\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__10336__A1 _01256_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07840_ _02536_ _02546_ vssd1 vssd1 vccd1 vccd1 _02547_ sky130_fd_sc_hd__nor2_1
XANTENNA__09780__S _04238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07752__A2 _01577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07771_ _02475_ _02477_ vssd1 vssd1 vccd1 vccd1 _02478_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09510_ _04046_ vssd1 vssd1 vccd1 vccd1 _04047_ sky130_fd_sc_hd__buf_4
X_06722_ genblk1\[4\].osc.clkdiv_C.cnt\[3\] _01605_ vssd1 vssd1 vccd1 vccd1 _01609_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_78_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_149_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09441_ _03954_ _04003_ _04004_ vssd1 vssd1 vccd1 vccd1 _04005_ sky130_fd_sc_hd__a21o_1
XFILLER_0_78_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06653_ _01523_ _01547_ vssd1 vssd1 vccd1 vccd1 _01548_ sky130_fd_sc_hd__nor2_1
XFILLER_0_149_648 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_47_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_91_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07313__B _01439_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09372_ _03940_ vssd1 vssd1 vccd1 vccd1 _03941_ sky130_fd_sc_hd__buf_4
XFILLER_0_47_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06584_ genblk1\[3\].osc.clkdiv_C.cnt\[10\] _01231_ _01488_ _01490_ _01491_ vssd1
+ vssd1 vccd1 vccd1 _01492_ sky130_fd_sc_hd__a221o_1
XFILLER_0_115_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08323_ _03013_ _03029_ vssd1 vssd1 vccd1 vccd1 _03030_ sky130_fd_sc_hd__and2_1
XFILLER_0_86_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12261__A1 _01329_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_808 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_90_903 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08254_ genblk2\[6\].wave_shpr.div.fin_quo\[5\] _02733_ _02959_ _02261_ vssd1 vssd1
+ vccd1 vccd1 _02961_ sky130_fd_sc_hd__a31o_1
XFILLER_0_145_865 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_6_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_15_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_43_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07205_ _01954_ _01987_ _01988_ vssd1 vssd1 vccd1 vccd1 _01989_ sky130_fd_sc_hd__and3_1
XANTENNA__06491__A2 _01363_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__12013__A1 _03726_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08185_ genblk2\[3\].wave_shpr.div.fin_quo\[7\] _02539_ vssd1 vssd1 vccd1 vccd1 _02892_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_104_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08144__B _01576_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_132_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07136_ genblk1\[9\].osc.clkdiv_C.cnt\[15\] _01361_ vssd1 vssd1 vccd1 vccd1 _01936_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07067_ _01863_ _01872_ _01873_ _01884_ vssd1 vssd1 vccd1 vccd1 _01885_ sky130_fd_sc_hd__or4b_1
XANTENNA__06243__A2 _01197_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_11_760 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_771 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08160__A _01489_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06599__B _01249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07969_ _02650_ _02667_ _02675_ vssd1 vssd1 vccd1 vccd1 _02676_ sky130_fd_sc_hd__a21oi_2
X_09708_ _04166_ _04186_ _04187_ vssd1 vssd1 vccd1 vccd1 _04188_ sky130_fd_sc_hd__a21o_1
X_10980_ net609 _05051_ _05064_ net616 _05075_ vssd1 vssd1 vccd1 vccd1 _00649_ sky130_fd_sc_hd__a221o_1
XANTENNA__07504__A net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09639_ _04130_ _04131_ vssd1 vssd1 vccd1 vccd1 _04132_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12650_ clknet_leaf_10_clk genblk1\[5\].osc.clkdiv_C.next_cnt\[17\] net57 vssd1 vssd1
+ vccd1 vccd1 genblk1\[5\].osc.clkdiv_C.cnt\[17\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_84_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10566__A_N genblk2\[5\].wave_shpr.div.b1\[7\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_78_782 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08038__C _02365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11601_ _05397_ _05511_ vssd1 vssd1 vccd1 vccd1 _05512_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_155_629 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_136_810 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_136_821 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12581_ clknet_leaf_14_clk genblk1\[2\].osc.clkdiv_C.next_cnt\[2\] net70 vssd1 vssd1
+ vccd1 vccd1 genblk1\[2\].osc.clkdiv_C.cnt\[2\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_26_819 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_92_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_93_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11532_ _05450_ genblk1\[8\].osc.clkdiv_C.cnt\[10\] vssd1 vssd1 vccd1 vccd1 _05463_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_147_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_136_865 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_19_893 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_92_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_92_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_46_690 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12004__A1 _01500_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_108_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11463_ _05428_ vssd1 vssd1 vccd1 vccd1 _00779_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__08054__B _01223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13202_ clknet_leaf_8_clk _00525_ net55 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.b1\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_61_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_10414_ _03719_ vssd1 vssd1 vccd1 vccd1 _04676_ sky130_fd_sc_hd__buf_6
X_11394_ genblk2\[8\].wave_shpr.div.acc\[5\] genblk2\[8\].wave_shpr.div.b1\[5\] vssd1
+ vssd1 vccd1 vccd1 _05370_ sky130_fd_sc_hd__or2b_1
X_13133_ clknet_leaf_0_clk _00458_ net41 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.b1\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_103_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10345_ net1303 _04639_ _04637_ vssd1 vssd1 vccd1 vccd1 _04640_ sky130_fd_sc_hd__mux2_1
XFILLER_0_103_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12307__A2 _06009_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13064_ clknet_leaf_29_clk _00391_ net95 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.quo\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10276_ _04582_ _04586_ _04587_ vssd1 vssd1 vccd1 vccd1 _04588_ sky130_fd_sc_hd__a21o_1
XANTENNA__11515__B1 _05449_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12015_ _05811_ vssd1 vssd1 vccd1 vccd1 _00948_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__10105__A _04269_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06302__B _01263_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_136_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xmax_cap3 _03923_ vssd1 vssd1 vccd1 vccd1 net1352 sky130_fd_sc_hd__buf_1
X_12917_ clknet_leaf_35_clk _00248_ net105 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.acc\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11294__A2 _05279_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_152_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_2170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12848_ clknet_leaf_58_clk _00179_ net194 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.i\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_118_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12779_ clknet_leaf_41_clk _00112_ net116 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.b1\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__06972__B _01214_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_124_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_43_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_813 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_841 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_43_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_153_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_9_69 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_25_874 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09775__S _04039_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_4_757 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold904 genblk2\[6\].wave_shpr.div.acc\[1\] vssd1 vssd1 vccd1 vccd1 net1122 sky130_fd_sc_hd__dlygate4sd3_1
Xhold915 genblk1\[0\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 net1133 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold926 genblk2\[4\].wave_shpr.div.acc\[24\] vssd1 vssd1 vccd1 vccd1 net1144 sky130_fd_sc_hd__dlygate4sd3_1
Xhold937 sig_norm.acc\[6\] vssd1 vssd1 vccd1 vccd1 net1155 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_10_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold948 genblk1\[2\].osc.clkdiv_C.cnt\[13\] vssd1 vssd1 vccd1 vccd1 net1166 sky130_fd_sc_hd__dlygate4sd3_1
X_09990_ genblk2\[3\].wave_shpr.div.b1\[3\] genblk2\[3\].wave_shpr.div.acc\[3\] vssd1
+ vssd1 vccd1 vccd1 _04386_ sky130_fd_sc_hd__and2b_1
Xhold959 genblk2\[6\].wave_shpr.div.i\[3\] vssd1 vssd1 vccd1 vccd1 net1177 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_122_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08941_ _03540_ _03550_ vssd1 vssd1 vccd1 vccd1 _03633_ sky130_fd_sc_hd__or2_1
XFILLER_0_86_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11506__B1 _05446_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08872_ sig_norm.acc\[0\] vssd1 vssd1 vccd1 vccd1 _03578_ sky130_fd_sc_hd__inv_2
XFILLER_0_19_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07823_ _02469_ _02528_ _02529_ vssd1 vssd1 vccd1 vccd1 _02530_ sky130_fd_sc_hd__o21ai_1
X_07754_ _02460_ vssd1 vssd1 vccd1 vccd1 _02461_ sky130_fd_sc_hd__clkbuf_2
X_06705_ _01489_ _01196_ vssd1 vssd1 vccd1 vccd1 _01595_ sky130_fd_sc_hd__nor2_4
XFILLER_0_67_708 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_07685_ _02390_ _02391_ _01995_ _02016_ vssd1 vssd1 vccd1 vccd1 _02392_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__08139__B _02364_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_91_clk clknet_4_9_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_91_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__08150__A2 _01234_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_149_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09424_ genblk2\[1\].wave_shpr.div.b1\[9\] genblk2\[1\].wave_shpr.div.acc\[9\] vssd1
+ vssd1 vccd1 vccd1 _03988_ sky130_fd_sc_hd__and2b_1
XANTENNA_hold1002_A genblk1\[11\].osc.clkdiv_C.cnt\[17\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06636_ genblk1\[3\].osc.clkdiv_C.cnt\[7\] _01535_ _01524_ vssd1 vssd1 vccd1 vccd1
+ _01537_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_47_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09355_ net1032 _03903_ _03910_ _03929_ vssd1 vssd1 vccd1 vccd1 _00170_ sky130_fd_sc_hd__a22o_1
X_06567_ genblk1\[2\].osc.clkdiv_C.cnt\[15\] genblk1\[2\].osc.clkdiv_C.cnt\[14\] _01474_
+ vssd1 vssd1 vccd1 vccd1 _01478_ sky130_fd_sc_hd__and3_1
XFILLER_0_74_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08306_ _03012_ _02989_ vssd1 vssd1 vccd1 vccd1 _03013_ sky130_fd_sc_hd__xnor2_1
X_09286_ _03838_ vssd1 vssd1 vccd1 vccd1 _03877_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_35_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_19_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_7_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06498_ genblk1\[2\].osc.clkdiv_C.cnt\[2\] net36 vssd1 vssd1 vccd1 vccd1 _01424_
+ sky130_fd_sc_hd__nand2_1
XANTENNA_clkbuf_leaf_7_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_145_673 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_34_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_62_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08237_ _02939_ _02942_ _02943_ vssd1 vssd1 vccd1 vccd1 _02944_ sky130_fd_sc_hd__o21a_1
XFILLER_0_105_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_133_835 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08168_ _02872_ _02873_ _02874_ vssd1 vssd1 vccd1 vccd1 _02875_ sky130_fd_sc_hd__nand3_1
XFILLER_0_31_844 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11745__B1 _05624_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07119_ genblk1\[9\].osc.clkdiv_C.cnt\[10\] _01227_ vssd1 vssd1 vccd1 vccd1 _01919_
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__10624__S _04834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08099_ genblk1\[4\].osc.clkdiv_C.cnt\[13\] _01498_ _02805_ genblk1\[4\].osc.clkdiv_C.cnt\[12\]
+ vssd1 vssd1 vccd1 vccd1 _02806_ sky130_fd_sc_hd__o22a_1
XFILLER_0_100_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10130_ _04465_ genblk1\[3\].osc.clkdiv_C.cnt\[15\] vssd1 vssd1 vccd1 vccd1 _04476_
+ sky130_fd_sc_hd__and2_1
XANTENNA__06403__A genblk1\[1\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10061_ _03701_ vssd1 vssd1 vccd1 vccd1 _04440_ sky130_fd_sc_hd__buf_4
XFILLER_0_98_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13751_ clknet_leaf_74_clk _01062_ net212 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.acc\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_15_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10963_ net498 _05062_ _05064_ genblk2\[6\].wave_shpr.div.quo\[13\] _05066_ vssd1
+ vssd1 vccd1 vccd1 _00641_ sky130_fd_sc_hd__a221o_1
XANTENNA__08049__B _01355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_82_clk clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_82_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_85_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12702_ clknet_leaf_89_clk genblk1\[8\].osc.clkdiv_C.next_cnt\[15\] net173 vssd1
+ vssd1 vccd1 vccd1 genblk1\[8\].osc.clkdiv_C.cnt\[15\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_97_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13682_ clknet_leaf_42_clk _00995_ net190 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.acc\[20\]
+ sky130_fd_sc_hd__dfrtp_1
X_10894_ genblk2\[6\].wave_shpr.div.fin_quo\[7\] net1349 _00017_ vssd1 vssd1 vccd1
+ vccd1 _05031_ sky130_fd_sc_hd__mux2_1
X_12633_ clknet_leaf_16_clk genblk1\[5\].osc.clkdiv_C.next_cnt\[0\] net74 vssd1 vssd1
+ vccd1 vccd1 genblk1\[5\].osc.clkdiv_C.cnt\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_155_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_127_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_122_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_31_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10236__B1 _04454_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_53_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12564_ clknet_leaf_29_clk genblk1\[1\].osc.clkdiv_C.next_cnt\[3\] net96 vssd1 vssd1
+ vccd1 vccd1 genblk1\[1\].osc.clkdiv_C.cnt\[3\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_108_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_142_109 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11515_ genblk2\[8\].wave_shpr.div.quo\[11\] _05448_ _05449_ net469 _05453_ vssd1
+ vssd1 vccd1 vccd1 _00806_ sky130_fd_sc_hd__a221o_1
XFILLER_0_123_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12495_ clknet_leaf_104_clk _00057_ net153 vssd1 vssd1 vccd1 vccd1 sig_norm.quo\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_107 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11446_ genblk2\[8\].wave_shpr.div.fin_quo\[2\] genblk2\[8\].wave_shpr.div.quo\[1\]
+ _00021_ vssd1 vssd1 vccd1 vccd1 _05420_ sky130_fd_sc_hd__mux2_1
XFILLER_0_123_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_1_705 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_153 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_321 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11377_ _00018_ _05353_ net1181 vssd1 vssd1 vccd1 vccd1 _05355_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_150_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_0_237 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12315__A _03941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13116_ clknet_leaf_2_clk _00441_ net52 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.b1\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10328_ genblk2\[5\].wave_shpr.div.b1\[0\] _01735_ _04440_ vssd1 vssd1 vccd1 vccd1
+ _04632_ sky130_fd_sc_hd__mux2_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__09157__A1 _03804_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13047_ clknet_leaf_129_clk _00374_ net65 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.b1\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10259_ genblk2\[4\].wave_shpr.div.acc\[11\] genblk2\[4\].wave_shpr.div.b1\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04571_ sky130_fd_sc_hd__or2b_1
XFILLER_0_56_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_89_800 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08380__A2 _01209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_76_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_73_clk clknet_4_15_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_73_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_72_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07470_ _02196_ _02153_ genblk2\[8\].wave_shpr.div.busy vssd1 vssd1 vccd1 vccd1 _02199_
+ sky130_fd_sc_hd__and3b_1
XANTENNA__06983__A _01436_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06421_ _01336_ vssd1 vssd1 vccd1 vccd1 _01365_ sky130_fd_sc_hd__buf_8
XANTENNA__06694__A2 _01313_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07798__B genblk1\[0\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09140_ _03751_ _03786_ _03787_ vssd1 vssd1 vccd1 vccd1 _03788_ sky130_fd_sc_hd__a21o_1
X_06352_ genblk1\[0\].osc.clkdiv_C.cnt\[16\] genblk1\[0\].osc.clkdiv_C.cnt\[15\] _01295_
+ vssd1 vssd1 vccd1 vccd1 _01298_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_16_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_126_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_06283_ _01173_ _01187_ vssd1 vssd1 vccd1 vccd1 _01245_ sky130_fd_sc_hd__or2_2
XFILLER_0_114_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09071_ _03726_ net1084 _01302_ _03727_ _03728_ vssd1 vssd1 vccd1 vccd1 _00087_ sky130_fd_sc_hd__o221a_1
XFILLER_0_32_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08022_ _02709_ _02708_ _02728_ vssd1 vssd1 vccd1 vccd1 _02729_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_112_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_21_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07134__A2_N _01311_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold701 genblk2\[2\].wave_shpr.div.acc\[5\] vssd1 vssd1 vccd1 vccd1 net919 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold712 genblk2\[3\].wave_shpr.div.acc\[15\] vssd1 vssd1 vccd1 vccd1 net930 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold723 genblk2\[3\].wave_shpr.div.acc\[6\] vssd1 vssd1 vccd1 vccd1 net941 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_4_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold734 genblk2\[2\].wave_shpr.div.acc\[10\] vssd1 vssd1 vccd1 vccd1 net952 sky130_fd_sc_hd__dlygate4sd3_1
Xhold745 genblk2\[3\].wave_shpr.div.acc\[5\] vssd1 vssd1 vccd1 vccd1 net963 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold756 genblk2\[9\].wave_shpr.div.acc\[9\] vssd1 vssd1 vccd1 vccd1 net974 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07946__A2 _01574_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold767 genblk2\[11\].wave_shpr.div.acc\[4\] vssd1 vssd1 vccd1 vccd1 net985 sky130_fd_sc_hd__dlygate4sd3_1
Xhold778 PWM.counter\[3\] vssd1 vssd1 vccd1 vccd1 net996 sky130_fd_sc_hd__dlygate4sd3_1
X_09973_ genblk2\[3\].wave_shpr.div.acc\[9\] genblk2\[3\].wave_shpr.div.b1\[9\] vssd1
+ vssd1 vccd1 vccd1 _04369_ sky130_fd_sc_hd__or2b_1
Xhold789 genblk2\[11\].wave_shpr.div.b1\[0\] vssd1 vssd1 vccd1 vccd1 net1007 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07149__A2_N _01799_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08924_ net717 _02260_ _03621_ _03574_ vssd1 vssd1 vccd1 vccd1 _00047_ sky130_fd_sc_hd__a22o_1
X_08855_ _03498_ _03553_ _03554_ vssd1 vssd1 vccd1 vccd1 _03562_ sky130_fd_sc_hd__nor3_1
XANTENNA__11783__B genblk1\[9\].osc.clkdiv_C.cnt\[13\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06877__B _01249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07806_ genblk2\[0\].wave_shpr.div.fin_quo\[4\] _02512_ vssd1 vssd1 vccd1 vccd1 _02513_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_137_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08786_ genblk2\[2\].wave_shpr.div.fin_quo\[0\] genblk2\[2\].wave_shpr.div.fin_quo\[1\]
+ _03113_ _02224_ vssd1 vssd1 vccd1 vccd1 _03493_ sky130_fd_sc_hd__a31o_1
X_07737_ genblk1\[1\].osc.clkdiv_C.cnt\[8\] vssd1 vssd1 vccd1 vccd1 _02444_ sky130_fd_sc_hd__inv_2
Xclkbuf_leaf_64_clk clknet_4_13_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_64_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__08123__A2 _01224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_138_905 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_67_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06893__A _01308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07668_ genblk1\[10\].osc.clkdiv_C.cnt\[3\] _02374_ _02013_ genblk1\[10\].osc.clkdiv_C.cnt\[2\]
+ vssd1 vssd1 vccd1 vccd1 _02375_ sky130_fd_sc_hd__o22a_1
XFILLER_0_1_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_137_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_94_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09407_ genblk2\[1\].wave_shpr.div.acc\[0\] genblk2\[1\].wave_shpr.div.b1\[0\] vssd1
+ vssd1 vccd1 vccd1 _03971_ sky130_fd_sc_hd__or2b_1
X_06619_ genblk1\[3\].osc.clkdiv_C.cnt\[1\] genblk1\[3\].osc.clkdiv_C.cnt\[0\] vssd1
+ vssd1 vccd1 vccd1 _01526_ sky130_fd_sc_hd__or2_1
XFILLER_0_137_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_48_763 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07599_ _02261_ _02305_ vssd1 vssd1 vccd1 vccd1 _02306_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_48_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09338_ _03795_ _03747_ vssd1 vssd1 vccd1 vccd1 _03917_ sky130_fd_sc_hd__or2b_1
XFILLER_0_47_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07501__B net18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_152_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_62_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_51_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_63_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_118_695 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09269_ net715 _00000_ _03863_ net578 _03864_ vssd1 vssd1 vccd1 vccd1 _00149_ sky130_fd_sc_hd__o221a_1
XFILLER_0_133_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_106_857 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11300_ _05196_ _05298_ vssd1 vssd1 vccd1 vccd1 _05299_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_133_643 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12280_ _06001_ vssd1 vssd1 vccd1 vccd1 _01023_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_121_838 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11231_ _05074_ genblk1\[7\].osc.clkdiv_C.cnt\[2\] vssd1 vssd1 vccd1 vccd1 _05254_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_31_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07229__A _01229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11162_ _05221_ vssd1 vssd1 vccd1 vccd1 _05222_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_184 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06133__A net8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10113_ net514 _04461_ _04462_ net634 _04467_ vssd1 vssd1 vccd1 vccd1 _00390_ sky130_fd_sc_hd__a221o_1
X_11093_ genblk2\[6\].wave_shpr.div.i\[1\] genblk2\[6\].wave_shpr.div.i\[0\] vssd1
+ vssd1 vccd1 vccd1 _05157_ sky130_fd_sc_hd__nand2_1
X_10044_ net1100 vssd1 vssd1 vccd1 vccd1 _04431_ sky130_fd_sc_hd__inv_2
Xhold50 _00872_ vssd1 vssd1 vccd1 vccd1 net268 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06787__B _01658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08362__A2 _02539_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold61 sig_norm.i\[3\] vssd1 vssd1 vccd1 vccd1 net279 sky130_fd_sc_hd__dlygate4sd3_1
Xhold72 genblk2\[9\].wave_shpr.div.quo\[9\] vssd1 vssd1 vccd1 vccd1 net290 sky130_fd_sc_hd__dlygate4sd3_1
Xhold83 _00300_ vssd1 vssd1 vccd1 vccd1 net301 sky130_fd_sc_hd__dlygate4sd3_1
Xhold94 genblk2\[8\].wave_shpr.div.quo\[13\] vssd1 vssd1 vccd1 vccd1 net312 sky130_fd_sc_hd__dlygate4sd3_1
X_11995_ net1242 _02805_ _05802_ vssd1 vssd1 vccd1 vccd1 _05803_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_55_clk clknet_4_12_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_55_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_58_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13734_ clknet_leaf_46_clk net444 net119 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.quo\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_10946_ genblk2\[6\].wave_shpr.div.quo\[7\] _05052_ _05056_ net241 vssd1 vssd1 vccd1
+ vccd1 _00634_ sky130_fd_sc_hd__a22o_1
XFILLER_0_97_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_133_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_86_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13665_ clknet_leaf_43_clk _00978_ net123 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.acc\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10877_ genblk2\[6\].wave_shpr.div.acc\[23\] _05020_ vssd1 vssd1 vccd1 vccd1 _05021_
+ sky130_fd_sc_hd__or2_2
XFILLER_0_85_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12616_ clknet_leaf_18_clk genblk1\[4\].osc.clkdiv_C.next_cnt\[1\] net80 vssd1 vssd1
+ vccd1 vccd1 genblk1\[4\].osc.clkdiv_C.cnt\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_38_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13596_ clknet_leaf_77_clk net936 net208 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.acc\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06428__A2 _01304_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12547_ clknet_leaf_61_clk genblk1\[0\].osc.clkdiv_C.next_cnt\[4\] net186 vssd1 vssd1
+ vccd1 vccd1 genblk1\[0\].osc.clkdiv_C.cnt\[4\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_13_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12478_ clknet_leaf_108_clk _00040_ net152 vssd1 vssd1 vccd1 vccd1 sig_norm.acc\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_3 _01507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_630 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_22_652 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11429_ _05360_ _05403_ _05404_ vssd1 vssd1 vccd1 vccd1 _05405_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08242__B _02309_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11185__B2 _03687_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_21_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_10_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06970_ genblk1\[7\].osc.clkdiv_C.cnt\[5\] _01805_ _01801_ genblk1\[7\].osc.clkdiv_C.cnt\[1\]
+ vssd1 vssd1 vccd1 vccd1 _01806_ sky130_fd_sc_hd__o2bb2a_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08640_ _02216_ _02553_ genblk2\[7\].wave_shpr.div.fin_quo\[3\] vssd1 vssd1 vccd1
+ vccd1 _03347_ sky130_fd_sc_hd__and3_1
XANTENNA__10696__B1 _04856_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_107_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08571_ genblk2\[9\].wave_shpr.div.fin_quo\[0\] genblk2\[9\].wave_shpr.div.fin_quo\[1\]
+ _02303_ _02316_ vssd1 vssd1 vccd1 vccd1 _03278_ sky130_fd_sc_hd__a31o_1
XFILLER_0_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_46_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_46_clk sky130_fd_sc_hd__clkbuf_16
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_77_825 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_89_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07522_ _02227_ net286 _02229_ _02241_ vssd1 vssd1 vccd1 vccd1 _02242_ sky130_fd_sc_hd__o22a_1
XANTENNA__07602__A _02308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07453_ genblk2\[6\].wave_shpr.div.busy _02186_ vssd1 vssd1 vccd1 vccd1 _02187_ sky130_fd_sc_hd__and2_1
XFILLER_0_64_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_9_646 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06404_ genblk1\[1\].osc.clkdiv_C.cnt\[14\] _01327_ vssd1 vssd1 vccd1 vccd1 _01348_
+ sky130_fd_sc_hd__and2_1
XANTENNA__07321__B _01359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07384_ genblk1\[11\].osc.clkdiv_C.cnt\[13\] _02132_ vssd1 vssd1 vccd1 vccd1 _02135_
+ sky130_fd_sc_hd__or2_1
X_09123_ genblk2\[0\].wave_shpr.div.b1\[4\] genblk2\[0\].wave_shpr.div.acc\[4\] vssd1
+ vssd1 vccd1 vccd1 _03771_ sky130_fd_sc_hd__and2b_1
XFILLER_0_134_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_72_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_8_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_06335_ _01269_ _01286_ _01287_ vssd1 vssd1 vccd1 vccd1 genblk1\[0\].osc.clkdiv_C.next_cnt\[9\]
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_115_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_44_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_5_863 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_736 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09054_ _03714_ net727 _03715_ _03717_ vssd1 vssd1 vccd1 vccd1 _00081_ sky130_fd_sc_hd__o211a_1
X_06266_ _01194_ vssd1 vssd1 vccd1 vccd1 _01228_ sky130_fd_sc_hd__inv_2
XFILLER_0_4_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_373 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08005_ _02700_ _02703_ _02711_ vssd1 vssd1 vccd1 vccd1 _02712_ sky130_fd_sc_hd__a21boi_1
Xhold520 _00378_ vssd1 vssd1 vccd1 vccd1 net738 sky130_fd_sc_hd__dlygate4sd3_1
Xhold531 genblk2\[4\].wave_shpr.div.quo\[4\] vssd1 vssd1 vccd1 vccd1 net749 sky130_fd_sc_hd__dlygate4sd3_1
X_06197_ net1307 vssd1 vssd1 vccd1 vccd1 _01163_ sky130_fd_sc_hd__inv_2
Xhold542 modein.delay_in\[1\] vssd1 vssd1 vccd1 vccd1 net760 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__07919__A2 _01430_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_12_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
Xhold553 genblk2\[1\].wave_shpr.div.quo\[5\] vssd1 vssd1 vccd1 vccd1 net771 sky130_fd_sc_hd__dlygate4sd3_1
Xhold564 genblk2\[2\].wave_shpr.div.acc\[1\] vssd1 vssd1 vccd1 vccd1 net782 sky130_fd_sc_hd__dlygate4sd3_1
Xhold575 genblk2\[4\].wave_shpr.div.quo\[2\] vssd1 vssd1 vccd1 vccd1 net793 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_12_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold586 genblk2\[0\].wave_shpr.div.quo\[0\] vssd1 vssd1 vccd1 vccd1 net804 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold597 _00381_ vssd1 vssd1 vccd1 vccd1 net815 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08592__A2 _02527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09956_ genblk2\[2\].wave_shpr.div.i\[1\] genblk2\[2\].wave_shpr.div.i\[0\] genblk2\[2\].wave_shpr.div.i\[2\]
+ vssd1 vssd1 vccd1 vccd1 _04355_ sky130_fd_sc_hd__a21o_1
XANTENNA__10902__S _04848_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06888__A _01658_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_110_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08907_ _03609_ net1240 _01157_ vssd1 vssd1 vccd1 vccd1 _03610_ sky130_fd_sc_hd__mux2_1
XTAP_880 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09887_ net895 _04282_ _04289_ _04305_ vssd1 vssd1 vccd1 vccd1 _00326_ sky130_fd_sc_hd__a22o_1
XTAP_891 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08838_ _03542_ _03544_ vssd1 vssd1 vccd1 vccd1 _03545_ sky130_fd_sc_hd__and2_1
XTAP_2703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08769_ _03457_ _03459_ vssd1 vssd1 vccd1 vccd1 _03476_ sky130_fd_sc_hd__or2b_1
XTAP_2725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_37_clk clknet_4_7_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_37_clk sky130_fd_sc_hd__clkbuf_16
XTAP_2747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10800_ _04819_ _04855_ _04951_ _04858_ net1038 vssd1 vssd1 vccd1 vccd1 _00593_ sky130_fd_sc_hd__a32o_1
XTAP_2758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_11780_ genblk2\[9\].wave_shpr.div.quo\[20\] _05628_ _05629_ net362 _05639_ vssd1
+ vssd1 vccd1 vccd1 _00885_ sky130_fd_sc_hd__a221o_1
XANTENNA__07304__B1 _01925_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09844__A2 _04247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_68_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09203__S _03822_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_94_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10731_ _04791_ _04899_ vssd1 vssd1 vccd1 vccd1 _04900_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_95_666 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__10349__S _04637_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_82_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_36_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13450_ clknet_leaf_119_clk _00767_ net143 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.i\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_94_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_10662_ genblk2\[5\].wave_shpr.div.quo\[6\] _04853_ _04857_ net253 vssd1 vssd1 vccd1
+ vccd1 _00549_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_35_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__06128__A net13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_727 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_137_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12401_ _03941_ vssd1 vssd1 vccd1 vccd1 _06073_ sky130_fd_sc_hd__clkbuf_4
X_13381_ clknet_leaf_96_clk _00700_ net167 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.b1\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_10593_ _04820_ vssd1 vssd1 vccd1 vccd1 _04821_ sky130_fd_sc_hd__buf_4
XFILLER_0_91_883 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_118_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_50_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_91_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12332_ _03833_ _02128_ vssd1 vssd1 vccd1 vccd1 _06024_ sky130_fd_sc_hd__nor2_1
XFILLER_0_106_665 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06297__A2_N _01190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12263_ genblk2\[1\].wave_shpr.div.b1\[1\] _01263_ _05802_ vssd1 vssd1 vccd1 vccd1
+ _05992_ sky130_fd_sc_hd__mux2_1
XANTENNA__09873__S _04214_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11214_ _05247_ vssd1 vssd1 vccd1 vccd1 _05248_ sky130_fd_sc_hd__clkbuf_4
X_12194_ genblk2\[11\].wave_shpr.div.acc\[10\] genblk2\[11\].wave_shpr.div.b1\[10\]
+ vssd1 vssd1 vccd1 vccd1 _05932_ sky130_fd_sc_hd__or2b_1
XANTENNA__09780__A1 _01858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08583__A2 _02308_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102_893 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11145_ genblk2\[7\].wave_shpr.div.b1\[12\] genblk2\[7\].wave_shpr.div.acc\[12\]
+ vssd1 vssd1 vccd1 vccd1 _05205_ sky130_fd_sc_hd__and2b_1
XFILLER_0_37_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11076_ genblk2\[6\].wave_shpr.div.acc\[21\] genblk2\[6\].wave_shpr.div.acc\[20\]
+ _05019_ net1350 vssd1 vssd1 vccd1 vccd1 _05146_ sky130_fd_sc_hd__or4_1
XANTENNA_clkbuf_leaf_94_clk_A clknet_4_11_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10027_ genblk2\[3\].wave_shpr.div.fin_quo\[0\] _04420_ _04422_ vssd1 vssd1 vccd1
+ vccd1 _04423_ sky130_fd_sc_hd__mux2_1
XANTENNA__11209__A _02171_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_144_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06897__A2 _01367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_28_clk clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_28_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_86_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_53_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11978_ genblk2\[10\].wave_shpr.div.fin_quo\[6\] net1324 _00003_ vssd1 vssd1 vccd1
+ vccd1 _05794_ sky130_fd_sc_hd__mux2_1
XANTENNA__07422__A _02147_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13717_ clknet_leaf_36_clk _01028_ net105 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.b1\[13\]
+ sky130_fd_sc_hd__dfrtp_1
X_10929_ net758 vssd1 vssd1 vccd1 vccd1 _05049_ sky130_fd_sc_hd__inv_2
XANTENNA__11642__A2 _05448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13648_ clknet_leaf_38_clk net224 net126 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.quo\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_6_605 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_39_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_32_clk_A clknet_4_5_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_6_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_13579_ clknet_leaf_76_clk _00894_ net207 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.acc\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_137 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_42_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_81_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06120_ net365 _01088_ net395 vssd1 vssd1 vccd1 vccd1 _01093_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_81_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_2_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__13329__RESET_B net91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_41_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_42_769 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_124_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_152_793 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_484 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_112_635 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_47_clk_A clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_151_281 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__08023__A1 _01229_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09220__B1 _03840_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09810_ genblk2\[2\].wave_shpr.div.quo\[9\] _04253_ _04251_ net300 _04254_ vssd1
+ vssd1 vccd1 vccd1 _00300_ sky130_fd_sc_hd__a221o_1
XANTENNA__08574__A2 net33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_10_699 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__09084__A _03735_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09741_ genblk2\[2\].wave_shpr.div.fin_quo\[3\] net1329 _00009_ vssd1 vssd1 vccd1
+ vccd1 _04218_ sky130_fd_sc_hd__mux2_1
X_06953_ _01760_ _01789_ _01790_ vssd1 vssd1 vccd1 vccd1 _01791_ sky130_fd_sc_hd__and3b_1
XFILLER_0_94_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_105_clk_A clknet_4_10_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10669__B1 _04855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_118_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09672_ genblk2\[1\].wave_shpr.div.i\[3\] _02158_ _04151_ vssd1 vssd1 vccd1 vccd1
+ _04154_ sky130_fd_sc_hd__and3_1
X_06884_ _01241_ _01660_ vssd1 vssd1 vccd1 vccd1 _01738_ sky130_fd_sc_hd__nor2_2
X_08623_ _03328_ _03329_ vssd1 vssd1 vccd1 vccd1 _03330_ sky130_fd_sc_hd__nor2_1
Xclkbuf_leaf_19_clk clknet_4_6_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_19_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_11_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08554_ _03259_ _03260_ vssd1 vssd1 vccd1 vccd1 _03261_ sky130_fd_sc_hd__nor2_1
X_07505_ _02215_ net760 _02225_ vssd1 vssd1 vccd1 vccd1 _02226_ sky130_fd_sc_hd__o21a_1
XANTENNA__11094__B1 _05057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08485_ genblk2\[3\].wave_shpr.div.fin_quo\[3\] _03191_ vssd1 vssd1 vccd1 vccd1 _03192_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_677 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_147_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_58_880 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_76_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07436_ genblk2\[4\].wave_shpr.div.i\[2\] genblk2\[4\].wave_shpr.div.i\[3\] genblk2\[4\].wave_shpr.div.i\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02174_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_91_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07051__B _01183_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_716 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_107_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_91_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_73_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07367_ _02122_ vssd1 vssd1 vccd1 vccd1 genblk1\[11\].osc.clkdiv_C.next_cnt\[8\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_60_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09106_ genblk2\[0\].wave_shpr.div.acc\[9\] genblk2\[0\].wave_shpr.div.b1\[9\] vssd1
+ vssd1 vccd1 vccd1 _03754_ sky130_fd_sc_hd__or2b_1
XANTENNA__09259__A _03853_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06318_ genblk1\[0\].osc.clkdiv_C.cnt\[3\] _01274_ vssd1 vssd1 vccd1 vccd1 _01277_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__07065__A2 _01211_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07298_ net695 _02061_ vssd1 vssd1 vccd1 vccd1 genblk1\[10\].osc.clkdiv_C.next_cnt\[17\]
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_115_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_60_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09037_ _03704_ net861 _03705_ vssd1 vssd1 vccd1 vccd1 _00076_ sky130_fd_sc_hd__a21bo_1
X_06249_ _01182_ vssd1 vssd1 vccd1 vccd1 _01211_ sky130_fd_sc_hd__buf_4
XFILLER_0_32_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_102_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_13_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xhold350 _00648_ vssd1 vssd1 vccd1 vccd1 net568 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_102_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold361 _00148_ vssd1 vssd1 vccd1 vccd1 net579 sky130_fd_sc_hd__dlygate4sd3_1
Xhold372 genblk2\[10\].wave_shpr.div.acc\[18\] vssd1 vssd1 vccd1 vccd1 net590 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__09762__A1 _04230_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11728__S _00023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold383 _00128_ vssd1 vssd1 vccd1 vccd1 net601 sky130_fd_sc_hd__dlygate4sd3_1
Xhold394 sig_norm.acc\[7\] vssd1 vssd1 vccd1 vccd1 net612 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10632__S _04834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07773__B1 _01190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09939_ net968 _04315_ _04322_ _04344_ vssd1 vssd1 vccd1 vccd1 _00339_ sky130_fd_sc_hd__a22o_1
Xclkbuf_4_13_0_clk clknet_0_clk vssd1 vssd1 vccd1 vccd1 clknet_4_13_0_clk sky130_fd_sc_hd__clkbuf_8
X_12950_ clknet_leaf_125_clk _00279_ net71 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.b1\[6\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1050 genblk2\[9\].wave_shpr.div.b1\[4\] vssd1 vssd1 vccd1 vccd1 net1268 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__12634__RESET_B net74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold1061 genblk2\[5\].wave_shpr.div.b1\[12\] vssd1 vssd1 vccd1 vccd1 net1279 sky130_fd_sc_hd__dlygate4sd3_1
X_11901_ genblk2\[0\].wave_shpr.div.i\[1\] genblk2\[0\].wave_shpr.div.i\[0\] genblk2\[0\].wave_shpr.div.i\[2\]
+ vssd1 vssd1 vccd1 vccd1 _05726_ sky130_fd_sc_hd__and3_1
Xhold1072 genblk2\[3\].wave_shpr.div.b1\[3\] vssd1 vssd1 vccd1 vccd1 net1290 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12881_ clknet_leaf_91_clk net415 net146 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold1083 genblk2\[7\].wave_shpr.div.b1\[12\] vssd1 vssd1 vccd1 vccd1 net1301 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1094 genblk2\[1\].wave_shpr.div.quo\[1\] vssd1 vssd1 vccd1 vccd1 net1312 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_2522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11832_ _05589_ _05675_ vssd1 vssd1 vccd1 vccd1 _05676_ sky130_fd_sc_hd__xnor2_1
XTAP_2544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11085__B1 _05055_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11763_ net243 _05628_ _05629_ net481 _05630_ vssd1 vssd1 vccd1 vccd1 _00877_ sky130_fd_sc_hd__a221o_1
XTAP_2599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_23_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__08057__B _01223_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1876 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_10714_ _04785_ _04780_ vssd1 vssd1 vccd1 vccd1 _04887_ sky130_fd_sc_hd__or2b_1
X_13502_ clknet_leaf_87_clk _00819_ net180 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.quo\[24\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1887 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_138_565 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_1898 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11694_ genblk2\[9\].wave_shpr.div.b1\[7\] genblk2\[9\].wave_shpr.div.acc\[7\] vssd1
+ vssd1 vccd1 vccd1 _05586_ sky130_fd_sc_hd__and2b_1
X_13433_ clknet_leaf_82_clk _00752_ net201 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.acc\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__07896__B net136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10645_ genblk2\[6\].wave_shpr.div.b1\[15\] _01365_ _04848_ vssd1 vssd1 vccd1 vccd1
+ _04850_ sky130_fd_sc_hd__mux2_1
XFILLER_0_130_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_13364_ clknet_leaf_12_clk _00683_ net53 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.i\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_10576_ genblk2\[5\].wave_shpr.div.b1\[12\] genblk2\[5\].wave_shpr.div.acc\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04804_ sky130_fd_sc_hd__and2b_1
XFILLER_0_24_769 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_23_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12315_ _03941_ vssd1 vssd1 vccd1 vccd1 _06015_ sky130_fd_sc_hd__clkbuf_4
X_13295_ clknet_leaf_53_clk _00616_ net112 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.b1\[7\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_20_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__12337__B1 _03941_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12246_ _05983_ vssd1 vssd1 vccd1 vccd1 _01007_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_139_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__10899__B1 _04233_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12177_ _05816_ _05917_ _05918_ _05818_ net1090 vssd1 vssd1 vccd1 vccd1 _01003_ sky130_fd_sc_hd__a32o_1
X_11128_ genblk2\[7\].wave_shpr.div.b1\[3\] genblk2\[7\].wave_shpr.div.acc\[3\] vssd1
+ vssd1 vccd1 vccd1 _05188_ sky130_fd_sc_hd__and2b_1
XFILLER_0_3_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_155_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11059_ genblk2\[6\].wave_shpr.div.acc\[16\] _05133_ _05105_ vssd1 vssd1 vccd1 vccd1
+ _05134_ sky130_fd_sc_hd__mux2_1
XANTENNA__07136__B _01361_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_64_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_78_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xwire28 net1356 vssd1 vssd1 vccd1 vccd1 net28 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_99_780 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06975__B _01355_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_154_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_59_633 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_58_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__09778__S _04238_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_58_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08270_ _02366_ _02976_ vssd1 vssd1 vccd1 vccd1 _02977_ sky130_fd_sc_hd__nor2_1
XFILLER_0_73_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_80_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_129_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_104_63 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07221_ genblk1\[10\].osc.clkdiv_C.cnt\[8\] vssd1 vssd1 vccd1 vccd1 _02003_ sky130_fd_sc_hd__inv_2
XFILLER_0_104_85 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_61_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_82_680 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_89_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_07152_ _01919_ _01922_ _01927_ _01951_ vssd1 vssd1 vccd1 vccd1 _01952_ sky130_fd_sc_hd__and4_2
XANTENNA__09079__A _03708_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_758 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_131_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__06255__B1 _01215_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_70_875 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_07083_ genblk1\[8\].osc.clkdiv_C.cnt\[4\] _01892_ genblk1\[8\].osc.clkdiv_C.cnt\[5\]
+ vssd1 vssd1 vccd1 vccd1 _01896_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_112_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_8_clk clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 clknet_leaf_8_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__08547__A2 _02527_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_649 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xfanout104 net107 vssd1 vssd1 vccd1 vccd1 net104 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xfanout115 net118 vssd1 vssd1 vccd1 vccd1 net115 sky130_fd_sc_hd__clkbuf_4
Xfanout126 net127 vssd1 vssd1 vccd1 vccd1 net126 sky130_fd_sc_hd__buf_2
Xfanout137 net145 vssd1 vssd1 vccd1 vccd1 net137 sky130_fd_sc_hd__clkbuf_4
Xfanout148 net150 vssd1 vssd1 vccd1 vccd1 net148 sky130_fd_sc_hd__clkbuf_4
X_07985_ _02682_ _02690_ _02691_ vssd1 vssd1 vccd1 vccd1 _02692_ sky130_fd_sc_hd__o21ai_1
Xfanout159 net162 vssd1 vssd1 vccd1 vccd1 net159 sky130_fd_sc_hd__clkbuf_4
XANTENNA__06231__A _01181_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09724_ _04158_ _04202_ _04203_ vssd1 vssd1 vccd1 vccd1 _04204_ sky130_fd_sc_hd__a21o_1
XFILLER_0_38_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06936_ genblk1\[6\].osc.clkdiv_C.cnt\[11\] _01777_ vssd1 vssd1 vccd1 vccd1 _01779_
+ sky130_fd_sc_hd__and2_1
XANTENNA__07046__B _01328_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09655_ _04045_ _04141_ _04142_ _04048_ net448 vssd1 vssd1 vccd1 vccd1 _00257_ sky130_fd_sc_hd__a32o_1
X_06867_ genblk1\[5\].osc.clkdiv_C.cnt\[16\] _01721_ vssd1 vssd1 vccd1 vccd1 _01723_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_78_920 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_97_739 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06885__B _01209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08606_ _02891_ _03311_ _03312_ _02893_ vssd1 vssd1 vccd1 vccd1 _03313_ sky130_fd_sc_hd__a31o_1
XFILLER_0_145_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__09261__B genblk1\[0\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_1106 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09586_ _03981_ _04090_ vssd1 vssd1 vccd1 vccd1 _04091_ sky130_fd_sc_hd__xnor2_1
XTAP_1117 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_06798_ genblk1\[5\].osc.clkdiv_C.cnt\[6\] vssd1 vssd1 vccd1 vccd1 _01670_ sky130_fd_sc_hd__inv_2
XFILLER_0_77_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1128 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08537_ _03240_ _03242_ vssd1 vssd1 vccd1 vccd1 _03244_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_1139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__10814__B1 _04858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08468_ _03154_ _03173_ _03051_ _03174_ vssd1 vssd1 vccd1 vccd1 _03175_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_65_647 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07419_ genblk2\[2\].wave_shpr.div.i\[2\] genblk2\[2\].wave_shpr.div.i\[3\] genblk2\[2\].wave_shpr.div.i\[0\]
+ vssd1 vssd1 vccd1 vccd1 _02161_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_92_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_08399_ _03103_ _03104_ _03105_ vssd1 vssd1 vccd1 vccd1 _03106_ sky130_fd_sc_hd__or3b_1
XFILLER_0_107_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__08605__B _02467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_46_894 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10430_ _04587_ _04582_ vssd1 vssd1 vccd1 vccd1 _04687_ sky130_fd_sc_hd__or2b_1
XFILLER_0_33_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__08235__A1 _02592_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07038__A2 _01855_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_150_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10361_ net834 vssd1 vssd1 vccd1 vccd1 _04649_ sky130_fd_sc_hd__inv_2
XFILLER_0_103_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_103_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06125__B _01095_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_752 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12100_ net929 _05844_ _05850_ _05862_ vssd1 vssd1 vccd1 vccd1 _00982_ sky130_fd_sc_hd__a22o_1
X_13080_ clknet_leaf_125_clk _00407_ net63 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.acc\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10292_ genblk2\[4\].wave_shpr.div.b1\[11\] genblk2\[4\].wave_shpr.div.acc\[11\]
+ vssd1 vssd1 vccd1 vccd1 _04604_ sky130_fd_sc_hd__and2b_1
XFILLER_0_131_785 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12886__RESET_B net98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12031_ _05812_ vssd1 vssd1 vccd1 vccd1 _05818_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__09735__A1 _04214_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold180 genblk2\[10\].wave_shpr.div.quo\[10\] vssd1 vssd1 vccd1 vccd1 net398 sky130_fd_sc_hd__dlygate4sd3_1
Xhold191 genblk2\[1\].wave_shpr.div.b1\[17\] vssd1 vssd1 vccd1 vccd1 net409 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__08943__C1 _01155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06141__A net14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07210__A2 _01224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12933_ clknet_leaf_31_clk _00262_ net102 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.i\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12864_ clknet_leaf_129_clk _00195_ net64 vssd1 vssd1 vccd1 vccd1 genblk2\[2\].wave_shpr.div.b1\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11815_ _05662_ _05581_ vssd1 vssd1 vccd1 vccd1 _05663_ sky130_fd_sc_hd__xnor2_1
XTAP_2374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_841 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12795_ clknet_leaf_92_clk net601 net148 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_625 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_11746_ net649 _05623_ _05624_ net746 vssd1 vssd1 vccd1 vccd1 _00866_ sky130_fd_sc_hd__a22o_1
XFILLER_0_154_811 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_83_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_1695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_11677_ _05567_ _05568_ vssd1 vssd1 vccd1 vccd1 _05569_ sky130_fd_sc_hd__nand2_1
XFILLER_0_83_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_153_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_64_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_153_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_141_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13416_ clknet_leaf_119_clk net535 net141 vssd1 vssd1 vccd1 vccd1 genblk2\[7\].wave_shpr.div.quo\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_10628_ net1211 _01189_ _04834_ vssd1 vssd1 vccd1 vccd1 _04841_ sky130_fd_sc_hd__mux2_1
XFILLER_0_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_24_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_24_566 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_107_793 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_13347_ clknet_leaf_5_clk _00668_ net45 vssd1 vssd1 vccd1 vccd1 genblk2\[6\].wave_shpr.div.acc\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__11230__B1 _05248_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10559_ genblk2\[5\].wave_shpr.div.b1\[3\] genblk2\[5\].wave_shpr.div.acc\[3\] vssd1
+ vssd1 vccd1 vccd1 _04787_ sky130_fd_sc_hd__and2b_1
XFILLER_0_24_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13278_ clknet_leaf_11_clk _00599_ net56 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.i\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_121_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12229_ genblk2\[11\].wave_shpr.div.b1\[13\] genblk2\[11\].wave_shpr.div.acc\[13\]
+ vssd1 vssd1 vccd1 vccd1 _05967_ sky130_fd_sc_hd__and2b_1
XFILLER_0_20_783 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07147__A _01241_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07770_ genblk1\[0\].osc.clkdiv_C.cnt\[12\] _01240_ _02476_ vssd1 vssd1 vccd1 vccd1
+ _02477_ sky130_fd_sc_hd__a21bo_1
X_06721_ _01608_ vssd1 vssd1 vccd1 vccd1 genblk1\[4\].osc.clkdiv_C.next_cnt\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_78_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09440_ genblk2\[1\].wave_shpr.div.b1\[17\] genblk2\[1\].wave_shpr.div.acc\[17\]
+ vssd1 vssd1 vccd1 vccd1 _04004_ sky130_fd_sc_hd__and2b_1
X_06652_ genblk1\[3\].osc.clkdiv_C.cnt\[13\] genblk1\[3\].osc.clkdiv_C.cnt\[12\] _01543_
+ vssd1 vssd1 vccd1 vccd1 _01547_ sky130_fd_sc_hd__and3_1
XFILLER_0_149_638 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_115_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09371_ _02170_ genblk2\[11\].wave_shpr.div.busy _02211_ vssd1 vssd1 vccd1 vccd1
+ _03940_ sky130_fd_sc_hd__and3_1
XFILLER_0_59_463 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06583_ genblk1\[3\].osc.clkdiv_C.cnt\[5\] _01250_ vssd1 vssd1 vccd1 vccd1 _01491_
+ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_636 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08322_ _02419_ _03018_ _03022_ _03024_ _03028_ vssd1 vssd1 vccd1 vccd1 _03029_ sky130_fd_sc_hd__a32o_1
XANTENNA__09662__A0 _04046_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_7_711 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_74_444 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_7_722 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_145_833 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_46_157 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_62_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08253_ _02734_ _02959_ genblk2\[6\].wave_shpr.div.fin_quo\[5\] vssd1 vssd1 vccd1
+ vccd1 _02960_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_117_535 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_6_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_145_877 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_07204_ genblk1\[9\].osc.clkdiv_C.cnt\[16\] _01985_ vssd1 vssd1 vccd1 vccd1 _01988_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_27_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08184_ _02225_ _02885_ vssd1 vssd1 vccd1 vccd1 _02891_ sky130_fd_sc_hd__nand2_1
XFILLER_0_15_544 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__11221__B1 _05250_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07135_ genblk1\[9\].osc.clkdiv_C.cnt\[4\] _01311_ _01925_ genblk1\[9\].osc.clkdiv_C.cnt\[5\]
+ _01934_ vssd1 vssd1 vccd1 vccd1 _01935_ sky130_fd_sc_hd__o221a_1
XFILLER_0_42_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_70_672 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_43_897 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07066_ genblk1\[8\].osc.clkdiv_C.cnt\[16\] _01578_ _01870_ genblk1\[8\].osc.clkdiv_C.cnt\[11\]
+ _01883_ vssd1 vssd1 vccd1 vccd1 _01884_ sky130_fd_sc_hd__o221a_1
XFILLER_0_113_785 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_11_783 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_100_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07968_ _02672_ _02674_ vssd1 vssd1 vccd1 vccd1 _02675_ sky130_fd_sc_hd__or2_1
XANTENNA__06896__A _01342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09707_ genblk2\[2\].wave_shpr.div.b1\[7\] genblk2\[2\].wave_shpr.div.acc\[7\] vssd1
+ vssd1 vccd1 vccd1 _04187_ sky130_fd_sc_hd__and2b_1
X_06919_ genblk1\[6\].osc.clkdiv_C.cnt\[5\] genblk1\[6\].osc.clkdiv_C.cnt\[4\] _01765_
+ vssd1 vssd1 vccd1 vccd1 _01768_ sky130_fd_sc_hd__and3_1
X_07899_ _01181_ _01852_ _01245_ genblk1\[8\].osc.clkdiv_C.cnt\[13\] vssd1 vssd1 vccd1
+ vccd1 _02606_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__08153__B1 _01494_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09638_ _04005_ _04129_ genblk2\[1\].wave_shpr.div.acc\[18\] vssd1 vssd1 vccd1 vccd1
+ _04131_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_97_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09569_ _03973_ _04077_ vssd1 vssd1 vccd1 vccd1 _04078_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_78_794 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_65_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11600_ _05398_ _05363_ vssd1 vssd1 vccd1 vccd1 _05511_ sky130_fd_sc_hd__or2b_1
XFILLER_0_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_65_422 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12580_ clknet_leaf_14_clk genblk1\[2\].osc.clkdiv_C.next_cnt\[1\] net70 vssd1 vssd1
+ vccd1 vccd1 genblk1\[2\].osc.clkdiv_C.cnt\[1\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_136_833 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11531_ genblk2\[8\].wave_shpr.div.quo\[18\] _05454_ _05458_ net263 _05462_ vssd1
+ vssd1 vccd1 vccd1 _00813_ sky130_fd_sc_hd__a221o_1
XFILLER_0_135_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_135_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_53_639 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_34_831 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_505 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11462_ net1294 _01797_ _05237_ vssd1 vssd1 vccd1 vccd1 _05428_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06136__A net1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13201_ clknet_leaf_114_clk _00524_ net132 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.fin_quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__08759__A2 _02467_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10413_ net698 _04651_ _04654_ net665 _04675_ vssd1 vssd1 vccd1 vccd1 _00482_ sky130_fd_sc_hd__a221o_1
XFILLER_0_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_1_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11393_ genblk2\[8\].wave_shpr.div.acc\[6\] genblk2\[8\].wave_shpr.div.b1\[6\] vssd1
+ vssd1 vccd1 vccd1 _05369_ sky130_fd_sc_hd__or2b_1
X_13132_ clknet_leaf_3_clk _00457_ net46 vssd1 vssd1 vccd1 vccd1 genblk2\[5\].wave_shpr.div.b1\[16\]
+ sky130_fd_sc_hd__dfrtp_1
X_10344_ _01678_ vssd1 vssd1 vccd1 vccd1 _04639_ sky130_fd_sc_hd__inv_2
XFILLER_0_60_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__11188__S _05042_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_131_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13063_ clknet_leaf_29_clk _00390_ net95 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.quo\[15\]
+ sky130_fd_sc_hd__dfrtp_1
X_10275_ genblk2\[4\].wave_shpr.div.b1\[2\] genblk2\[4\].wave_shpr.div.acc\[2\] vssd1
+ vssd1 vccd1 vccd1 _04587_ sky130_fd_sc_hd__and2b_1
XANTENNA__07719__B1 _01209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12014_ _02171_ net1278 vssd1 vssd1 vccd1 vccd1 _05811_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xmax_cap4 net1354 vssd1 vssd1 vccd1 vccd1 net1353 sky130_fd_sc_hd__clkbuf_1
XANTENNA__11217__A _05249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12916_ clknet_leaf_35_clk _00247_ net105 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.acc\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_152_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_29_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_75_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_2160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12847_ clknet_leaf_58_clk _00178_ net211 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.i\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_2182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_139_671 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_1470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_12778_ clknet_leaf_41_clk _00111_ net123 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.b1\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_1481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_904 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_84_764 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11729_ _05617_ vssd1 vssd1 vccd1 vccd1 _00856_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_15 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_680 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_71_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_117_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_142_825 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_71_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_126_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_142_869 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold905 genblk2\[2\].wave_shpr.div.i\[3\] vssd1 vssd1 vccd1 vccd1 net1123 sky130_fd_sc_hd__dlygate4sd3_1
Xhold916 PWM.final_in\[0\] vssd1 vssd1 vccd1 vccd1 net1134 sky130_fd_sc_hd__dlygate4sd3_1
Xhold927 genblk1\[3\].osc.clkdiv_C.cnt\[9\] vssd1 vssd1 vccd1 vccd1 net1145 sky130_fd_sc_hd__dlygate4sd3_1
Xhold938 sig_norm.quo\[9\] vssd1 vssd1 vccd1 vccd1 net1156 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold949 genblk1\[2\].osc.clkdiv_C.cnt\[15\] vssd1 vssd1 vccd1 vccd1 net1167 sky130_fd_sc_hd__dlygate4sd3_1
X_08940_ _03632_ vssd1 vssd1 vccd1 vccd1 _00052_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_110_777 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_08871_ sig_norm.b1\[1\] sig_norm.acc\[1\] vssd1 vssd1 vccd1 vccd1 _03577_ sky130_fd_sc_hd__or2b_1
X_07822_ net7 net150 _02312_ vssd1 vssd1 vccd1 vccd1 _02529_ sky130_fd_sc_hd__and3_2
XFILLER_0_19_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07605__A net17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09092__A _01367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07753_ _02458_ _02459_ vssd1 vssd1 vccd1 vccd1 _02460_ sky130_fd_sc_hd__and2_1
XANTENNA__13596__RESET_B net208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06704_ genblk1\[4\].osc.clkdiv_C.cnt\[9\] _01592_ vssd1 vssd1 vccd1 vccd1 _01594_
+ sky130_fd_sc_hd__or2_1
X_07684_ _01179_ _01575_ genblk1\[10\].osc.clkdiv_C.cnt\[15\] vssd1 vssd1 vccd1 vccd1
+ _02391_ sky130_fd_sc_hd__mux2_1
XFILLER_0_126_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08139__C _02365_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09423_ _03963_ _03985_ _03986_ vssd1 vssd1 vccd1 vccd1 _03987_ sky130_fd_sc_hd__a21o_1
XANTENNA__06697__B1 _01304_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06635_ _01523_ _01535_ _01536_ vssd1 vssd1 vccd1 vccd1 genblk1\[3\].osc.clkdiv_C.next_cnt\[6\]
+ sky130_fd_sc_hd__nor3_1
XANTENNA__10966__A _04676_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09354_ genblk2\[0\].wave_shpr.div.acc\[20\] _03927_ vssd1 vssd1 vccd1 vccd1 _03929_
+ sky130_fd_sc_hd__xor2_1
X_06566_ net1207 _01474_ _01477_ vssd1 vssd1 vccd1 vccd1 genblk1\[2\].osc.clkdiv_C.next_cnt\[14\]
+ sky130_fd_sc_hd__o21a_1
XFILLER_0_59_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_47_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08305_ _02977_ _02983_ vssd1 vssd1 vccd1 vccd1 _03012_ sky130_fd_sc_hd__xnor2_1
XANTENNA__11442__A0 genblk2\[8\].wave_shpr.div.fin_quo\[0\] vssd1 vssd1 vccd1 vccd1
+ sky130_fd_sc_hd__diode_2
XFILLER_0_117_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_09285_ net1033 _03870_ _03840_ _03876_ vssd1 vssd1 vccd1 vccd1 _00153_ sky130_fd_sc_hd__a22o_1
XANTENNA__10177__S _04507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_75_797 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07110__A1 genblk1\[8\].osc.clkdiv_C.cnt\[14\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06497_ _01173_ _01191_ _01175_ vssd1 vssd1 vccd1 vccd1 _01423_ sky130_fd_sc_hd__nor3b_4
XFILLER_0_34_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_62_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__10796__A2 _04858_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_62_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_08236_ net9 _02744_ _02365_ vssd1 vssd1 vccd1 vccd1 _02943_ sky130_fd_sc_hd__and3_1
XFILLER_0_145_685 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__07661__A2 _01190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_43_650 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_144_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_31_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_08167_ genblk1\[3\].osc.clkdiv_C.cnt\[9\] _01231_ vssd1 vssd1 vccd1 vccd1 _02874_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_30_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__12478__RESET_B net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__11745__B2 _05613_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07118_ net691 _01917_ vssd1 vssd1 vccd1 vccd1 genblk1\[8\].osc.clkdiv_C.next_cnt\[17\]
+ sky130_fd_sc_hd__xnor2_1
XANTENNA__09267__A _03838_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_31_856 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08098_ _01440_ _01576_ vssd1 vssd1 vccd1 vccd1 _02805_ sky130_fd_sc_hd__nand2_2
XANTENNA__08602__C _02885_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_100_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07049_ genblk1\[8\].osc.clkdiv_C.cnt\[4\] _01866_ _01865_ genblk1\[8\].osc.clkdiv_C.cnt\[9\]
+ vssd1 vssd1 vccd1 vccd1 _01867_ sky130_fd_sc_hd__o22a_1
XFILLER_0_30_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06403__B _01327_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10060_ _04439_ vssd1 vssd1 vccd1 vccd1 _00365_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_100_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__11736__S _00023_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10962_ _05059_ genblk1\[6\].osc.clkdiv_C.cnt\[5\] vssd1 vssd1 vccd1 vccd1 _05066_
+ sky130_fd_sc_hd__and2_1
XANTENNA__07234__B _01359_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13750_ clknet_leaf_75_clk _01061_ net211 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.acc\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__13266__RESET_B net38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12701_ clknet_leaf_89_clk genblk1\[8\].osc.clkdiv_C.next_cnt\[14\] net172 vssd1
+ vssd1 vccd1 vccd1 genblk1\[8\].osc.clkdiv_C.cnt\[14\] sky130_fd_sc_hd__dfrtp_4
X_13681_ clknet_leaf_63_clk _00994_ net125 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.acc\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_10893_ _05030_ vssd1 vssd1 vccd1 vccd1 _00607_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_155_405 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12632_ clknet_leaf_18_clk genblk1\[4\].osc.clkdiv_C.next_cnt\[17\] net112 vssd1
+ vssd1 vccd1 vccd1 genblk1\[4\].osc.clkdiv_C.cnt\[17\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_155_449 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_12563_ clknet_leaf_30_clk genblk1\[1\].osc.clkdiv_C.next_cnt\[2\] net96 vssd1 vssd1
+ vccd1 vccd1 genblk1\[1\].osc.clkdiv_C.cnt\[2\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_31_39 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__07101__A1 genblk1\[8\].osc.clkdiv_C.cnt\[11\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_65_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__11984__A1 _03813_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_135_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_19_691 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_11514_ _04676_ _01879_ vssd1 vssd1 vccd1 vccd1 _05453_ sky130_fd_sc_hd__nor2_1
XFILLER_0_135_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_108_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_12494_ clknet_leaf_106_clk _00056_ net153 vssd1 vssd1 vccd1 vccd1 sig_norm.quo\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_135_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_150_121 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11445_ _05419_ vssd1 vssd1 vccd1 vccd1 _00770_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_124_869 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_40_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_150_165 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_21_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11376_ _05248_ _05352_ _05354_ _05251_ net801 vssd1 vssd1 vccd1 vccd1 _00766_ sky130_fd_sc_hd__a32o_1
XFILLER_0_0_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10327_ net1264 vssd1 vssd1 vccd1 vccd1 _00440_ sky130_fd_sc_hd__clkbuf_1
X_13115_ clknet_leaf_115_clk _00440_ net135 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.fin_quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_131_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07409__B _02153_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13046_ clknet_leaf_112_clk _00373_ net128 vssd1 vssd1 vccd1 vccd1 genblk2\[4\].wave_shpr.div.b1\[16\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_147_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_10258_ genblk2\[4\].wave_shpr.div.acc\[12\] genblk2\[4\].wave_shpr.div.b1\[12\]
+ vssd1 vssd1 vccd1 vccd1 _04570_ sky130_fd_sc_hd__or2b_1
X_10189_ _04402_ _04519_ vssd1 vssd1 vccd1 vccd1 _04520_ sky130_fd_sc_hd__xnor2_1
XANTENNA__09865__B1 _04252_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_72_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__06679__B1 _01242_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_48_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__06983__B _01334_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_06420_ genblk1\[1\].osc.clkdiv_C.cnt\[16\] _01363_ _01341_ vssd1 vssd1 vccd1 vccd1
+ _01364_ sky130_fd_sc_hd__o21a_1
XFILLER_0_9_828 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_146_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_56_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07798__C _01209_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_29_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_45_904 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_57_775 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__07160__A genblk1\[9\].osc.clkdiv_C.cnt\[2\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_06351_ genblk1\[0\].osc.clkdiv_C.cnt\[15\] _01295_ _01297_ vssd1 vssd1 vccd1 vccd1
+ genblk1\[0\].osc.clkdiv_C.next_cnt\[15\] sky130_fd_sc_hd__o21a_1
XFILLER_0_29_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_56_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09093__A1 _01367_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__09093__B2 _01342_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_112_41 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09070_ _03702_ _01996_ vssd1 vssd1 vccd1 vccd1 _03728_ sky130_fd_sc_hd__nand2_4
X_06282_ genblk1\[0\].osc.clkdiv_C.cnt\[16\] _01242_ vssd1 vssd1 vccd1 vccd1 _01244_
+ sky130_fd_sc_hd__nand2_1
XFILLER_0_114_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_112_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_154_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_4_533 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08021_ genblk1\[6\].osc.clkdiv_C.cnt\[15\] _01577_ _02704_ vssd1 vssd1 vccd1 vccd1
+ _02728_ sky130_fd_sc_hd__a21o_1
XFILLER_0_112_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_31_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_13_812 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold702 genblk2\[0\].wave_shpr.div.acc\[13\] vssd1 vssd1 vccd1 vccd1 net920 sky130_fd_sc_hd__dlygate4sd3_1
Xhold713 genblk2\[11\].wave_shpr.div.acc\[21\] vssd1 vssd1 vccd1 vccd1 net931 sky130_fd_sc_hd__dlygate4sd3_1
Xhold724 genblk2\[3\].wave_shpr.div.acc\[12\] vssd1 vssd1 vccd1 vccd1 net942 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_40_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold735 genblk2\[2\].wave_shpr.div.acc\[13\] vssd1 vssd1 vccd1 vccd1 net953 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__06504__A _01224_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold746 genblk2\[0\].wave_shpr.div.acc\[7\] vssd1 vssd1 vccd1 vccd1 net964 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_13_889 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xhold757 genblk2\[2\].wave_shpr.div.acc\[4\] vssd1 vssd1 vccd1 vccd1 net975 sky130_fd_sc_hd__dlygate4sd3_1
Xhold768 genblk2\[6\].wave_shpr.div.acc\[4\] vssd1 vssd1 vccd1 vccd1 net986 sky130_fd_sc_hd__dlygate4sd3_1
X_09972_ genblk2\[3\].wave_shpr.div.acc\[10\] genblk2\[3\].wave_shpr.div.b1\[10\]
+ vssd1 vssd1 vccd1 vccd1 _04368_ sky130_fd_sc_hd__or2b_1
XANTENNA__10026__A _04421_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_0_750 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xhold779 genblk2\[11\].wave_shpr.div.acc\[7\] vssd1 vssd1 vccd1 vccd1 net997 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10950__A2 _05057_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08923_ _03589_ _03602_ _03620_ vssd1 vssd1 vccd1 vccd1 _03621_ sky130_fd_sc_hd__o21ai_1
XANTENNA__09815__A _04247_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_41_3 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_08854_ _03500_ _03503_ _03501_ _03502_ vssd1 vssd1 vccd1 vccd1 _03561_ sky130_fd_sc_hd__o211ai_1
XANTENNA__06906__A1 _01675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10702__A2 _02183_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07805_ genblk2\[0\].wave_shpr.div.fin_quo\[3\] _02511_ vssd1 vssd1 vccd1 vccd1 _02512_
+ sky130_fd_sc_hd__or2_1
X_08785_ genblk2\[2\].wave_shpr.div.fin_quo\[0\] _03113_ genblk2\[2\].wave_shpr.div.fin_quo\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03492_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_137_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_07736_ _02441_ _02437_ _02439_ _02442_ vssd1 vssd1 vccd1 vccd1 _02443_ sky130_fd_sc_hd__o22a_1
XANTENNA__09856__B1 _04253_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08123__A3 _01249_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07667_ _01308_ _01187_ vssd1 vssd1 vccd1 vccd1 _02374_ sky130_fd_sc_hd__nor2_4
XFILLER_0_79_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_138_917 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__06893__B _01577_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_153_81 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_1_93 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_06618_ genblk1\[3\].osc.clkdiv_C.cnt\[1\] genblk1\[3\].osc.clkdiv_C.cnt\[0\] vssd1
+ vssd1 vccd1 vccd1 _01525_ sky130_fd_sc_hd__nand2_1
X_09406_ genblk2\[1\].wave_shpr.div.acc\[1\] genblk2\[1\].wave_shpr.div.b1\[1\] vssd1
+ vssd1 vccd1 vccd1 _03970_ sky130_fd_sc_hd__xnor2_1
X_07598_ genblk2\[9\].wave_shpr.div.fin_quo\[6\] _02304_ vssd1 vssd1 vccd1 vccd1 _02305_
+ sky130_fd_sc_hd__xor2_1
XFILLER_0_109_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_75_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_153_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_09337_ net1050 _03903_ _03910_ _03916_ vssd1 vssd1 vccd1 vccd1 _00165_ sky130_fd_sc_hd__a22o_1
X_06549_ genblk1\[2\].osc.clkdiv_C.cnt\[9\] _01464_ vssd1 vssd1 vccd1 vccd1 _01466_
+ sky130_fd_sc_hd__and2_1
XANTENNA__11966__A1 _05787_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_90_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_133_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_09268_ _02171_ genblk1\[0\].osc.clkdiv_C.cnt\[17\] vssd1 vssd1 vccd1 vccd1 _03864_
+ sky130_fd_sc_hd__or2_1
XANTENNA__07634__A2 _01190_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08219_ _02602_ _02924_ vssd1 vssd1 vccd1 vccd1 _02926_ sky130_fd_sc_hd__xor2_1
XFILLER_0_105_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09199_ net1292 _03827_ _03822_ vssd1 vssd1 vccd1 vccd1 _03828_ sky130_fd_sc_hd__mux2_1
XANTENNA__10635__S _04834_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_15_182 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11230_ genblk2\[7\].wave_shpr.div.quo\[10\] _05251_ _05248_ net302 _05253_ vssd1
+ vssd1 vccd1 vccd1 _00721_ sky130_fd_sc_hd__a221o_1
XFILLER_0_120_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11161_ _05219_ _05220_ vssd1 vssd1 vccd1 vccd1 _05221_ sky130_fd_sc_hd__or2_1
XFILLER_0_113_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_101_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__06133__B net9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10941__A2 _05052_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10112_ _04465_ genblk1\[3\].osc.clkdiv_C.cnt\[6\] vssd1 vssd1 vccd1 vccd1 _04467_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_101_574 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11092_ genblk2\[6\].wave_shpr.div.i\[1\] genblk2\[6\].wave_shpr.div.i\[0\] vssd1
+ vssd1 vccd1 vccd1 _05156_ sky130_fd_sc_hd__or2_1
X_10043_ _03732_ net1071 _03733_ vssd1 vssd1 vccd1 vccd1 _00357_ sky130_fd_sc_hd__o21a_1
Xhold40 _00228_ vssd1 vssd1 vccd1 vccd1 net258 sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 genblk2\[0\].wave_shpr.div.quo\[6\] vssd1 vssd1 vccd1 vccd1 net269 sky130_fd_sc_hd__buf_1
Xhold62 genblk2\[6\].wave_shpr.div.i\[4\] vssd1 vssd1 vccd1 vccd1 net280 sky130_fd_sc_hd__dlygate4sd3_1
Xhold73 _00875_ vssd1 vssd1 vccd1 vccd1 net291 sky130_fd_sc_hd__dlygate4sd3_1
Xhold84 genblk2\[7\].wave_shpr.div.quo\[9\] vssd1 vssd1 vccd1 vccd1 net302 sky130_fd_sc_hd__dlygate4sd3_1
Xhold95 genblk2\[6\].wave_shpr.div.quo\[19\] vssd1 vssd1 vccd1 vccd1 net313 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_98_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11994_ _03707_ vssd1 vssd1 vccd1 vccd1 _05802_ sky130_fd_sc_hd__clkbuf_8
X_13733_ clknet_leaf_45_clk net468 net121 vssd1 vssd1 vccd1 vccd1 genblk2\[11\].wave_shpr.div.quo\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10945_ net241 _05052_ _05056_ net742 vssd1 vssd1 vccd1 vccd1 _00633_ sky130_fd_sc_hd__a22o_1
XFILLER_0_85_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_98_697 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_42_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_13664_ clknet_leaf_43_clk _00977_ net124 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.acc\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_155_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_10876_ genblk2\[6\].wave_shpr.div.acc\[22\] genblk2\[6\].wave_shpr.div.acc\[21\]
+ genblk2\[6\].wave_shpr.div.acc\[20\] _05019_ vssd1 vssd1 vccd1 vccd1 _05020_ sky130_fd_sc_hd__or4_1
XFILLER_0_54_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_128_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_12615_ clknet_leaf_121_clk genblk1\[4\].osc.clkdiv_C.next_cnt\[0\] net81 vssd1 vssd1
+ vccd1 vccd1 genblk1\[4\].osc.clkdiv_C.cnt\[0\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_94_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_66_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_155_257 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_26_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_13595_ clknet_leaf_72_clk _00910_ net216 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.acc\[19\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_26_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__07625__A2 _01208_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12546_ clknet_leaf_61_clk genblk1\[0\].osc.clkdiv_C.next_cnt\[3\] net188 vssd1 vssd1
+ vccd1 vccd1 genblk1\[0\].osc.clkdiv_C.cnt\[3\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_108_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12477_ clknet_leaf_107_clk _00039_ net152 vssd1 vssd1 vccd1 vccd1 sig_norm.acc\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__12326__A _03689_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_4 _01507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_22_642 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11428_ genblk2\[8\].wave_shpr.div.b1\[15\] genblk2\[8\].wave_shpr.div.acc\[15\]
+ vssd1 vssd1 vccd1 vccd1 _05404_ sky130_fd_sc_hd__and2b_1
XFILLER_0_105_880 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_22_664 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_6_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_104_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_11359_ genblk2\[7\].wave_shpr.div.acc\[23\] _05219_ vssd1 vssd1 vccd1 vccd1 _05343_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_67_35 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_13029_ clknet_leaf_113_clk _00356_ net131 vssd1 vssd1 vccd1 vccd1 genblk2\[3\].wave_shpr.div.fin_quo\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__12061__A _02155_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_83_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_6_clk_A clknet_4_1_0_clk vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08570_ genblk2\[9\].wave_shpr.div.fin_quo\[0\] _02303_ genblk2\[9\].wave_shpr.div.fin_quo\[1\]
+ vssd1 vssd1 vccd1 vccd1 _03277_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_88_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07521_ _02228_ PWM.final_sample_in\[6\] _02231_ _02240_ vssd1 vssd1 vccd1 vccd1
+ _02241_ sky130_fd_sc_hd__o22a_1
XFILLER_0_16_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_107_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_88_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_9_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_07452_ genblk2\[6\].wave_shpr.div.i\[1\] _02185_ genblk2\[6\].wave_shpr.div.i\[4\]
+ vssd1 vssd1 vccd1 vccd1 _02186_ sky130_fd_sc_hd__or3b_1
XANTENNA__12000__S _05802_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_76_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_45_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06403_ genblk1\[1\].osc.clkdiv_C.cnt\[14\] _01327_ vssd1 vssd1 vccd1 vccd1 _01347_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_119_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_135_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_9_658 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_123_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_07383_ _02134_ vssd1 vssd1 vccd1 vccd1 genblk1\[11\].osc.clkdiv_C.next_cnt\[12\]
+ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_57_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_09122_ _03760_ _03768_ _03769_ vssd1 vssd1 vccd1 vccd1 _03770_ sky130_fd_sc_hd__a21o_1
XFILLER_0_72_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06334_ genblk1\[0\].osc.clkdiv_C.cnt\[9\] _01284_ vssd1 vssd1 vccd1 vccd1 _01287_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_72_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_09053_ _03716_ vssd1 vssd1 vccd1 vccd1 _03717_ sky130_fd_sc_hd__buf_8
X_06265_ _01224_ _01226_ vssd1 vssd1 vccd1 vccd1 _01227_ sky130_fd_sc_hd__nor2_8
XFILLER_0_89_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA_fanout212_A net213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_5_875 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_60_748 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_08004_ genblk1\[6\].osc.clkdiv_C.cnt\[11\] _01519_ _02708_ _02710_ vssd1 vssd1 vccd1
+ vccd1 _02711_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_5_897 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold510 genblk2\[0\].wave_shpr.div.quo\[3\] vssd1 vssd1 vccd1 vccd1 net728 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_103_839 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_06196_ _01161_ _01162_ vssd1 vssd1 vccd1 vccd1 PWM.next_counter\[3\] sky130_fd_sc_hd__nor2_1
XFILLER_0_13_653 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_4_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_12_141 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
Xhold521 genblk2\[6\].wave_shpr.div.i\[2\] vssd1 vssd1 vccd1 vccd1 net739 sky130_fd_sc_hd__dlygate4sd3_1
Xhold532 _00464_ vssd1 vssd1 vccd1 vccd1 net750 sky130_fd_sc_hd__dlygate4sd3_1
Xhold543 genblk2\[2\].wave_shpr.div.b1\[17\] vssd1 vssd1 vccd1 vccd1 net761 sky130_fd_sc_hd__dlygate4sd3_1
Xhold554 genblk2\[5\].wave_shpr.div.acc\[9\] vssd1 vssd1 vccd1 vccd1 net772 sky130_fd_sc_hd__dlygate4sd3_1
Xhold565 genblk2\[5\].wave_shpr.div.i\[3\] vssd1 vssd1 vccd1 vccd1 net783 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__10384__B1 _04655_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xhold576 genblk2\[3\].wave_shpr.div.quo\[0\] vssd1 vssd1 vccd1 vccd1 net794 sky130_fd_sc_hd__dlymetal6s2s_1
Xhold587 genblk2\[7\].wave_shpr.div.acc\[14\] vssd1 vssd1 vccd1 vccd1 net805 sky130_fd_sc_hd__dlygate4sd3_1
Xhold598 genblk2\[11\].wave_shpr.div.acc\[10\] vssd1 vssd1 vccd1 vccd1 net816 sky130_fd_sc_hd__dlygate4sd3_1
X_09955_ _04251_ _04353_ _04354_ _04253_ net1110 vssd1 vssd1 vccd1 vccd1 _00345_ sky130_fd_sc_hd__a32o_1
XANTENNA__06888__B _01675_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__10190__S _04507_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08906_ sig_norm.acc\[3\] _03596_ _03608_ vssd1 vssd1 vccd1 vccd1 _03609_ sky130_fd_sc_hd__o21a_1
XTAP_870 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_09886_ genblk2\[2\].wave_shpr.div.acc\[8\] _04304_ _04301_ vssd1 vssd1 vccd1 vccd1
+ _04305_ sky130_fd_sc_hd__mux2_1
XTAP_881 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_892 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__08349__A_N _02789_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_08837_ _02574_ _03543_ vssd1 vssd1 vccd1 vccd1 _03544_ sky130_fd_sc_hd__xnor2_2
XANTENNA__11884__B1 _03694_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_2704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08768_ _03455_ _03456_ _03459_ vssd1 vssd1 vccd1 vccd1 _03475_ sky130_fd_sc_hd__o21ba_1
XTAP_2726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_2748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__11636__B1 _05448_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_07719_ genblk1\[1\].osc.clkdiv_C.cnt\[15\] _01309_ _01209_ genblk1\[1\].osc.clkdiv_C.cnt\[14\]
+ vssd1 vssd1 vccd1 vccd1 _02426_ sky130_fd_sc_hd__o22ai_2
XTAP_2759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_08699_ _03401_ _03404_ _03405_ vssd1 vssd1 vccd1 vccd1 _03406_ sky130_fd_sc_hd__nand3b_2
X_10730_ _04792_ _04774_ vssd1 vssd1 vccd1 vccd1 _04899_ sky130_fd_sc_hd__or2b_1
XFILLER_0_137_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_36_701 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_83_829 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_10661_ net253 _04853_ _04857_ net729 vssd1 vssd1 vccd1 vccd1 _00548_ sky130_fd_sc_hd__a22o_1
XFILLER_0_76_881 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_126_909 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XANTENNA__12493__RESET_B net152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__06128__B net15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_12400_ _03942_ vssd1 vssd1 vccd1 vccd1 _06072_ sky130_fd_sc_hd__clkbuf_4
X_13380_ clknet_leaf_80_clk _00699_ net200 vssd1 vssd1 vccd1 vccd1 genblk2\[8\].wave_shpr.div.b1\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_10592_ _04818_ _04819_ vssd1 vssd1 vccd1 vccd1 _04820_ sky130_fd_sc_hd__or2_1
XFILLER_0_51_704 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_152_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_12331_ net483 _06014_ _06015_ net509 _06023_ vssd1 vssd1 vccd1 vccd1 _01052_ sky130_fd_sc_hd__a221o_1
XFILLER_0_51_737 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_51_748 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_90_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_121_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12262_ _05991_ vssd1 vssd1 vccd1 vccd1 _01015_ sky130_fd_sc_hd__clkbuf_1
X_11213_ _02170_ genblk2\[7\].wave_shpr.div.busy _02191_ vssd1 vssd1 vccd1 vccd1 _05247_
+ sky130_fd_sc_hd__and3_1
X_12193_ genblk2\[11\].wave_shpr.div.acc\[11\] genblk2\[11\].wave_shpr.div.b1\[11\]
+ vssd1 vssd1 vccd1 vccd1 _05931_ sky130_fd_sc_hd__or2b_1
XFILLER_0_102_861 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_11144_ _05170_ _05202_ _05203_ vssd1 vssd1 vccd1 vccd1 _05204_ sky130_fd_sc_hd__a21o_1
XFILLER_0_101_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_128_29 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_37_27 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
X_11075_ genblk2\[6\].wave_shpr.div.acc\[20\] _05019_ net1350 vssd1 vssd1 vccd1 vccd1
+ _05145_ sky130_fd_sc_hd__or3_1
XANTENNA__10127__B1 _04455_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_10026_ _04421_ vssd1 vssd1 vccd1 vccd1 _04422_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_53_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__08099__A2 _01498_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_11977_ _05793_ vssd1 vssd1 vccd1 vccd1 _00928_ sky130_fd_sc_hd__clkbuf_1
X_13716_ clknet_leaf_36_clk _01027_ net103 vssd1 vssd1 vccd1 vccd1 genblk2\[1\].wave_shpr.div.b1\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_129_725 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_10928_ _05048_ vssd1 vssd1 vccd1 vccd1 _00624_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_129_736 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_0_86_689 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_0_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_39_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__09048__A1 _03712_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_13647_ clknet_leaf_47_clk _00960_ net114 vssd1 vssd1 vccd1 vccd1 genblk2\[10\].wave_shpr.div.quo\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_10859_ _04973_ _05001_ _05002_ vssd1 vssd1 vccd1 vccd1 _05003_ sky130_fd_sc_hd__a21o_1
XFILLER_0_128_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_26_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_6_617 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_82_851 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__07059__B1 _01869_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_27_767 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_13578_ clknet_leaf_78_clk _00893_ net207 vssd1 vssd1 vccd1 vccd1 genblk2\[9\].wave_shpr.div.acc\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_109_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_14_406 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_5_149 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_81_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_12529_ clknet_leaf_59_clk _00081_ net187 vssd1 vssd1 vccd1 vccd1 genblk2\[0\].wave_shpr.div.b1\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_78_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_78_34 vssd1 vssd1 vccd1 vccd1 sky130_ef_sc_hd__decap_12
XFILLER_0_111_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_124_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_151_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_2_867 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_50_792 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__09220__B2 net804 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__08574__A3 _02350_ vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__07782__A1 genblk1\[0\].osc.clkdiv_C.cnt\[4\] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_09740_ _04217_ vssd1 vssd1 vccd1 vccd1 _00267_ sky130_fd_sc_hd__clkbuf_1
X_06952_ genblk1\[6\].osc.clkdiv_C.cnt\[16\] _01787_ vssd1 vssd1 vccd1 vccd1 _01790_
+ sky130_fd_sc_hd__nand2_1
.ends

