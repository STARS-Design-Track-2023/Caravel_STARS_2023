magic
tech sky130A
magscale 1 2
timestamp 1693970324
<< obsli1 >>
rect 1104 2159 34684 35377
<< obsm1 >>
rect 14 2128 34854 35408
<< metal2 >>
rect 1306 37217 1362 38017
rect 7746 37217 7802 38017
rect 13542 37217 13598 38017
rect 19982 37217 20038 38017
rect 26422 37217 26478 38017
rect 32862 37217 32918 38017
rect 18 0 74 800
rect 5814 0 5870 800
rect 12254 0 12310 800
rect 18694 0 18750 800
rect 24490 0 24546 800
rect 30930 0 30986 800
<< obsm2 >>
rect 20 37161 1250 37346
rect 1418 37161 7690 37346
rect 7858 37161 13486 37346
rect 13654 37161 19926 37346
rect 20094 37161 26366 37346
rect 26534 37161 32806 37346
rect 32974 37161 34850 37346
rect 20 856 34850 37161
rect 130 734 5758 856
rect 5926 734 12198 856
rect 12366 734 18638 856
rect 18806 734 24434 856
rect 24602 734 30874 856
rect 31042 734 34850 856
<< metal3 >>
rect 35073 34688 35873 34808
rect 0 32648 800 32768
rect 35073 27888 35873 28008
rect 0 25848 800 25968
rect 35073 21088 35873 21208
rect 0 19728 800 19848
rect 35073 14288 35873 14408
rect 0 12928 800 13048
rect 35073 8168 35873 8288
rect 0 6128 800 6248
rect 35073 1368 35873 1488
<< obsm3 >>
rect 798 34888 35082 35393
rect 798 34608 34993 34888
rect 798 32848 35082 34608
rect 880 32568 35082 32848
rect 798 28088 35082 32568
rect 798 27808 34993 28088
rect 798 26048 35082 27808
rect 880 25768 35082 26048
rect 798 21288 35082 25768
rect 798 21008 34993 21288
rect 798 19928 35082 21008
rect 880 19648 35082 19928
rect 798 14488 35082 19648
rect 798 14208 34993 14488
rect 798 13128 35082 14208
rect 880 12848 35082 13128
rect 798 8368 35082 12848
rect 798 8088 34993 8368
rect 798 6328 35082 8088
rect 880 6048 35082 6328
rect 798 1568 35082 6048
rect 798 1395 34993 1568
<< metal4 >>
rect 5141 2128 5461 35408
rect 9338 2128 9658 35408
rect 13535 2128 13855 35408
rect 17732 2128 18052 35408
rect 21929 2128 22249 35408
rect 26126 2128 26446 35408
rect 30323 2128 30643 35408
rect 34520 2128 34840 35408
<< obsm4 >>
rect 8339 13363 9141 17781
<< labels >>
rlabel metal3 s 35073 34688 35873 34808 6 clk
port 1 nsew signal input
rlabel metal3 s 0 32648 800 32768 6 en
port 2 nsew signal input
rlabel metal2 s 30930 0 30986 800 6 keypad_i[0]
port 3 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 keypad_i[10]
port 4 nsew signal input
rlabel metal3 s 0 19728 800 19848 6 keypad_i[11]
port 5 nsew signal input
rlabel metal2 s 7746 37217 7802 38017 6 keypad_i[12]
port 6 nsew signal input
rlabel metal2 s 13542 37217 13598 38017 6 keypad_i[13]
port 7 nsew signal input
rlabel metal2 s 32862 37217 32918 38017 6 keypad_i[14]
port 8 nsew signal input
rlabel metal3 s 35073 8168 35873 8288 6 keypad_i[1]
port 9 nsew signal input
rlabel metal2 s 24490 0 24546 800 6 keypad_i[2]
port 10 nsew signal input
rlabel metal2 s 18 0 74 800 6 keypad_i[3]
port 11 nsew signal input
rlabel metal2 s 5814 0 5870 800 6 keypad_i[4]
port 12 nsew signal input
rlabel metal3 s 0 12928 800 13048 6 keypad_i[5]
port 13 nsew signal input
rlabel metal3 s 35073 1368 35873 1488 6 keypad_i[6]
port 14 nsew signal input
rlabel metal2 s 12254 0 12310 800 6 keypad_i[7]
port 15 nsew signal input
rlabel metal3 s 35073 21088 35873 21208 6 keypad_i[8]
port 16 nsew signal input
rlabel metal3 s 35073 27888 35873 28008 6 keypad_i[9]
port 17 nsew signal input
rlabel metal2 s 19982 37217 20038 38017 6 n_rst
port 18 nsew signal input
rlabel metal2 s 26422 37217 26478 38017 6 pwm_o
port 19 nsew signal output
rlabel metal2 s 18694 0 18750 800 6 sound_series[0]
port 20 nsew signal output
rlabel metal3 s 0 25848 800 25968 6 sound_series[1]
port 21 nsew signal output
rlabel metal2 s 1306 37217 1362 38017 6 sound_series[2]
port 22 nsew signal output
rlabel metal3 s 35073 14288 35873 14408 6 sound_series[3]
port 23 nsew signal output
rlabel metal4 s 5141 2128 5461 35408 6 vccd1
port 24 nsew power bidirectional
rlabel metal4 s 13535 2128 13855 35408 6 vccd1
port 24 nsew power bidirectional
rlabel metal4 s 21929 2128 22249 35408 6 vccd1
port 24 nsew power bidirectional
rlabel metal4 s 30323 2128 30643 35408 6 vccd1
port 24 nsew power bidirectional
rlabel metal4 s 9338 2128 9658 35408 6 vssd1
port 25 nsew ground bidirectional
rlabel metal4 s 17732 2128 18052 35408 6 vssd1
port 25 nsew ground bidirectional
rlabel metal4 s 26126 2128 26446 35408 6 vssd1
port 25 nsew ground bidirectional
rlabel metal4 s 34520 2128 34840 35408 6 vssd1
port 25 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 35873 38017
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3646582
string GDS_FILE /home/designer-25/CUP/openlane/synth/runs/23_09_05_20_15/results/signoff/synth.magic.gds
string GDS_START 799820
<< end >>

