* NGSPICE file created from top8227.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_4 abstract view
.subckt sky130_fd_sc_hd__a31oi_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_2 abstract view
.subckt sky130_fd_sc_hd__a21boi_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_4 abstract view
.subckt sky130_fd_sc_hd__nand4b_4 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_2 abstract view
.subckt sky130_fd_sc_hd__a311oi_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4b_2 abstract view
.subckt sky130_fd_sc_hd__nand4b_2 A_N B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41oi_4 abstract view
.subckt sky130_fd_sc_hd__a41oi_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_1 abstract view
.subckt sky130_fd_sc_hd__o2111ai_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41ai_2 abstract view
.subckt sky130_fd_sc_hd__o41ai_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_1 abstract view
.subckt sky130_fd_sc_hd__o41a_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_2 abstract view
.subckt sky130_fd_sc_hd__a31oi_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_2 abstract view
.subckt sky130_fd_sc_hd__a221oi_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_4 abstract view
.subckt sky130_fd_sc_hd__mux2_4 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_2 abstract view
.subckt sky130_fd_sc_hd__o21ba_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_2 abstract view
.subckt sky130_fd_sc_hd__o22ai_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311oi_4 abstract view
.subckt sky130_fd_sc_hd__a311oi_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_2 abstract view
.subckt sky130_fd_sc_hd__or4bb_2 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_4 abstract view
.subckt sky130_fd_sc_hd__and4b_4 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_2 abstract view
.subckt sky130_fd_sc_hd__o311a_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_4 abstract view
.subckt sky130_fd_sc_hd__o221ai_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

.subckt top8227 M10ClkOut VGND VPWR addressBusHigh[0] addressBusHigh[1] addressBusHigh[2]
+ addressBusHigh[3] addressBusHigh[4] addressBusHigh[5] addressBusHigh[6] addressBusHigh[7]
+ addressBusLow[0] addressBusLow[1] addressBusLow[2] addressBusLow[3] addressBusLow[4]
+ addressBusLow[5] addressBusLow[6] addressBusLow[7] clk dataBusEnable dataBusInput[0]
+ dataBusInput[1] dataBusInput[2] dataBusInput[3] dataBusInput[4] dataBusInput[5]
+ dataBusInput[6] dataBusInput[7] dataBusOutput[0] dataBusOutput[1] dataBusOutput[2]
+ dataBusOutput[3] dataBusOutput[4] dataBusOutput[5] dataBusOutput[6] dataBusOutput[7]
+ dataBusSelect functionalClockOut interruptRequest nonMaskableInterrupt nrst readNotWrite
+ ready setOverflow sync
X_2037_ _0959_ net42 _0951_ _1241_ VGND VGND VPWR VPWR _1310_ sky130_fd_sc_hd__a211o_1
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3086_ clknet_4_8_0_clk _0078_ net63 VGND VGND VPWR VPWR internalDataflow.stackBusModule.busInputs\[43\]
+ sky130_fd_sc_hd__dfrtp_1
X_2106_ internalDataflow.addressLowBusModule.busInputs\[30\] _1377_ _1378_ internalDataflow.addressLowBusModule.busInputs\[38\]
+ VGND VGND VPWR VPWR _1379_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2939_ _0740_ _0741_ _0738_ VGND VGND VPWR VPWR _0752_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_67_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_383 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1606_ _0909_ _0865_ _0871_ VGND VGND VPWR VPWR _0913_ sky130_fd_sc_hd__a21oi_4
X_2724_ _0544_ _0567_ _0572_ VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__a21o_1
X_2655_ internalDataflow.accRegToDB\[1\] _0274_ _0511_ VGND VGND VPWR VPWR _0513_
+ sky130_fd_sc_hd__mux2_1
X_1537_ _0843_ VGND VGND VPWR VPWR _0844_ sky130_fd_sc_hd__clkbuf_4
X_2586_ _0290_ _0406_ _0452_ _0453_ _0455_ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__a32o_1
X_3138_ clknet_4_15_0_clk _0020_ net71 VGND VGND VPWR VPWR demux.state_machine.currentInstruction\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_3069_ clknet_4_9_0_clk _0061_ net63 VGND VGND VPWR VPWR internalDataflow.addressLowBusModule.busInputs\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_64_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2440_ _1008_ _0873_ _0327_ VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__a21oi_1
X_2371_ _0998_ _0253_ _0258_ VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__and3_1
XFILLER_0_42_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_4_12_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_12_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_6_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2707_ _0556_ VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__buf_2
X_2638_ net79 _0503_ _0281_ VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__a21o_1
X_2569_ net82 net45 _0436_ _0440_ VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__a211o_1
XFILLER_0_60_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1940_ _1061_ _1123_ _1157_ _1183_ VGND VGND VPWR VPWR _1220_ sky130_fd_sc_hd__or4_1
XFILLER_0_68_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1871_ _1150_ _0975_ _0972_ _1069_ _1153_ VGND VGND VPWR VPWR _1154_ sky130_fd_sc_hd__a221o_1
XFILLER_0_9_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2423_ internalDataflow.addressLowBusModule.busInputs\[23\] _1502_ _0127_ net9 _0122_
+ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__a221o_1
X_2354_ _0154_ _0241_ VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__and2_1
X_2285_ _1467_ _1479_ _0172_ VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2070_ _1182_ _1128_ _0910_ _1097_ VGND VGND VPWR VPWR _1343_ sky130_fd_sc_hd__or4_1
XFILLER_0_56_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2972_ _0999_ _0779_ _0781_ VGND VGND VPWR VPWR _0782_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1785_ _1068_ _1023_ VGND VGND VPWR VPWR _1069_ sky130_fd_sc_hd__nor2_4
X_1923_ _0882_ _1076_ VGND VGND VPWR VPWR _1204_ sky130_fd_sc_hd__nor2_1
X_1854_ _0866_ _0815_ VGND VGND VPWR VPWR _1138_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_161 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2406_ internalDataflow.addressLowBusModule.busInputs\[31\] _1377_ _1378_ internalDataflow.addressLowBusModule.busInputs\[39\]
+ VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__a22o_1
XFILLER_0_46_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2199_ _0873_ _0910_ _1471_ _1360_ _1006_ VGND VGND VPWR VPWR _1472_ sky130_fd_sc_hd__o32a_1
XFILLER_0_34_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2268_ _0147_ _0155_ VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__nand2_1
X_2337_ _0224_ _1366_ _1368_ _1350_ VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__or4_1
XFILLER_0_62_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold41 demux.state_machine.currentAddress\[9\] VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold30 net16 VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__dlygate4sd3_1
Xhold52 net22 VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_220 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1570_ _0876_ VGND VGND VPWR VPWR _0877_ sky130_fd_sc_hd__clkbuf_4
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2122_ _0936_ _0927_ _0847_ demux.state_machine.timeState\[0\] VGND VGND VPWR VPWR
+ _1395_ sky130_fd_sc_hd__a22o_1
X_2053_ _1323_ _1280_ _1324_ _1325_ VGND VGND VPWR VPWR _1326_ sky130_fd_sc_hd__a31oi_4
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2955_ _0665_ _0766_ _0544_ VGND VGND VPWR VPWR _0767_ sky130_fd_sc_hd__o21ai_1
X_1906_ _1065_ _1164_ _1184_ _1187_ VGND VGND VPWR VPWR _1188_ sky130_fd_sc_hd__or4_1
X_1768_ _0962_ _1026_ VGND VGND VPWR VPWR _1052_ sky130_fd_sc_hd__nor2_2
X_1837_ _0830_ _0885_ VGND VGND VPWR VPWR _1121_ sky130_fd_sc_hd__nor2_2
X_2886_ _0636_ _0702_ VGND VGND VPWR VPWR _0704_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1699_ _0879_ _0981_ _1000_ _0983_ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__a22o_1
XFILLER_0_12_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput31 net31 VGND VGND VPWR VPWR addressBusLow[7] sky130_fd_sc_hd__clkbuf_4
Xoutput20 net20 VGND VGND VPWR VPWR addressBusHigh[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput42 net42 VGND VGND VPWR VPWR readNotWrite sky130_fd_sc_hd__clkbuf_4
XFILLER_0_53_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1622_ _0926_ _0927_ _0928_ VGND VGND VPWR VPWR _0929_ sky130_fd_sc_hd__or3b_1
X_2671_ _0520_ _0324_ _0521_ VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_26_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2740_ _0585_ _0586_ VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__nor2_1
X_1553_ _0859_ VGND VGND VPWR VPWR _0860_ sky130_fd_sc_hd__buf_4
XTAP_189 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2036_ _1097_ _1248_ _1004_ VGND VGND VPWR VPWR _1309_ sky130_fd_sc_hd__o21ai_1
X_3085_ clknet_4_8_0_clk _0077_ net62 VGND VGND VPWR VPWR internalDataflow.stackBusModule.busInputs\[42\]
+ sky130_fd_sc_hd__dfrtp_1
X_2105_ net50 _1350_ _1303_ _1366_ VGND VGND VPWR VPWR _1378_ sky130_fd_sc_hd__and4b_2
XFILLER_0_72_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2938_ _0749_ _0750_ VGND VGND VPWR VPWR _0751_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2869_ _0691_ VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__clkbuf_1
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2723_ _0546_ _0570_ _0571_ _0555_ internalDataflow.addressLowBusModule.busInputs\[18\]
+ VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__a32o_1
XFILLER_0_13_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1536_ demux.state_machine.currentInstruction\[1\] demux.state_machine.currentInstruction\[2\]
+ demux.state_machine.currentInstruction\[3\] demux.state_machine.currentInstruction\[0\]
+ VGND VGND VPWR VPWR _0843_ sky130_fd_sc_hd__or4b_1
XFILLER_0_54_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1605_ _0826_ _0857_ VGND VGND VPWR VPWR _0912_ sky130_fd_sc_hd__nor2_4
X_2585_ _0158_ _0412_ _0410_ _0454_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__a211o_1
X_2654_ _0512_ VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3137_ clknet_4_4_0_clk internalDataflow.psr.processStatusReg.stat_buf_nxt\[6\] net60
+ VGND VGND VPWR VPWR demux.PSR_V sky130_fd_sc_hd__dfrtp_4
XFILLER_0_1_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2019_ branch_ff.branchForward _1290_ _1291_ _1261_ VGND VGND VPWR VPWR _1292_ sky130_fd_sc_hd__a211o_1
X_3068_ clknet_4_9_0_clk _0060_ net65 VGND VGND VPWR VPWR internalDataflow.addressLowBusModule.busInputs\[18\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_68_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2370_ _0255_ _0257_ _1439_ VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__or3b_1
XFILLER_0_46_104 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2706_ _0536_ VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__buf_2
XFILLER_0_6_278 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1519_ demux.state_machine.currentInstruction\[5\] _0820_ VGND VGND VPWR VPWR _0826_
+ sky130_fd_sc_hd__nand2b_4
X_2499_ _0134_ _0315_ _0372_ _0317_ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__a31o_2
X_2637_ net97 _0503_ _0241_ VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2568_ _0202_ _0407_ _0439_ _0361_ VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__o211a_1
XFILLER_0_65_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1870_ _1052_ _1133_ _1151_ _1066_ _1152_ VGND VGND VPWR VPWR _1153_ sky130_fd_sc_hd__a32o_1
XFILLER_0_28_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2353_ _0238_ _0239_ _0240_ VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__or3_4
XFILLER_0_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2422_ internalDataflow.addressLowBusModule.busInputs\[39\] net46 _0125_ internalDataflow.addressLowBusModule.busInputs\[31\]
+ VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__a22o_1
X_2284_ _0162_ _0169_ _0148_ VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__mux2_2
XFILLER_0_59_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1999_ _0868_ _1131_ _1271_ _1263_ VGND VGND VPWR VPWR _1272_ sky130_fd_sc_hd__o31a_1
XFILLER_0_34_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_11_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_11_0_clk sky130_fd_sc_hd__clkbuf_8
X_1922_ _1202_ _0976_ _1019_ _1087_ _1155_ VGND VGND VPWR VPWR _1203_ sky130_fd_sc_hd__a221o_1
XFILLER_0_56_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2971_ _1002_ _0929_ _1282_ _1102_ _0780_ VGND VGND VPWR VPWR _0781_ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1853_ _1033_ _1017_ _1133_ _1136_ VGND VGND VPWR VPWR _1137_ sky130_fd_sc_hd__a22o_1
X_1784_ _0965_ VGND VGND VPWR VPWR _1068_ sky130_fd_sc_hd__inv_2
XFILLER_0_24_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2405_ internalDataflow.stackBusModule.busInputs\[47\] _1373_ _1374_ internalDataflow.accRegToDB\[7\]
+ _1375_ VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__a221o_1
X_2336_ internalDataflow.stackBusModule.busInputs\[40\] VGND VGND VPWR VPWR _0224_
+ sky130_fd_sc_hd__inv_2
XFILLER_0_12_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2198_ _0913_ _1298_ _1248_ _1390_ VGND VGND VPWR VPWR _1471_ sky130_fd_sc_hd__or4b_1
XFILLER_0_27_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2267_ _0150_ _0153_ _0154_ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold20 demux.setInterruptFlag VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__dlygate4sd3_1
Xhold42 internalDataflow.stackBusModule.busInputs\[36\] VGND VGND VPWR VPWR net114
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold53 internalDataflow.addressHighBusModule.busInputs\[21\] VGND VGND VPWR VPWR
+ net125 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 internalDataflow.stackBusModule.busInputs\[45\] VGND VGND VPWR VPWR net103
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2121_ _0936_ _1144_ _0872_ _0875_ _1393_ VGND VGND VPWR VPWR _1394_ sky130_fd_sc_hd__a221o_1
X_2052_ _1310_ VGND VGND VPWR VPWR _1325_ sky130_fd_sc_hd__buf_4
XFILLER_0_16_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1905_ _1186_ VGND VGND VPWR VPWR _1187_ sky130_fd_sc_hd__inv_2
XFILLER_0_44_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2885_ _0636_ _0702_ VGND VGND VPWR VPWR _0703_ sky130_fd_sc_hd__nand2_1
X_2954_ _0755_ _0765_ VGND VGND VPWR VPWR _0766_ sky130_fd_sc_hd__nor2_1
X_1836_ _1052_ _1112_ _1113_ _1119_ VGND VGND VPWR VPWR _1120_ sky130_fd_sc_hd__a31o_1
X_1767_ _0819_ _0820_ VGND VGND VPWR VPWR _1051_ sky130_fd_sc_hd__and2b_1
X_1698_ _0982_ _0996_ _0962_ _0999_ VGND VGND VPWR VPWR _1000_ sky130_fd_sc_hd__o211a_2
XFILLER_0_4_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2319_ internalDataflow.addressLowBusModule.busInputs\[18\] _1315_ _0205_ _0206_
+ net48 VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__a2111o_1
Xoutput43 net43 VGND VGND VPWR VPWR sync sky130_fd_sc_hd__clkbuf_4
Xoutput21 net21 VGND VGND VPWR VPWR addressBusHigh[5] sky130_fd_sc_hd__clkbuf_4
Xoutput32 net32 VGND VGND VPWR VPWR dataBusOutput[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_53_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1621_ _0885_ _0855_ _0866_ VGND VGND VPWR VPWR _0928_ sky130_fd_sc_hd__a21o_1
X_1552_ _0813_ _0811_ _0810_ _0812_ VGND VGND VPWR VPWR _0859_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_41_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2670_ demux.nmi instructionLoader.interruptInjector.irqGenerated net43 instructionLoader.interruptInjector.resetDetected
+ VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__o22ai_4
XFILLER_0_1_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2104_ _1366_ _1341_ _1350_ VGND VGND VPWR VPWR _1377_ sky130_fd_sc_hd__and3_2
X_2035_ _1307_ VGND VGND VPWR VPWR _1308_ sky130_fd_sc_hd__inv_2
XFILLER_0_27_95 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3084_ clknet_4_2_0_clk _0076_ net59 VGND VGND VPWR VPWR internalDataflow.stackBusModule.busInputs\[41\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2868_ internalDataflow.addressLowBusModule.busInputs\[35\] _0194_ _0687_ VGND VGND
+ VPWR VPWR _0691_ sky130_fd_sc_hd__mux2_1
X_2937_ internalDataflow.addressHighBusModule.busInputs\[21\] _0558_ VGND VGND VPWR
+ VPWR _0750_ sky130_fd_sc_hd__nand2_1
XFILLER_0_68_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1819_ _0964_ _1017_ _1095_ _0974_ VGND VGND VPWR VPWR _1103_ sky130_fd_sc_hd__a31o_1
X_2799_ _1384_ _1487_ _0488_ _0641_ VGND VGND VPWR VPWR _0642_ sky130_fd_sc_hd__or4_1
XFILLER_0_25_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_94 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_116 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2722_ _0568_ _0569_ VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__or2_1
X_1535_ _0841_ _0836_ VGND VGND VPWR VPWR _0842_ sky130_fd_sc_hd__nor2_1
X_1604_ _0907_ _0908_ _0910_ VGND VGND VPWR VPWR _0911_ sky130_fd_sc_hd__or3_2
X_2584_ _1434_ _1460_ _0364_ _0408_ _0157_ VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__a32o_1
X_2653_ _0226_ _0249_ _0511_ VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__mux2_1
X_3067_ clknet_4_13_0_clk _0059_ net65 VGND VGND VPWR VPWR internalDataflow.addressLowBusModule.busInputs\[17\]
+ sky130_fd_sc_hd__dfrtp_4
X_3136_ clknet_4_12_0_clk internalDataflow.psr.processStatusReg.stat_buf_nxt\[3\]
+ net65 VGND VGND VPWR VPWR internalDataflow.dataBusModule.busInputs\[43\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_64_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2018_ _0912_ _1079_ _1003_ VGND VGND VPWR VPWR _1291_ sky130_fd_sc_hd__o21a_1
XFILLER_0_9_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2705_ _0554_ VGND VGND VPWR VPWR _0555_ sky130_fd_sc_hd__clkbuf_4
X_2636_ _0502_ VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__inv_2
XFILLER_0_57_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1518_ _0824_ VGND VGND VPWR VPWR _0825_ sky130_fd_sc_hd__buf_4
X_2498_ internalDataflow.dataBusModule.busInputs\[43\] _0320_ VGND VGND VPWR VPWR
+ _0382_ sky130_fd_sc_hd__and2_1
X_2567_ _0204_ _0412_ _0410_ _0438_ VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__a211o_1
XFILLER_0_69_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3119_ clknet_4_13_0_clk _0107_ net70 VGND VGND VPWR VPWR instructionLoader.interruptInjector.irqGenerated
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_52_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2352_ internalDataflow.addressLowBusModule.busInputs\[16\] _1502_ _0127_ net2 VGND
+ VGND VPWR VPWR _0240_ sky130_fd_sc_hd__a22o_1
X_2421_ _1468_ _1480_ _0308_ VGND VGND VPWR VPWR _0309_ sky130_fd_sc_hd__mux2_1
X_2283_ _1460_ _0170_ VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_414 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2619_ _1491_ _1150_ _1285_ _1259_ VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__a22o_1
X_1998_ _0818_ _0861_ _0901_ VGND VGND VPWR VPWR _1271_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_42_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1852_ _0958_ _1086_ _1134_ _1135_ VGND VGND VPWR VPWR _1136_ sky130_fd_sc_hd__a31o_1
XFILLER_0_56_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1921_ _0827_ _0882_ VGND VGND VPWR VPWR _1202_ sky130_fd_sc_hd__nor2_4
X_2970_ _1384_ _1260_ _1330_ VGND VGND VPWR VPWR _0780_ sky130_fd_sc_hd__or3_1
XFILLER_0_44_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1783_ _1066_ VGND VGND VPWR VPWR _1067_ sky130_fd_sc_hd__buf_2
XFILLER_0_71_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2404_ _0136_ _0291_ _0134_ VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__o21a_1
X_2266_ _1465_ VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__inv_2
X_2335_ _0216_ _0222_ VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__xor2_4
XFILLER_0_20_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2197_ _1469_ _1352_ _1001_ VGND VGND VPWR VPWR _1470_ sky130_fd_sc_hd__and3b_1
XFILLER_0_62_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold54 net32 VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__dlygate4sd3_1
Xhold32 internalDataflow.stackBusModule.busInputs\[33\] VGND VGND VPWR VPWR net104
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 internalDataflow.stackBusModule.busInputs\[34\] VGND VGND VPWR VPWR net93
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold43 net21 VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__dlygate4sd3_1
Xhold10 internalDataflow.addressLowBusModule.busInputs\[27\] VGND VGND VPWR VPWR net82
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_38_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_122 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2120_ _0831_ _0837_ _1244_ VGND VGND VPWR VPWR _1393_ sky130_fd_sc_hd__o21a_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2051_ _1005_ _0905_ VGND VGND VPWR VPWR _1324_ sky130_fd_sc_hd__nand2_2
XFILLER_0_29_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1835_ _0943_ _1066_ _1118_ VGND VGND VPWR VPWR _1119_ sky130_fd_sc_hd__a21bo_1
X_1904_ _0901_ _0852_ _0978_ _1185_ VGND VGND VPWR VPWR _1186_ sky130_fd_sc_hd__o31a_1
XFILLER_0_44_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2884_ _0605_ _0620_ _0621_ _0701_ VGND VGND VPWR VPWR _0702_ sky130_fd_sc_hd__and4_1
XFILLER_0_4_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2953_ _0557_ _0662_ VGND VGND VPWR VPWR _0765_ sky130_fd_sc_hd__xnor2_1
X_1766_ _0972_ _1048_ _1049_ _0939_ VGND VGND VPWR VPWR _1050_ sky130_fd_sc_hd__a22o_1
X_1697_ _0998_ VGND VGND VPWR VPWR _0999_ sky130_fd_sc_hd__buf_4
XFILLER_0_52_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2318_ internalDataflow.addressHighBusModule.busInputs\[18\] _1294_ _1314_ net4 VGND
+ VGND VPWR VPWR _0206_ sky130_fd_sc_hd__a22o_1
X_2249_ internalDataflow.stackBusModule.busInputs\[45\] _1373_ _1374_ internalDataflow.accRegToDB\[5\]
+ _1375_ VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__a221o_1
XFILLER_0_73_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_10_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_10_0_clk sky130_fd_sc_hd__clkbuf_8
Xoutput22 net22 VGND VGND VPWR VPWR addressBusHigh[6] sky130_fd_sc_hd__clkbuf_4
Xoutput33 net33 VGND VGND VPWR VPWR dataBusOutput[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1620_ _0841_ _0815_ VGND VGND VPWR VPWR _0927_ sky130_fd_sc_hd__nor2_4
X_1551_ _0834_ _0835_ VGND VGND VPWR VPWR _0858_ sky130_fd_sc_hd__or2b_1
XTAP_169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3083_ clknet_4_3_0_clk _0075_ net59 VGND VGND VPWR VPWR internalDataflow.stackBusModule.busInputs\[40\]
+ sky130_fd_sc_hd__dfrtp_1
X_2103_ internalDataflow.stackBusModule.busInputs\[46\] _1373_ _1374_ internalDataflow.accRegToDB\[6\]
+ _1375_ VGND VGND VPWR VPWR _1376_ sky130_fd_sc_hd__a221o_1
XFILLER_0_57_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2034_ _0941_ _1306_ VGND VGND VPWR VPWR _1307_ sky130_fd_sc_hd__or2_1
X_2798_ _0489_ _0637_ _0640_ VGND VGND VPWR VPWR _0641_ sky130_fd_sc_hd__or3_1
X_1818_ _0912_ VGND VGND VPWR VPWR _1102_ sky130_fd_sc_hd__clkbuf_4
X_2867_ _0690_ VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2936_ internalDataflow.addressHighBusModule.busInputs\[21\] _0557_ VGND VGND VPWR
+ VPWR _0749_ sky130_fd_sc_hd__or2_1
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1749_ _1026_ _1016_ _1036_ VGND VGND VPWR VPWR _1037_ sky130_fd_sc_hd__o21a_1
XFILLER_0_40_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2652_ _0345_ _0509_ _0510_ _0332_ VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__o31a_4
X_2721_ _0568_ _0569_ VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__nand2_1
XFILLER_0_14_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1534_ demux.state_machine.currentInstruction\[5\] demux.state_machine.currentInstruction\[4\]
+ VGND VGND VPWR VPWR _0841_ sky130_fd_sc_hd__or2_2
X_1603_ _0826_ _0909_ VGND VGND VPWR VPWR _0910_ sky130_fd_sc_hd__nor2_4
X_2583_ _0156_ _0410_ VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__nand2_1
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2017_ _0888_ net52 _0917_ VGND VGND VPWR VPWR _1290_ sky130_fd_sc_hd__a21oi_4
X_3135_ clknet_4_12_0_clk internalDataflow.psr.processStatusReg.stat_buf_nxt\[2\]
+ net70 VGND VGND VPWR VPWR instructionLoader.interruptInjector.processStatusRegIFlag
+ sky130_fd_sc_hd__dfrtp_2
X_3066_ clknet_4_9_0_clk _0058_ net65 VGND VGND VPWR VPWR internalDataflow.addressLowBusModule.busInputs\[16\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_70_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2919_ internalDataflow.addressHighBusModule.busInputs\[18\] _0556_ _0720_ VGND VGND
+ VPWR VPWR _0734_ sky130_fd_sc_hd__a21boi_2
XFILLER_0_72_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_320 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2635_ _0999_ _0497_ _0501_ VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__and3_4
XFILLER_0_42_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2704_ _0538_ _0553_ VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__and2_2
X_1517_ _0812_ _0813_ _0811_ _0810_ VGND VGND VPWR VPWR _0824_ sky130_fd_sc_hd__or4b_1
X_2497_ _0376_ _0379_ _0380_ VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__and3_1
XFILLER_0_4_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2566_ _0203_ _0437_ _0364_ _0171_ VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__a2bb2o_1
X_3118_ clknet_4_14_0_clk instructionLoader.interruptInjector.interruptRequest net71
+ VGND VGND VPWR VPWR instructionLoader.interruptInjector.irqSync.nextQ2 sky130_fd_sc_hd__dfrtp_1
X_3049_ clknet_4_0_0_clk _0041_ net57 VGND VGND VPWR VPWR internalDataflow.addressLowBusModule.busInputs\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2420_ _1257_ _0296_ _0307_ VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_24_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2351_ internalDataflow.addressLowBusModule.busInputs\[32\] net46 _0125_ internalDataflow.addressLowBusModule.busInputs\[24\]
+ VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__a22o_1
X_2282_ _0164_ _0169_ _1329_ VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__mux2_2
XFILLER_0_19_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1997_ _1266_ _1267_ _1269_ VGND VGND VPWR VPWR _1270_ sky130_fd_sc_hd__or3b_1
X_2618_ _1001_ _0848_ _1395_ _1396_ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__a211o_1
XFILLER_0_42_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2549_ _0216_ _0222_ _0408_ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__o21a_1
XFILLER_0_65_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1851_ _1012_ _0969_ _0956_ _1024_ VGND VGND VPWR VPWR _1135_ sky130_fd_sc_hd__o211a_1
X_1920_ _1200_ _0976_ _1054_ _1095_ _1158_ VGND VGND VPWR VPWR _1201_ sky130_fd_sc_hd__a221o_1
XFILLER_0_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1782_ _0974_ VGND VGND VPWR VPWR _1066_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2403_ _0156_ _0290_ VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2196_ _0888_ net53 VGND VGND VPWR VPWR _1469_ sky130_fd_sc_hd__and2_1
X_2265_ _0151_ _0152_ _0123_ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__o21a_4
X_2334_ _0218_ _0221_ _0154_ VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__mux2_2
XFILLER_0_62_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold22 branch_ff.branchForward VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__dlygate4sd3_1
Xhold11 internalDataflow.addressLowBusModule.busInputs\[31\] VGND VGND VPWR VPWR net83
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold55 net20 VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__dlygate4sd3_1
Xhold44 net36 VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 internalDataflow.stackBusModule.busInputs\[42\] VGND VGND VPWR VPWR net105
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_67_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2050_ _1005_ _0927_ VGND VGND VPWR VPWR _1323_ sky130_fd_sc_hd__nand2_1
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2952_ _0761_ _0763_ VGND VGND VPWR VPWR _0764_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1834_ _0974_ _0964_ _1115_ _1117_ VGND VGND VPWR VPWR _1118_ sky130_fd_sc_hd__or4_1
X_1903_ _1047_ _1087_ VGND VGND VPWR VPWR _1185_ sky130_fd_sc_hd__nand2_1
X_1765_ _0836_ _0978_ VGND VGND VPWR VPWR _1049_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2883_ _0312_ _0537_ VGND VGND VPWR VPWR _0701_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1696_ _0997_ VGND VGND VPWR VPWR _0998_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_73_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2179_ _1004_ _1237_ VGND VGND VPWR VPWR _1452_ sky130_fd_sc_hd__and2_1
X_2248_ _0134_ _0135_ VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__nand2_2
X_2317_ internalDataflow.accRegToDB\[2\] _1316_ _1318_ instructionLoader.interruptInjector.processStatusRegIFlag
+ VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__a22o_1
XFILLER_0_35_248 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput34 net34 VGND VGND VPWR VPWR dataBusOutput[2] sky130_fd_sc_hd__clkbuf_4
Xoutput23 net23 VGND VGND VPWR VPWR addressBusHigh[7] sky130_fd_sc_hd__buf_2
XFILLER_0_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1550_ _0812_ _0833_ _0834_ _0835_ VGND VGND VPWR VPWR _0857_ sky130_fd_sc_hd__nand4b_4
XFILLER_0_34_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3082_ clknet_4_13_0_clk _0074_ net70 VGND VGND VPWR VPWR demux.reset sky130_fd_sc_hd__dfrtp_4
X_2033_ _0876_ _0879_ _0912_ VGND VGND VPWR VPWR _1306_ sky130_fd_sc_hd__o21a_1
XTAP_159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2102_ _1370_ _1367_ VGND VGND VPWR VPWR _1375_ sky130_fd_sc_hd__nor2_2
XFILLER_0_49_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2935_ net132 _0555_ _0742_ _0743_ _0748_ VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1748_ net4 _0957_ VGND VGND VPWR VPWR _1036_ sky130_fd_sc_hd__nand2_1
X_1817_ _0907_ _0975_ _1048_ _1095_ VGND VGND VPWR VPWR _1101_ sky130_fd_sc_hd__a22o_1
X_2797_ demux.state_machine.timeState\[3\] _1079_ _0494_ _1102_ _0639_ VGND VGND VPWR
+ VPWR _0640_ sky130_fd_sc_hd__a221o_1
XFILLER_0_4_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2866_ internalDataflow.addressLowBusModule.busInputs\[34\] _0215_ _0687_ VGND VGND
+ VPWR VPWR _0690_ sky130_fd_sc_hd__mux2_1
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1679_ _0961_ VGND VGND VPWR VPWR _0981_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_63_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2651_ _0839_ _1058_ _1128_ _1008_ VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__o31a_1
X_1602_ _0810_ _0811_ _0812_ _0833_ VGND VGND VPWR VPWR _0909_ sky130_fd_sc_hd__nand4b_4
X_2720_ _0547_ _0550_ _0549_ VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__o21bai_2
XFILLER_0_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2582_ _0158_ _0289_ VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__or2_1
X_1533_ _0831_ _0837_ _0839_ VGND VGND VPWR VPWR _0840_ sky130_fd_sc_hd__or3_2
XFILLER_0_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2016_ _1278_ _1280_ _1281_ _1288_ VGND VGND VPWR VPWR _1289_ sky130_fd_sc_hd__a31o_2
X_3134_ clknet_4_12_0_clk internalDataflow.psr.processStatusReg.stat_buf_nxt\[1\]
+ net65 VGND VGND VPWR VPWR demux.PSR_Z sky130_fd_sc_hd__dfrtp_2
X_3065_ clknet_4_8_0_clk _0057_ net62 VGND VGND VPWR VPWR internalDataflow.accRegToDB\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2918_ _0731_ _0732_ VGND VGND VPWR VPWR _0733_ sky130_fd_sc_hd__nor2_1
X_2849_ _0679_ VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__clkbuf_1
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1516_ _0822_ VGND VGND VPWR VPWR _0823_ sky130_fd_sc_hd__inv_2
X_2634_ _0985_ _1244_ _1285_ _0987_ _0500_ VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2565_ _1131_ _0323_ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__nand2_1
X_2703_ _0542_ VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3117_ clknet_4_14_0_clk net74 net71 VGND VGND VPWR VPWR instructionLoader.interruptInjector.irqGeneratedFF.synchronizedIRQ
+ sky130_fd_sc_hd__dfrtp_1
X_2496_ _0134_ _0372_ _0378_ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__nand3_2
XFILLER_0_4_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3048_ clknet_4_1_0_clk _0040_ net60 VGND VGND VPWR VPWR internalDataflow.addressLowBusModule.busInputs\[30\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_5_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2350_ _1265_ _1303_ _1267_ _0122_ VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__and4_1
X_2281_ internalDataflow.addressHighBusModule.busInputs\[20\] _1294_ net134 _0168_
+ VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__a211o_1
XFILLER_0_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1996_ _1268_ _0832_ _0827_ _0858_ VGND VGND VPWR VPWR _1269_ sky130_fd_sc_hd__or4_1
XFILLER_0_27_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2617_ _1001_ _0911_ _1391_ _0934_ VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__a211o_1
XFILLER_0_42_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2548_ _0223_ _0412_ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__and2_1
X_2479_ _0909_ _0852_ _1076_ VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_65_246 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1850_ _1095_ VGND VGND VPWR VPWR _1134_ sky130_fd_sc_hd__inv_2
X_1781_ _1057_ _1061_ _1064_ VGND VGND VPWR VPWR _1065_ sky130_fd_sc_hd__or3_1
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2333_ internalDataflow.addressLowBusModule.busInputs\[18\] _1502_ _0127_ net4 _0220_
+ VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__a221o_4
XFILLER_0_20_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2402_ _0158_ _0289_ VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__nand2_1
X_2195_ _1467_ VGND VGND VPWR VPWR _1468_ sky130_fd_sc_hd__inv_2
X_2264_ internalDataflow.addressLowBusModule.busInputs\[21\] _1502_ _0127_ net7 _0122_
+ VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__a221o_1
XFILLER_0_47_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1979_ _1244_ _1247_ _1250_ _1001_ _1251_ VGND VGND VPWR VPWR _1252_ sky130_fd_sc_hd__a221o_1
Xhold12 demux.state_machine.timeState\[3\] VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__dlygate4sd3_1
Xhold23 branch_ff.branchBackward VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__dlygate4sd3_1
Xhold45 net37 VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__dlygate4sd3_1
Xhold56 internalDataflow.stackBusModule.busInputs\[41\] VGND VGND VPWR VPWR net128
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 internalDataflow.stackBusModule.busInputs\[35\] VGND VGND VPWR VPWR net106
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1902_ _1047_ _1059_ _1092_ _1180_ _1183_ VGND VGND VPWR VPWR _1184_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_32_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2951_ _0749_ _0752_ _0762_ VGND VGND VPWR VPWR _0763_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_55 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1764_ _0978_ _0964_ _1041_ VGND VGND VPWR VPWR _1048_ sky130_fd_sc_hd__and3_4
X_1833_ _1074_ _1116_ VGND VGND VPWR VPWR _1117_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2882_ _0696_ _0698_ VGND VGND VPWR VPWR _0700_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1695_ _0959_ net42 _0951_ VGND VGND VPWR VPWR _0997_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_12_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2316_ _0202_ _0203_ VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__nor2_2
X_2178_ _0982_ _1324_ VGND VGND VPWR VPWR _1451_ sky130_fd_sc_hd__nand2_1
X_2247_ _1461_ _0132_ VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__nand2_1
XFILLER_0_35_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput24 net24 VGND VGND VPWR VPWR addressBusLow[0] sky130_fd_sc_hd__clkbuf_4
Xoutput35 net35 VGND VGND VPWR VPWR dataBusOutput[3] sky130_fd_sc_hd__clkbuf_4
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3081_ clknet_4_14_0_clk _0073_ net71 VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__dfrtp_1
X_2032_ branch_ff.branchBackward _1290_ VGND VGND VPWR VPWR _1305_ sky130_fd_sc_hd__nand2_1
X_2101_ _1366_ _1342_ _1350_ VGND VGND VPWR VPWR _1374_ sky130_fd_sc_hd__and3b_2
X_2865_ _0689_ VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2934_ _0659_ _0746_ _0747_ VGND VGND VPWR VPWR _0748_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1747_ net78 _0977_ _1032_ _1035_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__a211o_1
X_1816_ _1065_ _1073_ _1093_ _1099_ VGND VGND VPWR VPWR _1100_ sky130_fd_sc_hd__or4_1
X_1678_ _0966_ _0972_ _0980_ VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__a21boi_1
X_2796_ _1007_ _0491_ _1084_ _0638_ VGND VGND VPWR VPWR _0639_ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_330 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1601_ _0829_ _0838_ VGND VGND VPWR VPWR _0908_ sky130_fd_sc_hd__nor2_1
X_1532_ _0827_ _0838_ VGND VGND VPWR VPWR _0839_ sky130_fd_sc_hd__nor2_2
X_2650_ _0868_ _0870_ _1202_ _1002_ VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__o31a_1
X_2581_ _0375_ _0381_ _0383_ _0321_ VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3133_ clknet_4_12_0_clk internalDataflow.psr.processStatusReg.stat_buf_nxt\[0\]
+ net65 VGND VGND VPWR VPWR demux.PSR_C sky130_fd_sc_hd__dfrtp_2
XFILLER_0_54_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2015_ _1284_ _1287_ VGND VGND VPWR VPWR _1288_ sky130_fd_sc_hd__nor2_1
X_3064_ clknet_4_8_0_clk _0056_ net63 VGND VGND VPWR VPWR internalDataflow.accRegToDB\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_2848_ net110 _0194_ _0675_ VGND VGND VPWR VPWR _0679_ sky130_fd_sc_hd__mux2_1
X_2917_ internalDataflow.addressHighBusModule.busInputs\[19\] _0556_ VGND VGND VPWR
+ VPWR _0732_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2779_ _0312_ _0622_ VGND VGND VPWR VPWR _0623_ sky130_fd_sc_hd__xor2_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_160 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2702_ _0547_ _0551_ VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1515_ _0815_ _0816_ _0818_ _0821_ VGND VGND VPWR VPWR _0822_ sky130_fd_sc_hd__a31o_2
X_2633_ _0498_ _1495_ _0499_ VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__or3b_1
X_2495_ _0134_ _0372_ _0378_ VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2564_ _0418_ _0433_ _0434_ _0435_ VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__o211a_1
X_3116_ clknet_4_15_0_clk instructionLoader.interruptInjector.nmiSync.in net71 VGND
+ VGND VPWR VPWR instructionLoader.interruptInjector.nmiSync.nextQ2 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3047_ clknet_4_1_0_clk _0039_ net60 VGND VGND VPWR VPWR internalDataflow.addressLowBusModule.busInputs\[29\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_60_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout70 net71 VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2280_ internalDataflow.accRegToDB\[4\] _1316_ _1314_ net6 _0167_ VGND VGND VPWR
+ VPWR _0168_ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_200 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2616_ _1406_ _1405_ VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__nand2_1
X_1995_ demux.state_machine.timeState\[0\] VGND VGND VPWR VPWR _1268_ sky130_fd_sc_hd__inv_2
XFILLER_0_15_358 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2478_ _0315_ _0318_ _0321_ _0361_ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__a31o_1
XFILLER_0_23_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2547_ net96 net45 _0417_ _0420_ VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__a22o_1
XFILLER_0_65_258 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1780_ _0842_ _0975_ _1048_ _1063_ VGND VGND VPWR VPWR _1064_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2332_ internalDataflow.addressLowBusModule.busInputs\[34\] net46 _0125_ internalDataflow.addressLowBusModule.busInputs\[26\]
+ _0219_ VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__a221o_1
X_2401_ _0182_ _0288_ _0179_ VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__a21o_1
XFILLER_0_46_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2194_ _1325_ _1466_ VGND VGND VPWR VPWR _1467_ sky130_fd_sc_hd__nor2_2
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2263_ internalDataflow.addressLowBusModule.busInputs\[37\] net46 _0125_ internalDataflow.addressLowBusModule.busInputs\[29\]
+ VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1978_ _0877_ _0915_ _0930_ _1004_ VGND VGND VPWR VPWR _1251_ sky130_fd_sc_hd__a22o_1
XFILLER_0_30_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold13 demux.state_machine.currentAddress\[3\] VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__dlygate4sd3_1
Xhold46 free_carry_ff.freeCarry VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__dlygate4sd3_1
Xhold57 internalDataflow.addressLowBusModule.busInputs\[30\] VGND VGND VPWR VPWR net129
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 internalDataflow.stackBusModule.busInputs\[44\] VGND VGND VPWR VPWR net107
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 internalDataflow.addressLowBusModule.busInputs\[25\] VGND VGND VPWR VPWR net96
+ sky130_fd_sc_hd__dlygate4sd3_1
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_16_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1901_ _0966_ _1063_ _1181_ _0974_ _1182_ VGND VGND VPWR VPWR _1183_ sky130_fd_sc_hd__a32o_1
X_1832_ _1055_ _1063_ VGND VGND VPWR VPWR _1116_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2881_ _0696_ _0698_ VGND VGND VPWR VPWR _0699_ sky130_fd_sc_hd__or2_1
XFILLER_0_29_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2950_ internalDataflow.addressHighBusModule.busInputs\[21\] _0557_ VGND VGND VPWR
+ VPWR _0762_ sky130_fd_sc_hd__and2_1
X_1763_ net76 _0977_ _1047_ VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__a21o_1
X_1694_ _0983_ _0985_ _0986_ _0990_ _0995_ VGND VGND VPWR VPWR _0996_ sky130_fd_sc_hd__a311oi_2
XFILLER_0_52_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2246_ _0133_ VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__buf_2
X_2315_ _0195_ _0201_ VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__nor2_1
X_2177_ _1439_ _1440_ _1445_ _1449_ VGND VGND VPWR VPWR _1450_ sky130_fd_sc_hd__a31o_1
XFILLER_0_18_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput36 net36 VGND VGND VPWR VPWR dataBusOutput[4] sky130_fd_sc_hd__clkbuf_4
Xoutput25 net25 VGND VGND VPWR VPWR addressBusLow[1] sky130_fd_sc_hd__clkbuf_4
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3080_ clknet_4_10_0_clk _0072_ net64 VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__dfrtp_1
X_2100_ _1366_ _1342_ _1369_ VGND VGND VPWR VPWR _1373_ sky130_fd_sc_hd__and3b_2
X_2031_ _1303_ _1292_ _1301_ VGND VGND VPWR VPWR _1304_ sky130_fd_sc_hd__a21boi_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1815_ _1096_ _1098_ VGND VGND VPWR VPWR _1099_ sky130_fd_sc_hd__or2_1
X_2795_ _0820_ VGND VGND VPWR VPWR _0638_ sky130_fd_sc_hd__inv_2
XFILLER_0_43_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2864_ internalDataflow.addressLowBusModule.busInputs\[33\] _0274_ _0687_ VGND VGND
+ VPWR VPWR _0689_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2933_ _0659_ _0746_ _0544_ VGND VGND VPWR VPWR _0747_ sky130_fd_sc_hd__o21ai_1
X_1746_ _0966_ _1033_ _1017_ _1019_ _1034_ VGND VGND VPWR VPWR _1035_ sky130_fd_sc_hd__a32o_1
X_1677_ demux.state_machine.currentAddress\[7\] _0958_ _0979_ VGND VGND VPWR VPWR
+ _0980_ sky130_fd_sc_hd__mux2_1
XFILLER_0_25_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2229_ _1501_ VGND VGND VPWR VPWR _1502_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_48_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1600_ _0857_ _0829_ VGND VGND VPWR VPWR _0907_ sky130_fd_sc_hd__nor2_1
X_1531_ _0833_ _0834_ _0835_ _0832_ VGND VGND VPWR VPWR _0838_ sky130_fd_sc_hd__nand4b_2
X_2580_ _0376_ _0379_ _0380_ _0383_ _0375_ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__a41oi_4
XFILLER_0_22_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_22_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3132_ clknet_4_5_0_clk _0019_ net69 VGND VGND VPWR VPWR demux.state_machine.timeState\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_38_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3063_ clknet_4_9_0_clk _0055_ net63 VGND VGND VPWR VPWR internalDataflow.accRegToDB\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2014_ _0985_ _1244_ _1286_ _0948_ VGND VGND VPWR VPWR _1287_ sky130_fd_sc_hd__a211o_1
XFILLER_0_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_323 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2778_ _0605_ _0620_ _0621_ VGND VGND VPWR VPWR _0622_ sky130_fd_sc_hd__and3_1
X_2847_ _0678_ VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2916_ internalDataflow.addressHighBusModule.busInputs\[19\] _0556_ VGND VGND VPWR
+ VPWR _0731_ sky130_fd_sc_hd__nor2_1
X_1729_ _1021_ VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2632_ demux.state_machine.currentAddress\[6\] _1441_ _0982_ VGND VGND VPWR VPWR
+ _0499_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_40_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2701_ _0549_ _0550_ VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__nor2_1
XFILLER_0_27_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1514_ _0819_ _0820_ VGND VGND VPWR VPWR _0821_ sky130_fd_sc_hd__nand2_4
XFILLER_0_49_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2494_ _0315_ _0377_ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__nand2_2
XFILLER_0_10_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2563_ _0204_ _0287_ VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__or2_1
X_3115_ clknet_4_15_0_clk net73 net71 VGND VGND VPWR VPWR instructionLoader.interruptInjector.nmiGeneratedFF.synchronizedNMI
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3046_ clknet_4_1_0_clk _0038_ net57 VGND VGND VPWR VPWR internalDataflow.addressLowBusModule.busInputs\[28\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xfanout71 net72 VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__buf_4
Xfanout60 net61 VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__buf_4
XFILLER_0_24_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1994_ demux.state_machine.timeState\[1\] _0891_ _1084_ VGND VGND VPWR VPWR _1267_
+ sky130_fd_sc_hd__and3_2
XFILLER_0_19_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2615_ net83 net45 _0482_ VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_15_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2477_ _0359_ _0360_ _1478_ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__o21ai_4
X_2546_ _0406_ _0419_ VGND VGND VPWR VPWR _0420_ sky130_fd_sc_hd__nand2_1
X_3029_ clknet_4_7_0_clk _0001_ net67 VGND VGND VPWR VPWR demux.state_machine.currentAddress\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_38_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_112 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2400_ _0204_ _0287_ _0202_ VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__a21o_1
XFILLER_0_21_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2331_ demux.nmi _1425_ _0122_ VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__and3b_1
X_2262_ _1467_ _1479_ _0149_ VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_384 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2193_ _1274_ _1453_ VGND VGND VPWR VPWR _1466_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1977_ _1121_ _0943_ _1131_ _1249_ VGND VGND VPWR VPWR _1250_ sky130_fd_sc_hd__or4_1
XFILLER_0_47_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2529_ _0261_ _0251_ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__and2b_1
XFILLER_0_15_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold14 demux.state_machine.currentAddress\[10\] VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__dlygate4sd3_1
Xhold25 net24 VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__dlygate4sd3_1
Xhold58 internalDataflow.addressHighBusModule.busInputs\[18\] VGND VGND VPWR VPWR
+ net130 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 net18 VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__dlygate4sd3_1
Xhold47 internalDataflow.addressHighBusModule.busInputs\[22\] VGND VGND VPWR VPWR
+ net119 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1831_ _1114_ net3 _1010_ _1053_ _1012_ VGND VGND VPWR VPWR _1115_ sky130_fd_sc_hd__o2111ai_1
X_1900_ _0866_ _0825_ VGND VGND VPWR VPWR _1182_ sky130_fd_sc_hd__nor2_1
XFILLER_0_44_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2880_ _0615_ _0617_ _0624_ _0697_ _0613_ VGND VGND VPWR VPWR _0698_ sky130_fd_sc_hd__a311o_1
XFILLER_0_29_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1762_ _1046_ VGND VGND VPWR VPWR _1047_ sky130_fd_sc_hd__clkbuf_4
X_1693_ _0991_ _0993_ _0994_ VGND VGND VPWR VPWR _0995_ sky130_fd_sc_hd__a21o_1
XFILLER_0_40_402 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2176_ _0982_ _1447_ _1448_ VGND VGND VPWR VPWR _1449_ sky130_fd_sc_hd__nor3_1
X_2245_ _1461_ _0132_ VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__or2_1
X_2314_ _0195_ _0201_ VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__and2_1
XFILLER_0_20_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput15 net15 VGND VGND VPWR VPWR M10ClkOut sky130_fd_sc_hd__buf_1
Xoutput37 net37 VGND VGND VPWR VPWR dataBusOutput[5] sky130_fd_sc_hd__clkbuf_4
Xoutput26 net26 VGND VGND VPWR VPWR addressBusLow[2] sky130_fd_sc_hd__clkbuf_4
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2030_ _0952_ VGND VGND VPWR VPWR _1303_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_27_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2932_ _0729_ _0744_ _0745_ VGND VGND VPWR VPWR _0746_ sky130_fd_sc_hd__and3_1
X_1814_ _1097_ _1067_ _1059_ _1069_ VGND VGND VPWR VPWR _1098_ sky130_fd_sc_hd__a22o_1
X_1745_ _0961_ _1023_ VGND VGND VPWR VPWR _1034_ sky130_fd_sc_hd__nor2_1
X_2794_ _1007_ _1400_ _1168_ VGND VGND VPWR VPWR _0637_ sky130_fd_sc_hd__o21a_1
X_2863_ _0688_ VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__inv_2
XFILLER_0_68_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1676_ _0978_ VGND VGND VPWR VPWR _0979_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_0_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2228_ _1484_ _1488_ _1490_ _1500_ VGND VGND VPWR VPWR _1501_ sky130_fd_sc_hd__and4_1
XFILLER_0_30_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2159_ internalDataflow.addressHighBusModule.busInputs\[22\] _1422_ _1424_ net8 _1431_
+ VGND VGND VPWR VPWR _1432_ sky130_fd_sc_hd__o221a_1
XFILLER_0_63_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1530_ _0827_ _0836_ VGND VGND VPWR VPWR _0837_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_11 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2013_ _0932_ _0991_ _1285_ demux.state_machine.currentAddress\[1\] VGND VGND VPWR
+ VPWR _1286_ sky130_fd_sc_hd__a22o_1
X_3131_ clknet_4_5_0_clk _0018_ net69 VGND VGND VPWR VPWR demux.state_machine.timeState\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_3062_ clknet_4_2_0_clk _0054_ net62 VGND VGND VPWR VPWR internalDataflow.accRegToDB\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_195 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2915_ _0656_ _0729_ VGND VGND VPWR VPWR _0730_ sky130_fd_sc_hd__xor2_1
X_1728_ _1015_ _1020_ VGND VGND VPWR VPWR _1021_ sky130_fd_sc_hd__and2b_1
XFILLER_0_60_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2777_ _0130_ _0153_ _0536_ VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__o21ai_1
X_2846_ net105 _0215_ _0675_ VGND VGND VPWR VPWR _0678_ sky130_fd_sc_hd__mux2_1
XFILLER_0_13_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1659_ _0961_ _0962_ VGND VGND VPWR VPWR _0963_ sky130_fd_sc_hd__nor2_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_195 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_46 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2631_ _1435_ _0993_ _1244_ demux.state_machine.currentAddress\[7\] _0994_ VGND VGND
+ VPWR VPWR _0498_ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2700_ _0548_ _0521_ _0533_ VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__and3_1
XFILLER_0_27_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2562_ _0204_ _0287_ _0361_ VGND VGND VPWR VPWR _0434_ sky130_fd_sc_hd__a21oi_1
X_1513_ demux.state_machine.currentInstruction\[4\] VGND VGND VPWR VPWR _0820_ sky130_fd_sc_hd__buf_4
X_2493_ _0317_ VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__inv_2
X_3114_ clknet_4_11_0_clk _0106_ net66 VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__dfrtp_1
X_3045_ clknet_4_0_0_clk _0037_ net57 VGND VGND VPWR VPWR internalDataflow.addressLowBusModule.busInputs\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2829_ net124 _0665_ _0645_ VGND VGND VPWR VPWR _0666_ sky130_fd_sc_hd__mux2_1
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout72 net12 VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_36_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout61 net12 VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__buf_2
XFILLER_0_32_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_316 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_10_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_257 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1993_ _1265_ _0871_ _0865_ VGND VGND VPWR VPWR _1266_ sky130_fd_sc_hd__nor3_1
XFILLER_0_15_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2614_ _0475_ _0481_ _0321_ VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2545_ _0367_ _0418_ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__xor2_1
X_2476_ _1462_ _1290_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__or2_2
X_3028_ clknet_4_7_0_clk _0012_ net68 VGND VGND VPWR VPWR demux.state_machine.currentAddress\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2192_ _1303_ _1464_ VGND VGND VPWR VPWR _1465_ sky130_fd_sc_hd__nand2_2
X_2261_ _0140_ _0145_ _0148_ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__mux2_2
X_2330_ _1467_ _1479_ _0217_ VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1976_ _0828_ _1248_ VGND VGND VPWR VPWR _1249_ sky130_fd_sc_hd__or2_2
XFILLER_0_47_249 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2528_ _0358_ _0360_ _0402_ _1478_ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__o31ai_2
XFILLER_0_30_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold26 pulse_slower.currentEnableState\[0\] VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__dlygate4sd3_1
Xhold48 internalDataflow.addressLowBusModule.busInputs\[22\] VGND VGND VPWR VPWR net120
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 net39 VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__dlygate4sd3_1
Xhold59 internalDataflow.stackBusModule.busInputs\[39\] VGND VGND VPWR VPWR net131
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold37 internalDataflow.stackBusModule.busInputs\[38\] VGND VGND VPWR VPWR net109
+ sky130_fd_sc_hd__dlygate4sd3_1
X_2459_ _0149_ _0172_ _0196_ _0217_ VGND VGND VPWR VPWR _0344_ sky130_fd_sc_hd__or4_1
XFILLER_0_38_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1761_ _0963_ _0964_ _1030_ VGND VGND VPWR VPWR _1046_ sky130_fd_sc_hd__and3_1
XFILLER_0_52_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1830_ net2 VGND VGND VPWR VPWR _1114_ sky130_fd_sc_hd__inv_2
X_1692_ _0932_ demux.state_machine.currentAddress\[5\] VGND VGND VPWR VPWR _0994_
+ sky130_fd_sc_hd__and2_1
XFILLER_0_40_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2313_ _0197_ _0200_ _0154_ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2175_ _0987_ demux.state_machine.currentAddress\[6\] _1283_ VGND VGND VPWR VPWR
+ _1448_ sky130_fd_sc_hd__o21a_1
XFILLER_0_32_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2244_ _1465_ _1483_ _0131_ VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__a21o_1
XFILLER_0_25_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1959_ net11 VGND VGND VPWR VPWR instructionLoader.interruptInjector.nmiSync.in sky130_fd_sc_hd__inv_2
XFILLER_0_22_90 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput38 net38 VGND VGND VPWR VPWR dataBusOutput[6] sky130_fd_sc_hd__clkbuf_4
Xoutput16 net16 VGND VGND VPWR VPWR addressBusHigh[0] sky130_fd_sc_hd__clkbuf_4
Xoutput27 net27 VGND VGND VPWR VPWR addressBusLow[3] sky130_fd_sc_hd__clkbuf_4
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2931_ _0557_ _0656_ VGND VGND VPWR VPWR _0745_ sky130_fd_sc_hd__or2_1
X_1744_ _1013_ VGND VGND VPWR VPWR _1033_ sky130_fd_sc_hd__inv_2
X_1813_ _0866_ _0861_ VGND VGND VPWR VPWR _1097_ sky130_fd_sc_hd__nor2_2
XFILLER_0_40_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2793_ _0231_ _0633_ _0634_ _0234_ _0635_ VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__a221o_2
X_2862_ _0684_ _0249_ _0687_ VGND VGND VPWR VPWR _0688_ sky130_fd_sc_hd__mux2_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1675_ _0963_ VGND VGND VPWR VPWR _0978_ sky130_fd_sc_hd__clkbuf_4
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2089_ _0875_ _0930_ _1266_ _1360_ _1361_ VGND VGND VPWR VPWR _1362_ sky130_fd_sc_hd__a2111o_1
X_2227_ _1498_ _1499_ _0960_ VGND VGND VPWR VPWR _1500_ sky130_fd_sc_hd__a21o_1
X_2158_ _1429_ _1430_ VGND VGND VPWR VPWR _1431_ sky130_fd_sc_hd__or2_2
XFILLER_0_23_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3130_ clknet_4_6_0_clk _0017_ net69 VGND VGND VPWR VPWR demux.state_machine.timeState\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_38_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2012_ demux.state_machine.timeState\[0\] _0896_ demux.state_machine.timeState\[4\]
+ VGND VGND VPWR VPWR _1285_ sky130_fd_sc_hd__or3_4
X_3061_ clknet_4_8_0_clk _0053_ net62 VGND VGND VPWR VPWR internalDataflow.accRegToDB\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_70_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2845_ _0677_ VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2914_ _0727_ _0728_ _0724_ VGND VGND VPWR VPWR _0729_ sky130_fd_sc_hd__a21oi_1
X_1727_ demux.state_machine.currentAddress\[11\] _1011_ _0979_ VGND VGND VPWR VPWR
+ _1020_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1658_ instructionLoader.interruptInjector.resetDetected net43 VGND VGND VPWR VPWR
+ _0962_ sky130_fd_sc_hd__nor2_2
X_2776_ _0129_ _0153_ _0176_ _0592_ _0536_ VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__a41o_1
XFILLER_0_13_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1589_ demux.state_machine.timeState\[2\] VGND VGND VPWR VPWR _0896_ sky130_fd_sc_hd__buf_2
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_58 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1512_ demux.state_machine.currentInstruction\[5\] VGND VGND VPWR VPWR _0819_ sky130_fd_sc_hd__buf_4
X_2630_ _0905_ _1441_ _0488_ _0490_ _0496_ VGND VGND VPWR VPWR _0497_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2492_ _0372_ _0373_ _0375_ VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__a21o_2
X_2561_ _0427_ _0432_ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__nor2_1
XFILLER_0_65_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3113_ clknet_4_5_0_clk _0105_ net69 VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3044_ clknet_4_0_0_clk _0036_ net57 VGND VGND VPWR VPWR internalDataflow.addressLowBusModule.busInputs\[26\]
+ sky130_fd_sc_hd__dfrtp_1
X_2828_ _1432_ _0632_ _0634_ _1321_ _0664_ VGND VGND VPWR VPWR _0665_ sky130_fd_sc_hd__a221o_2
XFILLER_0_41_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2759_ _0177_ _0604_ _0536_ VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__o21ai_2
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout62 net63 VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1992_ demux.state_machine.timeState\[6\] VGND VGND VPWR VPWR _1265_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_133 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2475_ _1474_ _0353_ _0354_ _0358_ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__or4_2
X_2613_ _0476_ _0477_ _0480_ VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__o21a_1
XFILLER_0_23_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2544_ _0288_ _0321_ _0369_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__or3_1
X_3027_ clknet_4_7_0_clk _0011_ net68 VGND VGND VPWR VPWR demux.state_machine.currentAddress\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2191_ _1001_ _0913_ _1462_ _1463_ VGND VGND VPWR VPWR _1464_ sky130_fd_sc_hd__a211o_1
X_2260_ _1257_ VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1975_ _0855_ _0860_ _0827_ VGND VGND VPWR VPWR _1248_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2458_ _0217_ _0333_ _0341_ _0343_ VGND VGND VPWR VPWR internalDataflow.psr.processStatusReg.stat_buf_nxt\[2\]
+ sky130_fd_sc_hd__a211o_1
X_2527_ _1452_ _1475_ _0354_ _0401_ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__or4_1
XFILLER_0_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold38 internalDataflow.stackBusModule.busInputs\[43\] VGND VGND VPWR VPWR net110
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_11_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold27 internalDataflow.stackBusModule.busInputs\[37\] VGND VGND VPWR VPWR net99
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 net35 VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__dlygate4sd3_1
Xhold49 net23 VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__dlygate4sd3_1
X_2389_ _1467_ _1479_ _0276_ VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1760_ _1045_ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__clkbuf_1
X_1691_ _0992_ VGND VGND VPWR VPWR _0993_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_52_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2312_ _0198_ _0199_ _0123_ VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__o21a_2
XFILLER_0_73_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2174_ _1273_ _0988_ _0945_ _1446_ VGND VGND VPWR VPWR _1447_ sky130_fd_sc_hd__a31o_1
X_2243_ _1465_ _0130_ VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__nor2_1
XFILLER_0_35_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput17 net17 VGND VGND VPWR VPWR addressBusHigh[1] sky130_fd_sc_hd__clkbuf_4
X_1889_ _1167_ _1170_ _1171_ VGND VGND VPWR VPWR _1172_ sky130_fd_sc_hd__or3_1
Xoutput28 net28 VGND VGND VPWR VPWR addressBusLow[4] sky130_fd_sc_hd__buf_2
X_1958_ _1235_ VGND VGND VPWR VPWR pulse_slower.nextEnableState\[1\] sky130_fd_sc_hd__clkbuf_1
Xoutput39 net39 VGND VGND VPWR VPWR dataBusOutput[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_3_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2861_ _0924_ _1362_ _0686_ _0332_ VGND VGND VPWR VPWR _0687_ sky130_fd_sc_hd__o31a_4
XFILLER_0_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2930_ _0557_ _0656_ VGND VGND VPWR VPWR _0744_ sky130_fd_sc_hd__nand2_1
X_1743_ net3 _0963_ _1010_ _1017_ VGND VGND VPWR VPWR _1032_ sky130_fd_sc_hd__and4_1
X_1674_ _0958_ _0966_ _0972_ _0977_ demux.state_machine.currentAddress\[6\] VGND VGND
+ VPWR VPWR _0009_ sky130_fd_sc_hd__a32o_1
X_1812_ _1094_ _0975_ _1069_ _1095_ VGND VGND VPWR VPWR _1096_ sky130_fd_sc_hd__a22o_1
X_2792_ _1430_ _0245_ _0246_ _0247_ _0632_ VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2226_ demux.state_machine.currentAddress\[5\] _0987_ _1384_ _1004_ VGND VGND VPWR
+ VPWR _1499_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_0_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2088_ demux.state_machine.timeState\[6\] _0891_ _1084_ VGND VGND VPWR VPWR _1361_
+ sky130_fd_sc_hd__and3_1
X_2157_ _1423_ _1418_ VGND VGND VPWR VPWR _1430_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_48_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_245 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3060_ clknet_4_8_0_clk _0052_ net62 VGND VGND VPWR VPWR internalDataflow.accRegToDB\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_10_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_56 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2011_ _0988_ demux.state_machine.currentAddress\[6\] _1283_ VGND VGND VPWR VPWR
+ _1284_ sky130_fd_sc_hd__o21a_1
XFILLER_0_70_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2844_ net128 _0274_ _0675_ VGND VGND VPWR VPWR _0677_ sky130_fd_sc_hd__mux2_1
X_2913_ _0537_ _0652_ VGND VGND VPWR VPWR _0728_ sky130_fd_sc_hd__or2_1
X_1726_ _0988_ _0977_ _1017_ _1019_ VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__a22o_1
X_1588_ demux.PSR_Z _0889_ _0892_ _0893_ _0894_ VGND VGND VPWR VPWR _0895_ sky130_fd_sc_hd__a2111oi_1
X_1657_ _0960_ VGND VGND VPWR VPWR _0961_ sky130_fd_sc_hd__buf_4
X_2775_ net120 _0555_ _0612_ _0544_ _0619_ VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__a221o_1
XFILLER_0_13_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2209_ _1257_ _1481_ _1322_ VGND VGND VPWR VPWR _1482_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_48_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1511_ _0817_ VGND VGND VPWR VPWR _0818_ sky130_fd_sc_hd__buf_4
X_2491_ _0371_ _0374_ VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__and2_2
XFILLER_0_10_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2560_ _0367_ _0425_ _0368_ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__mux2_1
XFILLER_0_65_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3112_ clknet_4_2_0_clk _0104_ net57 VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__dfrtp_1
X_3043_ clknet_4_0_0_clk _0035_ net57 VGND VGND VPWR VPWR internalDataflow.addressLowBusModule.busInputs\[25\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2758_ _0595_ VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__inv_2
XFILLER_0_5_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2827_ _1481_ _0654_ VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1709_ _1002_ _0981_ _1000_ _1008_ VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__a22o_1
X_2689_ demux.state_machine.currentAddress\[6\] demux.state_machine.currentAddress\[7\]
+ _0539_ _1273_ VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__o211a_1
XFILLER_0_41_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout63 net64 VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_19_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1991_ _0927_ _1143_ _1263_ VGND VGND VPWR VPWR _1264_ sky130_fd_sc_hd__o21a_1
X_2612_ _0315_ _0479_ _0407_ VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2474_ _1007_ _1249_ _1444_ _0356_ _0357_ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__a2111o_1
X_2543_ _0284_ _0410_ _0416_ _0406_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__a211o_1
X_3026_ clknet_4_7_0_clk _0010_ net68 VGND VGND VPWR VPWR demux.state_machine.currentAddress\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_46_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_91 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2190_ _1006_ _1102_ _1168_ _0983_ _1330_ VGND VGND VPWR VPWR _1463_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1974_ _1166_ _0910_ _1245_ _1246_ VGND VGND VPWR VPWR _1247_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2526_ _1121_ _1144_ _0873_ _1008_ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__o31a_1
XFILLER_0_46_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold17 negEdgeDetector.q1 VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__dlygate4sd3_1
Xhold39 net29 VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__dlygate4sd3_1
X_2457_ _1325_ _0342_ _0336_ instructionLoader.interruptInjector.processStatusRegIFlag
+ VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__o211a_1
X_2388_ _1257_ net44 _0266_ VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__a21oi_4
Xhold28 internalDataflow.stackBusModule.busInputs\[46\] VGND VGND VPWR VPWR net100
+ sky130_fd_sc_hd__dlygate4sd3_1
X_3009_ _0947_ _0996_ _0961_ VGND VGND VPWR VPWR _0803_ sky130_fd_sc_hd__a21o_1
XFILLER_0_34_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_69_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1690_ demux.state_machine.timeState\[0\] demux.state_machine.timeState\[4\] VGND
+ VGND VPWR VPWR _0992_ sky130_fd_sc_hd__and2b_1
XFILLER_0_52_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2242_ _0123_ _0129_ VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__and2_2
X_2311_ internalDataflow.addressLowBusModule.busInputs\[19\] _1502_ _0127_ _0957_
+ _0122_ VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__a221o_1
X_2173_ _1005_ demux.state_machine.currentAddress\[7\] _0993_ _0985_ VGND VGND VPWR
+ VPWR _1446_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1957_ pulse_slower.currentEnableState\[1\] net98 VGND VGND VPWR VPWR _1235_ sky130_fd_sc_hd__and2b_1
XFILLER_0_28_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1888_ _0880_ _0978_ _1047_ _1081_ VGND VGND VPWR VPWR _1171_ sky130_fd_sc_hd__a2bb2o_1
Xoutput29 net29 VGND VGND VPWR VPWR addressBusLow[5] sky130_fd_sc_hd__clkbuf_4
X_2509_ _0390_ _0391_ _0332_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__o21a_4
XFILLER_0_31_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput18 net18 VGND VGND VPWR VPWR addressBusHigh[2] sky130_fd_sc_hd__clkbuf_4
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1811_ _1012_ _0969_ net55 _0967_ VGND VGND VPWR VPWR _1095_ sky130_fd_sc_hd__and4bb_4
XFILLER_0_57_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2860_ _1008_ _1204_ _0685_ _0916_ VGND VGND VPWR VPWR _0686_ sky130_fd_sc_hd__a211o_1
XFILLER_0_43_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2791_ _1383_ _1386_ _1329_ VGND VGND VPWR VPWR _0634_ sky130_fd_sc_hd__and3_2
XFILLER_0_25_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1742_ net101 _0977_ _1031_ VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1673_ _0976_ VGND VGND VPWR VPWR _0977_ sky130_fd_sc_hd__clkbuf_4
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_25_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2225_ _1241_ _1290_ _1494_ _1497_ _1416_ VGND VGND VPWR VPWR _1498_ sky130_fd_sc_hd__o32ai_4
XFILLER_0_0_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2087_ _0896_ _0939_ _1084_ VGND VGND VPWR VPWR _1360_ sky130_fd_sc_hd__and3_1
X_2156_ _1425_ _1428_ VGND VGND VPWR VPWR _1429_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_390 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2989_ _0791_ VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_54_338 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2010_ _0993_ _1282_ VGND VGND VPWR VPWR _1283_ sky130_fd_sc_hd__and2b_1
XFILLER_0_54_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2912_ _0537_ _0652_ VGND VGND VPWR VPWR _0727_ sky130_fd_sc_hd__nand2_1
X_1725_ _1018_ VGND VGND VPWR VPWR _1019_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_53_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2774_ _0615_ _0617_ _0618_ VGND VGND VPWR VPWR _0619_ sky130_fd_sc_hd__o21a_1
X_2843_ _0676_ VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__inv_2
X_1587_ demux.PSR_V _0869_ _0852_ VGND VGND VPWR VPWR _0894_ sky130_fd_sc_hd__nor3_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1656_ _0959_ net42 _0951_ VGND VGND VPWR VPWR _0960_ sky130_fd_sc_hd__a21o_2
XFILLER_0_13_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2139_ demux.state_machine.timeState\[5\] _1079_ _1071_ _0879_ _1411_ VGND VGND VPWR
+ VPWR _1412_ sky130_fd_sc_hd__a221o_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2208_ _1372_ _1380_ VGND VGND VPWR VPWR _1481_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_360 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1510_ demux.state_machine.currentInstruction\[0\] demux.state_machine.currentInstruction\[2\]
+ demux.state_machine.currentInstruction\[3\] demux.state_machine.currentInstruction\[1\]
+ VGND VGND VPWR VPWR _0817_ sky130_fd_sc_hd__or4b_1
XFILLER_0_49_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2490_ _0158_ _0179_ _0370_ VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__or3_1
X_3042_ clknet_4_1_0_clk _0034_ net60 VGND VGND VPWR VPWR internalDataflow.addressLowBusModule.busInputs\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_3111_ clknet_4_0_0_clk _0103_ net57 VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1708_ _1007_ VGND VGND VPWR VPWR _1008_ sky130_fd_sc_hd__clkbuf_4
X_2688_ _1001_ _0933_ _1414_ VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_45_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2757_ _0601_ _0602_ VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__xnor2_1
X_2826_ _0663_ VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__clkbuf_1
X_1639_ _0926_ _0943_ _0944_ _0927_ _0945_ VGND VGND VPWR VPWR _0946_ sky130_fd_sc_hd__o41ai_2
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_36_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout64 net66 VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__buf_4
XFILLER_0_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_19_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1990_ _0932_ VGND VGND VPWR VPWR _1263_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2611_ _0378_ _0444_ _0437_ _0317_ _0478_ VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__o221a_1
X_2542_ _0216_ _0364_ _0412_ _0283_ _0415_ VGND VGND VPWR VPWR _0416_ sky130_fd_sc_hd__a221o_1
XFILLER_0_62_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2473_ _1273_ _1390_ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__nor2_1
X_3025_ clknet_4_7_0_clk _0009_ net68 VGND VGND VPWR VPWR demux.state_machine.currentAddress\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_46_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_168 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2809_ _0650_ VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1973_ _0847_ _0873_ _0877_ VGND VGND VPWR VPWR _1246_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_7_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2525_ _0400_ VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__clkbuf_1
Xhold29 demux.state_machine.currentAddress\[5\] VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__dlygate4sd3_1
Xhold18 instructionLoader.interruptInjector.irqGenerated VGND VGND VPWR VPWR net90
+ sky130_fd_sc_hd__dlygate4sd3_1
X_2456_ _1008_ _0846_ _0334_ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_39_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2387_ _1460_ _0274_ VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__and2_2
X_3008_ net94 _0801_ _0802_ _0385_ VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__a22o_1
XFILLER_0_19_400 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2172_ _1443_ _1444_ VGND VGND VPWR VPWR _1445_ sky130_fd_sc_hd__nor2_1
X_2241_ _0122_ _0126_ _0128_ VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__or3_2
X_2310_ internalDataflow.addressLowBusModule.busInputs\[35\] net46 _0125_ internalDataflow.addressLowBusModule.busInputs\[27\]
+ VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__a22o_1
X_1887_ _1168_ _0978_ _1169_ VGND VGND VPWR VPWR _1170_ sky130_fd_sc_hd__o21a_1
X_1956_ _1234_ VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2508_ _0910_ _1097_ _1002_ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__o21a_1
XFILLER_0_3_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput19 net19 VGND VGND VPWR VPWR addressBusHigh[3] sky130_fd_sc_hd__clkbuf_4
X_2439_ _1168_ _1094_ _0983_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__o21a_1
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_252 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap50 net51 VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_1
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1741_ _1026_ _1014_ _1024_ _0979_ VGND VGND VPWR VPWR _1031_ sky130_fd_sc_hd__o211a_1
X_1810_ _0871_ _0861_ VGND VGND VPWR VPWR _1094_ sky130_fd_sc_hd__nor2_2
XFILLER_0_25_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2790_ _1326_ _0632_ VGND VGND VPWR VPWR _0633_ sky130_fd_sc_hd__nor2_2
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1672_ _0975_ VGND VGND VPWR VPWR _0976_ sky130_fd_sc_hd__buf_2
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2224_ _0991_ _0993_ _1495_ _1496_ VGND VGND VPWR VPWR _1497_ sky130_fd_sc_hd__a211o_1
X_2155_ _1245_ _1426_ _1427_ VGND VGND VPWR VPWR _1428_ sky130_fd_sc_hd__and3_1
XFILLER_0_63_306 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2086_ _0915_ _1357_ _1249_ _1358_ _0876_ VGND VGND VPWR VPWR _1359_ sky130_fd_sc_hd__o41a_1
XFILLER_0_33_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1939_ _1056_ _1070_ _1098_ _1109_ VGND VGND VPWR VPWR _1219_ sky130_fd_sc_hd__or4_1
X_2988_ net87 _0308_ _0783_ VGND VGND VPWR VPWR _0791_ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2911_ net130 _0555_ _0720_ _0721_ _0726_ VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__a221o_1
X_1724_ net3 _0978_ _1010_ net2 VGND VGND VPWR VPWR _1018_ sky130_fd_sc_hd__and4b_1
XFILLER_0_53_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2773_ _0615_ _0617_ _0546_ VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_13_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2842_ _0224_ _0249_ _0675_ VGND VGND VPWR VPWR _0676_ sky130_fd_sc_hd__mux2_1
X_1586_ demux.PSR_C _0869_ _0825_ VGND VGND VPWR VPWR _0893_ sky130_fd_sc_hd__nor3_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1655_ _0950_ VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__inv_2
XFILLER_0_0_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2138_ _0912_ _1168_ demux.state_machine.timeState\[1\] VGND VGND VPWR VPWR _1411_
+ sky130_fd_sc_hd__o21a_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2207_ _1479_ VGND VGND VPWR VPWR _1480_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2069_ net135 _1341_ VGND VGND VPWR VPWR _1342_ sky130_fd_sc_hd__or2b_1
XFILLER_0_21_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3110_ clknet_4_11_0_clk _0102_ net66 VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3041_ clknet_4_4_0_clk pulse_slower.nextEnableState\[1\] net60 VGND VGND VPWR VPWR
+ pulse_slower.currentEnableState\[1\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2825_ net115 _0662_ _0645_ VGND VGND VPWR VPWR _0663_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1638_ _0896_ demux.state_machine.timeState\[4\] VGND VGND VPWR VPWR _0945_ sky130_fd_sc_hd__or2_2
XFILLER_0_41_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1707_ _1006_ VGND VGND VPWR VPWR _1007_ sky130_fd_sc_hd__clkbuf_4
X_2687_ _0522_ _0537_ VGND VGND VPWR VPWR _0538_ sky130_fd_sc_hd__nor2_2
X_2756_ _0587_ _0589_ _0585_ VGND VGND VPWR VPWR _0602_ sky130_fd_sc_hd__a21o_1
X_1569_ _0875_ VGND VGND VPWR VPWR _0876_ sky130_fd_sc_hd__clkbuf_4
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xfanout65 net66 VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__buf_4
XFILLER_0_17_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2472_ _1071_ _1285_ _1409_ _1102_ _0355_ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__a221o_1
X_2610_ _0259_ _0364_ VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2541_ _0275_ _0282_ _0408_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__o21a_1
XFILLER_0_55_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3024_ clknet_4_7_0_clk _0008_ net67 VGND VGND VPWR VPWR demux.state_machine.currentAddress\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_46_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2808_ net17 _0649_ _0645_ VGND VGND VPWR VPWR _0650_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2739_ internalDataflow.addressLowBusModule.busInputs\[20\] _0535_ VGND VGND VPWR
+ VPWR _0586_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1972_ _1003_ _0913_ VGND VGND VPWR VPWR _1245_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2455_ _0981_ _0340_ VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__nor2_1
X_2524_ net131 _0305_ _0392_ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold19 net19 VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__dlygate4sd3_1
X_2386_ _1326_ _0266_ _0271_ _0273_ VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_46_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3007_ _0968_ internalDataflow.addressLowBusModule.busInputs\[23\] _0905_ _0323_
+ VGND VGND VPWR VPWR _0802_ sky130_fd_sc_hd__and4_1
XFILLER_0_19_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2171_ _1005_ _0910_ _1384_ VGND VGND VPWR VPWR _1444_ sky130_fd_sc_hd__a21o_1
X_2240_ internalDataflow.addressLowBusModule.busInputs\[22\] _1502_ _0127_ net8 VGND
+ VGND VPWR VPWR _0128_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1886_ _0964_ _1017_ _1087_ _0975_ VGND VGND VPWR VPWR _1169_ sky130_fd_sc_hd__a31o_1
X_1955_ _1225_ _1226_ _1231_ _1233_ VGND VGND VPWR VPWR _1234_ sky130_fd_sc_hd__or4_1
XFILLER_0_31_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2507_ _0831_ _1108_ _1008_ VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__o21a_1
XFILLER_0_51_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2438_ _0866_ _0844_ _0324_ _0325_ demux.PSR_V VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__o311a_1
XFILLER_0_11_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2369_ _0868_ _1143_ _0256_ demux.PSR_C _1006_ VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__o311a_1
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1671_ _0974_ VGND VGND VPWR VPWR _0975_ sky130_fd_sc_hd__buf_2
X_1740_ _0987_ _0977_ _1019_ _1030_ VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_128 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2223_ _1273_ demux.state_machine.currentAddress\[1\] _0945_ _0993_ _0985_ VGND VGND
+ VPWR VPWR _1496_ sky130_fd_sc_hd__a32o_1
X_2085_ _0943_ _1166_ VGND VGND VPWR VPWR _1358_ sky130_fd_sc_hd__or2_2
X_2154_ _1259_ _1079_ _1003_ VGND VGND VPWR VPWR _1427_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_63_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2987_ _0790_ VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_33_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1938_ _1120_ _1141_ _1167_ _1196_ VGND VGND VPWR VPWR _1218_ sky130_fd_sc_hd__or4_1
X_1869_ _0821_ _0860_ VGND VGND VPWR VPWR _1152_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2841_ _0674_ VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2910_ _0553_ _0725_ VGND VGND VPWR VPWR _0726_ sky130_fd_sc_hd__nor2_1
X_1723_ _0954_ _1016_ _0956_ VGND VGND VPWR VPWR _1017_ sky130_fd_sc_hd__o21ai_4
X_1654_ net13 VGND VGND VPWR VPWR _0959_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2772_ _0587_ _0589_ _0599_ _0616_ _0585_ VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__a311o_1
X_1585_ demux.PSR_V _0890_ _0891_ VGND VGND VPWR VPWR _0892_ sky130_fd_sc_hd__and3_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2206_ _1470_ _1472_ _1475_ _1476_ _1478_ VGND VGND VPWR VPWR _1479_ sky130_fd_sc_hd__o41a_2
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2137_ _0899_ _1409_ _0905_ VGND VGND VPWR VPWR _1410_ sky130_fd_sc_hd__o21ai_2
X_2068_ _0959_ net42 net51 _1241_ _0951_ VGND VGND VPWR VPWR _1341_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_14_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3040_ clknet_4_4_0_clk pulse_slower.nextEnableState\[0\] net60 VGND VGND VPWR VPWR
+ pulse_slower.currentEnableState\[0\] sky130_fd_sc_hd__dfrtp_1
X_2824_ _0141_ _0632_ _0633_ _0140_ _0661_ VGND VGND VPWR VPWR _0662_ sky130_fd_sc_hd__a221o_2
X_1637_ _0827_ _0855_ VGND VGND VPWR VPWR _0944_ sky130_fd_sc_hd__nor2_2
XFILLER_0_53_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1706_ _1005_ VGND VGND VPWR VPWR _1006_ sky130_fd_sc_hd__buf_2
XFILLER_0_30_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2686_ _0536_ VGND VGND VPWR VPWR _0537_ sky130_fd_sc_hd__inv_2
X_2755_ _0599_ _0600_ VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__nand2_1
X_1568_ demux.state_machine.timeState\[4\] VGND VGND VPWR VPWR _0875_ sky130_fd_sc_hd__clkbuf_4
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_207 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout66 net12 VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_32_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_387 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2471_ _0847_ _0868_ _1006_ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__o21a_1
XFILLER_0_23_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2540_ net80 _0403_ _0405_ _0406_ _0414_ VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__a221o_1
X_3023_ clknet_4_6_0_clk _0007_ net67 VGND VGND VPWR VPWR demux.state_machine.currentAddress\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_73_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2807_ _0647_ _0633_ _0634_ _0265_ _0648_ VGND VGND VPWR VPWR _0649_ sky130_fd_sc_hd__a221o_2
X_2738_ internalDataflow.addressLowBusModule.busInputs\[20\] _0535_ VGND VGND VPWR
+ VPWR _0585_ sky130_fd_sc_hd__and2_1
X_2669_ _0939_ _0940_ VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__nand2_1
XFILLER_0_41_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1971_ _1243_ VGND VGND VPWR VPWR _1244_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_55_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2454_ _0982_ _0334_ VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__nand2_1
X_2385_ net47 _1431_ _0272_ _1329_ VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__a31o_1
X_2523_ _0399_ VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__clkbuf_1
Xinput1 dataBusEnable VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_1
X_3006_ _0905_ _0323_ VGND VGND VPWR VPWR _0801_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2170_ _1005_ _1102_ _1267_ _1442_ VGND VGND VPWR VPWR _1443_ sky130_fd_sc_hd__a211o_1
X_1954_ _1154_ _1176_ _1205_ _1232_ VGND VGND VPWR VPWR _1233_ sky130_fd_sc_hd__or4_1
XFILLER_0_28_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1885_ _0829_ _0865_ VGND VGND VPWR VPWR _1168_ sky130_fd_sc_hd__nor2_4
XFILLER_0_43_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2368_ _1121_ _1200_ _0853_ _1174_ VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__or4_1
XFILLER_0_47_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2437_ _1325_ _0319_ VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__or2_2
XFILLER_0_11_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2506_ internalDataflow.stackBusModule.busInputs\[32\] VGND VGND VPWR VPWR _0389_
+ sky130_fd_sc_hd__inv_2
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2299_ _1382_ _1329_ _1387_ VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__a21o_1
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap52 net53 VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__buf_1
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1670_ _0973_ VGND VGND VPWR VPWR _0974_ sky130_fd_sc_hd__buf_2
XFILLER_0_25_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2222_ _1273_ demux.state_machine.currentAddress\[12\] _1491_ VGND VGND VPWR VPWR
+ _1495_ sky130_fd_sc_hd__and3_1
XFILLER_0_0_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2153_ _1102_ _0930_ _1001_ VGND VGND VPWR VPWR _1426_ sky130_fd_sc_hd__o21ai_1
X_2084_ _0847_ _0873_ VGND VGND VPWR VPWR _1357_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1937_ _1078_ _1129_ VGND VGND VPWR VPWR _1217_ sky130_fd_sc_hd__or2_1
X_2986_ net38 _1482_ _0783_ VGND VGND VPWR VPWR _0790_ sky130_fd_sc_hd__mux2_1
X_1868_ _0999_ _1041_ VGND VGND VPWR VPWR _1151_ sky130_fd_sc_hd__and2_1
X_1799_ _1079_ _0978_ _1082_ VGND VGND VPWR VPWR _1083_ sky130_fd_sc_hd__o21a_1
XFILLER_0_62_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2840_ _0332_ _0673_ VGND VGND VPWR VPWR _0674_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2771_ internalDataflow.addressLowBusModule.busInputs\[21\] _0535_ VGND VGND VPWR
+ VPWR _0616_ sky130_fd_sc_hd__and2_1
X_1653_ _0954_ _0956_ net4 _0957_ VGND VGND VPWR VPWR _0958_ sky130_fd_sc_hd__and4b_2
X_1722_ net4 _0957_ VGND VGND VPWR VPWR _1016_ sky130_fd_sc_hd__or2_2
X_1584_ _0819_ _0820_ VGND VGND VPWR VPWR _0891_ sky130_fd_sc_hd__nor2_4
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2205_ _0998_ _1477_ VGND VGND VPWR VPWR _1478_ sky130_fd_sc_hd__and2_2
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2136_ _1004_ _0877_ _0879_ VGND VGND VPWR VPWR _1409_ sky130_fd_sc_hd__or3_1
X_2067_ _1336_ _1337_ _1338_ _1339_ VGND VGND VPWR VPWR _1340_ sky130_fd_sc_hd__nor4_1
X_2969_ _1297_ _1254_ VGND VGND VPWR VPWR _0779_ sky130_fd_sc_hd__or2b_1
XFILLER_0_29_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_300 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1705_ _1004_ VGND VGND VPWR VPWR _1005_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2823_ _0145_ _0634_ VGND VGND VPWR VPWR _0661_ sky130_fd_sc_hd__and2_1
X_2754_ internalDataflow.addressLowBusModule.busInputs\[21\] _0558_ VGND VGND VPWR
+ VPWR _0600_ sky130_fd_sc_hd__nand2_1
X_1567_ _0868_ _0870_ _0872_ _0873_ VGND VGND VPWR VPWR _0874_ sky130_fd_sc_hd__or4_1
X_1636_ _0827_ _0885_ VGND VGND VPWR VPWR _0943_ sky130_fd_sc_hd__nor2_1
X_2685_ _0535_ VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__clkbuf_4
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_219 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2119_ _0875_ _0911_ _1389_ _1391_ _0934_ VGND VGND VPWR VPWR _1392_ sky130_fd_sc_hd__a2111o_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout67 net72 VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_4
X_3099_ clknet_4_13_0_clk _0091_ net66 VGND VGND VPWR VPWR internalDataflow.addressHighBusModule.busInputs\[16\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_17_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2470_ _1168_ _1441_ _1330_ _1267_ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__a211o_1
X_3022_ clknet_4_7_0_clk _0006_ net67 VGND VGND VPWR VPWR demux.state_machine.currentAddress\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2806_ _1431_ _0272_ _0632_ VGND VGND VPWR VPWR _0648_ sky130_fd_sc_hd__and3_1
X_2668_ _0519_ VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__clkbuf_1
X_2737_ _0584_ VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__clkbuf_1
X_1619_ _0885_ _0844_ _0882_ _0830_ VGND VGND VPWR VPWR _0926_ sky130_fd_sc_hd__a31oi_2
X_2599_ _0465_ _0466_ _0383_ _0467_ _0376_ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__o2111a_1
XFILLER_0_5_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_288 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1970_ demux.state_machine.timeState\[0\] demux.state_machine.timeState\[4\] VGND
+ VGND VPWR VPWR _1243_ sky130_fd_sc_hd__or2_1
XFILLER_0_55_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2522_ net109 _1434_ _0392_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_119 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2453_ _0196_ _0333_ _0339_ VGND VGND VPWR VPWR internalDataflow.psr.processStatusReg.stat_buf_nxt\[3\]
+ sky130_fd_sc_hd__a21o_1
X_2384_ internalDataflow.addressHighBusModule.busInputs\[17\] _1422_ _1424_ net3 VGND
+ VGND VPWR VPWR _0272_ sky130_fd_sc_hd__o22a_1
Xinput2 dataBusInput[0] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_4
X_3005_ _0800_ VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1884_ _1166_ _1067_ _1069_ _1113_ VGND VGND VPWR VPWR _1167_ sky130_fd_sc_hd__a22o_1
X_1953_ _1072_ _1096_ _1101_ _1124_ VGND VGND VPWR VPWR _1232_ sky130_fd_sc_hd__or4_1
XFILLER_0_43_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2505_ _0236_ _0333_ _0352_ _0385_ _0388_ VGND VGND VPWR VPWR internalDataflow.psr.processStatusReg.stat_buf_nxt\[0\]
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_11_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2436_ _0323_ VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__inv_2
X_2367_ _0254_ _1274_ _1440_ VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__or3b_1
XFILLER_0_37_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2298_ _1257_ _0185_ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__nor2_1
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_372 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2221_ _1491_ _0913_ _0930_ _0876_ _1493_ VGND VGND VPWR VPWR _1494_ sky130_fd_sc_hd__a221o_1
X_2152_ _1267_ _1361_ _1303_ VGND VGND VPWR VPWR _1425_ sky130_fd_sc_hd__o21a_1
X_2083_ _0897_ _0904_ _1352_ _1355_ VGND VGND VPWR VPWR _1356_ sky130_fd_sc_hd__a31o_1
XFILLER_0_17_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1936_ _1048_ _1087_ _1177_ _1191_ _1215_ VGND VGND VPWR VPWR _1216_ sky130_fd_sc_hd__a2111o_1
X_1867_ _0830_ _0860_ VGND VGND VPWR VPWR _1150_ sky130_fd_sc_hd__nor2_4
XFILLER_0_31_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2985_ _0789_ VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__clkbuf_1
X_1798_ _0964_ _1017_ _1081_ _1066_ VGND VGND VPWR VPWR _1082_ sky130_fd_sc_hd__a31o_1
XFILLER_0_3_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2419_ _1257_ _0304_ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1721_ net85 _0977_ _1011_ _1015_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2770_ _0613_ _0614_ VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1652_ net5 VGND VGND VPWR VPWR _0957_ sky130_fd_sc_hd__clkbuf_4
X_1583_ _0832_ _0833_ _0834_ _0835_ VGND VGND VPWR VPWR _0890_ sky130_fd_sc_hd__and4b_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2204_ demux.state_machine.currentAddress\[6\] _1283_ _1285_ _0988_ _1287_ VGND VGND
+ VPWR VPWR _1477_ sky130_fd_sc_hd__a221o_1
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2135_ _0873_ _1244_ VGND VGND VPWR VPWR _1408_ sky130_fd_sc_hd__nand2_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2066_ _0847_ _0856_ _1202_ _1237_ _1263_ VGND VGND VPWR VPWR _1339_ sky130_fd_sc_hd__o41a_1
XFILLER_0_29_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1919_ _0871_ _0882_ VGND VGND VPWR VPWR _1200_ sky130_fd_sc_hd__nor2_1
XFILLER_0_56_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2899_ _0708_ _0715_ _0553_ VGND VGND VPWR VPWR _0716_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2968_ _0778_ VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_54_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_45_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2822_ _0660_ VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1704_ _1003_ VGND VGND VPWR VPWR _1004_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2684_ _0534_ VGND VGND VPWR VPWR _0535_ sky130_fd_sc_hd__buf_2
XFILLER_0_5_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2753_ internalDataflow.addressLowBusModule.busInputs\[21\] _0535_ VGND VGND VPWR
+ VPWR _0599_ sky130_fd_sc_hd__or2_1
X_1635_ _0912_ _0936_ _0920_ _0938_ _0941_ VGND VGND VPWR VPWR _0942_ sky130_fd_sc_hd__a221oi_2
X_1566_ _0869_ _0861_ VGND VGND VPWR VPWR _0873_ sky130_fd_sc_hd__nor2_4
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_60 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2118_ _0937_ _1390_ VGND VGND VPWR VPWR _1391_ sky130_fd_sc_hd__nor2_1
X_3098_ clknet_4_2_0_clk _0090_ net58 VGND VGND VPWR VPWR internalDataflow.addressLowBusModule.busInputs\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2049_ _1257_ _1321_ VGND VGND VPWR VPWR _1322_ sky130_fd_sc_hd__nor2_1
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xfanout68 net72 VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__buf_2
XFILLER_0_71_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xfanout57 net61 VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_32_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3021_ clknet_4_7_0_clk _0005_ net68 VGND VGND VPWR VPWR demux.state_machine.currentAddress\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_25_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_74 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2805_ net44 VGND VGND VPWR VPWR _0647_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_106 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1618_ _0914_ _0919_ _0922_ _0924_ VGND VGND VPWR VPWR _0925_ sky130_fd_sc_hd__or4_1
X_2667_ internalDataflow.accRegToDB\[7\] _0305_ _0511_ VGND VGND VPWR VPWR _0519_
+ sky130_fd_sc_hd__mux2_1
X_2736_ _0583_ internalDataflow.addressLowBusModule.busInputs\[19\] _0554_ VGND VGND
+ VPWR VPWR _0584_ sky130_fd_sc_hd__mux2_1
X_1549_ _0855_ _0825_ _0821_ VGND VGND VPWR VPWR _0856_ sky130_fd_sc_hd__a21oi_1
X_2598_ _1466_ _0325_ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2521_ _0398_ VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__clkbuf_1
X_2452_ _0335_ _0337_ _0338_ VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__mux2_1
X_2383_ _0187_ _0270_ VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__nor2_1
X_3004_ _0385_ net118 _0799_ VGND VGND VPWR VPWR _0800_ sky130_fd_sc_hd__mux2_1
Xinput3 dataBusInput[1] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_4
XFILLER_0_61_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2719_ internalDataflow.addressLowBusModule.busInputs\[18\] _0535_ VGND VGND VPWR
+ VPWR _0568_ sky130_fd_sc_hd__xor2_1
XFILLER_0_10_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_256 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1952_ _1050_ _1227_ _1230_ VGND VGND VPWR VPWR _1231_ sky130_fd_sc_hd__or3_1
X_1883_ _0866_ _0865_ VGND VGND VPWR VPWR _1166_ sky130_fd_sc_hd__nor2_1
XFILLER_0_43_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_212 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2435_ _1273_ _1325_ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__nor2_4
X_2504_ _0335_ _0386_ _0387_ VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2366_ _1071_ _1244_ _1285_ _1168_ _1444_ VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__a221o_1
XFILLER_0_2_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2297_ internalDataflow.addressLowBusModule.busInputs\[19\] _1315_ _0183_ _0184_
+ net48 VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_66_329 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap54 _0989_ VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__buf_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_65_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2220_ _0897_ _0912_ _1168_ demux.state_machine.timeState\[1\] _1492_ VGND VGND VPWR
+ VPWR _1493_ sky130_fd_sc_hd__a221o_1
X_2082_ _0876_ _1353_ _1354_ _0918_ _0916_ VGND VGND VPWR VPWR _1355_ sky130_fd_sc_hd__a2111o_1
X_2151_ _1423_ _1418_ VGND VGND VPWR VPWR _1424_ sky130_fd_sc_hd__nand2_2
XFILLER_0_48_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2984_ net117 _0149_ _0783_ VGND VGND VPWR VPWR _0789_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_343 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1797_ _0967_ _1010_ _1080_ VGND VGND VPWR VPWR _1081_ sky130_fd_sc_hd__a21boi_4
X_1866_ _1149_ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__clkbuf_1
X_1935_ _1214_ _0976_ _1019_ _1059_ VGND VGND VPWR VPWR _1215_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2418_ _1460_ _0305_ VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__nand2_1
X_2349_ _1467_ _1479_ _0236_ VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1651_ net55 VGND VGND VPWR VPWR _0956_ sky130_fd_sc_hd__clkbuf_4
X_1720_ net3 _0979_ _1014_ VGND VGND VPWR VPWR _1015_ sky130_fd_sc_hd__and3_1
XFILLER_0_5_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1582_ _0869_ _0860_ VGND VGND VPWR VPWR _0889_ sky130_fd_sc_hd__nor2_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2134_ _1403_ _1405_ _1406_ VGND VGND VPWR VPWR _1407_ sky130_fd_sc_hd__and3b_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2203_ _1384_ _1266_ _1267_ _1306_ VGND VGND VPWR VPWR _1476_ sky130_fd_sc_hd__or4_1
X_2065_ _0868_ _1143_ _1131_ _1271_ _1263_ VGND VGND VPWR VPWR _1338_ sky130_fd_sc_hd__o41a_1
XFILLER_0_28_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2967_ _0777_ internalDataflow.addressHighBusModule.busInputs\[23\] _0554_ VGND VGND
+ VPWR VPWR _0778_ sky130_fd_sc_hd__mux2_1
XFILLER_0_69_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1849_ _0967_ _0969_ _1013_ VGND VGND VPWR VPWR _1133_ sky130_fd_sc_hd__or3_2
X_1918_ _1199_ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__clkbuf_1
X_2898_ _0713_ _0714_ VGND VGND VPWR VPWR _0715_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2821_ net127 _0659_ _0645_ VGND VGND VPWR VPWR _0660_ sky130_fd_sc_hd__mux2_1
X_1703_ _0932_ VGND VGND VPWR VPWR _1003_ sky130_fd_sc_hd__buf_4
X_1634_ _0832_ _0939_ _0940_ demux.state_machine.timeState\[4\] VGND VGND VPWR VPWR
+ _0941_ sky130_fd_sc_hd__and4b_2
XFILLER_0_41_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2683_ _0521_ _0533_ VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2752_ _0590_ _0591_ _0598_ VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__o21ai_1
X_1565_ _0871_ _0818_ VGND VGND VPWR VPWR _0872_ sky130_fd_sc_hd__nor2_1
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2117_ _0882_ _0861_ _0830_ VGND VGND VPWR VPWR _1390_ sky130_fd_sc_hd__a21o_1
X_3097_ clknet_4_0_0_clk _0089_ net59 VGND VGND VPWR VPWR internalDataflow.addressLowBusModule.busInputs\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2048_ internalDataflow.addressHighBusModule.busInputs\[22\] _1294_ net134 _1320_
+ VGND VGND VPWR VPWR _1321_ sky130_fd_sc_hd__a211o_1
Xfanout69 net72 VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__clkbuf_4
Xfanout58 net59 VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_55_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3020_ clknet_4_6_0_clk _0004_ net67 VGND VGND VPWR VPWR demux.state_machine.currentAddress\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_25_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2804_ _0646_ VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__clkbuf_1
X_1617_ _0897_ _0923_ VGND VGND VPWR VPWR _0924_ sky130_fd_sc_hd__and2_1
X_2597_ _0378_ _0372_ _0134_ VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__and3b_1
XFILLER_0_26_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2666_ _0518_ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__clkbuf_1
X_2735_ _0544_ _0575_ _0581_ _0582_ VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__a22o_1
X_1548_ _0854_ VGND VGND VPWR VPWR _0855_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_74 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2451_ _0842_ _0908_ _0323_ VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_23_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_66 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_99 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2520_ net99 _0146_ _0392_ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__mux2_1
Xinput4 dataBusInput[2] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_4
X_3003_ _0529_ _1437_ _0961_ _1281_ VGND VGND VPWR VPWR _0799_ sky130_fd_sc_hd__a211o_1
X_2382_ _1375_ _0267_ _0268_ _0269_ _1372_ VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__o41ai_2
XFILLER_0_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2718_ _0221_ _0566_ VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__xor2_1
XFILLER_0_6_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2649_ _0508_ VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1882_ _1140_ _1162_ _1163_ _1164_ VGND VGND VPWR VPWR _1165_ sky130_fd_sc_hd__or4_1
X_1951_ _0831_ _0977_ _0966_ _1229_ _1170_ VGND VGND VPWR VPWR _1230_ sky130_fd_sc_hd__a221o_1
XFILLER_0_43_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2503_ _0907_ _0921_ _0323_ VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_51_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2434_ net14 VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__inv_2
X_2365_ _1006_ _0987_ free_carry_ff.freeCarry _0252_ _1364_ VGND VGND VPWR VPWR _0253_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2296_ internalDataflow.addressHighBusModule.busInputs\[19\] _1294_ _1314_ net5 VGND
+ VGND VPWR VPWR _0184_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xmax_cap44 _0270_ VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__clkbuf_2
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_33_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2081_ demux.state_machine.timeState\[4\] demux.state_machine.timeState\[6\] demux.state_machine.timeState\[1\]
+ _1051_ _0890_ VGND VGND VPWR VPWR _1354_ sky130_fd_sc_hd__o311a_1
X_2150_ _1407_ _1408_ _1410_ _1421_ VGND VGND VPWR VPWR _1423_ sky130_fd_sc_hd__a31o_1
X_1934_ _0816_ _1076_ VGND VGND VPWR VPWR _1214_ sky130_fd_sc_hd__nor2_1
X_2983_ _0788_ VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1796_ _1012_ _0969_ _1010_ VGND VGND VPWR VPWR _1080_ sky130_fd_sc_hd__o21ai_1
X_1865_ _1100_ _1111_ _1148_ VGND VGND VPWR VPWR _1149_ sky130_fd_sc_hd__or3_1
XFILLER_0_12_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2417_ _0301_ _0304_ _1329_ VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__mux2_4
X_2348_ _0148_ _0231_ _0235_ VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__o21a_2
X_2279_ internalDataflow.addressLowBusModule.busInputs\[20\] _1315_ _0166_ _1318_
+ VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1581_ demux.PSR_N _0880_ _0883_ _0886_ _0887_ VGND VGND VPWR VPWR _0888_ sky130_fd_sc_hd__o2111a_2
X_1650_ demux.nmi instructionLoader.interruptInjector.resetDetected instructionLoader.interruptInjector.irqGenerated
+ VGND VGND VPWR VPWR _0955_ sky130_fd_sc_hd__nor3_1
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2202_ _1006_ _1358_ _1473_ _1474_ VGND VGND VPWR VPWR _1475_ sky130_fd_sc_hd__a211o_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2133_ _0937_ _0928_ VGND VGND VPWR VPWR _1406_ sky130_fd_sc_hd__or2_1
XFILLER_0_48_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2064_ _1152_ _0913_ _1094_ _1263_ VGND VGND VPWR VPWR _1337_ sky130_fd_sc_hd__o31a_1
XFILLER_0_71_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1917_ _1111_ _1160_ _1188_ _1198_ VGND VGND VPWR VPWR _1199_ sky130_fd_sc_hd__or4_1
XFILLER_0_44_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2897_ _0709_ _0700_ _0712_ VGND VGND VPWR VPWR _0714_ sky130_fd_sc_hd__and3_1
X_2966_ _0772_ _0776_ _0553_ VGND VGND VPWR VPWR _0777_ sky130_fd_sc_hd__mux2_1
X_1779_ _1062_ VGND VGND VPWR VPWR _1063_ sky130_fd_sc_hd__buf_2
X_1848_ _1131_ _0974_ _1018_ _1081_ VGND VGND VPWR VPWR _1132_ sky130_fd_sc_hd__a22o_1
XFILLER_0_8_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_62_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2820_ _0169_ _0634_ _0658_ VGND VGND VPWR VPWR _0659_ sky130_fd_sc_hd__a21o_2
X_2751_ internalDataflow.addressLowBusModule.busInputs\[20\] _0555_ _0597_ _0553_
+ VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__o2bb2a_1
X_1564_ _0830_ VGND VGND VPWR VPWR _0871_ sky130_fd_sc_hd__buf_4
X_1633_ _0835_ _0834_ VGND VGND VPWR VPWR _0940_ sky130_fd_sc_hd__and2b_1
X_2682_ _0483_ _0524_ _0528_ _0532_ VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__o31a_2
X_1702_ _1001_ VGND VGND VPWR VPWR _1002_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_26_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2116_ _0912_ _1168_ demux.state_machine.timeState\[5\] VGND VGND VPWR VPWR _1389_
+ sky130_fd_sc_hd__o21a_1
X_2047_ net8 _1314_ _1315_ internalDataflow.addressLowBusModule.busInputs\[22\] _1319_
+ VGND VGND VPWR VPWR _1320_ sky130_fd_sc_hd__a221o_1
X_3096_ clknet_4_3_0_clk _0088_ net59 VGND VGND VPWR VPWR internalDataflow.addressLowBusModule.busInputs\[37\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_44_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2949_ _0759_ _0760_ VGND VGND VPWR VPWR _0761_ sky130_fd_sc_hd__and2_1
Xfanout59 net61 VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_55_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_203 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2803_ net102 _0636_ _0645_ VGND VGND VPWR VPWR _0646_ sky130_fd_sc_hd__mux2_1
X_2734_ _0576_ _0577_ _0580_ _0553_ VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__o31a_1
X_1616_ _0871_ _0855_ VGND VGND VPWR VPWR _0923_ sky130_fd_sc_hd__nor2_1
X_1547_ demux.state_machine.currentInstruction\[1\] _0811_ _0810_ _0813_ VGND VGND
+ VPWR VPWR _0854_ sky130_fd_sc_hd__or4bb_1
X_2596_ _0134_ _0372_ _0378_ VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_1_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2665_ internalDataflow.accRegToDB\[6\] _1434_ _0511_ VGND VGND VPWR VPWR _0518_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3148_ clknet_4_1_0_clk VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__buf_2
XFILLER_0_5_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3079_ clknet_4_10_0_clk _0071_ net64 VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_20_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2450_ internalDataflow.dataBusModule.busInputs\[43\] _0336_ VGND VGND VPWR VPWR
+ _0337_ sky130_fd_sc_hd__and2_1
X_2381_ internalDataflow.addressLowBusModule.busInputs\[25\] _1377_ _1378_ internalDataflow.addressLowBusModule.busInputs\[33\]
+ VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__a22o_1
XFILLER_0_11_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput5 dataBusInput[3] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_2
X_3002_ _0798_ VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2717_ _0559_ _0561_ _0562_ _0537_ VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__o22a_1
XFILLER_0_14_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2648_ net31 _0312_ _0502_ VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2579_ _0321_ _0370_ _0441_ _0449_ VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__o31ai_1
XFILLER_0_73_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1950_ _1055_ _1181_ _1228_ VGND VGND VPWR VPWR _1229_ sky130_fd_sc_hd__a21o_1
X_1881_ _0889_ _1091_ _1047_ _1113_ VGND VGND VPWR VPWR _1164_ sky130_fd_sc_hd__a22o_1
X_2502_ _0352_ demux.PSR_C _0336_ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__and3b_1
XFILLER_0_47_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2364_ _0983_ _0917_ _0987_ _0993_ _0985_ VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__a32o_1
X_2433_ internalDataflow.dataBusModule.busInputs\[43\] _0320_ VGND VGND VPWR VPWR
+ _0321_ sky130_fd_sc_hd__nand2_2
XFILLER_0_66_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2295_ internalDataflow.accRegToDB\[3\] _1316_ _1318_ internalDataflow.dataBusModule.busInputs\[43\]
+ VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__a22o_1
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_69_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap56 _0947_ VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__buf_1
XFILLER_0_68_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_4_9_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_9_0_clk sky130_fd_sc_hd__clkbuf_8
X_2080_ _1051_ _1084_ _1122_ _0939_ VGND VGND VPWR VPWR _1353_ sky130_fd_sc_hd__a22o_1
X_1933_ _1213_ VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2982_ net116 _0172_ _0783_ VGND VGND VPWR VPWR _0788_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1864_ _1126_ _1130_ _1147_ VGND VGND VPWR VPWR _1148_ sky130_fd_sc_hd__or3_1
X_1795_ _0920_ VGND VGND VPWR VPWR _1079_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2278_ _0983_ _1079_ _0165_ _1260_ VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__a31o_1
XFILLER_0_35_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2416_ internalDataflow.addressLowBusModule.busInputs\[23\] _1315_ _0303_ net48 VGND
+ VGND VPWR VPWR _0304_ sky130_fd_sc_hd__a211o_1
X_2347_ _1256_ _0234_ VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__or2_1
XFILLER_0_62_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1580_ _0819_ _0855_ _0820_ demux.PSR_C VGND VGND VPWR VPWR _0887_ sky130_fd_sc_hd__or4b_1
X_2132_ _0823_ _0828_ _1202_ _1404_ _1244_ VGND VGND VPWR VPWR _1405_ sky130_fd_sc_hd__o41ai_2
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2201_ _1264_ _1336_ VGND VGND VPWR VPWR _1474_ sky130_fd_sc_hd__or2_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2063_ _1263_ _1150_ _0941_ VGND VGND VPWR VPWR _1336_ sky130_fd_sc_hd__a21o_1
XFILLER_0_71_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1916_ _1099_ _1130_ _1192_ _1197_ VGND VGND VPWR VPWR _1198_ sky130_fd_sc_hd__or4_1
XFILLER_0_60_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1847_ _0830_ _0815_ VGND VGND VPWR VPWR _1131_ sky130_fd_sc_hd__nor2_4
X_2896_ _0709_ _0700_ _0712_ VGND VGND VPWR VPWR _0713_ sky130_fd_sc_hd__a21oi_1
X_2965_ _0537_ _0775_ VGND VGND VPWR VPWR _0776_ sky130_fd_sc_hd__xnor2_1
X_1778_ _0967_ _0969_ net55 _1012_ VGND VGND VPWR VPWR _1062_ sky130_fd_sc_hd__and4b_1
XFILLER_0_12_231 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1701_ _0877_ VGND VGND VPWR VPWR _1001_ sky130_fd_sc_hd__clkbuf_4
X_2681_ _0529_ _0499_ _0531_ _0961_ VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__a31oi_1
XFILLER_0_38_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2750_ _0593_ _0594_ _0596_ _0537_ VGND VGND VPWR VPWR _0597_ sky130_fd_sc_hd__o22a_1
X_1632_ _0820_ _0819_ VGND VGND VPWR VPWR _0939_ sky130_fd_sc_hd__and2b_2
X_1563_ _0844_ _0818_ _0869_ VGND VGND VPWR VPWR _0870_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_41_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3095_ clknet_4_2_0_clk _0087_ net58 VGND VGND VPWR VPWR internalDataflow.addressLowBusModule.busInputs\[36\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2115_ _1382_ _1328_ _1387_ VGND VGND VPWR VPWR _1388_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_71_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2046_ internalDataflow.accRegToDB\[6\] _1316_ _1318_ demux.PSR_V VGND VGND VPWR
+ VPWR _1319_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2879_ internalDataflow.addressLowBusModule.busInputs\[23\] _0536_ VGND VGND VPWR
+ VPWR _0697_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2948_ internalDataflow.addressHighBusModule.busInputs\[22\] _0558_ VGND VGND VPWR
+ VPWR _0760_ sky130_fd_sc_hd__or2_1
XFILLER_0_40_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2802_ _0644_ VGND VGND VPWR VPWR _0645_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_41_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2664_ _0517_ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_326 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2733_ _0576_ _0577_ _0580_ VGND VGND VPWR VPWR _0581_ sky130_fd_sc_hd__o21ai_1
X_1615_ demux.state_machine.timeState\[3\] _0920_ _0921_ _0875_ VGND VGND VPWR VPWR
+ _0922_ sky130_fd_sc_hd__a22o_1
X_1546_ _0821_ _0852_ VGND VGND VPWR VPWR _0853_ sky130_fd_sc_hd__nor2_1
X_2595_ _0382_ _0459_ _0463_ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__or3_1
XFILLER_0_5_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3078_ clknet_4_5_0_clk _0070_ net69 VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__dfrtp_1
X_3147_ clknet_4_9_0_clk _0117_ net65 VGND VGND VPWR VPWR demux.PSR_N sky130_fd_sc_hd__dfrtp_1
XFILLER_0_64_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2029_ _1262_ _1289_ _0960_ _1301_ VGND VGND VPWR VPWR _1302_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_9_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_72_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2380_ internalDataflow.stackBusModule.busInputs\[33\] _1371_ VGND VGND VPWR VPWR
+ _0268_ sky130_fd_sc_hd__and2_1
X_3001_ instructionLoader.interruptInjector.resetDetected _0981_ VGND VGND VPWR VPWR
+ _0798_ sky130_fd_sc_hd__and2_1
XFILLER_0_36_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput6 dataBusInput[4] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_61_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2716_ _0546_ _0552_ _0555_ internalDataflow.addressLowBusModule.busInputs\[17\]
+ _0565_ VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__a221o_1
X_2647_ _0507_ VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__clkbuf_1
X_1529_ _0832_ _0833_ _0834_ _0835_ VGND VGND VPWR VPWR _0836_ sky130_fd_sc_hd__nand4_4
X_2578_ internalDataflow.addressLowBusModule.busInputs\[28\] net45 _0448_ _0382_ VGND
+ VGND VPWR VPWR _0449_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_37_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1880_ _1034_ _1052_ _1113_ _1091_ _0872_ VGND VGND VPWR VPWR _1163_ sky130_fd_sc_hd__a32o_1
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2501_ _0362_ _0365_ _0381_ _0384_ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_24_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2432_ _1325_ _0319_ VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__nor2_1
X_2363_ _1465_ _0237_ _0242_ _0250_ VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__a211o_1
X_2294_ _0181_ VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__inv_2
XFILLER_0_59_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_34_218 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xmax_cap46 _0119_ VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__buf_2
XFILLER_0_69_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1863_ _1140_ _1141_ _1142_ _1146_ VGND VGND VPWR VPWR _1147_ sky130_fd_sc_hd__or4_1
XFILLER_0_71_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1932_ _1207_ _1210_ _1212_ VGND VGND VPWR VPWR _1213_ sky130_fd_sc_hd__or3_1
XFILLER_0_33_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2981_ _0787_ VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1794_ _0966_ _1059_ _1075_ _1067_ _1077_ VGND VGND VPWR VPWR _1078_ sky130_fd_sc_hd__a32o_1
XFILLER_0_58_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2415_ internalDataflow.addressHighBusModule.busInputs\[23\] _1294_ _1314_ _1012_
+ _0302_ VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__a221o_1
XFILLER_0_24_273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2277_ demux.reset demux.setInterruptFlag demux.nmi VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__nor3_1
X_2346_ internalDataflow.addressLowBusModule.busInputs\[16\] _1315_ _0232_ _0233_
+ net134 VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_28_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_298 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2131_ _0863_ _0867_ _1097_ _0876_ VGND VGND VPWR VPWR _1404_ sky130_fd_sc_hd__o31a_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2200_ _1006_ _1455_ VGND VGND VPWR VPWR _1473_ sky130_fd_sc_hd__and2_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2062_ _0959_ net42 _1332_ _1334_ _0951_ VGND VGND VPWR VPWR _1335_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_28_55 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2964_ internalDataflow.addressHighBusModule.busInputs\[23\] _0774_ VGND VGND VPWR
+ VPWR _0775_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1915_ _1193_ _1196_ VGND VGND VPWR VPWR _1197_ sky130_fd_sc_hd__or2_1
X_1777_ _1058_ _0974_ _1034_ _1060_ VGND VGND VPWR VPWR _1061_ sky130_fd_sc_hd__a22o_1
X_1846_ _1127_ _0976_ _1047_ _1055_ _1129_ VGND VGND VPWR VPWR _1130_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2895_ _0710_ _0711_ VGND VGND VPWR VPWR _0712_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2329_ _0148_ _0212_ _0208_ VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__o21ba_2
XFILLER_0_62_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_8_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_8_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_62_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_408 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1700_ demux.state_machine.timeState\[5\] _0981_ _1000_ demux.state_machine.timeState\[1\]
+ VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__a22o_1
X_1631_ _0917_ _0937_ demux.reset VGND VGND VPWR VPWR _0938_ sky130_fd_sc_hd__a21oi_1
X_2680_ _1005_ _0530_ demux.state_machine.currentAddress\[7\] VGND VGND VPWR VPWR
+ _0531_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_41_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1562_ _0841_ VGND VGND VPWR VPWR _0869_ sky130_fd_sc_hd__clkbuf_4
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2045_ _1317_ _1302_ VGND VGND VPWR VPWR _1318_ sky130_fd_sc_hd__and2_2
X_2114_ _1326_ _1383_ _1386_ VGND VGND VPWR VPWR _1387_ sky130_fd_sc_hd__nor3_2
X_3094_ clknet_4_2_0_clk _0086_ net58 VGND VGND VPWR VPWR internalDataflow.addressLowBusModule.busInputs\[35\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2947_ internalDataflow.addressHighBusModule.busInputs\[22\] _0557_ VGND VGND VPWR
+ VPWR _0759_ sky130_fd_sc_hd__nand2_1
X_1829_ _1012_ _0967_ _0969_ _1010_ VGND VGND VPWR VPWR _1113_ sky130_fd_sc_hd__and4_2
XFILLER_0_44_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2878_ internalDataflow.addressHighBusModule.busInputs\[16\] _0536_ VGND VGND VPWR
+ VPWR _0696_ sky130_fd_sc_hd__xor2_1
XFILLER_0_4_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_279 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2801_ _0999_ _0642_ _0643_ VGND VGND VPWR VPWR _0644_ sky130_fd_sc_hd__and3_1
XFILLER_0_46_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1614_ _0869_ _0838_ VGND VGND VPWR VPWR _0921_ sky130_fd_sc_hd__nor2_2
XFILLER_0_41_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_88 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2594_ _0410_ _0460_ _0461_ _0462_ _0361_ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__o311a_1
XFILLER_0_1_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2663_ internalDataflow.accRegToDB\[5\] _0146_ _0511_ VGND VGND VPWR VPWR _0517_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2732_ _0578_ _0579_ VGND VGND VPWR VPWR _0580_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1545_ _0851_ VGND VGND VPWR VPWR _0852_ sky130_fd_sc_hd__buf_4
XFILLER_0_1_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3146_ clknet_4_4_0_clk _0116_ net60 VGND VGND VPWR VPWR branch_ff.branchBackward
+ sky130_fd_sc_hd__dfrtp_2
X_2028_ net13 _0950_ _1297_ _1300_ pulse_slower.nextEnableState\[0\] VGND VGND VPWR
+ VPWR _1301_ sky130_fd_sc_hd__o2111a_1
X_3077_ clknet_4_10_0_clk _0069_ net64 VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_198 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput7 dataBusInput[5] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__buf_2
X_3000_ demux.nmi _0341_ _0797_ net77 VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__a22o_1
XFILLER_0_6_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2715_ _0553_ _0564_ VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__nor2_1
X_2646_ net123 _0130_ _0502_ VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2577_ _0442_ _0443_ _0447_ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__a21oi_1
X_1528_ _0811_ VGND VGND VPWR VPWR _0835_ sky130_fd_sc_hd__clkbuf_4
X_3129_ clknet_4_6_0_clk _0016_ net67 VGND VGND VPWR VPWR demux.state_machine.timeState\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_37_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2431_ _0868_ _1143_ _1007_ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__o21ai_2
X_2500_ _0382_ _0383_ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2362_ _0243_ _0249_ VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__nor2_1
X_2293_ _0179_ _0180_ VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__nand2b_2
XFILLER_0_59_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2629_ _1079_ _0492_ _0493_ _1102_ _0495_ VGND VGND VPWR VPWR _0496_ sky130_fd_sc_hd__a221o_1
Xmax_cap47 _1387_ VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_65_311 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2980_ net88 _0196_ _0783_ VGND VGND VPWR VPWR _0787_ sky130_fd_sc_hd__mux2_1
Xinput10 interruptRequest VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_1
X_1862_ _1143_ _1091_ _0972_ _1019_ _1145_ VGND VGND VPWR VPWR _1146_ sky130_fd_sc_hd__a221o_1
X_1931_ _1064_ _1126_ _1129_ _1211_ VGND VGND VPWR VPWR _1212_ sky130_fd_sc_hd__or4_1
X_1793_ _0815_ _1076_ VGND VGND VPWR VPWR _1077_ sky130_fd_sc_hd__nor2_2
XFILLER_0_24_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2414_ internalDataflow.accRegToDB\[7\] _1316_ _1318_ demux.PSR_N VGND VGND VPWR
+ VPWR _0302_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_285 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2345_ demux.PSR_C _1317_ _1302_ _1294_ internalDataflow.addressHighBusModule.busInputs\[16\]
+ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__a32o_1
X_2276_ _1388_ _0162_ _0163_ _1387_ VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__a22o_1
XFILLER_0_47_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2130_ _1392_ _1394_ _1398_ _1402_ VGND VGND VPWR VPWR _1403_ sky130_fd_sc_hd__or4_1
X_2061_ _1003_ _1333_ _1241_ VGND VGND VPWR VPWR _1334_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_67 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1914_ _1194_ _1195_ VGND VGND VPWR VPWR _1196_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_55 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2963_ _0773_ _0763_ _0759_ VGND VGND VPWR VPWR _0774_ sky130_fd_sc_hd__o21a_1
X_1776_ _1052_ _1059_ VGND VGND VPWR VPWR _1060_ sky130_fd_sc_hd__and2_1
X_1845_ _1128_ _1091_ _1048_ _1059_ VGND VGND VPWR VPWR _1129_ sky130_fd_sc_hd__a22o_1
X_2894_ internalDataflow.addressHighBusModule.busInputs\[17\] _0556_ VGND VGND VPWR
+ VPWR _0711_ sky130_fd_sc_hd__and2_1
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2328_ _1460_ _0215_ VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__and2_2
XFILLER_0_67_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2259_ _1460_ _0146_ VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__and2_1
XFILLER_0_62_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1630_ demux.state_machine.timeState\[2\] demux.state_machine.timeState\[6\] VGND
+ VGND VPWR VPWR _0937_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1561_ _0829_ _0852_ VGND VGND VPWR VPWR _0868_ sky130_fd_sc_hd__nor2_4
XFILLER_0_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2113_ _0982_ _1295_ _1385_ _0998_ VGND VGND VPWR VPWR _1386_ sky130_fd_sc_hd__o211a_2
X_2044_ _0952_ _1292_ VGND VGND VPWR VPWR _1317_ sky130_fd_sc_hd__and2_1
X_3093_ clknet_4_2_0_clk _0085_ net58 VGND VGND VPWR VPWR internalDataflow.addressLowBusModule.busInputs\[34\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_29_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2877_ _0695_ VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__clkbuf_1
X_2946_ net125 _0555_ _0753_ _0546_ _0758_ VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__a221o_1
X_1759_ net113 _1044_ _0979_ VGND VGND VPWR VPWR _1045_ sky130_fd_sc_hd__mux2_1
X_1828_ _0961_ _1074_ VGND VGND VPWR VPWR _1112_ sky130_fd_sc_hd__nor2_1
XFILLER_0_25_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2800_ _0985_ _1283_ _1441_ _0987_ _0500_ VGND VGND VPWR VPWR _0643_ sky130_fd_sc_hd__a221o_1
XFILLER_0_26_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2731_ internalDataflow.addressLowBusModule.busInputs\[19\] _0535_ VGND VGND VPWR
+ VPWR _0579_ sky130_fd_sc_hd__and2_1
X_1544_ _0812_ _0813_ _0810_ _0811_ VGND VGND VPWR VPWR _0851_ sky130_fd_sc_hd__or4bb_1
X_1613_ _0869_ _0909_ VGND VGND VPWR VPWR _0920_ sky130_fd_sc_hd__nor2_2
XFILLER_0_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2593_ _0134_ _0410_ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__nand2_1
X_2662_ _0516_ VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_7_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_7_0_clk sky130_fd_sc_hd__clkbuf_8
X_3145_ clknet_4_6_0_clk _0115_ net67 VGND VGND VPWR VPWR demux.isAddressing sky130_fd_sc_hd__dfstp_1
XFILLER_0_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2027_ _1241_ _1299_ _1258_ VGND VGND VPWR VPWR _1300_ sky130_fd_sc_hd__or3_1
X_3076_ clknet_4_2_0_clk _0068_ net58 VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_283 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2929_ _0740_ _0741_ _0546_ VGND VGND VPWR VPWR _0743_ sky130_fd_sc_hd__o21a_1
XFILLER_0_17_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_11_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xinput8 dataBusInput[6] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__buf_2
XFILLER_0_42_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2714_ _0560_ _0563_ VGND VGND VPWR VPWR _0564_ sky130_fd_sc_hd__xnor2_1
X_1527_ _0810_ VGND VGND VPWR VPWR _0834_ sky130_fd_sc_hd__buf_4
X_2645_ _0506_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__clkbuf_1
X_2576_ _0179_ _0407_ _0445_ _0446_ VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__o22a_1
X_3128_ clknet_4_5_0_clk _0015_ net69 VGND VGND VPWR VPWR demux.state_machine.timeState\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_3059_ clknet_4_8_0_clk _0051_ net62 VGND VGND VPWR VPWR internalDataflow.accRegToDB\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2430_ _0292_ _0317_ VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__or2_1
X_2361_ _1329_ _0244_ _0248_ _0235_ _1327_ VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__o32ai_4
XFILLER_0_11_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2292_ _0171_ _0178_ VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__or2_1
XFILLER_0_42_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2628_ _0983_ _0494_ _0913_ VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__o21a_1
X_2559_ _0431_ VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap48 _1312_ VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_65_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_242 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1930_ _0921_ _0977_ _1048_ _1081_ _1187_ VGND VGND VPWR VPWR _1211_ sky130_fd_sc_hd__a221o_1
XFILLER_0_33_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput11 nonMaskableInterrupt VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_1
X_1861_ _1144_ _1066_ _1054_ _1087_ VGND VGND VPWR VPWR _1145_ sky130_fd_sc_hd__a22o_1
XFILLER_0_56_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1792_ _0821_ VGND VGND VPWR VPWR _1076_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_58_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2344_ net2 _1313_ _1302_ _1316_ internalDataflow.accRegToDB\[0\] VGND VGND VPWR
+ VPWR _0232_ sky130_fd_sc_hd__a32o_1
X_2413_ _0300_ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2275_ internalDataflow.addressHighBusModule.busInputs\[20\] _1422_ _1424_ _0954_
+ _1431_ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__o221a_1
XFILLER_0_62_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_267 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_370 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_359 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2060_ _1138_ _1058_ _0867_ _1204_ VGND VGND VPWR VPWR _1333_ sky130_fd_sc_hd__or4_1
XFILLER_0_44_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1913_ _0958_ _0966_ _0970_ _1066_ _0933_ VGND VGND VPWR VPWR _1195_ sky130_fd_sc_hd__a32o_1
XFILLER_0_56_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2893_ internalDataflow.addressHighBusModule.busInputs\[17\] _0536_ VGND VGND VPWR
+ VPWR _0710_ sky130_fd_sc_hd__nor2_1
XFILLER_0_8_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2962_ internalDataflow.addressHighBusModule.busInputs\[22\] _0557_ VGND VGND VPWR
+ VPWR _0773_ sky130_fd_sc_hd__nor2_1
X_1775_ _0967_ _1014_ VGND VGND VPWR VPWR _1059_ sky130_fd_sc_hd__and2b_2
X_1844_ _0857_ _1076_ VGND VGND VPWR VPWR _1128_ sky130_fd_sc_hd__nor2_1
XFILLER_0_4_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2327_ _1326_ _0208_ _0214_ _1329_ VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__o2bb2a_2
X_2258_ _0142_ _0145_ _1329_ VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__mux2_2
XFILLER_0_67_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2189_ _1006_ _0905_ VGND VGND VPWR VPWR _1462_ sky130_fd_sc_hd__and2_1
XFILLER_0_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1560_ _0865_ _0860_ _0866_ VGND VGND VPWR VPWR _0867_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_53_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2112_ _0983_ _0905_ _1352_ _1384_ VGND VGND VPWR VPWR _1385_ sky130_fd_sc_hd__a31o_1
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2043_ _1301_ _1262_ _1289_ VGND VGND VPWR VPWR _1316_ sky130_fd_sc_hd__and3_2
X_3092_ clknet_4_2_0_clk _0084_ net58 VGND VGND VPWR VPWR internalDataflow.addressLowBusModule.busInputs\[33\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1827_ _1106_ _1107_ _1110_ VGND VGND VPWR VPWR _1111_ sky130_fd_sc_hd__or3_1
XFILLER_0_44_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2876_ internalDataflow.addressLowBusModule.busInputs\[39\] _0305_ _0687_ VGND VGND
+ VPWR VPWR _0695_ sky130_fd_sc_hd__mux2_1
X_2945_ _0756_ _0757_ _0553_ VGND VGND VPWR VPWR _0758_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1758_ net3 _1010_ _1042_ _1043_ _0964_ VGND VGND VPWR VPWR _1044_ sky130_fd_sc_hd__a32o_1
X_1689_ demux.state_machine.currentAddress\[11\] demux.state_machine.currentAddress\[3\]
+ demux.state_machine.currentAddress\[7\] VGND VGND VPWR VPWR _0991_ sky130_fd_sc_hd__or3_2
XFILLER_0_25_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2661_ internalDataflow.accRegToDB\[4\] _0170_ _0511_ VGND VGND VPWR VPWR _0516_
+ sky130_fd_sc_hd__mux2_1
X_2730_ internalDataflow.addressLowBusModule.busInputs\[19\] _0558_ VGND VGND VPWR
+ VPWR _0578_ sky130_fd_sc_hd__nor2_1
X_1543_ _0830_ _0836_ VGND VGND VPWR VPWR _0850_ sky130_fd_sc_hd__nor2_1
X_1612_ _0876_ _0915_ _0916_ _0918_ VGND VGND VPWR VPWR _0919_ sky130_fd_sc_hd__a211o_1
XFILLER_0_41_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2592_ _1460_ _0305_ _0364_ _0408_ _0135_ VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__a32o_1
XFILLER_0_22_340 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3075_ clknet_4_13_0_clk _0067_ net70 VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__dfrtp_2
X_3144_ clknet_4_4_0_clk _0114_ net60 VGND VGND VPWR VPWR branch_ff.branchForward
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_49_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2026_ _1189_ _1298_ _1263_ VGND VGND VPWR VPWR _1299_ sky130_fd_sc_hd__o21a_1
XFILLER_0_9_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2859_ _1489_ VGND VGND VPWR VPWR _0685_ sky130_fd_sc_hd__inv_2
X_2928_ _0740_ _0741_ VGND VGND VPWR VPWR _0742_ sky130_fd_sc_hd__nand2_1
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xinput9 dataBusInput[7] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_2
XFILLER_0_52_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2644_ net111 _0153_ _0502_ VGND VGND VPWR VPWR _0506_ sky130_fd_sc_hd__mux2_1
X_2713_ _0561_ _0562_ VGND VGND VPWR VPWR _0563_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1526_ _0813_ VGND VGND VPWR VPWR _0833_ sky130_fd_sc_hd__buf_4
X_2575_ _0147_ _0364_ _0408_ _0180_ _0410_ VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__a221o_1
X_3127_ clknet_4_6_0_clk _0014_ net69 VGND VGND VPWR VPWR demux.state_machine.timeState\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_3058_ clknet_4_3_0_clk _0050_ net63 VGND VGND VPWR VPWR internalDataflow.accRegToDB\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_2009_ demux.state_machine.timeState\[0\] _0896_ VGND VGND VPWR VPWR _1282_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_6_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_6_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_51_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2360_ _1430_ _0245_ _0246_ _0247_ _1387_ VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__o2111a_1
X_2291_ _0171_ _0178_ VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__and2_1
XFILLER_0_63_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2627_ _1001_ _0491_ VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1509_ _0812_ _0813_ _0810_ _0811_ VGND VGND VPWR VPWR _0816_ sky130_fd_sc_hd__or4_2
X_2489_ _0136_ _0156_ _0371_ VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__nand3_1
X_2558_ _0430_ internalDataflow.addressLowBusModule.busInputs\[26\] net45 VGND VGND
+ VPWR VPWR _0431_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xmax_cap49 net135 VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__buf_1
XFILLER_0_33_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_17_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1860_ _0871_ _0844_ VGND VGND VPWR VPWR _1144_ sky130_fd_sc_hd__nor2_2
XFILLER_0_56_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput12 nrst VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_71_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1791_ _1074_ VGND VGND VPWR VPWR _1075_ sky130_fd_sc_hd__inv_2
XFILLER_0_3_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2412_ _0296_ _0299_ net47 VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__mux2_1
X_2274_ _0159_ _0161_ _1372_ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__o21a_1
X_2343_ _0228_ _0230_ _1372_ VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__o21a_1
XFILLER_0_59_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1989_ _1258_ _1261_ _0948_ VGND VGND VPWR VPWR _1262_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_7_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_21_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1912_ _0853_ _0974_ _0972_ _1088_ VGND VGND VPWR VPWR _1194_ sky130_fd_sc_hd__a22o_1
X_1843_ _0901_ _0855_ VGND VGND VPWR VPWR _1127_ sky130_fd_sc_hd__nor2_1
X_2892_ internalDataflow.addressHighBusModule.busInputs\[16\] _0536_ VGND VGND VPWR
+ VPWR _0709_ sky130_fd_sc_hd__nand2_1
X_2961_ _0669_ _0771_ VGND VGND VPWR VPWR _0772_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_69_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1774_ _0821_ _0861_ VGND VGND VPWR VPWR _1058_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2326_ _1388_ _0212_ _0213_ net47 VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__a22o_1
X_2257_ internalDataflow.addressHighBusModule.busInputs\[21\] _1294_ _0143_ _0144_
+ VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__a211o_1
XFILLER_0_47_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2188_ _1434_ _1460_ VGND VGND VPWR VPWR _1461_ sky130_fd_sc_hd__nand2_1
XFILLER_0_62_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_382 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold1 instructionLoader.interruptInjector.nmiSync.nextQ2 VGND VGND VPWR VPWR net73
+ sky130_fd_sc_hd__dlygate4sd3_1
X_2111_ _1241_ VGND VGND VPWR VPWR _1384_ sky130_fd_sc_hd__clkbuf_4
X_2042_ _1262_ _1289_ _1304_ VGND VGND VPWR VPWR _1315_ sky130_fd_sc_hd__a21boi_4
X_3091_ clknet_4_3_0_clk _0083_ net61 VGND VGND VPWR VPWR internalDataflow.addressLowBusModule.busInputs\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1826_ _0923_ _0976_ _1069_ _1081_ _1109_ VGND VGND VPWR VPWR _1110_ sky130_fd_sc_hd__a221o_1
XFILLER_0_25_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2875_ _0694_ VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__clkbuf_1
X_2944_ _0662_ _0755_ VGND VGND VPWR VPWR _0757_ sky130_fd_sc_hd__or2_1
XFILLER_0_17_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1757_ _1013_ _1017_ _1040_ VGND VGND VPWR VPWR _1043_ sky130_fd_sc_hd__a21o_1
X_1688_ _0987_ _0988_ demux.state_machine.currentAddress\[6\] net54 VGND VGND VPWR
+ VPWR _0990_ sky130_fd_sc_hd__o31a_1
X_2309_ _1467_ _1479_ _0196_ VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__mux2_1
XFILLER_0_67_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1611_ _0917_ _0871_ _0815_ VGND VGND VPWR VPWR _0918_ sky130_fd_sc_hd__nor3_1
XFILLER_0_41_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2660_ _0515_ VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__clkbuf_1
X_1542_ _0823_ _0828_ _0840_ _0848_ VGND VGND VPWR VPWR _0849_ sky130_fd_sc_hd__or4_1
X_2591_ _0136_ _0444_ VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_352 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3143_ clknet_4_15_0_clk _0025_ net72 VGND VGND VPWR VPWR demux.state_machine.currentInstruction\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_2025_ _0885_ _0865_ _1076_ VGND VGND VPWR VPWR _1298_ sky130_fd_sc_hd__a21oi_2
X_3074_ clknet_4_10_0_clk _0066_ net64 VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_9_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2927_ _0731_ _0734_ _0732_ VGND VGND VPWR VPWR _0741_ sky130_fd_sc_hd__o21bai_2
X_1809_ _1078_ _1083_ _1089_ _1092_ VGND VGND VPWR VPWR _1093_ sky130_fd_sc_hd__or4_1
X_2789_ _1383_ _1386_ VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__nand2_4
X_2858_ internalDataflow.addressLowBusModule.busInputs\[32\] VGND VGND VPWR VPWR _0684_
+ sky130_fd_sc_hd__inv_2
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_182 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2643_ _0505_ VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__clkbuf_1
X_2712_ _0281_ _0241_ VGND VGND VPWR VPWR _0562_ sky130_fd_sc_hd__nor2_1
XFILLER_0_14_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2574_ _0181_ _0444_ VGND VGND VPWR VPWR _0445_ sky130_fd_sc_hd__nor2_1
X_1525_ _0812_ VGND VGND VPWR VPWR _0832_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3126_ clknet_4_6_0_clk _0013_ net67 VGND VGND VPWR VPWR demux.state_machine.timeState\[0\]
+ sky130_fd_sc_hd__dfstp_2
X_2008_ _1003_ _0904_ _1241_ VGND VGND VPWR VPWR _1281_ sky130_fd_sc_hd__a21oi_2
X_3057_ clknet_4_13_0_clk _0049_ net70 VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_5_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2290_ _0173_ _0177_ _0154_ VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__mux2_1
XFILLER_0_27_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2626_ _1007_ _0936_ _1400_ VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__or3_1
XFILLER_0_56_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2557_ _0424_ _0429_ _0382_ VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__mux2_1
X_1508_ _0814_ VGND VGND VPWR VPWR _0815_ sky130_fd_sc_hd__buf_4
XFILLER_0_37_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2488_ _0156_ _0371_ _0136_ VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__a21o_2
X_3109_ clknet_4_12_0_clk _0101_ net70 VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1790_ _0957_ _0954_ _1022_ _1039_ VGND VGND VPWR VPWR _1074_ sky130_fd_sc_hd__a211o_1
Xinput13 ready VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_2
X_2411_ _0297_ _1422_ _1424_ _0968_ _0298_ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__o221a_1
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2273_ internalDataflow.stackBusModule.busInputs\[36\] _1371_ _0160_ VGND VGND VPWR
+ VPWR _0161_ sky130_fd_sc_hd__a21o_1
X_2342_ internalDataflow.stackBusModule.busInputs\[32\] _1371_ _1378_ internalDataflow.addressLowBusModule.busInputs\[32\]
+ _0229_ VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1988_ _0897_ _1079_ _1260_ _0833_ VGND VGND VPWR VPWR _1261_ sky130_fd_sc_hd__a22o_1
XFILLER_0_23_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2609_ _0292_ _0378_ _0361_ VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__a21o_1
Xclkbuf_4_5_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_5_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_21_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2960_ _0755_ _0765_ _0769_ _0770_ VGND VGND VPWR VPWR _0771_ sky130_fd_sc_hd__or4_1
X_1773_ _1050_ _1056_ VGND VGND VPWR VPWR _1057_ sky130_fd_sc_hd__or2_1
X_1911_ _0868_ _0976_ _1019_ _1113_ VGND VGND VPWR VPWR _1193_ sky130_fd_sc_hd__a22o_1
X_1842_ _1120_ _1124_ _1125_ VGND VGND VPWR VPWR _1126_ sky130_fd_sc_hd__or3_1
XFILLER_0_37_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2891_ _0649_ _0707_ VGND VGND VPWR VPWR _0708_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_29_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2187_ _1459_ VGND VGND VPWR VPWR _1460_ sky130_fd_sc_hd__buf_2
XFILLER_0_19_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2256_ internalDataflow.accRegToDB\[5\] _1316_ _1314_ net7 _1318_ VGND VGND VPWR
+ VPWR _0144_ sky130_fd_sc_hd__a221o_1
X_2325_ internalDataflow.addressHighBusModule.busInputs\[18\] _1422_ _1424_ net4 _1431_
+ VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__o221a_1
XFILLER_0_62_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_53_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_166 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_380 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold2 instructionLoader.interruptInjector.irqSync.nextQ2 VGND VGND VPWR VPWR net74
+ sky130_fd_sc_hd__dlygate4sd3_1
X_2041_ _1313_ _1302_ VGND VGND VPWR VPWR _1314_ sky130_fd_sc_hd__and2_2
X_2110_ _1325_ _1382_ VGND VGND VPWR VPWR _1383_ sky130_fd_sc_hd__or2_2
X_3090_ clknet_4_8_0_clk _0082_ net62 VGND VGND VPWR VPWR internalDataflow.stackBusModule.busInputs\[47\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_72_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2943_ _0662_ _0755_ VGND VGND VPWR VPWR _0756_ sky130_fd_sc_hd__nand2_1
X_1756_ _1012_ _0969_ _1010_ _1024_ _1041_ VGND VGND VPWR VPWR _1042_ sky130_fd_sc_hd__a41o_1
X_1825_ _1108_ _1067_ _1055_ _1069_ VGND VGND VPWR VPWR _1109_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2874_ internalDataflow.addressLowBusModule.busInputs\[38\] _1434_ _0687_ VGND VGND
+ VPWR VPWR _0694_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1687_ _0932_ _0896_ _0875_ demux.state_machine.timeState\[6\] VGND VGND VPWR VPWR
+ _0989_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_29_80 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2308_ _1257_ _0191_ _0186_ VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__a21oi_4
X_2239_ _0120_ _1500_ _0124_ VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__nor3b_4
XFILLER_0_35_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_41_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1610_ demux.state_machine.timeState\[4\] VGND VGND VPWR VPWR _0917_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2590_ _0136_ _0291_ _0458_ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3142_ clknet_4_15_0_clk _0024_ net72 VGND VGND VPWR VPWR demux.state_machine.currentInstruction\[4\]
+ sky130_fd_sc_hd__dfrtp_1
X_1541_ _0842_ _0845_ _0846_ _0847_ VGND VGND VPWR VPWR _0848_ sky130_fd_sc_hd__or4_2
XFILLER_0_5_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2024_ _1214_ _1296_ _0948_ VGND VGND VPWR VPWR _1297_ sky130_fd_sc_hd__a21o_1
X_3073_ clknet_4_13_0_clk _0065_ net70 VGND VGND VPWR VPWR internalDataflow.addressLowBusModule.busInputs\[23\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_64_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2857_ _0683_ VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2926_ _0738_ _0739_ VGND VGND VPWR VPWR _0740_ sky130_fd_sc_hd__and2_1
XFILLER_0_17_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1808_ _0966_ _1080_ _1090_ _1091_ _0873_ VGND VGND VPWR VPWR _1092_ sky130_fd_sc_hd__a32o_1
X_1739_ _1016_ _1029_ VGND VGND VPWR VPWR _1030_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2788_ _0631_ VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_342 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_39_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2711_ _0281_ _0241_ VGND VGND VPWR VPWR _0561_ sky130_fd_sc_hd__and2_1
X_1524_ _0830_ _0816_ VGND VGND VPWR VPWR _0831_ sky130_fd_sc_hd__nor2_2
X_2642_ net28 _0177_ _0502_ VGND VGND VPWR VPWR _0505_ sky130_fd_sc_hd__mux2_1
X_2573_ _1202_ _0323_ VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__nand2_1
X_3125_ clknet_4_4_0_clk _0113_ net69 VGND VGND VPWR VPWR free_carry_ff.freeCarry
+ sky130_fd_sc_hd__dfrtp_1
X_2007_ _1003_ _0840_ _1150_ _0897_ _1279_ VGND VGND VPWR VPWR _1280_ sky130_fd_sc_hd__a221oi_4
XFILLER_0_26_92 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3056_ clknet_4_0_0_clk _0048_ net57 VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_18_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2909_ _0652_ _0724_ VGND VGND VPWR VPWR _0725_ sky130_fd_sc_hd__xor2_1
XFILLER_0_20_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2625_ demux.state_machine.timeState\[3\] _1285_ _0491_ VGND VGND VPWR VPWR _0492_
+ sky130_fd_sc_hd__or3_1
X_1507_ _0810_ _0811_ _0812_ _0813_ VGND VGND VPWR VPWR _0814_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_42_278 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2556_ _0368_ _0428_ VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__xnor2_1
X_2487_ _0179_ _0370_ _0158_ VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_49_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3108_ clknet_4_8_0_clk _0100_ net64 VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_65_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3039_ clknet_4_8_0_clk _0033_ net62 VGND VGND VPWR VPWR internalDataflow.stackBusModule.busInputs\[39\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_33_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput14 setOverflow VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__dlymetal6s2s_1
X_2410_ _1429_ _1422_ _1424_ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__nand3_1
X_2341_ internalDataflow.addressLowBusModule.busInputs\[24\] _1366_ _1341_ _1350_
+ VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__and4_1
X_2272_ internalDataflow.addressLowBusModule.busInputs\[28\] _1377_ _1378_ internalDataflow.addressLowBusModule.busInputs\[36\]
+ VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1987_ _0932_ _1259_ VGND VGND VPWR VPWR _1260_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2608_ _0292_ _0378_ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__nor2_1
X_2539_ _0261_ _0407_ _0411_ _0413_ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__o22a_1
XFILLER_0_3_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1910_ _1189_ _0976_ _1069_ _1087_ _1191_ VGND VGND VPWR VPWR _1192_ sky130_fd_sc_hd__a221o_1
XFILLER_0_29_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2890_ _0702_ _0706_ VGND VGND VPWR VPWR _0707_ sky130_fd_sc_hd__nand2_1
X_1772_ _1051_ _1049_ _1054_ _1055_ _1032_ VGND VGND VPWR VPWR _1056_ sky130_fd_sc_hd__a221o_1
X_1841_ _0891_ _1122_ _1091_ _1047_ _1063_ VGND VGND VPWR VPWR _1125_ sky130_fd_sc_hd__a32o_1
XFILLER_0_56_167 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2324_ _0209_ _0210_ _0211_ _1372_ VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__o31a_1
X_2186_ _0998_ _1438_ _1450_ _1458_ VGND VGND VPWR VPWR _1459_ sky130_fd_sc_hd__and4_1
X_2255_ internalDataflow.addressLowBusModule.busInputs\[21\] _1315_ net48 VGND VGND
+ VPWR VPWR _0143_ sky130_fd_sc_hd__a21o_1
XFILLER_0_47_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_392 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2040_ _1303_ _1292_ VGND VGND VPWR VPWR _1313_ sky130_fd_sc_hd__nand2_1
Xhold3 net26 VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_72_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_71_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2942_ _0746_ _0754_ VGND VGND VPWR VPWR _0755_ sky130_fd_sc_hd__nand2_1
X_2873_ _0693_ VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_318 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1755_ net86 _0977_ _1019_ _1041_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__a22o_1
X_1686_ demux.state_machine.currentAddress\[12\] VGND VGND VPWR VPWR _0988_ sky130_fd_sc_hd__buf_2
X_1824_ _0855_ _1076_ VGND VGND VPWR VPWR _1108_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_4_4_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_4_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2238_ internalDataflow.addressLowBusModule.busInputs\[38\] net46 _0125_ internalDataflow.addressLowBusModule.busInputs\[30\]
+ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__a22o_1
X_2307_ _1460_ _0194_ VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__and2_1
XFILLER_0_67_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2169_ _1071_ _1285_ _1441_ _1168_ VGND VGND VPWR VPWR _1442_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1540_ _0826_ _0818_ VGND VGND VPWR VPWR _0847_ sky130_fd_sc_hd__nor2_4
XFILLER_0_22_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3141_ clknet_4_15_0_clk _0023_ net72 VGND VGND VPWR VPWR demux.state_machine.currentInstruction\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_2023_ _0988_ net54 _1295_ _0995_ VGND VGND VPWR VPWR _1296_ sky130_fd_sc_hd__a211o_1
X_3072_ clknet_4_12_0_clk _0064_ net65 VGND VGND VPWR VPWR internalDataflow.addressLowBusModule.busInputs\[22\]
+ sky130_fd_sc_hd__dfrtp_4
X_1807_ _1066_ VGND VGND VPWR VPWR _1091_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_60_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2856_ internalDataflow.stackBusModule.busInputs\[47\] _0305_ _0675_ VGND VGND VPWR
+ VPWR _0683_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2925_ internalDataflow.addressHighBusModule.busInputs\[20\] _0556_ VGND VGND VPWR
+ VPWR _0739_ sky130_fd_sc_hd__or2_1
X_1738_ _0954_ _0956_ VGND VGND VPWR VPWR _1029_ sky130_fd_sc_hd__nand2_1
X_1669_ _0961_ _0962_ VGND VGND VPWR VPWR _0973_ sky130_fd_sc_hd__or2_1
X_2787_ _0630_ internalDataflow.addressLowBusModule.busInputs\[23\] _0554_ VGND VGND
+ VPWR VPWR _0631_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_354 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_48_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2710_ _0241_ _0558_ _0559_ VGND VGND VPWR VPWR _0560_ sky130_fd_sc_hd__a21o_1
X_1523_ _0829_ VGND VGND VPWR VPWR _0830_ sky130_fd_sc_hd__clkbuf_8
X_2641_ _0504_ VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__clkbuf_1
X_2572_ _0181_ _0366_ _0361_ VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__a21oi_1
X_3124_ clknet_4_12_0_clk _0112_ net70 VGND VGND VPWR VPWR instructionLoader.interruptInjector.resetDetected
+ sky130_fd_sc_hd__dfstp_2
X_3055_ clknet_4_4_0_clk _0047_ net69 VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__dfrtp_1
X_2006_ _0932_ _0926_ VGND VGND VPWR VPWR _1279_ sky130_fd_sc_hd__and2_1
XFILLER_0_26_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2839_ _1002_ _0867_ _0672_ _1008_ VGND VGND VPWR VPWR _0673_ sky130_fd_sc_hd__a22o_1
XFILLER_0_45_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2908_ _0707_ _0722_ _0723_ VGND VGND VPWR VPWR _0724_ sky130_fd_sc_hd__or3_1
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2624_ _0879_ _1400_ VGND VGND VPWR VPWR _0491_ sky130_fd_sc_hd__or2_1
XFILLER_0_30_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1506_ demux.state_machine.currentInstruction\[0\] VGND VGND VPWR VPWR _0813_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_2_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2555_ _0288_ _0369_ _0426_ _0427_ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__or4_1
X_2486_ _0366_ _0369_ _0181_ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__a21oi_1
X_3107_ clknet_4_0_0_clk _0099_ net57 VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__dfrtp_1
X_3038_ clknet_4_3_0_clk _0032_ net58 VGND VGND VPWR VPWR internalDataflow.stackBusModule.busInputs\[38\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_68_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2271_ internalDataflow.stackBusModule.busInputs\[44\] _1373_ _1374_ internalDataflow.accRegToDB\[4\]
+ _1375_ VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__a221o_1
X_2340_ _1371_ _1367_ _0225_ _0227_ VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_59_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1986_ _0832_ _0939_ _0940_ VGND VGND VPWR VPWR _1259_ sky130_fd_sc_hd__and3b_2
XFILLER_0_23_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2607_ _0376_ _0383_ _0473_ _0474_ VGND VGND VPWR VPWR _0475_ sky130_fd_sc_hd__a31o_1
X_2469_ _1097_ _1298_ _1358_ _1007_ VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__o31a_1
X_2538_ _0404_ _0412_ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__and2_1
XFILLER_0_65_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1840_ _1121_ _0975_ _0972_ _1054_ _1123_ VGND VGND VPWR VPWR _1124_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1771_ _0967_ _1014_ VGND VGND VPWR VPWR _1055_ sky130_fd_sc_hd__and2_2
XFILLER_0_69_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2323_ internalDataflow.addressLowBusModule.busInputs\[26\] _1377_ _1378_ internalDataflow.addressLowBusModule.busInputs\[34\]
+ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__a22o_1
X_2254_ _1388_ _0140_ _0141_ net47 VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__a22o_1
XFILLER_0_18_61 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2185_ _1451_ _1454_ _1457_ _1305_ VGND VGND VPWR VPWR _1458_ sky130_fd_sc_hd__or4b_1
XFILLER_0_34_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1969_ _0875_ _1237_ _1238_ _1239_ _1241_ VGND VGND VPWR VPWR _1242_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_35_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold4 demux.state_machine.currentAddress\[8\] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_39_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1823_ _0944_ _1067_ _1054_ _1063_ VGND VGND VPWR VPWR _1107_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2872_ internalDataflow.addressLowBusModule.busInputs\[37\] _0146_ _0687_ VGND VGND
+ VPWR VPWR _0693_ sky130_fd_sc_hd__mux2_1
X_2941_ _0537_ _0659_ VGND VGND VPWR VPWR _0754_ sky130_fd_sc_hd__xnor2_1
X_1754_ _0954_ _1040_ VGND VGND VPWR VPWR _1041_ sky130_fd_sc_hd__and2_2
X_1685_ demux.state_machine.currentAddress\[1\] VGND VGND VPWR VPWR _0987_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_40_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2237_ _0124_ _0121_ VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__nor2_2
X_2306_ _1326_ _0186_ _0193_ _1329_ VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_48_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2168_ _1003_ _0879_ _0945_ VGND VGND VPWR VPWR _1441_ sky130_fd_sc_hd__or3_2
XFILLER_0_0_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2099_ _1303_ _1330_ _1367_ _1371_ VGND VGND VPWR VPWR _1372_ sky130_fd_sc_hd__a211o_4
XFILLER_0_16_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3140_ clknet_4_15_0_clk _0022_ net72 VGND VGND VPWR VPWR demux.state_machine.currentInstruction\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_3071_ clknet_4_11_0_clk _0063_ net65 VGND VGND VPWR VPWR internalDataflow.addressLowBusModule.busInputs\[21\]
+ sky130_fd_sc_hd__dfrtp_4
X_2022_ _0897_ _0985_ _0986_ net54 demux.state_machine.currentAddress\[1\] VGND VGND
+ VPWR VPWR _1295_ sky130_fd_sc_hd__a32o_1
XFILLER_0_9_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1806_ _0967_ _0958_ _1024_ VGND VGND VPWR VPWR _1090_ sky130_fd_sc_hd__a21o_1
XFILLER_0_60_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2786_ _0544_ _0623_ _0628_ _0629_ VGND VGND VPWR VPWR _0630_ sky130_fd_sc_hd__a22o_1
XFILLER_0_25_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2855_ _0682_ VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__clkbuf_1
X_2924_ internalDataflow.addressHighBusModule.busInputs\[20\] _0556_ VGND VGND VPWR
+ VPWR _0738_ sky130_fd_sc_hd__nand2_1
XFILLER_0_17_138 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1737_ _1028_ VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__clkbuf_1
X_1668_ _0971_ VGND VGND VPWR VPWR _0972_ sky130_fd_sc_hd__buf_2
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1599_ _0879_ _0900_ _0905_ VGND VGND VPWR VPWR _0906_ sky130_fd_sc_hd__o21a_1
XFILLER_0_13_366 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_63_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xclkbuf_4_3_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_3_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2640_ net122 _0200_ _0502_ VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__mux2_1
X_1522_ demux.state_machine.currentInstruction\[4\] _0819_ VGND VGND VPWR VPWR _0829_
+ sky130_fd_sc_hd__nand2b_4
XFILLER_0_22_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2571_ _0182_ _0288_ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__nand2_1
X_3054_ clknet_4_14_0_clk _0046_ net70 VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__dfrtp_1
X_3123_ clknet_4_14_0_clk _0111_ net71 VGND VGND VPWR VPWR instructionLoader.interruptInjector.nmiGeneratedFF.nmiRunning
+ sky130_fd_sc_hd__dfrtp_1
X_2005_ _1264_ _1270_ _1272_ _1277_ VGND VGND VPWR VPWR _1278_ sky130_fd_sc_hd__nor4_1
XFILLER_0_26_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2907_ _0556_ _0649_ VGND VGND VPWR VPWR _0723_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_269 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2838_ _0837_ _1152_ _1190_ VGND VGND VPWR VPWR _0672_ sky130_fd_sc_hd__or3_1
XFILLER_0_33_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2769_ internalDataflow.addressLowBusModule.busInputs\[22\] _0536_ VGND VGND VPWR
+ VPWR _0614_ sky130_fd_sc_hd__nor2_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xwire2 _1335_ VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__buf_1
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_247 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_63_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2623_ _1384_ _1486_ _0489_ VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__or3_1
XFILLER_0_27_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2554_ _0367_ _0425_ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1505_ demux.state_machine.currentInstruction\[1\] VGND VGND VPWR VPWR _0812_ sky130_fd_sc_hd__buf_2
XFILLER_0_2_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2485_ _0204_ _0287_ _0367_ _0368_ VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__o22ai_2
X_3037_ clknet_4_3_0_clk _0031_ net59 VGND VGND VPWR VPWR internalDataflow.stackBusModule.busInputs\[37\]
+ sky130_fd_sc_hd__dfrtp_1
X_3106_ clknet_4_9_0_clk _0098_ net63 VGND VGND VPWR VPWR internalDataflow.addressHighBusModule.busInputs\[23\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_73_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_18_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2270_ _0156_ _0157_ VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_100 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1985_ _0897_ _0912_ _0920_ _0876_ VGND VGND VPWR VPWR _1258_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2537_ _1007_ _1303_ _1202_ VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__and3_2
X_2606_ _0465_ _0466_ VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_54_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2468_ _1274_ _1454_ _0332_ VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__o21a_1
X_2399_ _0223_ _0285_ _0286_ VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__a21o_1
XFILLER_0_65_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xwire51 _1340_ VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__buf_1
XFILLER_0_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1770_ _0998_ _1052_ _1053_ VGND VGND VPWR VPWR _1054_ sky130_fd_sc_hd__and3_2
XFILLER_0_60_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2184_ _1307_ _1330_ _1456_ VGND VGND VPWR VPWR _1457_ sky130_fd_sc_hd__or3_1
X_2322_ internalDataflow.stackBusModule.busInputs\[34\] _1371_ VGND VGND VPWR VPWR
+ _0210_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2253_ internalDataflow.addressHighBusModule.busInputs\[21\] _1422_ _1424_ net7 _1431_
+ VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__o221a_1
X_1899_ _0954_ _1010_ _1040_ VGND VGND VPWR VPWR _1181_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_62_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1968_ _1240_ VGND VGND VPWR VPWR _1241_ sky130_fd_sc_hd__buf_4
XFILLER_0_47_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_47_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_114 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold5 instructionLoader.interruptInjector.nmiGeneratedFF.nmiRunning VGND VGND VPWR
+ VPWR net77 sky130_fd_sc_hd__dlygate4sd3_1
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_71_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2940_ _0751_ _0752_ VGND VGND VPWR VPWR _0753_ sky130_fd_sc_hd__xnor2_1
X_1753_ _1039_ _0957_ _0956_ VGND VGND VPWR VPWR _1040_ sky130_fd_sc_hd__and3_1
X_1822_ _0972_ _1047_ _1101_ _1105_ VGND VGND VPWR VPWR _1106_ sky130_fd_sc_hd__a211o_1
XFILLER_0_44_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2871_ _0692_ VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1684_ _0932_ _0875_ VGND VGND VPWR VPWR _0986_ sky130_fd_sc_hd__nor2_1
XFILLER_0_52_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2167_ _0930_ _1358_ _1005_ VGND VGND VPWR VPWR _1440_ sky130_fd_sc_hd__o21ai_1
X_2236_ _1484_ _1488_ _0118_ VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_17_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2305_ _0187_ _0191_ _0192_ net47 VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_35_117 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2098_ _1370_ VGND VGND VPWR VPWR _1371_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_43_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2021_ _1293_ VGND VGND VPWR VPWR _1294_ sky130_fd_sc_hd__buf_2
X_3070_ clknet_4_11_0_clk _0062_ net65 VGND VGND VPWR VPWR internalDataflow.addressLowBusModule.busInputs\[20\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_17_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2923_ _0737_ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1736_ demux.state_machine.currentAddress\[0\] _1027_ _0979_ VGND VGND VPWR VPWR
+ _1028_ sky130_fd_sc_hd__mux2_1
X_1805_ _1084_ _1085_ _0975_ _1087_ _1088_ VGND VGND VPWR VPWR _1089_ sky130_fd_sc_hd__a32o_1
XFILLER_0_40_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2785_ _0626_ _0627_ _0544_ VGND VGND VPWR VPWR _0629_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2854_ net100 _1434_ _0675_ VGND VGND VPWR VPWR _0682_ sky130_fd_sc_hd__mux2_1
X_1667_ _0967_ _0970_ VGND VGND VPWR VPWR _0971_ sky130_fd_sc_hd__and2_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1598_ _0904_ VGND VGND VPWR VPWR _0905_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_378 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2219_ demux.state_machine.timeState\[5\] _0945_ _1084_ _0891_ VGND VGND VPWR VPWR
+ _1492_ sky130_fd_sc_hd__o211a_1
XFILLER_0_63_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_48_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2570_ _0181_ _0366_ _0369_ VGND VGND VPWR VPWR _0441_ sky130_fd_sc_hd__and3_1
X_1521_ _0815_ _0825_ _0827_ VGND VGND VPWR VPWR _0828_ sky130_fd_sc_hd__a21oi_1
X_3122_ clknet_4_5_0_clk _0110_ net69 VGND VGND VPWR VPWR negEdgeDetector.q1 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2004_ _0897_ _0913_ _1274_ _1276_ VGND VGND VPWR VPWR _1277_ sky130_fd_sc_hd__a211o_1
X_3053_ clknet_4_8_0_clk _0045_ net62 VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2906_ _0556_ _0649_ VGND VGND VPWR VPWR _0722_ sky130_fd_sc_hd__and2_1
XFILLER_0_9_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1719_ _0969_ _1013_ VGND VGND VPWR VPWR _1014_ sky130_fd_sc_hd__nor2_1
X_2837_ instructionLoader.interruptInjector.resetDetected _0999_ _0671_ demux.reset
+ VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__a22o_1
X_2699_ _0521_ _0533_ _0548_ VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__a21oi_1
X_2768_ internalDataflow.addressLowBusModule.busInputs\[22\] _0535_ VGND VGND VPWR
+ VPWR _0613_ sky130_fd_sc_hd__and2_1
XFILLER_0_67_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_42 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2622_ _0877_ _0921_ _1244_ _0839_ _1399_ VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__a221o_1
X_1504_ demux.state_machine.currentInstruction\[3\] VGND VGND VPWR VPWR _0811_ sky130_fd_sc_hd__buf_2
XFILLER_0_42_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2553_ _0367_ _0425_ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__and2_1
XFILLER_0_12_64 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3105_ clknet_4_10_0_clk _0097_ net64 VGND VGND VPWR VPWR internalDataflow.addressHighBusModule.busInputs\[22\]
+ sky130_fd_sc_hd__dfrtp_4
X_2484_ _0223_ _0285_ VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__xor2_4
XFILLER_0_65_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3036_ clknet_4_2_0_clk _0030_ net58 VGND VGND VPWR VPWR internalDataflow.stackBusModule.busInputs\[36\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_351 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_2_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_2_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_18_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1984_ _1256_ VGND VGND VPWR VPWR _1257_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_15_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2467_ _0276_ _0236_ _0349_ _0351_ VGND VGND VPWR VPWR internalDataflow.psr.processStatusReg.stat_buf_nxt\[1\]
+ sky130_fd_sc_hd__o31ai_1
XFILLER_0_30_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2605_ _0425_ _0469_ VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__or2_1
X_2536_ _0275_ _0364_ _0408_ _0251_ _0410_ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__a221o_1
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2398_ _0216_ _0222_ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__and2_1
X_3019_ clknet_4_7_0_clk _0000_ net68 VGND VGND VPWR VPWR demux.state_machine.currentAddress\[0\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_65_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2321_ internalDataflow.stackBusModule.busInputs\[42\] _1373_ _1374_ internalDataflow.accRegToDB\[2\]
+ _1375_ VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2183_ _1357_ _1249_ _1455_ _1004_ VGND VGND VPWR VPWR _1456_ sky130_fd_sc_hd__o31a_1
X_2252_ _0137_ _0139_ _1372_ VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__o21a_1
XFILLER_0_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1967_ demux.isAddressing _0947_ VGND VGND VPWR VPWR _1240_ sky130_fd_sc_hd__and2_1
X_1898_ _0901_ _0825_ _0978_ VGND VGND VPWR VPWR _1180_ sky130_fd_sc_hd__nor3_1
XFILLER_0_50_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2519_ _0397_ VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_46_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_126 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold6 demux.state_machine.currentAddress\[2\] VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_71_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2870_ internalDataflow.addressLowBusModule.busInputs\[36\] _0170_ _0687_ VGND VGND
+ VPWR VPWR _0692_ sky130_fd_sc_hd__mux2_1
X_1752_ net4 VGND VGND VPWR VPWR _1039_ sky130_fd_sc_hd__inv_2
X_1821_ _0890_ _0891_ _0976_ _1104_ VGND VGND VPWR VPWR _1105_ sky130_fd_sc_hd__a31o_1
X_1683_ _0984_ VGND VGND VPWR VPWR _0985_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_40_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2304_ internalDataflow.addressHighBusModule.busInputs\[19\] _1422_ _1424_ _0957_
+ _1431_ VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__o221a_1
X_2166_ branch_ff.branchForward _1290_ VGND VGND VPWR VPWR _1439_ sky130_fd_sc_hd__nand2_1
X_2235_ _1425_ _0122_ VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__nand2b_2
X_2097_ _1366_ _1368_ _1369_ VGND VGND VPWR VPWR _1370_ sky130_fd_sc_hd__and3b_1
XFILLER_0_63_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2999_ demux.nmi _0671_ VGND VGND VPWR VPWR _0797_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_287 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_66_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2020_ _0952_ _1262_ _1289_ _1292_ VGND VGND VPWR VPWR _1293_ sky130_fd_sc_hd__and4_1
XFILLER_0_45_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2853_ _0681_ VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_15_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2922_ _0736_ internalDataflow.addressHighBusModule.busInputs\[19\] _0554_ VGND VGND
+ VPWR VPWR _0737_ sky130_fd_sc_hd__mux2_1
X_1735_ _1023_ _1025_ _1026_ VGND VGND VPWR VPWR _1027_ sky130_fd_sc_hd__a21oi_1
X_1804_ _1034_ _1052_ VGND VGND VPWR VPWR _1088_ sky130_fd_sc_hd__and2_2
X_1666_ _0968_ _0969_ _0956_ VGND VGND VPWR VPWR _0970_ sky130_fd_sc_hd__and3_1
XFILLER_0_40_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2784_ _0626_ _0627_ VGND VGND VPWR VPWR _0628_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1597_ _0902_ _0903_ VGND VGND VPWR VPWR _0904_ sky130_fd_sc_hd__nand2_2
XFILLER_0_0_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2218_ _0917_ _0937_ VGND VGND VPWR VPWR _1491_ sky130_fd_sc_hd__nand2_1
X_2149_ _1407_ _1408_ _1410_ _1418_ _1421_ VGND VGND VPWR VPWR _1422_ sky130_fd_sc_hd__a311o_4
XFILLER_0_63_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1520_ _0826_ VGND VGND VPWR VPWR _0827_ sky130_fd_sc_hd__buf_4
XFILLER_0_42_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3121_ clknet_4_13_0_clk _0109_ net70 VGND VGND VPWR VPWR demux.setInterruptFlag
+ sky130_fd_sc_hd__dfrtp_1
X_2003_ _0896_ _0939_ _1275_ VGND VGND VPWR VPWR _1276_ sky130_fd_sc_hd__and3_1
X_3052_ clknet_4_1_0_clk _0044_ net61 VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_45_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2836_ instructionLoader.interruptInjector.processStatusRegIFlag demux.setInterruptFlag
+ _0961_ VGND VGND VPWR VPWR _0671_ sky130_fd_sc_hd__or3_1
X_2905_ _0711_ _0719_ _0718_ _0546_ VGND VGND VPWR VPWR _0721_ sky130_fd_sc_hd__o31a_1
XFILLER_0_9_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1718_ _1012_ net55 VGND VGND VPWR VPWR _1013_ sky130_fd_sc_hd__nand2_2
X_2698_ internalDataflow.addressLowBusModule.busInputs\[17\] VGND VGND VPWR VPWR _0548_
+ sky130_fd_sc_hd__inv_2
X_2767_ _0130_ _0611_ VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__xor2_1
XFILLER_0_13_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1649_ net6 VGND VGND VPWR VPWR _0954_ sky130_fd_sc_hd__buf_4
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_18 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1503_ demux.state_machine.currentInstruction\[2\] VGND VGND VPWR VPWR _0810_ sky130_fd_sc_hd__clkbuf_2
X_2621_ _0483_ _0484_ _0485_ _0487_ VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__or4_1
X_2552_ _1466_ _0325_ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2483_ _0262_ _0283_ VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__xor2_4
XFILLER_0_37_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3035_ clknet_4_2_0_clk _0029_ net58 VGND VGND VPWR VPWR internalDataflow.stackBusModule.busInputs\[35\]
+ sky130_fd_sc_hd__dfrtp_1
X_3104_ clknet_4_10_0_clk _0096_ net64 VGND VGND VPWR VPWR internalDataflow.addressHighBusModule.busInputs\[21\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_73_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_140 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2819_ _0163_ _0632_ _0633_ _0162_ VGND VGND VPWR VPWR _0658_ sky130_fd_sc_hd__a22o_1
XTAP_190 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_322 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1983_ _1242_ _1252_ _1255_ _0998_ VGND VGND VPWR VPWR _1256_ sky130_fd_sc_hd__o211a_1
X_2604_ net129 net45 _0464_ _0472_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2466_ _0276_ _0333_ _0348_ _0350_ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__o2bb2a_1
X_2535_ _0409_ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__buf_2
XFILLER_0_64_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xwire53 _0895_ VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__dlymetal6s2s_1
X_3018_ _0809_ VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__clkbuf_1
X_2397_ _0262_ _0283_ _0284_ VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__a21o_2
XFILLER_0_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2251_ internalDataflow.stackBusModule.busInputs\[37\] _1371_ _0138_ VGND VGND VPWR
+ VPWR _0139_ sky130_fd_sc_hd__a21o_1
X_2320_ _1257_ _0207_ VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__nor2_1
X_2182_ _1161_ _1131_ _0915_ VGND VGND VPWR VPWR _1455_ sky130_fd_sc_hd__or3_1
Xclkbuf_4_1_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_1_0_clk sky130_fd_sc_hd__clkbuf_8
X_1966_ _0844_ _0815_ _0818_ _0901_ _0917_ VGND VGND VPWR VPWR _1239_ sky130_fd_sc_hd__a311oi_2
XFILLER_0_34_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1897_ _1179_ VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_71 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2449_ _0332_ _0327_ VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__nand2_1
X_2518_ net114 _0170_ _0392_ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_263 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold7 net25 VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_71_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1820_ _1102_ _0978_ _1103_ VGND VGND VPWR VPWR _1104_ sky130_fd_sc_hd__o21a_1
XFILLER_0_29_127 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1751_ net81 _0979_ _1038_ VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__o21a_1
X_1682_ demux.state_machine.currentAddress\[4\] demux.state_machine.currentAddress\[10\]
+ VGND VGND VPWR VPWR _0984_ sky130_fd_sc_hd__or2_1
XFILLER_0_52_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2234_ _1502_ _0119_ _0121_ VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__nor3b_4
X_2303_ _0188_ _0190_ _1372_ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_48_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2165_ _1006_ _1436_ _1437_ VGND VGND VPWR VPWR _1438_ sky130_fd_sc_hd__a21bo_1
X_2096_ _0997_ _1346_ _1349_ _1335_ VGND VGND VPWR VPWR _1369_ sky130_fd_sc_hd__a31o_1
X_1949_ _1029_ _1036_ _1133_ _1011_ VGND VGND VPWR VPWR _1228_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_63_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2998_ _0796_ VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_16_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1803_ _0967_ _1086_ VGND VGND VPWR VPWR _1087_ sky130_fd_sc_hd__nor2_2
XFILLER_0_45_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2783_ _0615_ _0617_ _0613_ VGND VGND VPWR VPWR _0627_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_25_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2852_ net103 _0146_ _0675_ VGND VGND VPWR VPWR _0681_ sky130_fd_sc_hd__mux2_1
X_2921_ _0730_ _0735_ _0553_ VGND VGND VPWR VPWR _0736_ sky130_fd_sc_hd__mux2_1
X_1734_ net3 _0956_ VGND VGND VPWR VPWR _1026_ sky130_fd_sc_hd__nand2_2
X_1665_ net8 VGND VGND VPWR VPWR _0969_ sky130_fd_sc_hd__buf_2
X_1596_ _0885_ _0855_ _0860_ _0852_ _0901_ VGND VGND VPWR VPWR _0903_ sky130_fd_sc_hd__a41o_1
XFILLER_0_40_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2217_ _1427_ _1489_ _1310_ VGND VGND VPWR VPWR _1490_ sky130_fd_sc_hd__a21o_1
XFILLER_0_22_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2079_ branch_ff.branchForward branch_ff.branchBackward VGND VGND VPWR VPWR _1352_
+ sky130_fd_sc_hd__or2_1
X_2148_ _1384_ _1419_ _1420_ _0960_ VGND VGND VPWR VPWR _1421_ sky130_fd_sc_hd__a31o_1
XFILLER_0_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_341 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3120_ clknet_4_14_0_clk _0108_ net71 VGND VGND VPWR VPWR demux.nmi sky130_fd_sc_hd__dfrtp_4
X_3051_ clknet_4_0_0_clk _0043_ net57 VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dfrtp_1
X_2002_ _0835_ _0834_ _0833_ _0832_ VGND VGND VPWR VPWR _1275_ sky130_fd_sc_hd__and4b_1
XFILLER_0_9_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2835_ _0670_ VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2766_ _0605_ _0609_ _0610_ VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__and3_1
X_2904_ _0711_ _0718_ _0719_ VGND VGND VPWR VPWR _0720_ sky130_fd_sc_hd__o21ai_1
X_1717_ net9 VGND VGND VPWR VPWR _1012_ sky130_fd_sc_hd__clkbuf_4
X_1579_ demux.PSR_Z _0869_ _0885_ VGND VGND VPWR VPWR _0886_ sky130_fd_sc_hd__or3_1
X_1648_ _0953_ VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_2
X_2697_ internalDataflow.addressLowBusModule.busInputs\[16\] VGND VGND VPWR VPWR _0547_
+ sky130_fd_sc_hd__inv_2
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2620_ _1001_ _1094_ _1394_ _0486_ VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__a211o_1
XFILLER_0_42_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2551_ _0421_ _0422_ _0423_ _0368_ _0361_ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__o32a_1
X_2482_ _0204_ _0287_ _0202_ VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__a21oi_1
X_3034_ clknet_4_8_0_clk _0028_ net62 VGND VGND VPWR VPWR internalDataflow.stackBusModule.busInputs\[34\]
+ sky130_fd_sc_hd__dfrtp_1
X_3103_ clknet_4_10_0_clk _0095_ net64 VGND VGND VPWR VPWR internalDataflow.addressHighBusModule.busInputs\[20\]
+ sky130_fd_sc_hd__dfrtp_4
X_2749_ _0177_ _0595_ VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_5_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2818_ _0657_ VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__clkbuf_1
XTAP_191 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1982_ _1253_ _1254_ VGND VGND VPWR VPWR _1255_ sky130_fd_sc_hd__nand2_1
XFILLER_0_23_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2534_ _1007_ _1303_ _1271_ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__and3_1
X_2603_ _0470_ _0321_ _0471_ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__or3b_1
XFILLER_0_15_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2465_ demux.PSR_Z _0336_ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__nand2_1
X_2396_ _0275_ _0282_ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__and2_1
XFILLER_0_38_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3017_ demux.PSR_N _0308_ _0808_ VGND VGND VPWR VPWR _0809_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_69_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2250_ internalDataflow.addressLowBusModule.busInputs\[29\] _1377_ _1378_ internalDataflow.addressLowBusModule.busInputs\[37\]
+ VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__a22o_1
X_2181_ _1264_ _1279_ _1452_ _1453_ VGND VGND VPWR VPWR _1454_ sky130_fd_sc_hd__or4_1
XFILLER_0_34_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1965_ _0844_ _0882_ _0852_ _0871_ _0917_ VGND VGND VPWR VPWR _1238_ sky130_fd_sc_hd__a311oi_2
XFILLER_0_43_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1896_ _1100_ _1178_ VGND VGND VPWR VPWR _1179_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2517_ _0396_ VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_52_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2448_ _0982_ _0334_ _0819_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__a21o_1
X_2379_ internalDataflow.stackBusModule.busInputs\[41\] _1373_ _1374_ internalDataflow.accRegToDB\[1\]
+ VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xhold8 internalDataflow.addressLowBusModule.busInputs\[24\] VGND VGND VPWR VPWR net80
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1750_ _1029_ _1037_ _0979_ VGND VGND VPWR VPWR _1038_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_29_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1681_ _0897_ VGND VGND VPWR VPWR _0983_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_40_348 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2164_ _0987_ _0993_ _0982_ VGND VGND VPWR VPWR _1437_ sky130_fd_sc_hd__a21oi_1
X_2233_ _0120_ _1500_ VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__or2_1
X_2302_ internalDataflow.stackBusModule.busInputs\[35\] _1371_ _0189_ VGND VGND VPWR
+ VPWR _0190_ sky130_fd_sc_hd__a21o_1
XFILLER_0_61_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2095_ net135 _1341_ VGND VGND VPWR VPWR _1368_ sky130_fd_sc_hd__and2b_1
X_1879_ _1161_ _1067_ _1019_ _1095_ _1142_ VGND VGND VPWR VPWR _1162_ sky130_fd_sc_hd__a221o_1
X_1948_ _1061_ _1132_ _1145_ _1163_ VGND VGND VPWR VPWR _1227_ sky130_fd_sc_hd__or4_1
XFILLER_0_63_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2997_ net14 net89 _0981_ VGND VGND VPWR VPWR _0796_ sky130_fd_sc_hd__mux2_1
XFILLER_0_43_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_378 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xclkbuf_4_0_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_0_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_66_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2920_ _0733_ _0734_ VGND VGND VPWR VPWR _0735_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1802_ _1022_ _1012_ _0969_ VGND VGND VPWR VPWR _1086_ sky130_fd_sc_hd__or3b_1
X_1733_ _1013_ _1024_ VGND VGND VPWR VPWR _1025_ sky130_fd_sc_hd__nand2_1
XFILLER_0_57_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_45_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2782_ _0624_ _0625_ VGND VGND VPWR VPWR _0626_ sky130_fd_sc_hd__nand2_1
X_2851_ _0680_ VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_17_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1595_ _0857_ _0882_ _0825_ _0865_ _0901_ VGND VGND VPWR VPWR _0902_ sky130_fd_sc_hd__a41o_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1664_ net9 VGND VGND VPWR VPWR _0968_ sky130_fd_sc_hd__inv_2
XFILLER_0_0_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2216_ _1003_ demux.state_machine.timeState\[1\] _1102_ VGND VGND VPWR VPWR _1489_
+ sky130_fd_sc_hd__o21ai_2
X_2147_ demux.state_machine.currentAddress\[7\] _0985_ _1004_ VGND VGND VPWR VPWR
+ _1420_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_15_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2078_ _1336_ _1337_ _0982_ VGND VGND VPWR VPWR _1351_ sky130_fd_sc_hd__o21a_1
XFILLER_0_8_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_8_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2001_ _0815_ _0818_ _0825_ _0866_ _1273_ VGND VGND VPWR VPWR _1274_ sky130_fd_sc_hd__a311oi_4
X_3050_ clknet_4_4_0_clk _0042_ net60 VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__dfrtp_1
XFILLER_0_42_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2903_ internalDataflow.addressHighBusModule.busInputs\[18\] _0556_ VGND VGND VPWR
+ VPWR _0719_ sky130_fd_sc_hd__xor2_1
X_1716_ _0957_ _0954_ _1010_ net4 VGND VGND VPWR VPWR _1011_ sky130_fd_sc_hd__and4b_1
XFILLER_0_60_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2834_ net121 _0669_ _0645_ VGND VGND VPWR VPWR _0670_ sky130_fd_sc_hd__mux2_1
X_2696_ _0538_ _0543_ VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__nor2_4
X_2765_ _0153_ _0558_ VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__nand2_1
X_1578_ _0884_ VGND VGND VPWR VPWR _0885_ sky130_fd_sc_hd__clkbuf_4
X_1647_ _0878_ _0906_ _0935_ _0952_ VGND VGND VPWR VPWR _0953_ sky130_fd_sc_hd__o31a_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_150 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_44_292 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2550_ _0195_ _0364_ _0410_ _0286_ _0406_ VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__a221o_1
XFILLER_0_50_273 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2481_ _0250_ _0364_ VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3033_ clknet_4_2_0_clk _0027_ net58 VGND VGND VPWR VPWR internalDataflow.stackBusModule.busInputs\[33\]
+ sky130_fd_sc_hd__dfrtp_1
X_3102_ clknet_4_11_0_clk _0094_ net64 VGND VGND VPWR VPWR internalDataflow.addressHighBusModule.busInputs\[19\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_58_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_96 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_204 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2679_ _0877_ _0933_ VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__and2_1
X_2748_ _0200_ _0221_ _0522_ _0562_ VGND VGND VPWR VPWR _0595_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_5_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2817_ net91 _0656_ _0645_ VGND VGND VPWR VPWR _0657_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_192 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1981_ _1077_ _1173_ _0995_ VGND VGND VPWR VPWR _1254_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2533_ _1007_ _0332_ _1131_ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__and3_2
X_2602_ _0376_ _0469_ _0468_ _0450_ VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__a211o_1
XFILLER_0_23_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_6 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2464_ _1482_ _0344_ _0308_ _0348_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__or4b_1
X_2395_ _0275_ _0282_ VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__xor2_4
Xwire55 _0955_ VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_2
X_3016_ _0806_ _0347_ _0807_ _0332_ VGND VGND VPWR VPWR _0808_ sky130_fd_sc_hd__o31a_1
XFILLER_0_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2180_ _1004_ _0868_ VGND VGND VPWR VPWR _1453_ sky130_fd_sc_hd__and2_1
XFILLER_0_18_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_129 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1895_ _1160_ _1165_ _1172_ _1177_ VGND VGND VPWR VPWR _1178_ sky130_fd_sc_hd__or4_1
X_1964_ _0909_ _0885_ _0865_ _0852_ _0821_ VGND VGND VPWR VPWR _1237_ sky130_fd_sc_hd__a41oi_4
XFILLER_0_43_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2447_ demux.state_machine.timeState\[5\] demux.setInterruptFlag _1079_ VGND VGND
+ VPWR VPWR _0334_ sky130_fd_sc_hd__and3_1
X_2516_ net106 _0194_ _0392_ VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2378_ _1257_ _0265_ VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_143 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xhold9 demux.state_machine.currentAddress\[4\] VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_69_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1680_ _0948_ VGND VGND VPWR VPWR _0982_ sky130_fd_sc_hd__buf_4
X_2301_ internalDataflow.addressLowBusModule.busInputs\[27\] _1377_ _1378_ internalDataflow.addressLowBusModule.busInputs\[35\]
+ VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__a22o_1
X_2163_ _0988_ demux.state_machine.currentAddress\[4\] demux.state_machine.currentAddress\[10\]
+ _1435_ VGND VGND VPWR VPWR _1436_ sky130_fd_sc_hd__or4_1
X_2232_ _1427_ _1489_ _1310_ VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_0_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2094_ _1342_ _1350_ _1366_ VGND VGND VPWR VPWR _1367_ sky130_fd_sc_hd__mux2_1
X_1947_ _1110_ _1193_ _1194_ _1215_ VGND VGND VPWR VPWR _1226_ sky130_fd_sc_hd__or4_1
X_1878_ _0901_ _0818_ VGND VGND VPWR VPWR _1161_ sky130_fd_sc_hd__nor2_2
X_2996_ _0341_ _0795_ VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_162 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2850_ net107 _0170_ _0675_ VGND VGND VPWR VPWR _0680_ sky130_fd_sc_hd__mux2_1
XFILLER_0_15_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1663_ net7 VGND VGND VPWR VPWR _0967_ sky130_fd_sc_hd__clkbuf_4
X_1732_ _0957_ _0954_ _0956_ net4 VGND VGND VPWR VPWR _1024_ sky130_fd_sc_hd__and4bb_2
X_1801_ _0819_ _0820_ VGND VGND VPWR VPWR _1085_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2781_ internalDataflow.addressLowBusModule.busInputs\[23\] _0558_ VGND VGND VPWR
+ VPWR _0625_ sky130_fd_sc_hd__nand2_1
XFILLER_0_25_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_56_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1594_ _0869_ VGND VGND VPWR VPWR _0901_ sky130_fd_sc_hd__buf_4
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_210 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2215_ _1403_ _1487_ _1406_ _1405_ VGND VGND VPWR VPWR _1488_ sky130_fd_sc_hd__or4bb_2
X_2146_ demux.state_machine.currentAddress\[6\] _1283_ VGND VGND VPWR VPWR _1419_
+ sky130_fd_sc_hd__nand2_1
X_2077_ _0998_ _1346_ _1349_ net49 VGND VGND VPWR VPWR _1350_ sky130_fd_sc_hd__a31oi_4
XFILLER_0_48_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2979_ _0786_ VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2000_ _1268_ VGND VGND VPWR VPWR _1273_ sky130_fd_sc_hd__buf_4
XFILLER_0_45_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2902_ _0709_ _0700_ _0710_ VGND VGND VPWR VPWR _0718_ sky130_fd_sc_hd__a21oi_1
X_2833_ _0667_ _0632_ _0634_ _0304_ _0668_ VGND VGND VPWR VPWR _0669_ sky130_fd_sc_hd__a221o_2
X_1715_ _0956_ VGND VGND VPWR VPWR _1010_ sky130_fd_sc_hd__clkbuf_4
X_1646_ net13 _0950_ pulse_slower.nextEnableState\[0\] _0948_ VGND VGND VPWR VPWR
+ _0952_ sky130_fd_sc_hd__o211a_1
X_2695_ _0538_ _0545_ VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__xnor2_1
X_2764_ _0153_ _0176_ _0592_ _0558_ VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__a31o_1
XFILLER_0_5_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1577_ _0812_ _0810_ _0811_ _0813_ VGND VGND VPWR VPWR _0884_ sky130_fd_sc_hd__or4bb_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2129_ _0879_ _0912_ _0922_ _1399_ _1401_ VGND VGND VPWR VPWR _1402_ sky130_fd_sc_hd__a2111o_1
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2480_ _1121_ _1144_ _0363_ _0323_ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__o31a_4
XFILLER_0_50_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_10_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3101_ clknet_4_11_0_clk _0093_ net66 VGND VGND VPWR VPWR internalDataflow.addressHighBusModule.busInputs\[18\]
+ sky130_fd_sc_hd__dfrtp_4
X_3032_ clknet_4_3_0_clk _0026_ net60 VGND VGND VPWR VPWR internalDataflow.stackBusModule.busInputs\[32\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_58_385 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2816_ _0185_ _0634_ _0655_ VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__a21o_1
X_1629_ _0896_ demux.state_machine.timeState\[6\] VGND VGND VPWR VPWR _0936_ sky130_fd_sc_hd__or2_4
X_2678_ _1005_ _0985_ VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__nand2_1
X_2747_ _0177_ _0592_ VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_193 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_377 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1980_ _0988_ _0993_ _0948_ VGND VGND VPWR VPWR _1253_ sky130_fd_sc_hd__a21oi_1
X_2463_ _1359_ _0347_ _0332_ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__o21a_1
X_2532_ _1271_ _0323_ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__nand2_2
X_2601_ _0450_ _0468_ _0469_ _0376_ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__o211a_1
XFILLER_0_2_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3015_ _1002_ _0847_ _0328_ VGND VGND VPWR VPWR _0807_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2394_ _0277_ _0281_ _0154_ VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__mux2_2
XFILLER_0_58_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xwire45 _0403_ VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__buf_2
XFILLER_0_73_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_52_325 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1894_ _0847_ _0976_ _1019_ _1063_ _1176_ VGND VGND VPWR VPWR _1177_ sky130_fd_sc_hd__a221o_1
XFILLER_0_50_54 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1963_ _1236_ VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__buf_1
XFILLER_0_28_344 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2446_ _0332_ _0327_ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__and2_1
X_2515_ _0395_ VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2377_ internalDataflow.addressLowBusModule.busInputs\[17\] _1315_ _0263_ _0264_
+ net48 VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_34_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_61_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_155 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_369 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2231_ _1484_ _1488_ _1490_ _0118_ VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__a211oi_2
X_2300_ internalDataflow.stackBusModule.busInputs\[43\] _1373_ _1374_ internalDataflow.accRegToDB\[3\]
+ _1375_ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__a221o_1
X_2162_ demux.state_machine.currentAddress\[11\] demux.state_machine.currentAddress\[3\]
+ VGND VGND VPWR VPWR _1435_ sky130_fd_sc_hd__or2_1
XFILLER_0_45_98 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2093_ _1351_ _1365_ _0998_ VGND VGND VPWR VPWR _1366_ sky130_fd_sc_hd__o21a_2
X_2995_ _0999_ _1022_ net92 VGND VGND VPWR VPWR _0795_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_28_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1877_ _1154_ _1155_ _1157_ _1159_ VGND VGND VPWR VPWR _1160_ sky130_fd_sc_hd__or4_1
X_1946_ _1192_ _1201_ _1217_ VGND VGND VPWR VPWR _1225_ sky130_fd_sc_hd__or3_1
XFILLER_0_43_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2429_ _0306_ _0314_ VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__and2_1
XFILLER_0_66_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1800_ _0834_ _0835_ _0832_ _0833_ VGND VGND VPWR VPWR _1084_ sky130_fd_sc_hd__and4b_4
XFILLER_0_15_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1731_ net4 _0954_ _1022_ _0957_ VGND VGND VPWR VPWR _1023_ sky130_fd_sc_hd__or4b_2
X_1662_ _0965_ VGND VGND VPWR VPWR _0966_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_40_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_40_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2780_ internalDataflow.addressLowBusModule.busInputs\[23\] _0535_ VGND VGND VPWR
+ VPWR _0624_ sky130_fd_sc_hd__or2_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2214_ _0905_ _1485_ _1486_ VGND VGND VPWR VPWR _1487_ sky130_fd_sc_hd__a21o_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1593_ _0877_ _0888_ net53 _0899_ VGND VGND VPWR VPWR _0900_ sky130_fd_sc_hd__a31o_1
XFILLER_0_0_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2076_ _1347_ _1348_ demux.state_machine.currentAddress\[3\] _0948_ VGND VGND VPWR
+ VPWR _1349_ sky130_fd_sc_hd__a211o_2
XFILLER_0_56_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2145_ _1384_ _1381_ _1412_ _1417_ _0998_ VGND VGND VPWR VPWR _1418_ sky130_fd_sc_hd__o311a_2
XFILLER_0_48_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1929_ _1057_ _1073_ _1106_ _1209_ VGND VGND VPWR VPWR _1210_ sky130_fd_sc_hd__or4_1
X_2978_ net34 _0217_ _0783_ VGND VGND VPWR VPWR _0786_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_291 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_60_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2901_ _0717_ VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__clkbuf_1
X_2832_ _0296_ _0654_ VGND VGND VPWR VPWR _0668_ sky130_fd_sc_hd__nor2_1
X_2763_ net133 _0555_ _0603_ _0546_ _0608_ VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__a221o_1
XFILLER_0_18_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1714_ _1008_ _0999_ _1009_ net84 VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__o22a_1
X_1576_ _0819_ _0882_ _0820_ demux.PSR_N VGND VGND VPWR VPWR _0883_ sky130_fd_sc_hd__or4b_1
X_1645_ _0951_ VGND VGND VPWR VPWR pulse_slower.nextEnableState\[0\] sky130_fd_sc_hd__inv_2
X_2694_ internalDataflow.addressLowBusModule.busInputs\[16\] _0241_ _0544_ VGND VGND
+ VPWR VPWR _0545_ sky130_fd_sc_hd__mux2_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2128_ _0839_ _1243_ _1400_ _1071_ _1240_ VGND VGND VPWR VPWR _1401_ sky130_fd_sc_hd__a221o_1
X_2059_ _1173_ _0995_ _1331_ _1273_ VGND VGND VPWR VPWR _1332_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_36_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_412 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3031_ clknet_4_7_0_clk _0003_ net67 VGND VGND VPWR VPWR demux.state_machine.currentAddress\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_37_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3100_ clknet_4_13_0_clk _0092_ net66 VGND VGND VPWR VPWR internalDataflow.addressHighBusModule.busInputs\[17\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_58_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2746_ _0176_ _0592_ _0558_ VGND VGND VPWR VPWR _0593_ sky130_fd_sc_hd__a21o_1
XFILLER_0_14_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2815_ _0191_ _0654_ _0632_ _0192_ VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_18_228 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1559_ _0827_ VGND VGND VPWR VPWR _0866_ sky130_fd_sc_hd__buf_4
X_2677_ _1392_ _0525_ _0490_ _0527_ VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__or4_1
X_1628_ _0877_ _0911_ _0925_ _0931_ _0934_ VGND VGND VPWR VPWR _0935_ sky130_fd_sc_hd__a2111o_1
XFILLER_0_41_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_361 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2600_ _0375_ _0372_ _0373_ VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__nand3_1
XFILLER_0_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2462_ _1008_ _0840_ _0345_ _0346_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__a211o_1
X_2393_ internalDataflow.addressLowBusModule.busInputs\[17\] _1502_ _0278_ _0280_
+ VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__a211o_2
X_2531_ _0361_ VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__inv_2
XFILLER_0_64_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3014_ _0915_ _1249_ _1358_ _1002_ VGND VGND VPWR VPWR _0806_ sky130_fd_sc_hd__o31a_1
XFILLER_0_61_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_389 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_275 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2729_ _0568_ _0569_ VGND VGND VPWR VPWR _0577_ sky130_fd_sc_hd__and2_1
XFILLER_0_56_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_367 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_381 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1962_ clknet_4_4_0_clk pulse_slower.nextEnableState\[0\] VGND VGND VPWR VPWR _1236_
+ sky130_fd_sc_hd__and2_2
XFILLER_0_28_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_70_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1893_ _1173_ _1091_ _1060_ _1112_ _1175_ VGND VGND VPWR VPWR _1176_ sky130_fd_sc_hd__a221o_1
XFILLER_0_50_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2445_ _1303_ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__clkbuf_4
X_2376_ net3 _1313_ _1302_ _1294_ internalDataflow.addressHighBusModule.busInputs\[17\]
+ VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__a32o_1
X_2514_ net93 _0215_ _0392_ VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2230_ _0961_ _1498_ VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_23 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2092_ _1356_ _1359_ _1363_ _1295_ _1364_ VGND VGND VPWR VPWR _1365_ sky130_fd_sc_hd__o32a_1
X_2161_ _1322_ _1326_ _1329_ _1433_ VGND VGND VPWR VPWR _1434_ sky130_fd_sc_hd__o2bb2a_2
X_1945_ _1224_ VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__clkbuf_1
X_2994_ demux.nmi _0792_ _0794_ VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_1876_ _0921_ _1067_ _1048_ _1081_ _1158_ VGND VGND VPWR VPWR _1159_ sky130_fd_sc_hd__a221o_1
XFILLER_0_43_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2428_ _0292_ _0315_ VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__nand2_1
X_2359_ internalDataflow.addressHighBusModule.busInputs\[16\] _1422_ VGND VGND VPWR
+ VPWR _0247_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1661_ _0963_ _0964_ VGND VGND VPWR VPWR _0965_ sky130_fd_sc_hd__and2_1
X_1730_ demux.nmi instructionLoader.interruptInjector.resetDetected instructionLoader.interruptInjector.irqGenerated
+ VGND VGND VPWR VPWR _1022_ sky130_fd_sc_hd__or3_4
X_1592_ _0897_ _0898_ VGND VGND VPWR VPWR _0899_ sky130_fd_sc_hd__and2_1
XFILLER_0_25_189 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2144_ demux.state_machine.currentAddress\[7\] _0993_ _0989_ _0988_ _1416_ VGND VGND
+ VPWR VPWR _1417_ sky130_fd_sc_hd__a221o_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2213_ _0891_ _1275_ _1244_ VGND VGND VPWR VPWR _1486_ sky130_fd_sc_hd__and3_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2075_ demux.state_machine.currentAddress\[5\] _1077_ demux.state_machine.currentAddress\[10\]
+ _1273_ VGND VGND VPWR VPWR _1348_ sky130_fd_sc_hd__a211o_1
XFILLER_0_48_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_71_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1928_ _1047_ _1095_ _1175_ _1208_ _1083_ VGND VGND VPWR VPWR _1209_ sky130_fd_sc_hd__a2111o_1
X_1859_ _0901_ _0844_ VGND VGND VPWR VPWR _1143_ sky130_fd_sc_hd__nor2_2
XFILLER_0_44_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2977_ _0785_ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2900_ _0716_ internalDataflow.addressHighBusModule.busInputs\[17\] _0554_ VGND VGND
+ VPWR VPWR _0717_ sky130_fd_sc_hd__mux2_1
X_1713_ _1000_ VGND VGND VPWR VPWR _1009_ sky130_fd_sc_hd__inv_2
XFILLER_0_26_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2831_ _0299_ VGND VGND VPWR VPWR _0667_ sky130_fd_sc_hd__inv_2
X_2762_ _0553_ _0607_ VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__nor2_1
XFILLER_0_5_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1575_ _0881_ VGND VGND VPWR VPWR _0882_ sky130_fd_sc_hd__buf_4
X_1644_ pulse_slower.currentEnableState\[1\] pulse_slower.currentEnableState\[0\]
+ VGND VGND VPWR VPWR _0951_ sky130_fd_sc_hd__or2_2
X_2693_ _0543_ VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__clkbuf_4
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2127_ demux.state_machine.timeState\[1\] demux.state_machine.timeState\[5\] VGND
+ VGND VPWR VPWR _1400_ sky130_fd_sc_hd__or2_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_13_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2058_ demux.state_machine.currentAddress\[11\] _0988_ demux.state_machine.currentAddress\[4\]
+ _0948_ VGND VGND VPWR VPWR _1331_ sky130_fd_sc_hd__nor4_1
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3030_ clknet_4_6_0_clk _0002_ net67 VGND VGND VPWR VPWR demux.state_machine.currentAddress\[11\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_73_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2676_ _1071_ _0491_ _0526_ _1079_ _1411_ VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__a221o_1
XFILLER_0_41_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2745_ _0200_ _0221_ _0561_ VGND VGND VPWR VPWR _0592_ sky130_fd_sc_hd__and3_1
XFILLER_0_26_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2814_ _1326_ _0632_ VGND VGND VPWR VPWR _0654_ sky130_fd_sc_hd__or2_1
X_1558_ _0864_ VGND VGND VPWR VPWR _0865_ sky130_fd_sc_hd__clkbuf_8
X_1627_ _0932_ _0933_ VGND VGND VPWR VPWR _0934_ sky130_fd_sc_hd__and2_1
XTAP_184 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_373 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_70_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_254 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2530_ _0404_ _0259_ VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__xor2_1
X_2461_ _1002_ _1353_ _1239_ _1238_ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__a211o_1
X_2392_ _1425_ _0122_ _0279_ net46 internalDataflow.addressLowBusModule.busInputs\[33\]
+ VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__a32o_1
XFILLER_0_11_416 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3013_ _0385_ _0805_ _0801_ net95 VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_3_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_335 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2659_ internalDataflow.accRegToDB\[3\] _0194_ _0511_ VGND VGND VPWR VPWR _0515_
+ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_14_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2728_ internalDataflow.addressLowBusModule.busInputs\[18\] _0535_ VGND VGND VPWR
+ VPWR _0576_ sky130_fd_sc_hd__and2_1
XFILLER_0_69_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_379 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_1892_ _1088_ _1095_ _1174_ _0975_ VGND VGND VPWR VPWR _1175_ sky130_fd_sc_hd__a22o_1
X_1961_ net1 _0950_ VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__nand2_1
XFILLER_0_7_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_413 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2513_ _0394_ VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2444_ _0316_ _0318_ _0320_ _0321_ _0331_ VGND VGND VPWR VPWR internalDataflow.psr.processStatusReg.stat_buf_nxt\[6\]
+ sky130_fd_sc_hd__a41o_1
X_2375_ demux.PSR_Z _1317_ _1302_ internalDataflow.accRegToDB\[1\] _1316_ VGND VGND
+ VPWR VPWR _0263_ sky130_fd_sc_hd__a32o_1
XFILLER_0_11_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_368 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_59 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_68 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_29_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2160_ _1372_ _1380_ _1388_ _1432_ net47 VGND VGND VPWR VPWR _1433_ sky130_fd_sc_hd__a32o_1
XFILLER_0_45_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2091_ _1253_ VGND VGND VPWR VPWR _1364_ sky130_fd_sc_hd__inv_2
Xmax_cap1 _1312_ VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__buf_1
X_1875_ _0908_ _1066_ _1048_ _1113_ VGND VGND VPWR VPWR _1158_ sky130_fd_sc_hd__a22o_1
X_1944_ _1206_ _1216_ _1217_ _1223_ VGND VGND VPWR VPWR _1224_ sky130_fd_sc_hd__or4_1
XFILLER_0_61_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2993_ demux.nmi instructionLoader.interruptInjector.nmiGeneratedFF.nmiRunning instructionLoader.interruptInjector.nmiGeneratedFF.synchronizedNMI
+ VGND VGND VPWR VPWR _0794_ sky130_fd_sc_hd__or3b_1
XFILLER_0_43_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2427_ _0306_ _0314_ VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__or2_2
Xclkbuf_4_15_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_15_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_43_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2358_ _1114_ _1423_ _1418_ VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__nand3_1
X_2289_ _0123_ _0176_ VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__and2_2
XFILLER_0_19_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_124 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1660_ net2 net3 _0956_ VGND VGND VPWR VPWR _0964_ sky130_fd_sc_hd__o21ai_4
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1591_ branch_ff.branchForward branch_ff.branchBackward VGND VGND VPWR VPWR _0898_
+ sky130_fd_sc_hd__nor2_1
XFILLER_0_21_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2143_ _1415_ VGND VGND VPWR VPWR _1416_ sky130_fd_sc_hd__inv_2
X_2212_ _0876_ _0888_ net53 _0936_ _1263_ VGND VGND VPWR VPWR _1485_ sky130_fd_sc_hd__a311o_1
XFILLER_0_72_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2074_ _1263_ demux.state_machine.currentAddress\[11\] demux.state_machine.currentAddress\[1\]
+ demux.state_machine.currentAddress\[7\] VGND VGND VPWR VPWR _1347_ sky130_fd_sc_hd__or4_1
XFILLER_0_8_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1858_ _0927_ _1066_ _1054_ _1081_ VGND VGND VPWR VPWR _1142_ sky130_fd_sc_hd__a22o_1
X_1927_ _0901_ _0882_ _0979_ VGND VGND VPWR VPWR _1208_ sky130_fd_sc_hd__nor3_1
XFILLER_0_44_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2976_ net33 _0276_ _0783_ VGND VGND VPWR VPWR _0785_ sky130_fd_sc_hd__mux2_1
XFILLER_0_16_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1789_ _1070_ _1072_ VGND VGND VPWR VPWR _1073_ sky130_fd_sc_hd__or2_1
XFILLER_0_39_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_403 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2830_ _0666_ VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__clkbuf_1
X_1712_ demux.state_machine.timeState\[1\] _0981_ _1000_ _0879_ VGND VGND VPWR VPWR
+ _0014_ sky130_fd_sc_hd__a22o_1
X_1643_ _0942_ _0946_ _0822_ _0949_ VGND VGND VPWR VPWR _0950_ sky130_fd_sc_hd__a31oi_4
X_2692_ _0542_ VGND VGND VPWR VPWR _0543_ sky130_fd_sc_hd__inv_2
X_2761_ _0153_ _0606_ VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__xor2_1
XFILLER_0_5_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_305 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_1 _0652_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1574_ demux.state_machine.currentInstruction\[1\] _0813_ demux.state_machine.currentInstruction\[2\]
+ demux.state_machine.currentInstruction\[3\] VGND VGND VPWR VPWR _0881_ sky130_fd_sc_hd__or4b_1
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2126_ _0936_ _1121_ _0868_ _1243_ VGND VGND VPWR VPWR _1399_ sky130_fd_sc_hd__a22o_1
X_2057_ _0891_ _1084_ _1285_ VGND VGND VPWR VPWR _1330_ sky130_fd_sc_hd__and3_2
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2959_ _0558_ _0665_ VGND VGND VPWR VPWR _0770_ sky130_fd_sc_hd__nor2_1
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2813_ _0653_ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__clkbuf_1
X_1626_ _0827_ _0852_ VGND VGND VPWR VPWR _0933_ sky130_fd_sc_hd__nor2_2
X_2675_ demux.state_machine.timeState\[5\] demux.state_machine.timeState\[3\] VGND
+ VGND VPWR VPWR _0526_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2744_ _0587_ _0589_ _0538_ _0544_ VGND VGND VPWR VPWR _0591_ sky130_fd_sc_hd__a211o_1
X_1557_ _0813_ _0810_ _0811_ _0812_ VGND VGND VPWR VPWR _0864_ sky130_fd_sc_hd__or4bb_1
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2109_ branch_ff.branchBackward _1290_ _1381_ VGND VGND VPWR VPWR _1382_ sky130_fd_sc_hd__a21oi_2
X_3089_ clknet_4_3_0_clk _0081_ net59 VGND VGND VPWR VPWR internalDataflow.stackBusModule.busInputs\[46\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2460_ _0983_ _1150_ _1237_ _1002_ _0918_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__a221o_1
XFILLER_0_23_266 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2391_ demux.nmi demux.reset VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__or2b_1
XFILLER_0_64_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3012_ _0968_ internalDataflow.addressLowBusModule.busInputs\[23\] _0801_ VGND VGND
+ VPWR VPWR _0805_ sky130_fd_sc_hd__or3_1
XFILLER_0_3_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1609_ _0820_ _0825_ _0896_ _0819_ VGND VGND VPWR VPWR _0916_ sky130_fd_sc_hd__and4bb_1
X_2589_ _0136_ _0291_ _0406_ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__o21ai_1
X_2658_ _0514_ VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2727_ _0200_ _0574_ VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__xor2_1
XFILLER_0_69_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1960_ net10 VGND VGND VPWR VPWR instructionLoader.interruptInjector.interruptRequest
+ sky130_fd_sc_hd__inv_2
X_1891_ _1076_ _0865_ VGND VGND VPWR VPWR _1174_ sky130_fd_sc_hd__nor2_1
XFILLER_0_59_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2443_ _0322_ net89 _0999_ _0330_ VGND VGND VPWR VPWR _0331_ sky130_fd_sc_hd__a31o_1
XFILLER_0_3_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2512_ net104 _0274_ _0392_ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2374_ _0251_ _0259_ _0261_ VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__a21o_2
XFILLER_0_61_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2090_ _0924_ _1242_ _1362_ VGND VGND VPWR VPWR _1363_ sky130_fd_sc_hd__or3_1
XFILLER_0_45_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_280 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2992_ net90 _0792_ _0793_ VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_28_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1943_ _1218_ _1219_ _1222_ VGND VGND VPWR VPWR _1223_ sky130_fd_sc_hd__or3_1
X_1874_ _1156_ _0974_ _1063_ _1088_ VGND VGND VPWR VPWR _1157_ sky130_fd_sc_hd__a22o_1
XFILLER_0_61_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2426_ _1465_ _0309_ _0313_ VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__a21o_1
XFILLER_0_10_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2357_ _1325_ _1428_ _1425_ VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__o21bai_1
X_2288_ _0122_ _0174_ _0175_ VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__or3_2
XFILLER_0_62_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_136 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_1590_ _0896_ VGND VGND VPWR VPWR _0897_ sky130_fd_sc_hd__buf_4
XFILLER_0_0_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2073_ _1003_ _1343_ _1345_ _1241_ VGND VGND VPWR VPWR _1346_ sky130_fd_sc_hd__a22o_2
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2142_ _1263_ _1414_ _1241_ VGND VGND VPWR VPWR _1415_ sky130_fd_sc_hd__o21a_1
X_2211_ _1384_ _1419_ _1420_ _0960_ VGND VGND VPWR VPWR _1484_ sky130_fd_sc_hd__a31oi_2
XFILLER_0_72_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2975_ _0784_ VGND VGND VPWR VPWR _0099_ sky130_fd_sc_hd__clkbuf_1
X_1857_ _0845_ _1067_ _1048_ _1055_ VGND VGND VPWR VPWR _1141_ sky130_fd_sc_hd__a22o_1
XFILLER_0_71_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1926_ _1172_ _1197_ _1201_ _1206_ VGND VGND VPWR VPWR _1207_ sky130_fd_sc_hd__or4_1
X_1788_ _0966_ _0972_ _1017_ _1067_ _1071_ VGND VGND VPWR VPWR _1072_ sky130_fd_sc_hd__a32o_1
XFILLER_0_21_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2409_ internalDataflow.addressHighBusModule.busInputs\[23\] VGND VGND VPWR VPWR
+ _0297_ sky130_fd_sc_hd__inv_2
XFILLER_0_62_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold60 internalDataflow.addressHighBusModule.busInputs\[20\] VGND VGND VPWR VPWR
+ net132 sky130_fd_sc_hd__dlygate4sd3_1
Xclkbuf_4_14_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_14_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_53_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1642_ _0932_ _0822_ _0948_ VGND VGND VPWR VPWR _0949_ sky130_fd_sc_hd__o21ai_2
X_2691_ _0982_ _0540_ _0541_ _1290_ _0999_ VGND VGND VPWR VPWR _0542_ sky130_fd_sc_hd__o221ai_4
X_1711_ _0983_ _0981_ _1000_ _1002_ VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__a22o_1
XANTENNA_2 _0961_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2760_ _0593_ _0605_ VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__nand2_1
XFILLER_0_5_317 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1573_ _0869_ _0865_ VGND VGND VPWR VPWR _0880_ sky130_fd_sc_hd__or2_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2125_ _0875_ _0848_ _1395_ _1396_ _1397_ VGND VGND VPWR VPWR _1398_ sky130_fd_sc_hd__a2111o_1
X_2056_ _1328_ VGND VGND VPWR VPWR _1329_ sky130_fd_sc_hd__clkbuf_4
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1909_ _1190_ _1091_ _1055_ _1088_ VGND VGND VPWR VPWR _1191_ sky130_fd_sc_hd__a22o_1
XFILLER_0_44_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2958_ _0557_ _0665_ VGND VGND VPWR VPWR _0769_ sky130_fd_sc_hd__and2_1
XFILLER_0_17_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2889_ _0312_ _0636_ VGND VGND VPWR VPWR _0706_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_35_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2812_ net108 _0652_ _0645_ VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__mux2_1
X_2743_ _0587_ _0589_ VGND VGND VPWR VPWR _0590_ sky130_fd_sc_hd__nor2_1
X_2674_ _1394_ _1398_ VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__or2_1
X_1625_ demux.state_machine.timeState\[0\] VGND VGND VPWR VPWR _0932_ sky130_fd_sc_hd__clkbuf_4
X_1556_ _0850_ _0853_ _0856_ _0862_ VGND VGND VPWR VPWR _0863_ sky130_fd_sc_hd__or4b_1
XFILLER_0_5_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2108_ _1102_ _0944_ _1004_ VGND VGND VPWR VPWR _1381_ sky130_fd_sc_hd__o21a_1
X_2039_ _1302_ _1294_ _1304_ _1311_ VGND VGND VPWR VPWR _1312_ sky130_fd_sc_hd__nor4_1
X_3088_ clknet_4_9_0_clk _0080_ net63 VGND VGND VPWR VPWR internalDataflow.stackBusModule.busInputs\[45\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_17_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_55_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3011_ _0804_ VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__clkbuf_1
X_2390_ internalDataflow.addressLowBusModule.busInputs\[25\] _0125_ _0127_ net3 VGND
+ VGND VPWR VPWR _0278_ sky130_fd_sc_hd__a22o_1
XFILLER_0_3_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_156 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2726_ _0221_ _0537_ _0561_ _0573_ VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__a31o_1
XFILLER_0_6_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1539_ _0826_ _0816_ VGND VGND VPWR VPWR _0846_ sky130_fd_sc_hd__nor2_1
X_1608_ _0882_ _0861_ _0866_ VGND VGND VPWR VPWR _0915_ sky130_fd_sc_hd__a21oi_2
X_2657_ internalDataflow.accRegToDB\[2\] _0215_ _0511_ VGND VGND VPWR VPWR _0514_
+ sky130_fd_sc_hd__mux2_1
X_2588_ _0450_ _0451_ _0457_ VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_69_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_215 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1890_ _1076_ _0818_ VGND VGND VPWR VPWR _1173_ sky130_fd_sc_hd__nor2_1
XFILLER_0_55_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2442_ _1482_ _0326_ _0329_ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__mux2_1
X_2373_ _0154_ _0237_ _0260_ _0250_ VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__o211a_1
X_2511_ _0393_ VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__inv_2
XFILLER_0_38_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_70 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_19_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2709_ _0522_ _0557_ VGND VGND VPWR VPWR _0559_ sky130_fd_sc_hd__and2_1
XFILLER_0_6_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1942_ _1107_ _1139_ _1220_ _1221_ VGND VGND VPWR VPWR _1222_ sky130_fd_sc_hd__or4_1
XFILLER_0_56_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2991_ instructionLoader.interruptInjector.processStatusRegIFlag demux.setInterruptFlag
+ instructionLoader.interruptInjector.irqGenerated instructionLoader.interruptInjector.irqGeneratedFF.synchronizedIRQ
+ VGND VGND VPWR VPWR _0793_ sky130_fd_sc_hd__or4b_1
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1873_ _0866_ _0860_ VGND VGND VPWR VPWR _1156_ sky130_fd_sc_hd__nor2_1
XFILLER_0_24_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_234 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2425_ _1465_ _0312_ VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__nor2_1
X_2356_ _0228_ _0230_ _1372_ _1388_ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__o211a_1
X_2287_ internalDataflow.addressLowBusModule.busInputs\[20\] _1502_ _0127_ net6 VGND
+ VGND VPWR VPWR _0175_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_57_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_310 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2210_ _1468_ _1480_ _1482_ VGND VGND VPWR VPWR _1483_ sky130_fd_sc_hd__mux2_1
XFILLER_0_0_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2072_ _1273_ _1344_ VGND VGND VPWR VPWR _1345_ sky130_fd_sc_hd__nand2_1
X_2141_ _0875_ _1413_ demux.state_machine.currentAddress\[6\] VGND VGND VPWR VPWR
+ _1414_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1925_ _1203_ _1205_ VGND VGND VPWR VPWR _1206_ sky130_fd_sc_hd__or2_1
X_2974_ net126 _0236_ _0783_ VGND VGND VPWR VPWR _0784_ sky130_fd_sc_hd__mux2_1
X_1856_ _1132_ _1139_ VGND VGND VPWR VPWR _1140_ sky130_fd_sc_hd__or2_1
X_1787_ _0830_ _0909_ VGND VGND VPWR VPWR _1071_ sky130_fd_sc_hd__nor2_4
XFILLER_0_24_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2408_ _1372_ _0295_ VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__nand2_2
X_2339_ _0226_ _1366_ _1368_ _1369_ VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__or4_1
XFILLER_0_39_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_47_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_49 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold50 net27 VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__dlygate4sd3_1
Xhold61 internalDataflow.addressLowBusModule.busInputs\[21\] VGND VGND VPWR VPWR net133
+ sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_53_232 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_3 _0968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_1641_ demux.isAddressing net56 VGND VGND VPWR VPWR _0948_ sky130_fd_sc_hd__nand2_4
X_1710_ net84 _0981_ _1000_ demux.state_machine.timeState\[5\] VGND VGND VPWR VPWR
+ _0016_ sky130_fd_sc_hd__a22o_1
X_2690_ _0934_ _1385_ _1412_ VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__or3_1
X_1572_ demux.state_machine.timeState\[6\] VGND VGND VPWR VPWR _0879_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_41_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2124_ _1259_ _0945_ _1150_ _0936_ VGND VGND VPWR VPWR _1397_ sky130_fd_sc_hd__a22o_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2055_ _1256_ _1327_ VGND VGND VPWR VPWR _1328_ sky130_fd_sc_hd__nor2_1
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_1839_ _1122_ _1085_ _0974_ _1081_ _1088_ VGND VGND VPWR VPWR _1123_ sky130_fd_sc_hd__a32o_1
X_1908_ _1076_ _0825_ VGND VGND VPWR VPWR _1190_ sky130_fd_sc_hd__nor2_1
X_2888_ _0546_ _0699_ _0700_ _0705_ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__a31o_1
X_2957_ net119 _0555_ _0764_ _0546_ _0768_ VGND VGND VPWR VPWR _0097_ sky130_fd_sc_hd__a221o_1
XFILLER_0_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput40 net40 VGND VGND VPWR VPWR dataBusSelect sky130_fd_sc_hd__clkbuf_4
XFILLER_0_53_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2811_ _0213_ _0632_ _0633_ _0212_ _0651_ VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__a221o_2
X_2742_ _0568_ _0569_ _0588_ _0579_ _0576_ VGND VGND VPWR VPWR _0589_ sky130_fd_sc_hd__a311o_1
X_1624_ _0929_ _0930_ _0879_ VGND VGND VPWR VPWR _0931_ sky130_fd_sc_hd__o21a_1
X_1555_ _0857_ _0858_ _0860_ _0861_ _0821_ VGND VGND VPWR VPWR _0862_ sky130_fd_sc_hd__a41o_1
X_2673_ _1005_ _0936_ _0523_ _0905_ VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__o31a_1
XFILLER_0_27_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3087_ clknet_4_2_0_clk _0079_ net59 VGND VGND VPWR VPWR internalDataflow.stackBusModule.busInputs\[44\]
+ sky130_fd_sc_hd__dfrtp_1
X_2107_ internalDataflow.stackBusModule.busInputs\[38\] _1371_ _1376_ _1379_ VGND
+ VGND VPWR VPWR _1380_ sky130_fd_sc_hd__a211o_1
X_2038_ _1305_ _1308_ _1309_ _1310_ VGND VGND VPWR VPWR _1311_ sky130_fd_sc_hd__a31o_1
XFILLER_0_11_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_4_13_0_clk clknet_0_clk VGND VGND VPWR VPWR clknet_4_13_0_clk sky130_fd_sc_hd__clkbuf_8
XFILLER_0_23_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3010_ _0979_ _0803_ demux.isAddressing VGND VGND VPWR VPWR _0804_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_371 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2725_ _0221_ _0559_ _0562_ VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__and3b_1
X_2656_ _0513_ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_59_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1538_ _0826_ _0844_ VGND VGND VPWR VPWR _0845_ sky130_fd_sc_hd__nor2_1
X_1607_ _0912_ _0913_ demux.state_machine.timeState\[5\] VGND VGND VPWR VPWR _0914_
+ sky130_fd_sc_hd__o21a_1
X_2587_ net112 net45 _0456_ _0321_ VGND VGND VPWR VPWR _0457_ sky130_fd_sc_hd__a22oi_1
X_3139_ clknet_4_15_0_clk _0021_ net71 VGND VGND VPWR VPWR demux.state_machine.currentInstruction\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_49_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2510_ _0389_ _0249_ _0392_ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2441_ _1325_ _0328_ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__or2_1
X_2372_ _1465_ _0241_ VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__or2_1
XFILLER_0_24_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_393 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2708_ _0557_ VGND VGND VPWR VPWR _0558_ sky130_fd_sc_hd__clkbuf_4
X_2639_ net75 _0503_ _0221_ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__a21o_1
XFILLER_0_37_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_171 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1872_ _0839_ _0975_ _1018_ _1055_ VGND VGND VPWR VPWR _1155_ sky130_fd_sc_hd__a22o_1
X_1941_ _0846_ _1091_ _1104_ _1153_ VGND VGND VPWR VPWR _1221_ sky130_fd_sc_hd__a211o_1
X_2990_ _0981_ _0340_ VGND VGND VPWR VPWR _0792_ sky130_fd_sc_hd__or2_1
XFILLER_0_9_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2424_ _0310_ _0311_ _0123_ VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__o21a_2
X_2355_ _1460_ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__inv_2
X_2286_ internalDataflow.addressLowBusModule.busInputs\[36\] net46 _0125_ internalDataflow.addressLowBusModule.busInputs\[28\]
+ VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_293 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2140_ _0896_ demux.state_machine.timeState\[6\] VGND VGND VPWR VPWR _1413_ sky130_fd_sc_hd__and2b_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2071_ _0987_ _1077_ _0876_ VGND VGND VPWR VPWR _1344_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_29_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_1855_ _0966_ _1116_ _1137_ _1066_ _1138_ VGND VGND VPWR VPWR _1139_ sky130_fd_sc_hd__a32o_1
X_1924_ _1060_ _1151_ _1204_ _1091_ _1089_ VGND VGND VPWR VPWR _1205_ sky130_fd_sc_hd__a221o_1
X_2973_ _0782_ VGND VGND VPWR VPWR _0783_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_16_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_1786_ _0910_ _1067_ _1063_ _1069_ VGND VGND VPWR VPWR _1070_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2269_ _0147_ _0155_ VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__or2_1
X_2407_ internalDataflow.stackBusModule.busInputs\[39\] _1371_ _0293_ _0294_ VGND
+ VGND VPWR VPWR _0295_ sky130_fd_sc_hd__a211o_1
X_2338_ internalDataflow.accRegToDB\[0\] VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold40 internalDataflow.addressLowBusModule.busInputs\[29\] VGND VGND VPWR VPWR net112
+ sky130_fd_sc_hd__dlygate4sd3_1
Xhold51 net30 VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1640_ demux.state_machine.currentAddress\[8\] demux.state_machine.currentAddress\[0\]
+ demux.state_machine.currentAddress\[2\] demux.state_machine.currentAddress\[9\]
+ VGND VGND VPWR VPWR _0947_ sky130_fd_sc_hd__nor4_2
XFILLER_0_67_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_1571_ _0849_ _0863_ _0867_ _0874_ _0877_ VGND VGND VPWR VPWR _0878_ sky130_fd_sc_hd__o41a_1
XFILLER_0_41_417 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2123_ _0870_ _1131_ _1243_ VGND VGND VPWR VPWR _1396_ sky130_fd_sc_hd__o21a_1
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_2054_ _1323_ _1280_ _1324_ _1325_ VGND VGND VPWR VPWR _1327_ sky130_fd_sc_hd__a31o_1
XFILLER_0_8_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_16_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_1838_ _0832_ _0834_ _0835_ _0833_ VGND VGND VPWR VPWR _1122_ sky130_fd_sc_hd__and4bb_1
X_1907_ _0871_ _0825_ VGND VGND VPWR VPWR _1189_ sky130_fd_sc_hd__nor2_1
XFILLER_0_32_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2887_ _0544_ _0703_ _0704_ _0555_ internalDataflow.addressHighBusModule.busInputs\[16\]
+ VGND VGND VPWR VPWR _0705_ sky130_fd_sc_hd__a32o_1
XFILLER_0_29_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2956_ _0665_ _0766_ _0767_ VGND VGND VPWR VPWR _0768_ sky130_fd_sc_hd__a21oi_1
X_1769_ _1017_ _1040_ VGND VGND VPWR VPWR _1053_ sky130_fd_sc_hd__nor2_1
XFILLER_0_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput41 net41 VGND VGND VPWR VPWR functionalClockOut sky130_fd_sc_hd__buf_1
Xoutput30 net30 VGND VGND VPWR VPWR addressBusLow[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_336 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2672_ _1469_ _0898_ _0877_ VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__o21a_1
XFILLER_0_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_2810_ _0207_ _0634_ VGND VGND VPWR VPWR _0651_ sky130_fd_sc_hd__and2_1
X_2741_ internalDataflow.addressLowBusModule.busInputs\[19\] _0534_ VGND VGND VPWR
+ VPWR _0588_ sky130_fd_sc_hd__or2_1
X_1623_ _0860_ _0861_ _0830_ VGND VGND VPWR VPWR _0930_ sky130_fd_sc_hd__a21oi_4
X_1554_ _0835_ _0834_ _0833_ _0832_ VGND VGND VPWR VPWR _0861_ sky130_fd_sc_hd__nand4b_4
XTAP_155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

