* NGSPICE file created from z23.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_2 abstract view
.subckt sky130_fd_sc_hd__or3b_2 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_1 abstract view
.subckt sky130_fd_sc_hd__o2111a_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_2 abstract view
.subckt sky130_fd_sc_hd__dfstp_2 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_1 abstract view
.subckt sky130_fd_sc_hd__dfrtp_1 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_8 abstract view
.subckt sky130_fd_sc_hd__nor2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_2 abstract view
.subckt sky130_fd_sc_hd__dfrtp_2 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlygate4sd3_1 abstract view
.subckt sky130_fd_sc_hd__dlygate4sd3_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_1 abstract view
.subckt sky130_fd_sc_hd__or4b_1 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_1 abstract view
.subckt sky130_fd_sc_hd__and4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221a_1 abstract view
.subckt sky130_fd_sc_hd__o221a_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_4 abstract view
.subckt sky130_fd_sc_hd__o21a_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_4 abstract view
.subckt sky130_fd_sc_hd__o22a_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4_2 abstract view
.subckt sky130_fd_sc_hd__and4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_4 abstract view
.subckt sky130_fd_sc_hd__o41a_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_4 abstract view
.subckt sky130_fd_sc_hd__a21bo_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_4 abstract view
.subckt sky130_fd_sc_hd__or4b_4 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_4 abstract view
.subckt sky130_fd_sc_hd__or3b_4 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_4 abstract view
.subckt sky130_fd_sc_hd__o2111a_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_2 abstract view
.subckt sky130_fd_sc_hd__and4bb_2 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_4 abstract view
.subckt sky130_fd_sc_hd__a22oi_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_2 abstract view
.subckt sky130_fd_sc_hd__nand2b_2 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_4 abstract view
.subckt sky130_fd_sc_hd__nor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_1 abstract view
.subckt sky130_fd_sc_hd__and4b_1 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_1 abstract view
.subckt sky130_fd_sc_hd__o311a_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_4 abstract view
.subckt sky130_fd_sc_hd__or4bb_4 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_8 abstract view
.subckt sky130_fd_sc_hd__nand2_8 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_1 abstract view
.subckt sky130_fd_sc_hd__a2111oi_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_4 abstract view
.subckt sky130_fd_sc_hd__and3b_4 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o41a_2 abstract view
.subckt sky130_fd_sc_hd__o41a_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_1 abstract view
.subckt sky130_fd_sc_hd__dfstp_1 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_2 abstract view
.subckt sky130_fd_sc_hd__nor4_2 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4_1 abstract view
.subckt sky130_fd_sc_hd__nor4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2b_2 abstract view
.subckt sky130_fd_sc_hd__nor2b_2 A B_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_4 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_4 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_4 abstract view
.subckt sky130_fd_sc_hd__o211a_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_2 abstract view
.subckt sky130_fd_sc_hd__nor3b_2 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_4 abstract view
.subckt sky130_fd_sc_hd__nor3b_4 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_2 abstract view
.subckt sky130_fd_sc_hd__nor4b_2 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_2 abstract view
.subckt sky130_fd_sc_hd__a311o_2 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_4 abstract view
.subckt sky130_fd_sc_hd__a22o_4 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_2 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_4 abstract view
.subckt sky130_fd_sc_hd__o31a_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_4 abstract view
.subckt sky130_fd_sc_hd__or2b_4 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4bb_1 abstract view
.subckt sky130_fd_sc_hd__or4bb_1 A B C_N D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_4 abstract view
.subckt sky130_fd_sc_hd__nor3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32a_1 abstract view
.subckt sky130_fd_sc_hd__o32a_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_1 abstract view
.subckt sky130_fd_sc_hd__o31ai_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_4 abstract view
.subckt sky130_fd_sc_hd__nand3b_4 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_4 abstract view
.subckt sky130_fd_sc_hd__a41o_4 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4b_2 abstract view
.subckt sky130_fd_sc_hd__and4b_2 A_N B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_4 abstract view
.subckt sky130_fd_sc_hd__a2111o_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2b_4 abstract view
.subckt sky130_fd_sc_hd__nand2b_4 A_N B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_4 abstract view
.subckt sky130_fd_sc_hd__a2111oi_4 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux4_1 abstract view
.subckt sky130_fd_sc_hd__mux4_1 A0 A1 A2 A3 S0 S1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_2 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_2 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_1 abstract view
.subckt sky130_fd_sc_hd__o22ai_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o311a_4 abstract view
.subckt sky130_fd_sc_hd__o311a_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfxtp_1 abstract view
.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_2 abstract view
.subckt sky130_fd_sc_hd__a21bo_2 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31oi_1 abstract view
.subckt sky130_fd_sc_hd__a31oi_1 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_4 abstract view
.subckt sky130_fd_sc_hd__a21o_4 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_4 abstract view
.subckt sky130_fd_sc_hd__o21bai_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_2 abstract view
.subckt sky130_fd_sc_hd__and3b_2 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_2 abstract view
.subckt sky130_fd_sc_hd__a32o_2 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_2 abstract view
.subckt sky130_fd_sc_hd__or4_2 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_4 abstract view
.subckt sky130_fd_sc_hd__a31o_4 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111oi_2 abstract view
.subckt sky130_fd_sc_hd__a2111oi_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_4 abstract view
.subckt sky130_fd_sc_hd__and4bb_4 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111a_2 abstract view
.subckt sky130_fd_sc_hd__o2111a_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_1 abstract view
.subckt sky130_fd_sc_hd__o221ai_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_1 abstract view
.subckt sky130_fd_sc_hd__a41o_1 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3b_1 abstract view
.subckt sky130_fd_sc_hd__nor3b_1 A B C_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2111ai_2 abstract view
.subckt sky130_fd_sc_hd__o2111ai_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_2 abstract view
.subckt sky130_fd_sc_hd__o31a_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor4b_1 abstract view
.subckt sky130_fd_sc_hd__nor4b_1 A B C D_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a41o_2 abstract view
.subckt sky130_fd_sc_hd__a41o_2 A1 A2 A3 A4 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

.subckt z23 VGND VPWR clk interrupt_gpio_in keypad_input[0] keypad_input[10] keypad_input[11]
+ keypad_input[12] keypad_input[13] keypad_input[14] keypad_input[15] keypad_input[1]
+ keypad_input[2] keypad_input[3] keypad_input[4] keypad_input[5] keypad_input[6]
+ keypad_input[7] keypad_input[8] keypad_input[9] memory_address_out[0] memory_address_out[10]
+ memory_address_out[11] memory_address_out[12] memory_address_out[13] memory_address_out[14]
+ memory_address_out[15] memory_address_out[1] memory_address_out[2] memory_address_out[3]
+ memory_address_out[4] memory_address_out[5] memory_address_out[6] memory_address_out[7]
+ memory_address_out[8] memory_address_out[9] memory_data_in[0] memory_data_in[1]
+ memory_data_in[2] memory_data_in[3] memory_data_in[4] memory_data_in[5] memory_data_in[6]
+ memory_data_in[7] memory_data_out[0] memory_data_out[1] memory_data_out[2] memory_data_out[3]
+ memory_data_out[4] memory_data_out[5] memory_data_out[6] memory_data_out[7] memory_wr
+ nrst programmable_gpio_in[0] programmable_gpio_in[1] programmable_gpio_in[2] programmable_gpio_in[3]
+ programmable_gpio_in[4] programmable_gpio_in[5] programmable_gpio_in[6] programmable_gpio_in[7]
+ programmable_gpio_out[0] programmable_gpio_out[1] programmable_gpio_out[2] programmable_gpio_out[3]
+ programmable_gpio_out[4] programmable_gpio_out[5] programmable_gpio_out[6] programmable_gpio_out[7]
+ programmable_gpio_wr[0] programmable_gpio_wr[1] programmable_gpio_wr[2] programmable_gpio_wr[3]
+ programmable_gpio_wr[4] programmable_gpio_wr[5] programmable_gpio_wr[6] programmable_gpio_wr[7]
+ ss0[0] ss0[1] ss0[2] ss0[3] ss0[4] ss0[5] ss0[6] ss0[7] ss1[0] ss1[1] ss1[2] ss1[3]
+ ss1[4] ss1[5] ss1[6] ss1[7] ss2[0] ss2[1] ss2[2] ss2[3] ss2[4] ss2[5] ss2[6] ss2[7]
+ ss3[0] ss3[1] ss3[2] ss3[3] ss3[4] ss3[5] ss3[6] ss3[7] ss4[0] ss4[1] ss4[2] ss4[3]
+ ss4[4] ss4[5] ss4[6] ss4[7] ss5[0] ss5[1] ss5[2] ss5[3] ss5[4] ss5[5] ss5[6] ss5[7]
+ ss6[0] ss6[1] ss6[2] ss6[3] ss6[4] ss6[5] ss6[6] ss6[7] ss7[0] ss7[1] ss7[2] ss7[3]
+ ss7[4] ss7[5] ss7[6] ss7[7]
XTAP_199 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5417__A0 _1194_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3155_ cu.id.alu_opcode\[0\] VGND VGND VPWR VPWR _2892_ sky130_fd_sc_hd__clkbuf_4
X_3086_ _2752_ _2822_ ih.t.count\[9\] VGND VGND VPWR VPWR _2824_ sky130_fd_sc_hd__a21oi_1
XANTENNA__5968__A1 _2486_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout162_A net163 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3988_ _0588_ _1059_ _0606_ _1061_ VGND VGND VPWR VPWR _1062_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_91_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5727_ _2518_ mc.cl.next_data\[2\] _2111_ VGND VGND VPWR VPWR _2524_ sky130_fd_sc_hd__and3_1
XANTENNA__5485__B _2284_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_9_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5658_ net91 _1329_ VGND VGND VPWR VPWR _2471_ sky130_fd_sc_hd__or2_1
X_4609_ _1652_ mc.cc.count\[3\] mc.cc.enable_edge_detector.prev_data VGND VGND VPWR
+ VPWR _1653_ sky130_fd_sc_hd__or3b_2
X_5589_ _2169_ _2398_ _2405_ _2136_ VGND VGND VPWR VPWR _2406_ sky130_fd_sc_hd__o211a_1
XFILLER_0_4_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4829__B cu.pc.pc_o\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3643__B _0663_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5350__S _2215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output56_A net56 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4960_ _1799_ _1942_ _1948_ _1949_ VGND VGND VPWR VPWR _1950_ sky130_fd_sc_hd__a22o_1
XFILLER_0_80_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4891_ _2920_ cu.pc.pc_o\[7\] VGND VGND VPWR VPWR _1886_ sky130_fd_sc_hd__nand2_1
XFILLER_0_58_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3911_ _0973_ _0329_ _0379_ VGND VGND VPWR VPWR _0987_ sky130_fd_sc_hd__nor3_1
XFILLER_0_80_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3842_ _0917_ VGND VGND VPWR VPWR _0918_ sky130_fd_sc_hd__buf_2
XFILLER_0_39_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5512_ net67 _1638_ _2279_ net66 VGND VGND VPWR VPWR _2332_ sky130_fd_sc_hd__a22o_1
XANTENNA__3820__B_N _0895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3594__D1 _0576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3773_ cu.reg_file.reg_a\[5\] _0625_ _0628_ cu.reg_file.reg_mem\[13\] _0848_ VGND
+ VGND VPWR VPWR _0849_ sky130_fd_sc_hd__a221o_1
XFILLER_0_14_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5886__A0 _1189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5443_ _2139_ _2247_ VGND VGND VPWR VPWR _2272_ sky130_fd_sc_hd__nand2_1
X_5374_ _2230_ VGND VGND VPWR VPWR _0161_ sky130_fd_sc_hd__clkbuf_1
X_4325_ cu.reg_file.reg_sp\[3\] _0993_ _1344_ cu.id.cb_opcode_y\[0\] _1324_ VGND VGND
+ VPWR VPWR _1390_ sky130_fd_sc_hd__a221o_1
XFILLER_0_10_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4256_ _1323_ VGND VGND VPWR VPWR _1324_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_38_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5260__S _1666_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3207_ _2897_ _2932_ _2935_ _2937_ _2943_ VGND VGND VPWR VPWR _2944_ sky130_fd_sc_hd__o2111a_1
X_4187_ _1234_ _1182_ _1023_ VGND VGND VPWR VPWR _1257_ sky130_fd_sc_hd__o21a_1
X_3138_ cu.id.opcode\[6\] VGND VGND VPWR VPWR _2875_ sky130_fd_sc_hd__clkbuf_4
XTAP_1129 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1118 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1107 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3069_ _2756_ _2806_ ih.t.count\[15\] VGND VGND VPWR VPWR _2807_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_9_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_92_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_clkbuf_leaf_31_clk_A clknet_2_1__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_339 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5565__C1 _1661_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5580__A2 _2147_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3591__B2 cu.reg_file.reg_h\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3591__A1 cu.reg_file.reg_sp\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5345__S _2206_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3654__A _0566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5090_ cu.reg_file.reg_d\[4\] _2047_ _2039_ VGND VGND VPWR VPWR _2048_ sky130_fd_sc_hd__mux2_1
X_4110_ _1013_ _1182_ _1023_ VGND VGND VPWR VPWR _1184_ sky130_fd_sc_hd__o21ai_2
X_4041_ _0607_ _1114_ _0632_ VGND VGND VPWR VPWR _1115_ sky130_fd_sc_hd__o21a_1
XANTENNA__5080__S _2035_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3646__A2 _0663_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5992_ clknet_leaf_33_clk _0030_ net161 VGND VGND VPWR VPWR cu.pc.pc_o\[14\] sky130_fd_sc_hd__dfrtp_4
X_4943_ _1932_ _1933_ VGND VGND VPWR VPWR _1934_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_74_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4874_ cu.pc.pc_o\[5\] _1870_ _1815_ VGND VGND VPWR VPWR _1871_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3825_ _0737_ _0752_ _0898_ _0900_ VGND VGND VPWR VPWR _0901_ sky130_fd_sc_hd__a31o_1
XFILLER_0_34_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5020__A1 _1263_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3756_ cu.reg_file.reg_mem\[15\] _0640_ _0830_ _0831_ VGND VGND VPWR VPWR _0832_
+ sky130_fd_sc_hd__a211oi_4
XFILLER_0_42_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3582__B2 cu.reg_file.reg_a\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3582__A1 cu.reg_file.reg_b\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5426_ _2022_ net69 _2260_ VGND VGND VPWR VPWR _2261_ sky130_fd_sc_hd__mux2_1
X_3687_ _0762_ VGND VGND VPWR VPWR _0763_ sky130_fd_sc_hd__inv_2
XFILLER_0_2_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5357_ _2220_ VGND VGND VPWR VPWR _0154_ sky130_fd_sc_hd__clkbuf_1
X_5288_ _1369_ _2179_ VGND VGND VPWR VPWR _2180_ sky130_fd_sc_hd__and2_4
X_4308_ _1373_ VGND VGND VPWR VPWR _1374_ sky130_fd_sc_hd__clkbuf_4
X_4239_ _0343_ _1295_ _1298_ _1299_ _1306_ VGND VGND VPWR VPWR _1307_ sky130_fd_sc_hd__a221o_1
XANTENNA__4826__C cu.pc.pc_o\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_69_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4842__B cu.pc.pc_o\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3458__B _0501_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5011__A1 _1213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3573__B2 cu.reg_file.reg_e\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_68_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5002__A1 _1623_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4590_ _1415_ _1630_ _1633_ VGND VGND VPWR VPWR _1634_ sky130_fd_sc_hd__or3_2
XFILLER_0_9_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3610_ _0464_ _0487_ _0482_ cu.reg_file.reg_l\[3\] VGND VGND VPWR VPWR _0686_ sky130_fd_sc_hd__o211a_1
X_3541_ _0616_ VGND VGND VPWR VPWR _0617_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_386 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6260_ clknet_leaf_21_clk _0242_ net190 VGND VGND VPWR VPWR ih.t.timer_max\[8\] sky130_fd_sc_hd__dfstp_2
XANTENNA__5688__A2_N _1643_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3472_ _0371_ _0376_ VGND VGND VPWR VPWR _0548_ sky130_fd_sc_hd__or2_2
XFILLER_0_10_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6191_ clknet_leaf_23_clk _0224_ net192 VGND VGND VPWR VPWR mc.cl.next_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_5211_ _0619_ ih.gpio_interrupt_mask\[0\] _2127_ VGND VGND VPWR VPWR _2128_ sky130_fd_sc_hd__mux2_1
X_5142_ _2081_ cu.reg_file.reg_h\[6\] _2069_ VGND VGND VPWR VPWR _2082_ sky130_fd_sc_hd__mux2_1
XANTENNA__4927__B _1521_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5073_ _2034_ _1792_ VGND VGND VPWR VPWR _2035_ sky130_fd_sc_hd__nor2_8
X_4024_ _1032_ _1095_ _1097_ _0770_ VGND VGND VPWR VPWR _1098_ sky130_fd_sc_hd__o22a_1
XFILLER_0_47_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5975_ clknet_leaf_32_clk _0012_ net161 VGND VGND VPWR VPWR cu.alu_f\[5\] sky130_fd_sc_hd__dfrtp_1
X_4926_ _2920_ _1521_ VGND VGND VPWR VPWR _1918_ sky130_fd_sc_hd__or2_1
XFILLER_0_47_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4857_ _1853_ _1854_ VGND VGND VPWR VPWR _1855_ sky130_fd_sc_hd__xnor2_1
XANTENNA__3278__B _2936_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_15_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3808_ cu.reg_file.reg_b\[2\] _0426_ _0429_ cu.reg_file.reg_d\[2\] VGND VGND VPWR
+ VPWR _0884_ sky130_fd_sc_hd__a22o_1
XANTENNA__5493__B _1648_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4752__B1 _0350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4788_ _2953_ _0339_ VGND VGND VPWR VPWR _1790_ sky130_fd_sc_hd__nor2_2
XFILLER_0_70_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3739_ _0813_ _0814_ VGND VGND VPWR VPWR _0815_ sky130_fd_sc_hd__nand2_1
XFILLER_0_42_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5409_ _1075_ net134 _2248_ VGND VGND VPWR VPWR _2251_ sky130_fd_sc_hd__mux2_1
XANTENNA__4268__C1 _1335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4853__A _0374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3794__A1 cu.reg_file.reg_a\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3794__B2 cu.reg_file.reg_mem\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5535__A2 _2194_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xwire144 _0985_ VGND VGND VPWR VPWR net144 sky130_fd_sc_hd__buf_1
XANTENNA__3546__B2 cu.reg_file.reg_l\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5299__A1 net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_507 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4763__A _1739_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5578__B _1330_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3379__A _0298_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2972_ net10 VGND VGND VPWR VPWR _2711_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5760_ cu.reg_file.reg_sp\[3\] _2534_ VGND VGND VPWR VPWR _2549_ sky130_fd_sc_hd__and2_1
X_4711_ ih.t.count\[25\] ih.t.count\[26\] _1723_ VGND VGND VPWR VPWR _1726_ sky130_fd_sc_hd__and3_1
X_5691_ mc.cl.next_data\[11\] _2359_ _2490_ _2499_ VGND VGND VPWR VPWR _2500_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__3785__A1 cu.id.imm_i\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4642_ ih.t.count\[0\] ih.t.count\[1\] ih.t.count\[2\] ih.t.count\[3\] VGND VGND
+ VPWR VPWR _1680_ sky130_fd_sc_hd__a31o_1
XFILLER_0_71_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4573_ _2702_ _1052_ _1623_ _2697_ VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__a22o_1
XANTENNA__4734__B1 _2878_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6312_ clknet_leaf_36_clk _0005_ net158 VGND VGND VPWR VPWR cu.id.state\[1\] sky130_fd_sc_hd__dfrtp_1
X_3524_ _0599_ VGND VGND VPWR VPWR _0600_ sky130_fd_sc_hd__inv_2
X_6243_ clknet_leaf_23_clk ih.t.next_count\[31\] net192 VGND VGND VPWR VPWR ih.t.count\[31\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__4938__A cu.pc.pc_o\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3455_ _0530_ VGND VGND VPWR VPWR _0531_ sky130_fd_sc_hd__buf_2
X_6174_ clknet_leaf_19_clk _0208_ net185 VGND VGND VPWR VPWR cu.reg_file.reg_mem\[10\]
+ sky130_fd_sc_hd__dfrtp_2
X_3386_ _0455_ _0461_ VGND VGND VPWR VPWR _0462_ sky130_fd_sc_hd__nand2_1
X_5125_ _2070_ VGND VGND VPWR VPWR _0072_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5056_ cu.reg_file.reg_c\[0\] _2022_ _2025_ VGND VGND VPWR VPWR _2026_ sky130_fd_sc_hd__mux2_1
XANTENNA__5462__A1 _2085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4007_ _1076_ _1077_ _1080_ _0517_ VGND VGND VPWR VPWR _1081_ sky130_fd_sc_hd__o31a_1
XFILLER_0_67_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5958_ cu.id.imm_i\[10\] _2391_ _2686_ VGND VGND VPWR VPWR _2689_ sky130_fd_sc_hd__mux2_1
X_4909_ _1900_ _1901_ _1798_ VGND VGND VPWR VPWR _1903_ sky130_fd_sc_hd__a21oi_1
XANTENNA__3776__B2 cu.reg_file.reg_d\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3776__A1 cu.reg_file.reg_b\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4973__A0 cu.pc.pc_o\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5889_ _2651_ VGND VGND VPWR VPWR _0255_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4740__A3 _0968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold30 ih.t.count\[7\] VGND VGND VPWR VPWR net226 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_26_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4583__A _1561_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_38_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4716__B1 _1687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3519__B2 _0340_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_5 _1188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output86_A net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_315 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_304 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3662__A _2950_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5141__A0 _1624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4477__B _1530_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6108__RESET_B net195 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_326 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3240_ _0308_ _0315_ VGND VGND VPWR VPWR _0316_ sky130_fd_sc_hd__nor2_1
XANTENNA__5692__B2 _1646_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3171_ cu.id.opcode\[7\] cu.id.opcode\[6\] VGND VGND VPWR VPWR _2908_ sky130_fd_sc_hd__and2b_2
XTAP_359 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5444__A1 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3207__B1 _2935_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5812_ _1623_ _2594_ _2545_ VGND VGND VPWR VPWR _2595_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5743_ _2533_ VGND VGND VPWR VPWR _2534_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_29_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3758__A1 cu.reg_file.reg_d\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3758__B2 cu.reg_file.reg_h\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2955_ mc.rw.state\[2\] _2695_ mc.rw.state\[0\] VGND VGND VPWR VPWR _2696_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5674_ cu.reg_file.reg_mem\[7\] _2486_ _1739_ VGND VGND VPWR VPWR _2487_ sky130_fd_sc_hd__mux2_1
XANTENNA__4707__B1 _1687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4625_ _1666_ VGND VGND VPWR VPWR _1667_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_25_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4556_ _1296_ _1607_ _1608_ VGND VGND VPWR VPWR _1609_ sky130_fd_sc_hd__a21o_1
X_3507_ _0321_ _0322_ _0328_ _0334_ VGND VGND VPWR VPWR _0583_ sky130_fd_sc_hd__or4_4
XANTENNA__5263__S _1666_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4487_ cu.reg_file.reg_h\[3\] _1316_ _1312_ cu.reg_file.reg_b\[3\] _1543_ VGND VGND
+ VPWR VPWR _1544_ sky130_fd_sc_hd__a221o_1
XANTENNA__5132__A0 _1222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6226_ clknet_leaf_11_clk ih.t.next_count\[14\] net177 VGND VGND VPWR VPWR ih.t.count\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_3438_ _0384_ _0392_ VGND VGND VPWR VPWR _0514_ sky130_fd_sc_hd__nand2_1
X_6157_ clknet_leaf_17_clk _0191_ net172 VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__dfrtp_4
XTAP_871 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_860 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4486__A2 _1321_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3369_ cu.id.cb_opcode_y\[0\] _0361_ _0444_ _0343_ _0322_ VGND VGND VPWR VPWR _0445_
+ sky130_fd_sc_hd__a221o_1
XTAP_893 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_882 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5108_ _2059_ VGND VGND VPWR VPWR _0066_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5499__A _2180_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5435__A1 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6088_ clknet_leaf_19_clk _0122_ net190 VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__dfrtp_4
X_5039_ _2013_ VGND VGND VPWR VPWR _0043_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3945__C_N _0986_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3749__A1 cu.reg_file.reg_d\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3749__B2 cu.reg_file.reg_h\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5371__A0 _1075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput42 net42 VGND VGND VPWR VPWR memory_address_out[1] sky130_fd_sc_hd__clkbuf_4
XANTENNA__4578__A _0516_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput75 net75 VGND VGND VPWR VPWR programmable_gpio_wr[7] sky130_fd_sc_hd__clkbuf_4
Xoutput64 net64 VGND VGND VPWR VPWR programmable_gpio_out[4] sky130_fd_sc_hd__clkbuf_4
Xoutput53 net53 VGND VGND VPWR VPWR memory_data_out[2] sky130_fd_sc_hd__buf_2
Xoutput97 net97 VGND VGND VPWR VPWR ss2[5] sky130_fd_sc_hd__clkbuf_4
Xoutput86 net86 VGND VGND VPWR VPWR ss1[2] sky130_fd_sc_hd__clkbuf_4
XANTENNA__5674__A1 _2486_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5426__A1 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output124_A net124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5348__S _2215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5362__A0 _1261_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4165__A1 _0387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4410_ cu.pc.pc_o\[7\] _1322_ _1315_ cu.reg_file.reg_e\[7\] _1470_ VGND VGND VPWR
+ VPWR _1471_ sky130_fd_sc_hd__a221o_1
XFILLER_0_78_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5390_ _1075_ net126 _2237_ VGND VGND VPWR VPWR _2240_ sky130_fd_sc_hd__mux2_1
X_4341_ _1382_ _1398_ _1399_ _1405_ VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__a31o_2
XANTENNA__5083__S _2035_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3912__A1 _2936_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4272_ cu.reg_file.reg_c\[1\] _1281_ _1338_ VGND VGND VPWR VPWR _1339_ sky130_fd_sc_hd__a21oi_1
X_6011_ clknet_leaf_4_clk _0049_ net170 VGND VGND VPWR VPWR cu.reg_file.reg_c\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_3223_ _2902_ _2884_ VGND VGND VPWR VPWR _0299_ sky130_fd_sc_hd__and2_1
XANTENNA__5417__A1 net138 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3154_ _2888_ _2889_ _2890_ VGND VGND VPWR VPWR _2891_ sky130_fd_sc_hd__and3_1
X_3085_ ih.t.count\[9\] _2752_ _2822_ VGND VGND VPWR VPWR _2823_ sky130_fd_sc_hd__and3_1
XFILLER_0_89_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout155_A net163 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3987_ _1060_ _0588_ _0599_ VGND VGND VPWR VPWR _1061_ sky130_fd_sc_hd__and3_1
XFILLER_0_91_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5726_ net19 _2519_ _2523_ VGND VGND VPWR VPWR _0220_ sky130_fd_sc_hd__a21o_1
XFILLER_0_45_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3600__B1 _0498_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5657_ net99 _2193_ _2469_ VGND VGND VPWR VPWR _2470_ sky130_fd_sc_hd__a21o_1
XFILLER_0_60_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4608_ mc.cc.count\[2\] mc.cc.count\[1\] mc.cc.count\[0\] VGND VGND VPWR VPWR _1652_
+ sky130_fd_sc_hd__or3_1
X_5588_ ih.gpio_interrupt_mask\[3\] _2326_ _2404_ _2125_ _2327_ VGND VGND VPWR VPWR
+ _2405_ sky130_fd_sc_hd__a221o_1
XFILLER_0_60_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4539_ _1296_ _1591_ _1592_ VGND VGND VPWR VPWR _1593_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5105__A0 cu.reg_file.reg_e\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5656__A1 net131 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5656__B2 net139 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6209_ clknet_leaf_4_clk net7 net171 VGND VGND VPWR VPWR ih.ih.ih.prev_data\[14\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_690 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_5_clk_A clknet_2_2__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5895__A1 _0618_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output49_A net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4890_ _2920_ cu.pc.pc_o\[7\] VGND VGND VPWR VPWR _1885_ sky130_fd_sc_hd__nor2_1
X_3910_ _0526_ net144 VGND VGND VPWR VPWR _0986_ sky130_fd_sc_hd__nand2_4
XANTENNA__4490__B _1545_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5078__S _2039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3841_ _0401_ _0916_ VGND VGND VPWR VPWR _0917_ sky130_fd_sc_hd__nand2_1
XANTENNA__4386__A1 cu.reg_file.reg_c\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3772_ cu.pc.pc_o\[13\] _0740_ _0846_ _0847_ VGND VGND VPWR VPWR _0848_ sky130_fd_sc_hd__a211o_1
X_5511_ net64 _2277_ _2179_ net65 VGND VGND VPWR VPWR _2331_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5335__A0 _1075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6194__RESET_B net162 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4138__A1 _0916_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5442_ _2271_ VGND VGND VPWR VPWR _0188_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_73_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5373_ _1188_ net119 _2226_ VGND VGND VPWR VPWR _2230_ sky130_fd_sc_hd__mux2_1
XFILLER_0_22_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4649__C _1672_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4324_ cu.reg_file.reg_l\[3\] _1317_ VGND VGND VPWR VPWR _1389_ sky130_fd_sc_hd__and2_1
X_4255_ _1268_ _1302_ VGND VGND VPWR VPWR _1323_ sky130_fd_sc_hd__nand2_4
XFILLER_0_38_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3206_ _2940_ _2942_ VGND VGND VPWR VPWR _2943_ sky130_fd_sc_hd__nor2_1
X_4186_ _1127_ _1236_ _1238_ _1255_ VGND VGND VPWR VPWR _1256_ sky130_fd_sc_hd__a31o_2
X_3137_ cu.id.alu_opcode\[1\] cu.id.alu_opcode\[0\] cu.id.alu_opcode\[3\] VGND VGND
+ VPWR VPWR _2874_ sky130_fd_sc_hd__and3_2
XTAP_1119 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1108 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3068_ ih.t.timer_max\[15\] _2755_ VGND VGND VPWR VPWR _2806_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_432 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5574__A0 cu.reg_file.reg_mem\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5709_ net8 _1650_ _2488_ _2513_ VGND VGND VPWR VPWR _0213_ sky130_fd_sc_hd__a31o_1
XANTENNA__5326__A0 _1261_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5877__A1 _1667_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4065__B1 _0652_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4591__A _1455_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3812__B1 _0624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4368__B2 _0373_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4368__A1 cu.reg_file.reg_sp\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3591__A2 _0413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4540__A1 cu.pc.pc_o\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4040_ _0610_ _1111_ _1112_ _1113_ VGND VGND VPWR VPWR _1114_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_91_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5991_ clknet_leaf_33_clk _0029_ net161 VGND VGND VPWR VPWR cu.pc.pc_o\[13\] sky130_fd_sc_hd__dfrtp_4
X_4942_ _1918_ _1923_ _1919_ VGND VGND VPWR VPWR _1933_ sky130_fd_sc_hd__a21bo_1
XANTENNA__3803__B1 _0624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4873_ _1862_ _1869_ _1809_ VGND VGND VPWR VPWR _1870_ sky130_fd_sc_hd__mux2_1
XANTENNA__5556__B1 _2247_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3824_ _0892_ _0895_ _0898_ _0899_ VGND VGND VPWR VPWR _0900_ sky130_fd_sc_hd__a2bb2o_1
X_3755_ cu.reg_file.reg_b\[7\] _0426_ _0429_ cu.reg_file.reg_d\[7\] VGND VGND VPWR
+ VPWR _0831_ sky130_fd_sc_hd__a22o_1
X_3686_ _0694_ _0701_ VGND VGND VPWR VPWR _0762_ sky130_fd_sc_hd__xor2_1
XANTENNA__3582__A2 _0502_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5425_ _2139_ _2180_ VGND VGND VPWR VPWR _2260_ sky130_fd_sc_hd__nand2_1
XFILLER_0_64_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5356_ _1190_ net112 _2215_ VGND VGND VPWR VPWR _2220_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5271__S _2170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5287_ _1329_ _1354_ VGND VGND VPWR VPWR _2179_ sky130_fd_sc_hd__nor2_2
X_4307_ _1306_ _1362_ _1367_ VGND VGND VPWR VPWR _1373_ sky130_fd_sc_hd__o21a_1
XANTENNA__3580__A cu.pc.pc_o\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4238_ _1305_ VGND VGND VPWR VPWR _1306_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4169_ _0829_ _0838_ _1060_ VGND VGND VPWR VPWR _1239_ sky130_fd_sc_hd__mux2_1
XFILLER_0_92_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3474__B _0384_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4522__B2 cu.reg_file.reg_d\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4522__A1 cu.pc.pc_o\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4586__A _1434_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5538__B1 _2225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4210__B1 _0293_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5356__S _2215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3540_ _0518_ _0568_ _0571_ _0615_ VGND VGND VPWR VPWR _0616_ sky130_fd_sc_hd__or4b_1
XFILLER_0_24_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_24_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5210_ _2126_ VGND VGND VPWR VPWR _2127_ sky130_fd_sc_hd__buf_2
X_3471_ _0399_ _0546_ VGND VGND VPWR VPWR _0547_ sky130_fd_sc_hd__nor2_2
XFILLER_0_24_398 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6190_ clknet_leaf_20_clk _0223_ net189 VGND VGND VPWR VPWR mc.cl.next_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_50_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5141_ _1624_ _1126_ _2066_ VGND VGND VPWR VPWR _2081_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5072_ _1790_ _0348_ _0351_ VGND VGND VPWR VPWR _2034_ sky130_fd_sc_hd__or3_2
X_4023_ _0918_ _1096_ VGND VGND VPWR VPWR _1097_ sky130_fd_sc_hd__and2_1
XFILLER_0_79_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5974_ clknet_leaf_32_clk _0011_ net161 VGND VGND VPWR VPWR cu.alu_f\[4\] sky130_fd_sc_hd__dfrtp_1
X_4925_ _1521_ _1907_ VGND VGND VPWR VPWR _1917_ sky130_fd_sc_hd__xor2_1
X_4856_ _1841_ _1844_ _1842_ VGND VGND VPWR VPWR _1854_ sky130_fd_sc_hd__o21a_1
XFILLER_0_51_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_30_clk_A clknet_2_3__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_34_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3807_ cu.reg_file.reg_sp\[10\] _0636_ _0748_ cu.reg_file.reg_h\[2\] VGND VGND VPWR
+ VPWR _0883_ sky130_fd_sc_hd__a22o_1
XANTENNA__5266__S _1666_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4787_ _0343_ _1299_ VGND VGND VPWR VPWR _1789_ sky130_fd_sc_hd__xor2_1
XFILLER_0_15_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3738_ _0801_ _0812_ _0798_ VGND VGND VPWR VPWR _0814_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_30_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_42_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3669_ cu.pc.pc_o\[8\] _0740_ _0742_ _0744_ VGND VGND VPWR VPWR _0745_ sky130_fd_sc_hd__a211o_1
X_5408_ _2250_ VGND VGND VPWR VPWR _0175_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4504__B2 cu.reg_file.reg_b\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4504__A1 cu.reg_file.reg_h\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5339_ _1190_ net104 _2206_ VGND VGND VPWR VPWR _2211_ sky130_fd_sc_hd__mux2_1
XANTENNA__4853__B cu.pc.pc_o\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5940__A0 _0341_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3932__B _0986_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_508 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_519 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3482__A1 _0547_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3379__B _2923_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2971_ net4 VGND VGND VPWR VPWR _2710_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4710_ net215 _1723_ _1725_ VGND VGND VPWR VPWR ih.t.next_count\[25\] sky130_fd_sc_hd__a21oi_1
X_5690_ ih.t.timer_max\[27\] _2151_ _2320_ ih.t.timer_max\[11\] VGND VGND VPWR VPWR
+ _2499_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_44_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4641_ ih.t.count\[0\] ih.t.count\[1\] ih.t.count\[2\] ih.t.count\[3\] VGND VGND
+ VPWR VPWR _1679_ sky130_fd_sc_hd__and4_1
XANTENNA__5086__S _2035_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4572_ _0516_ _1230_ VGND VGND VPWR VPWR _1623_ sky130_fd_sc_hd__nor2_8
X_6311_ clknet_leaf_36_clk _0004_ net158 VGND VGND VPWR VPWR cu.id.state\[0\] sky130_fd_sc_hd__dfrtp_1
X_3523_ _0598_ VGND VGND VPWR VPWR _0599_ sky130_fd_sc_hd__clkbuf_4
X_6242_ clknet_leaf_23_clk ih.t.next_count\[30\] net192 VGND VGND VPWR VPWR ih.t.count\[30\]
+ sky130_fd_sc_hd__dfrtp_2
X_3454_ _0519_ _0529_ VGND VGND VPWR VPWR _0530_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4938__B _1521_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4498__B1 _1284_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6173_ clknet_leaf_19_clk _0207_ net184 VGND VGND VPWR VPWR cu.reg_file.reg_mem\[9\]
+ sky130_fd_sc_hd__dfrtp_4
X_3385_ _2896_ _0324_ _2912_ _0346_ _2949_ VGND VGND VPWR VPWR _0461_ sky130_fd_sc_hd__o221a_1
X_5124_ _2067_ cu.reg_file.reg_h\[0\] _2069_ VGND VGND VPWR VPWR _2070_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout185_A net196 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4954__A _1233_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5055_ _2002_ _2024_ _2951_ VGND VGND VPWR VPWR _2025_ sky130_fd_sc_hd__o21a_4
X_4006_ _0817_ _1078_ _1079_ _0810_ VGND VGND VPWR VPWR _1080_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5957_ _2688_ VGND VGND VPWR VPWR _0286_ sky130_fd_sc_hd__clkbuf_1
X_4908_ _1900_ _1901_ VGND VGND VPWR VPWR _1902_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3776__A2 _0426_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5888_ _1191_ ih.t.timer_max\[5\] _2645_ VGND VGND VPWR VPWR _2651_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4839_ cu.pc.pc_o\[3\] _1826_ VGND VGND VPWR VPWR _1838_ sky130_fd_sc_hd__and2_1
XFILLER_0_62_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold20 ih.t.count\[28\] VGND VGND VPWR VPWR net216 sky130_fd_sc_hd__dlygate4sd3_1
Xhold31 ih.t.count\[6\] VGND VGND VPWR VPWR net227 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_42_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_93_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3519__A2 _0361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_6 _1188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5634__S _2351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_305 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_output79_A net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_327 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_316 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5141__A1 _1126_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3170_ cu.id.alu_opcode\[0\] cu.id.alu_opcode\[3\] cu.id.alu_opcode\[1\] VGND VGND
+ VPWR VPWR _2907_ sky130_fd_sc_hd__and3b_1
XANTENNA__4774__A _2948_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5811_ _2592_ _2593_ VGND VGND VPWR VPWR _2594_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_17_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5742_ _0296_ _0469_ VGND VGND VPWR VPWR _2533_ sky130_fd_sc_hd__or2_1
XANTENNA__3758__A2 _0488_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2954_ mc.rw.state\[1\] VGND VGND VPWR VPWR _2695_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5673_ _2482_ _2483_ _2485_ _1641_ VGND VGND VPWR VPWR _2486_ sky130_fd_sc_hd__o22a_4
X_4624_ _1665_ VGND VGND VPWR VPWR _1666_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_32_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4555_ cu.id.imm_i\[15\] _1294_ _1297_ cu.pc.pc_o\[15\] _1489_ VGND VGND VPWR VPWR
+ _1608_ sky130_fd_sc_hd__a221o_1
XANTENNA__4949__A cu.pc.pc_o\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3506_ _0341_ _0443_ _0336_ VGND VGND VPWR VPWR _0582_ sky130_fd_sc_hd__a21o_1
X_4486_ cu.pc.pc_o\[11\] _1321_ _1314_ cu.reg_file.reg_d\[3\] _1542_ VGND VGND VPWR
+ VPWR _1543_ sky130_fd_sc_hd__a221o_1
X_6225_ clknet_leaf_11_clk ih.t.next_count\[13\] net177 VGND VGND VPWR VPWR ih.t.count\[13\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__5132__A1 _1089_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3437_ alu.Cin _0512_ _0510_ VGND VGND VPWR VPWR _0513_ sky130_fd_sc_hd__a21o_1
X_6156_ clknet_leaf_16_clk _0190_ net181 VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__dfrtp_1
XTAP_861 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3368_ _0442_ _0437_ _0443_ VGND VGND VPWR VPWR _0444_ sky130_fd_sc_hd__a21o_1
XTAP_894 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_883 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_872 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5107_ cu.reg_file.reg_e\[2\] _1074_ _2056_ VGND VGND VPWR VPWR _2059_ sky130_fd_sc_hd__mux2_1
XANTENNA__5499__B _2193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6087_ clknet_leaf_5_clk _0121_ net168 VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__dfrtp_4
X_3299_ _0373_ _0374_ VGND VGND VPWR VPWR _0375_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5038_ cu.reg_file.reg_b\[3\] _2012_ _2006_ VGND VGND VPWR VPWR _2013_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3749__A2 _0488_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5371__A1 net118 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput43 net43 VGND VGND VPWR VPWR memory_address_out[2] sky130_fd_sc_hd__buf_2
Xoutput76 net76 VGND VGND VPWR VPWR ss0[0] sky130_fd_sc_hd__clkbuf_4
Xoutput65 net65 VGND VGND VPWR VPWR programmable_gpio_out[5] sky130_fd_sc_hd__clkbuf_4
Xoutput54 net54 VGND VGND VPWR VPWR memory_data_out[3] sky130_fd_sc_hd__clkbuf_4
XANTENNA__5123__A1 _2066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput87 net87 VGND VGND VPWR VPWR ss1[3] sky130_fd_sc_hd__clkbuf_4
Xoutput98 net98 VGND VGND VPWR VPWR ss2[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6241__RESET_B net194 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5584__A_N _1400_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3437__A1 alu.Cin VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_73_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5362__A1 net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4340_ _1400_ _1403_ _1404_ _1371_ VGND VGND VPWR VPWR _1405_ sky130_fd_sc_hd__a22o_1
X_4271_ cu.reg_file.reg_e\[1\] _1283_ _1285_ cu.reg_file.reg_l\[1\] _1337_ VGND VGND
+ VPWR VPWR _1338_ sky130_fd_sc_hd__a221o_1
XFILLER_0_94_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6010_ clknet_leaf_6_clk _0048_ net164 VGND VGND VPWR VPWR cu.reg_file.reg_c\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_3222_ _2892_ VGND VGND VPWR VPWR _0298_ sky130_fd_sc_hd__inv_2
X_3153_ cu.id.alu_opcode\[3\] cu.id.alu_opcode\[1\] VGND VGND VPWR VPWR _2890_ sky130_fd_sc_hd__and2b_1
X_3084_ ih.t.timer_max\[9\] _2751_ VGND VGND VPWR VPWR _2822_ sky130_fd_sc_hd__nand2_1
XANTENNA__3428__A1 _2948_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3986_ _0575_ VGND VGND VPWR VPWR _1060_ sky130_fd_sc_hd__clkbuf_4
X_5725_ _2518_ mc.cl.next_data\[1\] _2111_ VGND VGND VPWR VPWR _2523_ sky130_fd_sc_hd__and3_1
XFILLER_0_57_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3600__A1 cu.reg_file.reg_h\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_72_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5656_ net131 _2235_ _2246_ net139 VGND VGND VPWR VPWR _2469_ sky130_fd_sc_hd__a22o_1
X_4607_ mc.rw.state\[2\] mc.rw.state\[1\] mc.rw.state\[0\] VGND VGND VPWR VPWR _1651_
+ sky130_fd_sc_hd__nor3_1
XFILLER_0_72_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5587_ mc.cl.next_data\[3\] _2313_ net141 _2403_ VGND VGND VPWR VPWR _2404_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4398__B _1455_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4538_ cu.id.imm_i\[14\] _1295_ _1298_ cu.pc.pc_o\[14\] _1489_ VGND VGND VPWR VPWR
+ _1592_ sky130_fd_sc_hd__a221o_1
XFILLER_0_13_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4469_ cu.reg_file.reg_sp\[10\] _0992_ _1344_ cu.id.imm_i\[10\] _1324_ VGND VGND
+ VPWR VPWR _1527_ sky130_fd_sc_hd__a221o_1
XANTENNA__5105__A1 _1051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6208_ clknet_leaf_5_clk net6 net169 VGND VGND VPWR VPWR ih.ih.ih.prev_data\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__4864__B1 cu.pc.pc_o\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6139_ clknet_leaf_19_clk _0173_ net184 VGND VGND VPWR VPWR net131 sky130_fd_sc_hd__dfrtp_4
XTAP_691 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_680 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5041__A0 cu.reg_file.reg_b\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4304__C1 _1369_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_488 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5032__A0 cu.reg_file.reg_b\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3840_ _0774_ _0775_ VGND VGND VPWR VPWR _0916_ sky130_fd_sc_hd__and2_2
XFILLER_0_6_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3771_ cu.reg_file.reg_b\[5\] _0743_ _0624_ cu.reg_file.reg_sp\[13\] VGND VGND VPWR
+ VPWR _0847_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5510_ net68 _1648_ _2137_ _2274_ VGND VGND VPWR VPWR _2330_ sky130_fd_sc_hd__a31o_1
XFILLER_0_81_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5441_ _2022_ net74 _2270_ VGND VGND VPWR VPWR _2271_ sky130_fd_sc_hd__mux2_1
X_5372_ _2229_ VGND VGND VPWR VPWR _0160_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5099__A0 cu.reg_file.reg_d\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4323_ cu.id.cb_opcode_y\[0\] _1295_ _1298_ cu.pc.pc_o\[3\] _1305_ VGND VGND VPWR
+ VPWR _1388_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4254_ _1321_ VGND VGND VPWR VPWR _1322_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__3649__B2 cu.reg_file.reg_h\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3649__A1 cu.reg_file.reg_sp\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3205_ _2902_ _2936_ _2885_ _2941_ VGND VGND VPWR VPWR _2942_ sky130_fd_sc_hd__and4_2
X_4185_ _0387_ _1234_ _1254_ VGND VGND VPWR VPWR _1255_ sky130_fd_sc_hd__and3_1
X_3136_ _2745_ _2869_ _2871_ net140 net203 VGND VGND VPWR VPWR _0000_ sky130_fd_sc_hd__a32o_1
XFILLER_0_96_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3067_ ih.t.count\[16\] _2804_ VGND VGND VPWR VPWR _2805_ sky130_fd_sc_hd__xnor2_1
XTAP_1109 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5271__A0 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_18_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5574__A1 _2391_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5708_ _2512_ _1643_ cu.reg_file.reg_mem\[15\] _1646_ VGND VGND VPWR VPWR _2513_
+ sky130_fd_sc_hd__a2bb2o_1
X_3969_ _0611_ VGND VGND VPWR VPWR _1044_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5326__A1 net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5639_ net106 _2204_ _2452_ _1401_ VGND VGND VPWR VPWR _2453_ sky130_fd_sc_hd__a22o_1
XANTENNA__5877__A2 _2180_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4837__A0 cu.pc.pc_o\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4591__B _1473_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3812__A1 cu.reg_file.reg_b\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3812__B2 cu.reg_file.reg_sp\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5014__A0 _1191_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4368__A2 _0993_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5565__B2 ih.t.timer_max\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3000__B net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_514 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3951__A _2951_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output61_A net61 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5990_ clknet_leaf_28_clk _0028_ net188 VGND VGND VPWR VPWR cu.pc.pc_o\[12\] sky130_fd_sc_hd__dfstp_2
XFILLER_0_59_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5089__S _2035_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4941_ _2920_ cu.pc.pc_o\[11\] VGND VGND VPWR VPWR _1932_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3803__A1 cu.reg_file.reg_b\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3803__B2 cu.reg_file.reg_sp\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4872_ _1867_ _1868_ _1799_ VGND VGND VPWR VPWR _1869_ sky130_fd_sc_hd__mux2_1
XANTENNA__5005__A0 _1074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5556__A1 net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3823_ _0747_ _0751_ VGND VGND VPWR VPWR _0899_ sky130_fd_sc_hd__nor2_1
XANTENNA__5556__B2 net134 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_213 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_27_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3754_ cu.reg_file.reg_sp\[15\] _0636_ _0748_ cu.reg_file.reg_h\[7\] VGND VGND VPWR
+ VPWR _0830_ sky130_fd_sc_hd__a22o_1
X_3685_ _0758_ _0760_ VGND VGND VPWR VPWR _0761_ sky130_fd_sc_hd__nand2_1
XANTENNA__3845__B _0892_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5424_ _2259_ VGND VGND VPWR VPWR _0182_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5355_ _2219_ VGND VGND VPWR VPWR _0153_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5286_ _2178_ VGND VGND VPWR VPWR _0125_ sky130_fd_sc_hd__clkbuf_1
X_4306_ _1348_ VGND VGND VPWR VPWR _1372_ sky130_fd_sc_hd__inv_2
X_4237_ _1304_ VGND VGND VPWR VPWR _1305_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__3580__B _0501_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_4_clk_A clknet_2_0__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4168_ _1144_ _1160_ _1237_ VGND VGND VPWR VPWR _1238_ sky130_fd_sc_hd__nor3_1
X_3119_ _2797_ _2799_ _2800_ _2856_ VGND VGND VPWR VPWR _2857_ sky130_fd_sc_hd__or4_1
X_4099_ _0948_ _0959_ _0773_ VGND VGND VPWR VPWR _1173_ sky130_fd_sc_hd__o21a_1
XFILLER_0_81_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_65_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4867__A _0373_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4522__A2 _1321_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3797__B1 _0429_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4210__A1 _2877_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3470_ _0296_ _0528_ VGND VGND VPWR VPWR _0546_ sky130_fd_sc_hd__or2_2
XFILLER_0_86_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5140_ _2080_ VGND VGND VPWR VPWR _0077_ sky130_fd_sc_hd__clkbuf_1
X_5071_ _2033_ VGND VGND VPWR VPWR _0055_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5474__A0 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4022_ _0768_ _0772_ VGND VGND VPWR VPWR _1096_ sky130_fd_sc_hd__nand2_1
X_5973_ clknet_leaf_38_clk _0010_ net159 VGND VGND VPWR VPWR cu.alu_f\[3\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_87_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4924_ _1916_ VGND VGND VPWR VPWR _0025_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_59_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5529__A1 _1649_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4855_ _1851_ _1852_ VGND VGND VPWR VPWR _1853_ sky130_fd_sc_hd__and2b_1
XANTENNA__3004__A2 net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4786_ _1299_ VGND VGND VPWR VPWR _1788_ sky130_fd_sc_hd__inv_2
X_3806_ cu.id.imm_i\[10\] _0739_ _0881_ _0653_ VGND VGND VPWR VPWR _0882_ sky130_fd_sc_hd__a22o_2
X_3737_ _0801_ _0812_ _0798_ VGND VGND VPWR VPWR _0813_ sky130_fd_sc_hd__or3_1
XFILLER_0_70_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3668_ cu.reg_file.reg_b\[0\] _0743_ _0624_ cu.reg_file.reg_sp\[8\] VGND VGND VPWR
+ VPWR _0744_ sky130_fd_sc_hd__a22o_1
X_5407_ _1052_ net133 _2248_ VGND VGND VPWR VPWR _2250_ sky130_fd_sc_hd__mux2_1
XANTENNA__5701__A1 net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3599_ cu.reg_file.reg_l\[4\] _0621_ _0674_ VGND VGND VPWR VPWR _0675_ sky130_fd_sc_hd__a21o_1
X_5338_ _2210_ VGND VGND VPWR VPWR _0145_ sky130_fd_sc_hd__clkbuf_1
X_5269_ _1642_ VGND VGND VPWR VPWR _2169_ sky130_fd_sc_hd__buf_4
XANTENNA__5217__A0 _1188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5940__A1 _2391_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_509 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5920__S _2668_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4259__A1 cu.reg_file.reg_e\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2970_ net9 VGND VGND VPWR VPWR _2709_ sky130_fd_sc_hd__inv_2
XANTENNA__4431__A1 _1296_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5367__S _2226_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4640_ _1678_ VGND VGND VPWR VPWR ih.t.next_count\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_44_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4195__B1 _1263_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_491 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4571_ _2702_ _0619_ _1622_ _2697_ VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__a22o_1
X_6310_ clknet_leaf_30_clk _0292_ net183 VGND VGND VPWR VPWR cu.id.imm_i\[15\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__6202__D net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5989__RESET_B net188 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3522_ _0440_ _0589_ _0591_ _0593_ _0597_ VGND VGND VPWR VPWR _0598_ sky130_fd_sc_hd__o41a_4
X_6241_ clknet_leaf_22_clk ih.t.next_count\[29\] net194 VGND VGND VPWR VPWR ih.t.count\[29\]
+ sky130_fd_sc_hd__dfrtp_1
X_3453_ _0400_ _0528_ VGND VGND VPWR VPWR _0529_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6172_ clknet_leaf_19_clk _0206_ net183 VGND VGND VPWR VPWR cu.reg_file.reg_mem\[8\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__4498__B2 cu.reg_file.reg_h\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4498__A1 cu.reg_file.reg_b\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3384_ _0345_ _0450_ _0459_ VGND VGND VPWR VPWR _0460_ sky130_fd_sc_hd__or3b_2
X_5123_ _2066_ _2068_ _2951_ VGND VGND VPWR VPWR _2069_ sky130_fd_sc_hd__a21bo_4
XANTENNA__4954__B cu.pc.pc_o\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5054_ _2004_ _2023_ VGND VGND VPWR VPWR _2024_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4005_ _0817_ _0808_ _0776_ VGND VGND VPWR VPWR _1079_ sky130_fd_sc_hd__a21o_1
XANTENNA_fanout178_A net182 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5956_ cu.id.imm_i\[9\] _2372_ _2686_ VGND VGND VPWR VPWR _2688_ sky130_fd_sc_hd__mux2_1
X_5887_ _2650_ VGND VGND VPWR VPWR _0254_ sky130_fd_sc_hd__clkbuf_1
X_4907_ _1885_ _1888_ _1886_ VGND VGND VPWR VPWR _1901_ sky130_fd_sc_hd__o21a_1
XFILLER_0_47_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5277__S _2170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4838_ _1837_ VGND VGND VPWR VPWR _0018_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4769_ _1300_ _1644_ _1268_ VGND VGND VPWR VPWR _1776_ sky130_fd_sc_hd__o21a_1
XANTENNA__5922__A1 _2372_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold32 mc.cc.count\[1\] VGND VGND VPWR VPWR net228 sky130_fd_sc_hd__dlygate4sd3_1
Xhold21 ih.t.count\[16\] VGND VGND VPWR VPWR net217 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5438__A0 _2022_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold10 cu.id.is_halted VGND VGND VPWR VPWR net206 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4583__C _1598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4880__A _0387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3496__A alu.Cin VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4177__A0 _0663_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_7 _2496_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3943__B _0986_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4120__A _1144_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_306 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3662__C _0536_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_328 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5429__A0 _2022_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4774__B _0986_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5810_ _2583_ _2586_ _2584_ VGND VGND VPWR VPWR _2593_ sky130_fd_sc_hd__a21bo_1
XANTENNA__4404__A1 cu.reg_file.reg_e\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5741_ _1007_ _0981_ _0989_ _0994_ VGND VGND VPWR VPWR _2532_ sky130_fd_sc_hd__or4b_4
XANTENNA__4404__B2 cu.reg_file.reg_l\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5672_ _1649_ _2484_ VGND VGND VPWR VPWR _2485_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4623_ _0315_ _1658_ _1659_ VGND VGND VPWR VPWR _1665_ sky130_fd_sc_hd__or3b_4
XFILLER_0_44_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4554_ cu.reg_file.reg_b\[7\] net143 _1284_ cu.reg_file.reg_h\[7\] _1606_ VGND VGND
+ VPWR VPWR _1607_ sky130_fd_sc_hd__a221o_1
XANTENNA__3391__A1 _2923_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3505_ cu.reg_file.reg_l\[2\] _0422_ _0577_ _0579_ _0580_ VGND VGND VPWR VPWR _0581_
+ sky130_fd_sc_hd__a2111o_1
XANTENNA__4668__C _1672_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6224_ clknet_leaf_11_clk ih.t.next_count\[12\] net177 VGND VGND VPWR VPWR ih.t.count\[12\]
+ sky130_fd_sc_hd__dfrtp_1
X_4485_ cu.reg_file.reg_sp\[11\] _0992_ _1343_ cu.id.imm_i\[11\] _1324_ VGND VGND
+ VPWR VPWR _1542_ sky130_fd_sc_hd__a221o_1
X_3436_ _0395_ _0400_ VGND VGND VPWR VPWR _0512_ sky130_fd_sc_hd__nor2_2
XFILLER_0_0_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6155_ clknet_leaf_8_clk _0189_ net168 VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__dfrtp_2
XTAP_862 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4965__A _1233_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3367_ _0328_ _0334_ VGND VGND VPWR VPWR _0443_ sky130_fd_sc_hd__or2_1
X_6086_ clknet_leaf_9_clk _0120_ net174 VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__dfrtp_1
XTAP_895 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_884 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_873 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5106_ _2058_ VGND VGND VPWR VPWR _0065_ sky130_fd_sc_hd__clkbuf_1
X_5037_ _1187_ _1222_ _2002_ VGND VGND VPWR VPWR _2012_ sky130_fd_sc_hd__mux2_1
X_3298_ cu.id.cb_opcode_y\[1\] VGND VGND VPWR VPWR _0374_ sky130_fd_sc_hd__buf_4
XFILLER_0_94_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5939_ _2678_ VGND VGND VPWR VPWR _0278_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_63_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4205__A _0359_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_23_409 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput44 net44 VGND VGND VPWR VPWR memory_address_out[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_9_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput55 net55 VGND VGND VPWR VPWR memory_data_out[4] sky130_fd_sc_hd__clkbuf_4
Xoutput66 net66 VGND VGND VPWR VPWR programmable_gpio_out[6] sky130_fd_sc_hd__clkbuf_4
Xoutput77 net77 VGND VGND VPWR VPWR ss0[1] sky130_fd_sc_hd__buf_2
Xoutput99 net99 VGND VGND VPWR VPWR ss2[7] sky130_fd_sc_hd__buf_2
Xoutput88 net88 VGND VGND VPWR VPWR ss1[4] sky130_fd_sc_hd__clkbuf_4
XANTENNA__3003__B net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4115__A _1187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output91_A net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4270_ cu.reg_file.reg_a\[1\] _1276_ _1287_ cu.reg_file.reg_sp\[1\] VGND VGND VPWR
+ VPWR _1337_ sky130_fd_sc_hd__a22o_1
X_3221_ _2925_ _2932_ _2904_ VGND VGND VPWR VPWR _0297_ sky130_fd_sc_hd__o21ai_2
X_3152_ cu.id.opcode\[0\] cu.id.opcode\[2\] cu.id.opcode\[1\] VGND VGND VPWR VPWR
+ _2889_ sky130_fd_sc_hd__and3_1
X_3083_ ih.t.count\[10\] _2820_ VGND VGND VPWR VPWR _2821_ sky130_fd_sc_hd__xnor2_1
XANTENNA__3428__A2 _0501_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3985_ _0603_ VGND VGND VPWR VPWR _1059_ sky130_fd_sc_hd__inv_2
X_5724_ net18 _2519_ _2522_ VGND VGND VPWR VPWR _0219_ sky130_fd_sc_hd__a21o_1
XFILLER_0_17_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3600__A2 _0495_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5655_ _2468_ VGND VGND VPWR VPWR _0204_ sky130_fd_sc_hd__clkbuf_1
X_4606_ _1649_ VGND VGND VPWR VPWR _1650_ sky130_fd_sc_hd__clkbuf_4
X_5586_ _1666_ _2401_ _2402_ VGND VGND VPWR VPWR _2403_ sky130_fd_sc_hd__o21a_1
XFILLER_0_13_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4537_ cu.reg_file.reg_b\[6\] _1281_ _1285_ cu.reg_file.reg_h\[6\] _1590_ VGND VGND
+ VPWR VPWR _1591_ sky130_fd_sc_hd__a221o_1
XFILLER_0_40_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4468_ _1521_ _1485_ _1525_ VGND VGND VPWR VPWR _1526_ sky130_fd_sc_hd__o21a_1
XFILLER_0_68_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6207_ clknet_leaf_5_clk net5 net172 VGND VGND VPWR VPWR ih.ih.ih.prev_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3419_ net146 _0473_ _0479_ _0463_ _0458_ VGND VGND VPWR VPWR _0495_ sky130_fd_sc_hd__o2111a_4
X_4399_ _1455_ _1459_ _1460_ _1371_ VGND VGND VPWR VPWR _1461_ sky130_fd_sc_hd__a22o_1
X_6138_ clknet_leaf_27_clk _0172_ net187 VGND VGND VPWR VPWR net130 sky130_fd_sc_hd__dfrtp_4
XANTENNA__4864__A1 cu.pc.pc_o\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_670 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_681 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6069_ clknet_leaf_17_clk _0103_ net172 VGND VGND VPWR VPWR ih.gpio_interrupt_mask\[2\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__6039__RESET_B net161 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5813__A0 cu.reg_file.reg_sp\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4589__B _1401_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3355__A1 cu.reg_file.reg_c\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3355__B2 cu.reg_file.reg_e\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5501__C1 _1660_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3014__A ih.t.timer_max\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5804__A0 _1622_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4771__C _1646_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5583__A2 _2193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3770_ cu.reg_file.reg_d\[5\] _0488_ _0741_ cu.reg_file.reg_h\[5\] VGND VGND VPWR
+ VPWR _0846_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5440_ _2139_ _2236_ VGND VGND VPWR VPWR _2270_ sky130_fd_sc_hd__nand2_1
XANTENNA__5375__S _2226_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5371_ _1075_ net118 _2226_ VGND VGND VPWR VPWR _2229_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6210__D net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4322_ _1271_ _1386_ VGND VGND VPWR VPWR _1387_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4253_ _1319_ _1320_ VGND VGND VPWR VPWR _1321_ sky130_fd_sc_hd__nor2_2
X_3204_ cu.id.opcode\[2\] cu.id.opcode\[1\] _2875_ _2876_ VGND VGND VPWR VPWR _2941_
+ sky130_fd_sc_hd__and4bb_2
XANTENNA__3649__A2 _0413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4184_ _0701_ _1245_ _1253_ VGND VGND VPWR VPWR _1254_ sky130_fd_sc_hd__a21o_1
XFILLER_0_38_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3135_ net1 _2872_ _2870_ VGND VGND VPWR VPWR _2873_ sky130_fd_sc_hd__nor3_1
X_3066_ ih.t.timer_max\[16\] _2756_ VGND VGND VPWR VPWR _2804_ sky130_fd_sc_hd__xor2_1
XANTENNA__6132__RESET_B net195 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5271__A1 _2085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout160_A net162 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3968_ _0599_ _0603_ _0606_ _1042_ VGND VGND VPWR VPWR _1043_ sky130_fd_sc_hd__o22a_1
XFILLER_0_45_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5707_ mc.cl.next_data\[15\] _2359_ _2490_ _2511_ VGND VGND VPWR VPWR _2512_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_45_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5285__S _2170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_45_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3899_ _0359_ _0973_ _0364_ _0974_ _0296_ VGND VGND VPWR VPWR _0975_ sky130_fd_sc_hd__a221o_1
X_5638_ net90 _1330_ VGND VGND VPWR VPWR _2452_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5569_ _2169_ _2379_ _2386_ _2136_ VGND VGND VPWR VPWR _2387_ sky130_fd_sc_hd__o211a_1
XFILLER_0_13_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3812__A2 _0743_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3567__A1_N _0576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5014__A1 _1209_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_301 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3951__B _0368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output54_A net54 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4940_ _1929_ _1930_ VGND VGND VPWR VPWR _1931_ sky130_fd_sc_hd__nor2_1
XANTENNA__3803__A2 _0743_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4871_ _1144_ _1862_ _1795_ VGND VGND VPWR VPWR _1868_ sky130_fd_sc_hd__mux2_1
XANTENNA__5005__A1 _1226_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6205__D net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3822_ _0896_ _0897_ VGND VGND VPWR VPWR _0898_ sky130_fd_sc_hd__nand2_2
XFILLER_0_39_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5556__A2 _2236_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3753_ cu.id.imm_i\[15\] _0739_ _0828_ _0653_ VGND VGND VPWR VPWR _0829_ sky130_fd_sc_hd__a22oi_4
X_3684_ _0714_ _0759_ VGND VGND VPWR VPWR _0760_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5423_ net68 _2085_ _2258_ VGND VGND VPWR VPWR _2259_ sky130_fd_sc_hd__mux2_1
XANTENNA__4516__B1 _1286_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5354_ _1188_ net111 _2215_ VGND VGND VPWR VPWR _2219_ sky130_fd_sc_hd__mux2_1
X_4305_ _2701_ VGND VGND VPWR VPWR _1371_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_49_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5285_ net83 _1260_ _2170_ VGND VGND VPWR VPWR _2178_ sky130_fd_sc_hd__mux2_1
XANTENNA__4819__A1 _0343_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4236_ _2946_ _1303_ VGND VGND VPWR VPWR _1304_ sky130_fd_sc_hd__nor2_2
XFILLER_0_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5492__A1 net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4167_ _0617_ _1050_ _1073_ _1089_ VGND VGND VPWR VPWR _1237_ sky130_fd_sc_hd__or4_1
X_3118_ _2802_ _2803_ _2855_ VGND VGND VPWR VPWR _2856_ sky130_fd_sc_hd__or3_1
XANTENNA__5244__A1 _1661_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4098_ _0916_ _0946_ _1171_ _1032_ _0918_ VGND VGND VPWR VPWR _1172_ sky130_fd_sc_hd__o221a_1
X_3049_ _2761_ _2785_ ih.t.count\[23\] VGND VGND VPWR VPWR _2787_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4213__A _1280_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4867__B cu.pc.pc_o\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4586__C _1473_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3797__B2 cu.reg_file.reg_d\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3797__A1 cu.reg_file.reg_b\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5538__A2 _2147_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4123__A _1126_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5070_ cu.reg_file.reg_c\[7\] _1260_ _2025_ VGND VGND VPWR VPWR _2033_ sky130_fd_sc_hd__mux2_1
XANTENNA__5474__A1 _2085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4021_ _1093_ _1094_ VGND VGND VPWR VPWR _1095_ sky130_fd_sc_hd__nor2_1
XANTENNA__3485__B1 _0492_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5972_ clknet_leaf_35_clk _0009_ net159 VGND VGND VPWR VPWR cu.alu_f\[2\] sky130_fd_sc_hd__dfrtp_1
X_4923_ cu.pc.pc_o\[9\] _1915_ _1815_ VGND VGND VPWR VPWR _1916_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3788__A1 cu.reg_file.reg_mem\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4732__S _0359_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4017__B _0773_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4854_ _0374_ cu.pc.pc_o\[4\] VGND VGND VPWR VPWR _1852_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4785_ net199 _1787_ VGND VGND VPWR VPWR _0001_ sky130_fd_sc_hd__nor2_1
X_3805_ cu.reg_file.reg_a\[2\] _0625_ _0628_ cu.reg_file.reg_mem\[10\] _0880_ VGND
+ VGND VPWR VPWR _0881_ sky130_fd_sc_hd__a221o_1
X_3736_ _0802_ _0804_ _0811_ VGND VGND VPWR VPWR _0812_ sky130_fd_sc_hd__or3_2
XFILLER_0_27_183 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4752__A3 _2935_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3667_ _0464_ _0480_ VGND VGND VPWR VPWR _0743_ sky130_fd_sc_hd__and2_2
X_5406_ _2249_ VGND VGND VPWR VPWR _0174_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5701__A2 _1650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3598_ cu.reg_file.reg_c\[4\] _0485_ _0489_ cu.reg_file.reg_e\[4\] VGND VGND VPWR
+ VPWR _0674_ sky130_fd_sc_hd__a22o_1
X_5337_ _1188_ net103 _2206_ VGND VGND VPWR VPWR _2210_ sky130_fd_sc_hd__mux2_1
X_5268_ _2168_ VGND VGND VPWR VPWR _0117_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5799__A cu.reg_file.reg_sp\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4219_ _1286_ VGND VGND VPWR VPWR _1287_ sky130_fd_sc_hd__clkbuf_4
X_5199_ net210 _2708_ _2119_ mc.cc.enable_edge_detector.prev_data VGND VGND VPWR VPWR
+ _0097_ sky130_fd_sc_hd__a22o_1
XFILLER_0_78_540 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5311__B _2194_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4976__B1 cu.pc.pc_o\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5153__A0 cu.reg_file.reg_l\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4118__A _1189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5392__A0 _1188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4570_ _0824_ _0819_ VGND VGND VPWR VPWR _1622_ sky130_fd_sc_hd__and2_4
XANTENNA__4195__A1 _0516_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4195__B2 _1027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3521_ _0293_ _0596_ _0440_ VGND VGND VPWR VPWR _0597_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_52_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5144__A0 _1263_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_3_clk_A clknet_2_0__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6240_ clknet_leaf_22_clk ih.t.next_count\[28\] net194 VGND VGND VPWR VPWR ih.t.count\[28\]
+ sky130_fd_sc_hd__dfrtp_2
X_3452_ _0527_ VGND VGND VPWR VPWR _0528_ sky130_fd_sc_hd__buf_2
X_3383_ _2889_ _0301_ _2933_ VGND VGND VPWR VPWR _0459_ sky130_fd_sc_hd__or3_1
X_6171_ clknet_leaf_37_clk _0205_ net159 VGND VGND VPWR VPWR cu.reg_file.reg_mem\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_5122_ _0352_ _1792_ _1790_ VGND VGND VPWR VPWR _2068_ sky130_fd_sc_hd__or3b_1
X_5053_ _0350_ _0358_ _0366_ VGND VGND VPWR VPWR _2023_ sky130_fd_sc_hd__or3_1
X_4004_ _0808_ _0810_ VGND VGND VPWR VPWR _1078_ sky130_fd_sc_hd__nor2_1
XFILLER_0_94_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5955_ _2687_ VGND VGND VPWR VPWR _0285_ sky130_fd_sc_hd__clkbuf_1
X_5886_ _1189_ ih.t.timer_max\[4\] _2645_ VGND VGND VPWR VPWR _2650_ sky130_fd_sc_hd__mux2_1
X_4906_ _1898_ _1899_ VGND VGND VPWR VPWR _1900_ sky130_fd_sc_hd__or2_1
XFILLER_0_90_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4837_ cu.pc.pc_o\[2\] _1836_ _1815_ VGND VGND VPWR VPWR _1837_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4768_ net206 _1775_ VGND VGND VPWR VPWR _0005_ sky130_fd_sc_hd__nor2_1
XFILLER_0_15_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4699_ _1717_ _1718_ VGND VGND VPWR VPWR ih.t.next_count\[21\] sky130_fd_sc_hd__nor2_1
XANTENNA__5293__S _2182_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3719_ _0788_ _0794_ VGND VGND VPWR VPWR _0795_ sky130_fd_sc_hd__nand2_1
XANTENNA__5135__A0 _1213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5686__B2 ih.t.timer_max\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold22 ih.t.count\[30\] VGND VGND VPWR VPWR net218 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5438__A1 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold11 cu.alu_f\[3\] VGND VGND VPWR VPWR net207 sky130_fd_sc_hd__dlygate4sd3_1
Xhold33 ih.t.count\[8\] VGND VGND VPWR VPWR net229 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__5610__A1 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4880__B cu.pc.pc_o\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_53_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_8 _2919_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4401__A _1455_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5126__A0 _1623_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5677__B2 ih.t.timer_max\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_329 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_307 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5429__A1 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5232__A _1364_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5601__A1 net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3612__B1 _0499_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5740_ _2530_ _1050_ _2116_ VGND VGND VPWR VPWR _2531_ sky130_fd_sc_hd__mux2_1
XTAP_1090 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_17_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5671_ net15 _2345_ _2369_ net8 VGND VGND VPWR VPWR _2484_ sky130_fd_sc_hd__a22o_1
X_4622_ _1653_ VGND VGND VPWR VPWR _1664_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4553_ cu.reg_file.reg_d\[7\] _1282_ _1286_ cu.reg_file.reg_sp\[15\] VGND VGND VPWR
+ VPWR _1606_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4484_ cu.pc.pc_o\[11\] _1485_ _1540_ VGND VGND VPWR VPWR _1541_ sky130_fd_sc_hd__o21a_1
X_3504_ cu.reg_file.reg_mem\[2\] _0418_ _0419_ cu.reg_file.reg_h\[2\] VGND VGND VPWR
+ VPWR _0580_ sky130_fd_sc_hd__a22o_1
XANTENNA__5117__A0 cu.reg_file.reg_e\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6223_ clknet_leaf_11_clk ih.t.next_count\[11\] net176 VGND VGND VPWR VPWR ih.t.count\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_3435_ alu.Cin _0510_ VGND VGND VPWR VPWR _0511_ sky130_fd_sc_hd__nand2_1
XANTENNA__4340__A1 _1400_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6154_ clknet_leaf_9_clk _0188_ net175 VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__dfrtp_4
XTAP_852 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4965__B cu.pc.pc_o\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3366_ _0321_ VGND VGND VPWR VPWR _0442_ sky130_fd_sc_hd__inv_2
XANTENNA_fanout190_A net194 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6085_ clknet_leaf_9_clk _0119_ net174 VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__dfrtp_1
XTAP_885 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_874 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5105_ cu.reg_file.reg_e\[1\] _1051_ _2056_ VGND VGND VPWR VPWR _2058_ sky130_fd_sc_hd__mux2_1
X_3297_ cu.id.cb_opcode_y\[2\] VGND VGND VPWR VPWR _0373_ sky130_fd_sc_hd__clkbuf_4
XTAP_896 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5036_ _2011_ VGND VGND VPWR VPWR _0042_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5938_ _0340_ _2372_ _2666_ VGND VGND VPWR VPWR _2678_ sky130_fd_sc_hd__mux2_1
XANTENNA__3603__B1 _0492_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5869_ _2161_ ih.t.timer_max\[12\] _2636_ VGND VGND VPWR VPWR _2641_ sky130_fd_sc_hd__mux2_1
XANTENNA__5356__A0 _1190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5659__A1 net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5659__B2 _1401_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput45 net45 VGND VGND VPWR VPWR memory_address_out[4] sky130_fd_sc_hd__clkbuf_4
Xoutput56 net56 VGND VGND VPWR VPWR memory_data_out[5] sky130_fd_sc_hd__clkbuf_4
Xoutput67 net67 VGND VGND VPWR VPWR programmable_gpio_out[7] sky130_fd_sc_hd__clkbuf_4
Xoutput89 net89 VGND VGND VPWR VPWR ss1[5] sky130_fd_sc_hd__clkbuf_4
Xoutput78 net78 VGND VGND VPWR VPWR ss0[2] sky130_fd_sc_hd__clkbuf_4
XANTENNA__5052__A _0618_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4891__A _2920_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5926__S _2668_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output84_A net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3220_ _0295_ VGND VGND VPWR VPWR _0296_ sky130_fd_sc_hd__clkbuf_4
X_3151_ _2875_ _2876_ VGND VGND VPWR VPWR _2888_ sky130_fd_sc_hd__nor2_2
XFILLER_0_27_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3082_ ih.t.timer_max\[10\] _2752_ VGND VGND VPWR VPWR _2820_ sky130_fd_sc_hd__xor2_1
XANTENNA__6208__D net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4306__A _1348_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3984_ _0370_ _1052_ _1058_ VGND VGND VPWR VPWR _0008_ sky130_fd_sc_hd__a21o_1
X_5723_ _2518_ mc.cl.next_data\[0\] _2111_ VGND VGND VPWR VPWR _2522_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5654_ cu.reg_file.reg_mem\[6\] _2467_ _1739_ VGND VGND VPWR VPWR _2468_ sky130_fd_sc_hd__mux2_1
X_4605_ _1648_ VGND VGND VPWR VPWR _1649_ sky130_fd_sc_hd__buf_2
XFILLER_0_60_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5585_ ih.t.timer_max\[19\] _2150_ _2319_ ih.t.timer_max\[3\] _1661_ VGND VGND VPWR
+ VPWR _2402_ sky130_fd_sc_hd__a221o_1
XFILLER_0_13_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4536_ cu.reg_file.reg_d\[6\] _1283_ _1589_ VGND VGND VPWR VPWR _1590_ sky130_fd_sc_hd__a21bo_1
X_4467_ _1296_ _1523_ _1524_ VGND VGND VPWR VPWR _1525_ sky130_fd_sc_hd__a21o_1
XFILLER_0_40_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4398_ _1441_ _1455_ VGND VGND VPWR VPWR _1460_ sky130_fd_sc_hd__nor2_1
X_6206_ clknet_leaf_7_clk net4 net167 VGND VGND VPWR VPWR ih.ih.ih.prev_data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_3418_ _0482_ _0493_ VGND VGND VPWR VPWR _0494_ sky130_fd_sc_hd__and2_2
X_6137_ clknet_leaf_6_clk _0171_ net165 VGND VGND VPWR VPWR net129 sky130_fd_sc_hd__dfrtp_2
XTAP_660 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3349_ _0405_ _0412_ VGND VGND VPWR VPWR _0425_ sky130_fd_sc_hd__or2b_2
XTAP_693 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6068_ clknet_leaf_13_clk _0102_ net181 VGND VGND VPWR VPWR ih.gpio_interrupt_mask\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_5019_ _1998_ VGND VGND VPWR VPWR _0038_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_95_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output122_A net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3291__A1 _0350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_39_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3965__A _0710_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5370_ _2228_ VGND VGND VPWR VPWR _0159_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4543__A1 cu.reg_file.reg_h\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_134 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_22_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4543__B2 cu.reg_file.reg_b\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4321_ cu.reg_file.reg_c\[3\] _1281_ _1385_ VGND VGND VPWR VPWR _1386_ sky130_fd_sc_hd__a21oi_1
XANTENNA__4796__A _2948_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4252_ _0295_ _2914_ _0320_ _1310_ VGND VGND VPWR VPWR _1320_ sky130_fd_sc_hd__or4_1
XANTENNA__5404__B _2247_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3203_ _2938_ _2939_ VGND VGND VPWR VPWR _2940_ sky130_fd_sc_hd__nor2_2
XFILLER_0_38_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4183_ _0701_ _1252_ VGND VGND VPWR VPWR _1253_ sky130_fd_sc_hd__nor2_1
XFILLER_0_38_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3134_ _2745_ _2869_ VGND VGND VPWR VPWR _2872_ sky130_fd_sc_hd__or2b_1
X_3065_ ih.t.count\[17\] _2757_ _2801_ VGND VGND VPWR VPWR _2803_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6101__RESET_B net195 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_201 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3967_ _0599_ _1041_ VGND VGND VPWR VPWR _1042_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5706_ ih.t.timer_max\[31\] _2151_ _2320_ ih.t.timer_max\[15\] VGND VGND VPWR VPWR
+ _2511_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_70_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4782__A1 _0350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_30_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_30_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_60_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3898_ _0520_ VGND VGND VPWR VPWR _0974_ sky130_fd_sc_hd__inv_2
XFILLER_0_33_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5637_ net98 _2194_ _2450_ VGND VGND VPWR VPWR _2451_ sky130_fd_sc_hd__a21o_1
XFILLER_0_60_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5568_ ih.gpio_interrupt_mask\[2\] _2326_ _2385_ _2125_ _2327_ VGND VGND VPWR VPWR
+ _2386_ sky130_fd_sc_hd__a221o_1
X_4519_ _1296_ _1572_ _1573_ VGND VGND VPWR VPWR _1574_ sky130_fd_sc_hd__a21o_1
XFILLER_0_13_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5499_ _2180_ _2193_ VGND VGND VPWR VPWR _2319_ sky130_fd_sc_hd__or2_2
XTAP_490 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5330__A _2205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_21_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_21_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_36_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_538 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output47_A net47 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5789__A0 cu.reg_file.reg_sp\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4870_ _1865_ _1866_ VGND VGND VPWR VPWR _1867_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_24_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_86_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3821_ _0895_ _0892_ VGND VGND VPWR VPWR _0897_ sky130_fd_sc_hd__or2b_1
XANTENNA__5386__S _2237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_12_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_12_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_82_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3752_ cu.reg_file.reg_a\[7\] _0625_ _0628_ cu.reg_file.reg_mem\[15\] _0827_ VGND
+ VGND VPWR VPWR _0828_ sky130_fd_sc_hd__a221o_1
X_3683_ _0715_ _0711_ VGND VGND VPWR VPWR _0759_ sky130_fd_sc_hd__nand2b_2
X_5422_ _1306_ _2257_ _2137_ VGND VGND VPWR VPWR _2258_ sky130_fd_sc_hd__and3_1
XANTENNA__4516__A1 cu.reg_file.reg_d\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4516__B2 cu.reg_file.reg_sp\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5353_ _2218_ VGND VGND VPWR VPWR _0152_ sky130_fd_sc_hd__clkbuf_1
X_4304_ _2701_ _1354_ _1353_ _1369_ VGND VGND VPWR VPWR _1370_ sky130_fd_sc_hd__a211o_1
XFILLER_0_49_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5284_ _2177_ VGND VGND VPWR VPWR _0124_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4819__A2 _1299_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4235_ _1302_ VGND VGND VPWR VPWR _1303_ sky130_fd_sc_hd__inv_2
XANTENNA__5492__A2 _1633_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4166_ _1175_ _1200_ _1232_ _1235_ VGND VGND VPWR VPWR _1236_ sky130_fd_sc_hd__a31o_1
X_3117_ _2805_ _2807_ _2808_ _2854_ VGND VGND VPWR VPWR _2855_ sky130_fd_sc_hd__or4_1
XFILLER_0_65_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4097_ _0945_ _0946_ VGND VGND VPWR VPWR _1171_ sky130_fd_sc_hd__xor2_1
X_3048_ ih.t.count\[23\] _2761_ _2785_ VGND VGND VPWR VPWR _2786_ sky130_fd_sc_hd__and3_1
XFILLER_0_81_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4999_ _1984_ VGND VGND VPWR VPWR _1985_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_18_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4691__B1 _1670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3797__A2 _0426_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5934__S _2668_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4020_ _0801_ _0812_ VGND VGND VPWR VPWR _1094_ sky130_fd_sc_hd__and2_1
Xclkbuf_leaf_1_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_1_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__4682__B1 _1670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3485__B2 cu.reg_file.reg_d\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5564__A_N _1400_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5971_ clknet_leaf_35_clk _0008_ net159 VGND VGND VPWR VPWR cu.alu_f\[1\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_87_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4922_ _1909_ _1914_ _1809_ VGND VGND VPWR VPWR _1915_ sky130_fd_sc_hd__mux2_1
XANTENNA__3788__A2 _0640_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4853_ _0374_ cu.pc.pc_o\[4\] VGND VGND VPWR VPWR _1851_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_524 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4784_ _1000_ _1786_ cu.id.is_halted VGND VGND VPWR VPWR _1787_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3804_ cu.pc.pc_o\[10\] _0740_ _0878_ _0879_ VGND VGND VPWR VPWR _0880_ sky130_fd_sc_hd__a211o_1
XFILLER_0_15_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3735_ _0805_ _0808_ _0810_ VGND VGND VPWR VPWR _0811_ sky130_fd_sc_hd__or3_2
XFILLER_0_27_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5405_ _0619_ net132 _2248_ VGND VGND VPWR VPWR _2249_ sky130_fd_sc_hd__mux2_1
XFILLER_0_30_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3666_ cu.reg_file.reg_d\[0\] _0488_ _0741_ cu.reg_file.reg_h\[0\] VGND VGND VPWR
+ VPWR _0742_ sky130_fd_sc_hd__a22o_1
XFILLER_0_62_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3597_ _0374_ _0672_ _0294_ VGND VGND VPWR VPWR _0673_ sky130_fd_sc_hd__mux2_1
X_5336_ _2209_ VGND VGND VPWR VPWR _0144_ sky130_fd_sc_hd__clkbuf_1
X_5267_ ih.t.timer_max\[31\] _2167_ _2153_ VGND VGND VPWR VPWR _2168_ sky130_fd_sc_hd__mux2_1
X_4218_ _0295_ _0469_ VGND VGND VPWR VPWR _1286_ sky130_fd_sc_hd__nor2_4
X_5198_ mc.cc.count\[3\] _1652_ _2118_ VGND VGND VPWR VPWR _2119_ sky130_fd_sc_hd__o21ba_1
XANTENNA__4673__B1 _1670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4149_ _0941_ _1218_ VGND VGND VPWR VPWR _1219_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_552 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4976__A1 cu.pc.pc_o\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5153__A1 _1051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4664__B1 _1670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3467__A1 cu.reg_file.reg_sp\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3957__B _0528_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5392__A1 net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4195__A2 _1260_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3520_ _0594_ _0595_ VGND VGND VPWR VPWR _0596_ sky130_fd_sc_hd__nand2_1
XANTENNA__5144__A1 _1110_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3451_ _0521_ _0524_ _0525_ _0526_ VGND VGND VPWR VPWR _0527_ sky130_fd_sc_hd__and4b_1
X_3382_ net147 _0454_ _0457_ VGND VGND VPWR VPWR _0458_ sky130_fd_sc_hd__a21oi_4
X_6170_ clknet_2_1__leaf_clk _0204_ net161 VGND VGND VPWR VPWR cu.reg_file.reg_mem\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_5121_ _1622_ _0617_ _2066_ VGND VGND VPWR VPWR _2067_ sky130_fd_sc_hd__mux2_1
X_5052_ _0618_ VGND VGND VPWR VPWR _2022_ sky130_fd_sc_hd__buf_2
XFILLER_0_46_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4003_ _0764_ _1064_ VGND VGND VPWR VPWR _1077_ sky130_fd_sc_hd__nor2_1
XFILLER_0_87_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_75_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5954_ cu.id.imm_i\[8\] _2350_ _2686_ VGND VGND VPWR VPWR _2687_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5080__A0 _1051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5885_ _2649_ VGND VGND VPWR VPWR _0253_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4905_ cu.id.cb_opcode_x\[1\] cu.pc.pc_o\[8\] VGND VGND VPWR VPWR _1899_ sky130_fd_sc_hd__and2_1
XANTENNA__3630__B2 cu.reg_file.reg_mem\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4836_ _1828_ _1835_ _1809_ VGND VGND VPWR VPWR _1836_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_90_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4767_ _1483_ _1632_ _1643_ _1771_ _1774_ VGND VGND VPWR VPWR _1775_ sky130_fd_sc_hd__o311a_1
XFILLER_0_7_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5574__S _2351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4698_ net233 _1714_ _1687_ VGND VGND VPWR VPWR _1718_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3718_ _0664_ _0682_ _0793_ VGND VGND VPWR VPWR _0794_ sky130_fd_sc_hd__a21o_1
XFILLER_0_43_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3649_ cu.reg_file.reg_sp\[7\] _0413_ _0419_ cu.reg_file.reg_h\[7\] _0724_ VGND VGND
+ VPWR VPWR _0725_ sky130_fd_sc_hd__a221o_1
XANTENNA__5135__A1 _1160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5319_ _2199_ VGND VGND VPWR VPWR _0137_ sky130_fd_sc_hd__clkbuf_1
Xhold23 ih.t.count\[4\] VGND VGND VPWR VPWR net219 sky130_fd_sc_hd__dlygate4sd3_1
X_6299_ clknet_leaf_37_clk _0281_ net159 VGND VGND VPWR VPWR cu.id.cb_opcode_y\[1\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold12 cu.alu_f\[5\] VGND VGND VPWR VPWR net208 sky130_fd_sc_hd__dlygate4sd3_1
Xhold34 ih.t.count\[24\] VGND VGND VPWR VPWR net230 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3449__A1 _0359_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4219__A _1286_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2962__A _2697_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5610__A2 _1648_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3621__A1 cu.reg_file.reg_sp\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3621__B2 cu.reg_file.reg_h\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_19_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4889__A cu.pc.pc_o\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_9 clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5126__A1 _1050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3017__B ih.t.timer_max\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_319 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_308 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5062__A0 cu.reg_file.reg_c\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5601__A2 _1633_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3612__A1 cu.reg_file.reg_h\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1091 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1080 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5670_ net75 _1648_ _2137_ _2274_ VGND VGND VPWR VPWR _2483_ sky130_fd_sc_hd__a31o_1
XANTENNA__3612__B2 cu.reg_file.reg_a\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4621_ _1647_ _1663_ _2706_ VGND VGND VPWR VPWR mc.rw.next_state\[1\] sky130_fd_sc_hd__a21o_1
XFILLER_0_96_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5394__S _2237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4552_ _1382_ _1602_ _1603_ _1605_ VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__a31o_2
XFILLER_0_40_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4483_ _1296_ _1538_ _1539_ VGND VGND VPWR VPWR _1540_ sky130_fd_sc_hd__a21o_1
X_3503_ cu.reg_file.reg_sp\[2\] _0413_ _0415_ cu.reg_file.reg_d\[2\] _0578_ VGND VGND
+ VPWR VPWR _0579_ sky130_fd_sc_hd__a221o_1
XANTENNA__5117__A1 _1260_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6222_ clknet_leaf_11_clk ih.t.next_count\[10\] net176 VGND VGND VPWR VPWR ih.t.count\[10\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_12_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3434_ _0447_ net142 VGND VGND VPWR VPWR _0510_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_40_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6153_ clknet_leaf_8_clk _0187_ net169 VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__dfrtp_4
XTAP_853 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3365_ cu.reg_file.reg_l\[0\] _0422_ _0431_ _0434_ _0440_ VGND VGND VPWR VPWR _0441_
+ sky130_fd_sc_hd__a2111o_2
X_6084_ clknet_leaf_21_clk _0118_ net189 VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__dfrtp_1
XTAP_886 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_875 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5104_ _2057_ VGND VGND VPWR VPWR _0064_ sky130_fd_sc_hd__clkbuf_1
X_3296_ cu.id.cb_opcode_x\[1\] VGND VGND VPWR VPWR _0372_ sky130_fd_sc_hd__inv_2
XTAP_897 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5035_ cu.reg_file.reg_b\[2\] _2010_ _2006_ VGND VGND VPWR VPWR _2011_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout183_A net196 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5937_ _2677_ VGND VGND VPWR VPWR _0277_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3603__A1 cu.reg_file.reg_sp\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3603__B2 cu.reg_file.reg_d\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5868_ _2640_ VGND VGND VPWR VPWR _0245_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5356__A1 net112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4819_ _0343_ _1299_ _1818_ VGND VGND VPWR VPWR _1820_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5799_ cu.reg_file.reg_sp\[8\] _2535_ VGND VGND VPWR VPWR _2583_ sky130_fd_sc_hd__or2_1
XFILLER_0_35_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5659__A2 _2204_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput35 net35 VGND VGND VPWR VPWR memory_address_out[0] sky130_fd_sc_hd__clkbuf_4
Xoutput46 net46 VGND VGND VPWR VPWR memory_address_out[5] sky130_fd_sc_hd__clkbuf_4
Xoutput57 net57 VGND VGND VPWR VPWR memory_data_out[6] sky130_fd_sc_hd__buf_2
Xoutput68 net68 VGND VGND VPWR VPWR programmable_gpio_wr[0] sky130_fd_sc_hd__clkbuf_4
Xoutput79 net79 VGND VGND VPWR VPWR ss0[3] sky130_fd_sc_hd__clkbuf_4
XANTENNA__4619__A0 _1650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4891__B cu.pc.pc_o\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_2_clk_A clknet_2_0__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5044__A0 cu.reg_file.reg_b\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4555__C1 _1489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5942__S _2666_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5504__D1 _1417_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4858__A0 _1160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4248__B_N _1311_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3150_ _2883_ _2884_ _2885_ _2886_ VGND VGND VPWR VPWR _2887_ sky130_fd_sc_hd__and4_2
X_3081_ ih.t.count\[11\] _2753_ _2817_ VGND VGND VPWR VPWR _2819_ sky130_fd_sc_hd__and3_1
XANTENNA__5283__A0 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5035__A0 cu.reg_file.reg_b\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5586__A1 _1666_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5722_ _2869_ _2870_ _2873_ net204 VGND VGND VPWR VPWR _0218_ sky130_fd_sc_hd__a22o_1
X_3983_ cu.alu_f\[1\] _1023_ _1056_ _1057_ _1027_ VGND VGND VPWR VPWR _1058_ sky130_fd_sc_hd__o221a_1
XANTENNA__3597__A0 _0374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5653_ _2463_ _2464_ _2466_ _1641_ VGND VGND VPWR VPWR _2467_ sky130_fd_sc_hd__o22a_4
XFILLER_0_45_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5584_ _1400_ _2400_ VGND VGND VPWR VPWR _2401_ sky130_fd_sc_hd__and2b_1
XFILLER_0_72_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4604_ _1485_ VGND VGND VPWR VPWR _1648_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4535_ cu.reg_file.reg_sp\[14\] _1286_ VGND VGND VPWR VPWR _1589_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4466_ cu.id.imm_i\[10\] _1294_ _1297_ _1521_ _1489_ VGND VGND VPWR VPWR _1524_ sky130_fd_sc_hd__a221o_1
XFILLER_0_13_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4397_ _2701_ _1441_ _1353_ VGND VGND VPWR VPWR _1459_ sky130_fd_sc_hd__a21o_1
XFILLER_0_68_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5510__A1 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6205_ clknet_leaf_6_clk net3 net166 VGND VGND VPWR VPWR ih.ih.ih.prev_data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3417_ _0458_ _0486_ VGND VGND VPWR VPWR _0493_ sky130_fd_sc_hd__nor2_1
XANTENNA__4695__C _1672_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6136_ clknet_leaf_6_clk _0170_ net165 VGND VGND VPWR VPWR net128 sky130_fd_sc_hd__dfrtp_4
XTAP_661 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3348_ _0408_ _0407_ _0293_ VGND VGND VPWR VPWR _0424_ sky130_fd_sc_hd__a21o_1
XTAP_650 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_672 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6067_ clknet_leaf_16_clk _0101_ net181 VGND VGND VPWR VPWR ih.gpio_interrupt_mask\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_3279_ _0340_ _0341_ _0343_ VGND VGND VPWR VPWR _0355_ sky130_fd_sc_hd__a21bo_1
XANTENNA__5299__S _2182_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5018_ cu.reg_file.reg_a\[6\] _1997_ _1985_ VGND VGND VPWR VPWR _1998_ sky130_fd_sc_hd__mux2_1
XFILLER_0_95_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5577__A1 net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_469 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4304__A2 _1354_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3815__A1 cu.reg_file.reg_a\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output115_A net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5017__A0 _1193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3815__B2 cu.reg_file.reg_mem\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5002__S _0368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4240__A1 _0359_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5740__A1 _1050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4320_ cu.reg_file.reg_e\[3\] _1283_ _1285_ cu.reg_file.reg_l\[3\] _1384_ VGND VGND
+ VPWR VPWR _1385_ sky130_fd_sc_hd__a221o_1
XFILLER_0_59_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4251_ _1318_ VGND VGND VPWR VPWR _1319_ sky130_fd_sc_hd__inv_2
X_3202_ _2899_ cu.id.opcode\[1\] _2875_ _2876_ VGND VGND VPWR VPWR _2939_ sky130_fd_sc_hd__or4bb_4
XANTENNA__3503__B1 _0415_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3205__B _2936_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4182_ _1248_ _1251_ _0588_ VGND VGND VPWR VPWR _1252_ sky130_fd_sc_hd__mux2_1
X_3133_ _2870_ VGND VGND VPWR VPWR _2871_ sky130_fd_sc_hd__inv_2
XFILLER_0_89_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3064_ _2757_ _2801_ ih.t.count\[17\] VGND VGND VPWR VPWR _2802_ sky130_fd_sc_hd__a21oi_1
XANTENNA__3806__A1 cu.id.imm_i\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5008__A0 _1187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5559__B2 _1401_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3966_ _0447_ _0588_ VGND VGND VPWR VPWR _1041_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5705_ net7 _1650_ _2488_ _2510_ VGND VGND VPWR VPWR _0212_ sky130_fd_sc_hd__a31o_1
XANTENNA__4782__A2 _2948_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5636_ net130 _2236_ _2247_ net138 VGND VGND VPWR VPWR _2450_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3897_ _2885_ _2886_ VGND VGND VPWR VPWR _0973_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5567_ mc.cl.next_data\[2\] _2359_ _2324_ _2384_ VGND VGND VPWR VPWR _2385_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_41_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5498_ ih.t.timer_max\[0\] _2314_ _2317_ _1400_ VGND VGND VPWR VPWR _2318_ sky130_fd_sc_hd__o2bb2a_1
X_4518_ cu.id.imm_i\[13\] _1294_ _1297_ cu.pc.pc_o\[13\] _1488_ VGND VGND VPWR VPWR
+ _1573_ sky130_fd_sc_hd__a221o_1
X_4449_ cu.reg_file.reg_sp\[9\] _0993_ _1344_ cu.id.imm_i\[9\] _1324_ VGND VGND VPWR
+ VPWR _1508_ sky130_fd_sc_hd__a221o_1
X_6119_ clknet_leaf_7_clk _0153_ net167 VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__dfrtp_2
XTAP_480 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4470__A1 _1521_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4470__B2 cu.reg_file.reg_d\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2970__A net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4222__A1 cu.reg_file.reg_c\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5722__A1 _2869_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5486__A0 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3976__A _1050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3820_ _0892_ _0895_ VGND VGND VPWR VPWR _0896_ sky130_fd_sc_hd__or2b_1
X_3751_ cu.pc.pc_o\[15\] _0740_ _0825_ _0826_ VGND VGND VPWR VPWR _0827_ sky130_fd_sc_hd__a211o_1
XFILLER_0_54_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3682_ _0511_ _0712_ VGND VGND VPWR VPWR _0758_ sky130_fd_sc_hd__nor2_1
X_5421_ _1329_ _1372_ _1369_ VGND VGND VPWR VPWR _2257_ sky130_fd_sc_hd__and3_1
XANTENNA__4516__A2 _1282_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4600__A _1632_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5352_ _1075_ net110 _2215_ VGND VGND VPWR VPWR _2218_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4303_ _1368_ VGND VGND VPWR VPWR _1369_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5283_ net82 _1193_ _2170_ VGND VGND VPWR VPWR _2177_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4234_ _1300_ _1301_ VGND VGND VPWR VPWR _1302_ sky130_fd_sc_hd__and2b_1
XFILLER_0_4_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4165_ _0387_ _1234_ _0824_ VGND VGND VPWR VPWR _1235_ sky130_fd_sc_hd__a21oi_1
X_3116_ _2810_ _2811_ _2853_ VGND VGND VPWR VPWR _2854_ sky130_fd_sc_hd__or3_1
XANTENNA__5431__A _2139_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4096_ _0546_ _0733_ VGND VGND VPWR VPWR _1170_ sky130_fd_sc_hd__xor2_1
X_3047_ ih.t.timer_max\[22\] _2760_ ih.t.timer_max\[23\] VGND VGND VPWR VPWR _2785_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA_clkbuf_leaf_42_clk_A clknet_2_0__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4998_ _2951_ _0367_ _0352_ VGND VGND VPWR VPWR _1984_ sky130_fd_sc_hd__and3_1
X_3949_ _1023_ _1024_ alu.Cin _1021_ VGND VGND VPWR VPWR _1025_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_60_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4507__A2 _1545_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5619_ net105 _2205_ _2433_ _1401_ VGND VGND VPWR VPWR _2434_ sky130_fd_sc_hd__a22o_1
XANTENNA__5704__B2 _1646_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5640__B1 _2225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6063__RESET_B net195 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5950__S _2666_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3485__A2 _0502_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_509 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4434__A1 cu.pc.pc_o\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4434__B2 cu.reg_file.reg_d\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5970_ clknet_leaf_35_clk _0007_ net159 VGND VGND VPWR VPWR alu.Cin sky130_fd_sc_hd__dfrtp_4
XFILLER_0_87_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4921_ _1912_ _1913_ _1798_ VGND VGND VPWR VPWR _1914_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4852_ cu.pc.pc_o\[4\] _1838_ VGND VGND VPWR VPWR _1850_ sky130_fd_sc_hd__xor2_1
XFILLER_0_47_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3803_ cu.reg_file.reg_b\[2\] _0743_ _0624_ cu.reg_file.reg_sp\[10\] VGND VGND VPWR
+ VPWR _0879_ sky130_fd_sc_hd__a22o_1
XFILLER_0_55_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5934__A1 _2486_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_536 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4783_ _0986_ _0989_ _0994_ VGND VGND VPWR VPWR _1786_ sky130_fd_sc_hd__and3_1
XFILLER_0_7_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3734_ _0763_ _0809_ VGND VGND VPWR VPWR _0810_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_70_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3665_ _0464_ _0482_ VGND VGND VPWR VPWR _0741_ sky130_fd_sc_hd__and2_2
X_5404_ _2181_ _2247_ VGND VGND VPWR VPWR _2248_ sky130_fd_sc_hd__nand2_8
XFILLER_0_2_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3596_ ih.interrupt_source\[3\] ih.interrupt_source\[2\] VGND VGND VPWR VPWR _0672_
+ sky130_fd_sc_hd__or2_1
XFILLER_0_30_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5335_ _1075_ net102 _2206_ VGND VGND VPWR VPWR _2209_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5266_ _1110_ _1263_ _1666_ VGND VGND VPWR VPWR _2167_ sky130_fd_sc_hd__mux2_1
XFILLER_0_55_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4217_ _1284_ VGND VGND VPWR VPWR _1285_ sky130_fd_sc_hd__buf_2
X_5197_ mc.cc.count\[0\] _2708_ VGND VGND VPWR VPWR _2118_ sky130_fd_sc_hd__or2_1
X_4148_ _0939_ _0940_ VGND VGND VPWR VPWR _1218_ sky130_fd_sc_hd__or2_1
XFILLER_0_78_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4079_ _1060_ _0600_ VGND VGND VPWR VPWR _1153_ sky130_fd_sc_hd__nand2_1
XANTENNA__5622__B1 _2204_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4189__A0 _1194_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_199 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5684__A2_N _1643_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_214 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5916__A1 _1484_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3450_ _2925_ _2901_ _2912_ _2897_ _2935_ VGND VGND VPWR VPWR _0526_ sky130_fd_sc_hd__o221a_1
X_3381_ cu.id.starting_int_service _0382_ _0456_ _2896_ VGND VGND VPWR VPWR _0457_
+ sky130_fd_sc_hd__or4b_2
XFILLER_0_20_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5120_ _2065_ VGND VGND VPWR VPWR _2066_ sky130_fd_sc_hd__buf_4
X_5051_ _2021_ VGND VGND VPWR VPWR _0047_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4002_ _0761_ _0764_ _0772_ VGND VGND VPWR VPWR _1076_ sky130_fd_sc_hd__and3b_1
XFILLER_0_46_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4407__A1 cu.id.cb_opcode_x\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4407__B2 cu.pc.pc_o\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5953_ _2685_ VGND VGND VPWR VPWR _2686_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5080__A1 _1623_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5884_ _1187_ ih.t.timer_max\[3\] _2645_ VGND VGND VPWR VPWR _2649_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4904_ _2920_ cu.pc.pc_o\[8\] VGND VGND VPWR VPWR _1898_ sky130_fd_sc_hd__nor2_1
XANTENNA__3630__A2 _0498_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5907__A1 _1193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4835_ _1833_ _1834_ _1799_ VGND VGND VPWR VPWR _1835_ sky130_fd_sc_hd__mux2_1
XFILLER_0_28_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4766_ _1303_ _1772_ _1773_ _1765_ VGND VGND VPWR VPWR _1774_ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_355 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3717_ _0652_ _0663_ VGND VGND VPWR VPWR _0793_ sky130_fd_sc_hd__and2b_1
XFILLER_0_43_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4697_ ih.t.count\[21\] _1714_ VGND VGND VPWR VPWR _1717_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3648_ cu.reg_file.reg_d\[7\] _0415_ _0432_ cu.reg_file.reg_b\[7\] VGND VGND VPWR
+ VPWR _0724_ sky130_fd_sc_hd__a22o_1
X_3579_ cu.id.cb_opcode_y\[2\] _0654_ _0294_ VGND VGND VPWR VPWR _0655_ sky130_fd_sc_hd__mux2_1
X_5318_ _1188_ net95 _2195_ VGND VGND VPWR VPWR _2199_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6298_ clknet_leaf_41_clk _0280_ net152 VGND VGND VPWR VPWR cu.id.cb_opcode_y\[0\]
+ sky130_fd_sc_hd__dfrtp_4
Xhold13 cu.alu_f\[4\] VGND VGND VPWR VPWR net209 sky130_fd_sc_hd__dlygate4sd3_1
Xhold35 ih.t.count\[18\] VGND VGND VPWR VPWR net231 sky130_fd_sc_hd__dlygate4sd3_1
Xhold24 mc.cc.count\[3\] VGND VGND VPWR VPWR net220 sky130_fd_sc_hd__dlygate4sd3_1
X_5249_ ih.t.timer_max\[25\] _2155_ _2153_ VGND VGND VPWR VPWR _2156_ sky130_fd_sc_hd__mux2_1
XANTENNA__4934__S _1798_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2962__B _2702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3621__A2 _0413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_309 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5005__S _0368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4098__C1 _0918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5062__A1 _1187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3612__A2 _0495_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1092 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1081 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1070 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_8_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4620_ _1651_ _1662_ _2699_ VGND VGND VPWR VPWR _1663_ sky130_fd_sc_hd__a21o_1
XFILLER_0_72_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4573__B1 _1623_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4551_ _1402_ _1598_ _1604_ _1371_ VGND VGND VPWR VPWR _1605_ sky130_fd_sc_hd__a2bb2o_1
X_4482_ cu.id.imm_i\[11\] _1294_ _1297_ cu.pc.pc_o\[11\] _1489_ VGND VGND VPWR VPWR
+ _1539_ sky130_fd_sc_hd__a221o_1
X_3502_ cu.reg_file.reg_b\[2\] _0432_ _0433_ cu.reg_file.reg_a\[2\] VGND VGND VPWR
+ VPWR _0578_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6221_ clknet_leaf_11_clk ih.t.next_count\[9\] net176 VGND VGND VPWR VPWR ih.t.count\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_158 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3433_ _0491_ _0497_ _0506_ _0508_ VGND VGND VPWR VPWR _0509_ sky130_fd_sc_hd__o31ai_2
X_6152_ clknet_leaf_9_clk _0186_ net174 VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__dfrtp_4
XTAP_810 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5103_ cu.reg_file.reg_e\[0\] _2022_ _2056_ VGND VGND VPWR VPWR _2057_ sky130_fd_sc_hd__mux2_1
X_3364_ _0293_ _0362_ _0438_ _0439_ VGND VGND VPWR VPWR _0440_ sky130_fd_sc_hd__or4_4
X_6083_ clknet_leaf_21_clk _0117_ net189 VGND VGND VPWR VPWR ih.t.timer_max\[31\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_876 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_865 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3295_ _2950_ _0361_ VGND VGND VPWR VPWR _0371_ sky130_fd_sc_hd__nand2_2
XANTENNA__3224__A _0298_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_898 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_887 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5034_ _1074_ _1226_ _2002_ VGND VGND VPWR VPWR _2010_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5936_ _0343_ _2350_ _2666_ VGND VGND VPWR VPWR _2677_ sky130_fd_sc_hd__mux2_1
X_5867_ _2159_ ih.t.timer_max\[11\] _2636_ VGND VGND VPWR VPWR _2640_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4818_ _0343_ _1299_ _1818_ VGND VGND VPWR VPWR _1819_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5798_ _2582_ VGND VGND VPWR VPWR _0233_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_196 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4749_ _1739_ _1757_ _1483_ VGND VGND VPWR VPWR _1758_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput36 net36 VGND VGND VPWR VPWR memory_address_out[10] sky130_fd_sc_hd__clkbuf_4
Xoutput58 net58 VGND VGND VPWR VPWR memory_data_out[7] sky130_fd_sc_hd__clkbuf_4
Xoutput47 net47 VGND VGND VPWR VPWR memory_address_out[6] sky130_fd_sc_hd__clkbuf_4
Xoutput69 net69 VGND VGND VPWR VPWR programmable_gpio_wr[1] sky130_fd_sc_hd__clkbuf_4
XANTENNA__3134__A _2745_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2973__A net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3358__A1 cu.reg_file.reg_b\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3358__B2 cu.reg_file.reg_a\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_78_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3309__A _0359_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5504__C1 _1489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5524__A _1666_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3080_ _2753_ _2817_ ih.t.count\[11\] VGND VGND VPWR VPWR _2818_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5283__A1 _1193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3982_ _0298_ _1001_ _1002_ VGND VGND VPWR VPWR _1057_ sky130_fd_sc_hd__o21ai_1
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4794__A0 _0617_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5721_ net1 net197 _2872_ _2870_ _2521_ VGND VGND VPWR VPWR _0217_ sky130_fd_sc_hd__a2111oi_1
XANTENNA__4603__A _1646_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5652_ _1649_ _2465_ VGND VGND VPWR VPWR _2466_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5583_ ih.t.timer_max\[11\] _2193_ _2314_ ih.t.timer_max\[3\] _2399_ VGND VGND VPWR
+ VPWR _2400_ sky130_fd_sc_hd__a221o_1
X_4603_ _1646_ VGND VGND VPWR VPWR _1647_ sky130_fd_sc_hd__buf_2
XFILLER_0_72_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4534_ _1580_ _1582_ VGND VGND VPWR VPWR _1588_ sky130_fd_sc_hd__nand2_1
XFILLER_0_13_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5434__A _2139_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4465_ cu.reg_file.reg_b\[2\] net143 _1284_ cu.reg_file.reg_h\[2\] _1522_ VGND VGND
+ VPWR VPWR _1523_ sky130_fd_sc_hd__a221o_1
XFILLER_0_7_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4396_ _1419_ _1436_ _1456_ _1445_ VGND VGND VPWR VPWR _1458_ sky130_fd_sc_hd__nand4_1
XANTENNA__5510__A2 _1648_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6204_ clknet_leaf_5_clk net17 net171 VGND VGND VPWR VPWR ih.ih.ih.prev_data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
X_3416_ net146 _0473_ net145 _0463_ _0458_ VGND VGND VPWR VPWR _0492_ sky130_fd_sc_hd__o2111a_4
X_6135_ clknet_leaf_6_clk _0169_ net164 VGND VGND VPWR VPWR net127 sky130_fd_sc_hd__dfrtp_4
XANTENNA__3521__A1 _0293_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3347_ _0417_ VGND VGND VPWR VPWR _0423_ sky130_fd_sc_hd__inv_2
XTAP_640 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6066_ clknet_leaf_25_clk _0100_ net195 VGND VGND VPWR VPWR mc.cc.count\[3\] sky130_fd_sc_hd__dfrtp_1
XTAP_695 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3278_ _2883_ _2936_ VGND VGND VPWR VPWR _0354_ sky130_fd_sc_hd__or2_1
X_5017_ _1193_ _1624_ _0368_ VGND VGND VPWR VPWR _1997_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4482__C1 _1489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5577__A2 _2194_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5919_ cu.ir.idx\[0\] cu.ir.idx\[1\] VGND VGND VPWR VPWR _2668_ sky130_fd_sc_hd__nor2_4
XFILLER_0_90_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_63_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3760__A1 cu.pc.pc_o\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5017__A1 _1624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output108_A net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_81_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3751__A1 cu.pc.pc_o\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4250_ _2893_ _2901_ _2923_ _2936_ VGND VGND VPWR VPWR _1318_ sky130_fd_sc_hd__or4b_2
XANTENNA__4700__B1 _1670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3201_ cu.id.alu_opcode\[0\] _2894_ VGND VGND VPWR VPWR _2938_ sky130_fd_sc_hd__or2b_1
X_4181_ _1249_ _1250_ _0599_ VGND VGND VPWR VPWR _1251_ sky130_fd_sc_hd__mux2_1
XANTENNA__3503__A1 cu.reg_file.reg_sp\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3503__B2 cu.reg_file.reg_d\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3132_ ih.ih.int_f.prev_data ih.ih.int_f.data_in ih.input_handler_enable VGND VGND
+ VPWR VPWR _2870_ sky130_fd_sc_hd__and3b_4
X_3063_ ih.t.timer_max\[16\] _2756_ ih.t.timer_max\[17\] VGND VGND VPWR VPWR _2801_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_89_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5008__A1 _1222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5559__A2 _2205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3824__A2_N _0895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3965_ _0710_ VGND VGND VPWR VPWR _1040_ sky130_fd_sc_hd__inv_2
XFILLER_0_45_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5704_ _2509_ _1643_ cu.reg_file.reg_mem\[14\] _1646_ VGND VGND VPWR VPWR _2510_
+ sky130_fd_sc_hd__a2bb2o_1
X_3896_ _2935_ _0971_ VGND VGND VPWR VPWR _0972_ sky130_fd_sc_hd__nand2_1
XFILLER_0_45_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5635_ _2449_ VGND VGND VPWR VPWR _0203_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5566_ _1666_ _2382_ _2383_ VGND VGND VPWR VPWR _2384_ sky130_fd_sc_hd__o21a_1
XFILLER_0_79_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_clkbuf_2_1__f_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5497_ _2315_ _2316_ VGND VGND VPWR VPWR _2317_ sky130_fd_sc_hd__nor2_1
X_4517_ cu.reg_file.reg_b\[5\] net143 _1284_ cu.reg_file.reg_h\[5\] _1571_ VGND VGND
+ VPWR VPWR _1572_ sky130_fd_sc_hd__a221o_1
XANTENNA_clkbuf_leaf_1_clk_A clknet_2_0__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4448_ cu.reg_file.reg_h\[1\] _1316_ VGND VGND VPWR VPWR _1507_ sky130_fd_sc_hd__and2_1
XFILLER_0_13_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5495__B2 ih.t.timer_max\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4379_ _1404_ _1417_ _1434_ VGND VGND VPWR VPWR _1442_ sky130_fd_sc_hd__a21bo_1
X_6118_ clknet_leaf_7_clk _0152_ net167 VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__dfrtp_4
XTAP_470 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6049_ clknet_leaf_3_clk _0087_ net157 VGND VGND VPWR VPWR cu.reg_file.reg_l\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_95_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4470__A2 _1321_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3430__B1 _0499_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3981__B2 cu.alu_f\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5722__A2 _2870_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5486__A1 _0618_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4997__A0 _0618_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5948__S _2666_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3750_ cu.reg_file.reg_b\[7\] _0743_ _0624_ cu.reg_file.reg_sp\[15\] VGND VGND VPWR
+ VPWR _0826_ sky130_fd_sc_hd__a22o_1
X_3681_ _0664_ _0756_ VGND VGND VPWR VPWR _0757_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_27_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5420_ _2256_ VGND VGND VPWR VPWR _0181_ sky130_fd_sc_hd__clkbuf_1
X_5351_ _2217_ VGND VGND VPWR VPWR _0151_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4600__B _1643_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4302_ _1306_ _1362_ _1367_ VGND VGND VPWR VPWR _1368_ sky130_fd_sc_hd__o21ai_2
X_5282_ _2176_ VGND VGND VPWR VPWR _0123_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_50_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4233_ cu.id.state\[1\] VGND VGND VPWR VPWR _1301_ sky130_fd_sc_hd__buf_2
X_4164_ _1233_ _0371_ VGND VGND VPWR VPWR _1234_ sky130_fd_sc_hd__nor2_1
X_3115_ _2813_ _2815_ _2816_ _2852_ VGND VGND VPWR VPWR _2853_ sky130_fd_sc_hd__or4_1
XANTENNA__5431__B _2205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4095_ _0566_ _1110_ VGND VGND VPWR VPWR _1169_ sky130_fd_sc_hd__xnor2_1
X_3046_ _2762_ _2782_ ih.t.count\[24\] VGND VGND VPWR VPWR _2784_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_81_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4997_ _0618_ _1622_ _0368_ VGND VGND VPWR VPWR _1983_ sky130_fd_sc_hd__mux2_1
XFILLER_0_45_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3963__A1 _0918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3948_ _0572_ _1020_ VGND VGND VPWR VPWR _1024_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3879_ _0771_ _0954_ VGND VGND VPWR VPWR _0955_ sky130_fd_sc_hd__or2b_1
XANTENNA__4998__A _2951_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5165__A0 cu.reg_file.reg_l\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5618_ net89 _1330_ VGND VGND VPWR VPWR _2433_ sky130_fd_sc_hd__or2_1
XFILLER_0_5_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4510__B _1530_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4912__A0 cu.pc.pc_o\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5549_ net69 _1649_ _2137_ _2274_ VGND VGND VPWR VPWR _2368_ sky130_fd_sc_hd__a31o_1
XFILLER_0_41_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5640__A1 net114 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5640__B2 net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4903__A0 _1622_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3317__A _0384_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5008__S _0368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5631__A1 net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4434__A2 _1321_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4920_ _1623_ _1909_ _1794_ VGND VGND VPWR VPWR _1913_ sky130_fd_sc_hd__mux2_1
XANTENNA__5631__B2 net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4851_ _1849_ VGND VGND VPWR VPWR _0019_ sky130_fd_sc_hd__clkbuf_1
X_3802_ cu.reg_file.reg_d\[2\] _0488_ _0741_ cu.reg_file.reg_h\[2\] VGND VGND VPWR
+ VPWR _0878_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_548 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4782_ _0350_ _2948_ _1782_ net201 VGND VGND VPWR VPWR _0002_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3733_ _0759_ _0783_ _0784_ VGND VGND VPWR VPWR _0809_ sky130_fd_sc_hd__a21oi_1
X_3664_ _0501_ VGND VGND VPWR VPWR _0740_ sky130_fd_sc_hd__buf_4
X_5403_ _2246_ VGND VGND VPWR VPWR _2247_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_2_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3595_ _0576_ _0665_ _0667_ _0670_ VGND VGND VPWR VPWR _0671_ sky130_fd_sc_hd__o2bb2a_1
X_5334_ _2208_ VGND VGND VPWR VPWR _0143_ sky130_fd_sc_hd__clkbuf_1
X_5265_ _2166_ VGND VGND VPWR VPWR _0116_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5196_ _2117_ VGND VGND VPWR VPWR _0096_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4122__B2 _1192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4216_ _1279_ _1275_ VGND VGND VPWR VPWR _1284_ sky130_fd_sc_hd__nor2_2
X_4147_ _0951_ _1216_ VGND VGND VPWR VPWR _1217_ sky130_fd_sc_hd__nor2_1
X_4078_ _0558_ _0663_ _0822_ _0694_ VGND VGND VPWR VPWR _1152_ sky130_fd_sc_hd__a22o_1
X_3029_ ih.t.count\[31\] _2766_ VGND VGND VPWR VPWR _2767_ sky130_fd_sc_hd__xnor2_1
XANTENNA__5386__A0 _0619_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5138__A0 _1209_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5689__A1 net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4361__A1 _1415_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2976__A net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5861__A1 ih.t.timer_max\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3321__C1 _0387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_429 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5377__A0 _1192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_226 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5916__A2 _2351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5129__A0 _1226_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3380_ _0300_ _2911_ _0455_ VGND VGND VPWR VPWR _0456_ sky130_fd_sc_hd__o21ai_1
XANTENNA__5301__A0 _1192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5050_ cu.reg_file.reg_b\[7\] _2020_ _2006_ VGND VGND VPWR VPWR _2021_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_41_clk_A clknet_2_0__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4104__A1 _0547_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4001_ _1074_ VGND VGND VPWR VPWR _1075_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_79_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4606__A _1649_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5952_ _2663_ cu.ir.idx\[1\] VGND VGND VPWR VPWR _2685_ sky130_fd_sc_hd__and2_1
X_4903_ _1622_ _1896_ _1795_ VGND VGND VPWR VPWR _1897_ sky130_fd_sc_hd__mux2_1
XANTENNA__3615__B1 _0492_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5883_ _2648_ VGND VGND VPWR VPWR _0252_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_546 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4834_ _1073_ _1828_ _1795_ VGND VGND VPWR VPWR _1834_ sky130_fd_sc_hd__mux2_1
X_4765_ _1747_ _1763_ _1761_ VGND VGND VPWR VPWR _1773_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_28_484 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5437__A _2139_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3716_ _0733_ _0790_ _0729_ _0791_ VGND VGND VPWR VPWR _0792_ sky130_fd_sc_hd__o2bb2a_1
X_4696_ _1716_ VGND VGND VPWR VPWR ih.t.next_count\[20\] sky130_fd_sc_hd__clkbuf_1
X_3647_ _0293_ _0372_ _0634_ VGND VGND VPWR VPWR _0723_ sky130_fd_sc_hd__or3_1
XFILLER_0_11_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3578_ ih.interrupt_source\[3\] ih.interrupt_source\[1\] VGND VGND VPWR VPWR _0654_
+ sky130_fd_sc_hd__or2_1
X_5317_ _2198_ VGND VGND VPWR VPWR _0136_ sky130_fd_sc_hd__clkbuf_1
Xhold14 mc.cc.count\[0\] VGND VGND VPWR VPWR net210 sky130_fd_sc_hd__dlygate4sd3_1
X_6297_ clknet_leaf_42_clk _0279_ net152 VGND VGND VPWR VPWR cu.id.cb_opcode_z\[2\]
+ sky130_fd_sc_hd__dfrtp_1
Xhold25 _0099_ VGND VGND VPWR VPWR net221 sky130_fd_sc_hd__dlygate4sd3_1
Xhold36 ih.t.count\[27\] VGND VGND VPWR VPWR net232 sky130_fd_sc_hd__dlygate4sd3_1
X_5248_ _1050_ _1623_ _1667_ VGND VGND VPWR VPWR _2155_ sky130_fd_sc_hd__mux2_1
X_5179_ mc.cl.next_data\[12\] net22 mc.count VGND VGND VPWR VPWR _2105_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5347__A _2147_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_487 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output138_A net138 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5956__S _2686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4145__B _0779_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1082 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1071 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1060 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_365 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1093 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_89 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4573__A1 _2702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4161__A _0516_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_281 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4550_ _1585_ _1598_ VGND VGND VPWR VPWR _1604_ sky130_fd_sc_hd__xor2_1
XANTENNA__4573__B2 _2697_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4481_ cu.reg_file.reg_b\[3\] net143 _1284_ cu.reg_file.reg_h\[3\] _1537_ VGND VGND
+ VPWR VPWR _1538_ sky130_fd_sc_hd__a221o_1
XFILLER_0_25_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3501_ cu.reg_file.reg_c\[2\] _0427_ _0430_ cu.reg_file.reg_e\[2\] VGND VGND VPWR
+ VPWR _0577_ sky130_fd_sc_hd__a22o_1
X_6220_ clknet_leaf_11_clk ih.t.next_count\[8\] net176 VGND VGND VPWR VPWR ih.t.count\[8\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3432_ _0343_ _2949_ _0507_ VGND VGND VPWR VPWR _0508_ sky130_fd_sc_hd__a21o_1
XANTENNA__4325__A1 cu.reg_file.reg_sp\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4325__B2 cu.id.cb_opcode_y\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6151_ clknet_leaf_8_clk _0185_ net168 VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__dfrtp_4
XTAP_800 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3363_ net150 _2914_ _0318_ VGND VGND VPWR VPWR _0439_ sky130_fd_sc_hd__or3_1
XTAP_844 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5102_ _2035_ _2055_ _2951_ VGND VGND VPWR VPWR _2056_ sky130_fd_sc_hd__o21a_4
X_6082_ clknet_leaf_22_clk _0116_ net191 VGND VGND VPWR VPWR ih.t.timer_max\[30\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_877 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_866 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3294_ _0369_ VGND VGND VPWR VPWR _0370_ sky130_fd_sc_hd__buf_2
XTAP_899 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_888 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5033_ _2009_ VGND VGND VPWR VPWR _0041_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout169_A net182 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4336__A _1348_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3240__A _0308_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5935_ _2676_ VGND VGND VPWR VPWR _0276_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5866_ _2639_ VGND VGND VPWR VPWR _0244_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4817_ _0340_ cu.pc.pc_o\[1\] VGND VGND VPWR VPWR _1818_ sky130_fd_sc_hd__xor2_1
XFILLER_0_16_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5797_ cu.reg_file.reg_sp\[7\] _2581_ _2539_ VGND VGND VPWR VPWR _2582_ sky130_fd_sc_hd__mux2_1
X_4748_ _0371_ _1756_ VGND VGND VPWR VPWR _1757_ sky130_fd_sc_hd__nand2_1
X_4679_ ih.t.count\[15\] _1702_ VGND VGND VPWR VPWR _1705_ sky130_fd_sc_hd__and2_1
Xoutput37 net37 VGND VGND VPWR VPWR memory_address_out[11] sky130_fd_sc_hd__buf_2
Xoutput48 net48 VGND VGND VPWR VPWR memory_address_out[7] sky130_fd_sc_hd__buf_2
Xoutput59 net59 VGND VGND VPWR VPWR memory_wr sky130_fd_sc_hd__buf_2
XANTENNA__4945__S _1798_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3625__A1_N _0576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3000__A_N net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4246__A _1309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3150__A _2883_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4555__B2 cu.pc.pc_o\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3309__B _2893_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3818__B1 _0429_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4156__A _0516_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3981_ _1023_ _1054_ _1055_ cu.alu_f\[1\] VGND VGND VPWR VPWR _1056_ sky130_fd_sc_hd__o2bb2a_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5720_ net1 ih.interrupt_source\[3\] VGND VGND VPWR VPWR _2521_ sky130_fd_sc_hd__nor2_1
XFILLER_0_72_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_42_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_42_clk sky130_fd_sc_hd__clkbuf_16
X_5651_ net14 _2345_ _2369_ net7 VGND VGND VPWR VPWR _2465_ sky130_fd_sc_hd__a22o_1
XFILLER_0_17_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5582_ ih.t.timer_max\[27\] _2146_ _2204_ ih.t.timer_max\[19\] VGND VGND VPWR VPWR
+ _2399_ sky130_fd_sc_hd__a22o_1
X_4602_ _1645_ VGND VGND VPWR VPWR _1646_ sky130_fd_sc_hd__clkbuf_4
X_4533_ _1353_ _1579_ _1583_ _1584_ _1587_ VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__a221o_1
XFILLER_0_25_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5434__B _2147_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6203_ clknet_leaf_4_clk net16 net171 VGND VGND VPWR VPWR ih.ih.ih.prev_data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_4464_ cu.reg_file.reg_d\[2\] _1282_ _1286_ cu.reg_file.reg_sp\[10\] VGND VGND VPWR
+ VPWR _1522_ sky130_fd_sc_hd__a22o_1
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4395_ _1419_ _1436_ _1445_ _1456_ VGND VGND VPWR VPWR _1457_ sky130_fd_sc_hd__a31o_1
XFILLER_0_0_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3415_ cu.reg_file.reg_c\[0\] _0485_ _0489_ cu.reg_file.reg_e\[0\] _0490_ VGND VGND
+ VPWR VPWR _0491_ sky130_fd_sc_hd__a221o_1
X_6134_ clknet_leaf_6_clk _0168_ net165 VGND VGND VPWR VPWR net126 sky130_fd_sc_hd__dfrtp_2
XFILLER_0_0_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3346_ _0414_ _0421_ _0417_ VGND VGND VPWR VPWR _0422_ sky130_fd_sc_hd__a21oi_4
XTAP_630 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6065_ clknet_leaf_25_clk net221 net192 VGND VGND VPWR VPWR mc.cc.count\[2\] sky130_fd_sc_hd__dfrtp_1
XTAP_685 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_696 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3277_ _2892_ _0324_ VGND VGND VPWR VPWR _0353_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5016_ _1996_ VGND VGND VPWR VPWR _0037_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_67_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5918_ net201 _2667_ _1781_ VGND VGND VPWR VPWR _0268_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_48_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_33_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_33_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_90_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_48_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5849_ _2625_ _2626_ VGND VGND VPWR VPWR _2627_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_63_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4537__B2 cu.reg_file.reg_h\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4537__A1 cu.reg_file.reg_b\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3760__A2 _0740_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2984__A net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_39_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_24_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_24_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_81_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output82_A net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3751__A2 _0740_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3200_ _2936_ _2901_ _2898_ VGND VGND VPWR VPWR _2937_ sky130_fd_sc_hd__or3_2
X_4180_ _0694_ _1040_ _1060_ VGND VGND VPWR VPWR _1250_ sky130_fd_sc_hd__mux2_1
XANTENNA__3503__A2 _0413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3131_ _2768_ _2864_ _2867_ _2868_ VGND VGND VPWR VPWR _2869_ sky130_fd_sc_hd__or4b_4
X_3062_ ih.t.count\[18\] _2758_ _2798_ VGND VGND VPWR VPWR _2800_ sky130_fd_sc_hd__and3_1
XFILLER_0_54_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4464__B1 _1286_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_15_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_15_clk sky130_fd_sc_hd__clkbuf_16
X_3964_ _0570_ _0712_ VGND VGND VPWR VPWR _1039_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5703_ mc.cl.next_data\[14\] _2359_ _2490_ _2508_ VGND VGND VPWR VPWR _2509_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_57_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3895_ _2893_ _2896_ _2912_ _2923_ VGND VGND VPWR VPWR _0971_ sky130_fd_sc_hd__o22a_1
XFILLER_0_45_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4519__A1 _1296_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_357 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5634_ cu.reg_file.reg_mem\[5\] _2448_ _2351_ VGND VGND VPWR VPWR _2449_ sky130_fd_sc_hd__mux2_1
X_5565_ ih.t.timer_max\[18\] _2150_ _2319_ ih.t.timer_max\[2\] _1661_ VGND VGND VPWR
+ VPWR _2383_ sky130_fd_sc_hd__a221o_1
XFILLER_0_79_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5496_ ih.t.timer_max\[24\] _2146_ _2204_ ih.t.timer_max\[16\] VGND VGND VPWR VPWR
+ _2316_ sky130_fd_sc_hd__a22o_1
X_4516_ cu.reg_file.reg_d\[5\] _1282_ _1286_ cu.reg_file.reg_sp\[13\] VGND VGND VPWR
+ VPWR _1571_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4447_ cu.id.imm_i\[9\] _1295_ _1298_ cu.pc.pc_o\[9\] _1305_ VGND VGND VPWR VPWR
+ _1506_ sky130_fd_sc_hd__a221o_1
X_6117_ clknet_leaf_10_clk _0151_ net175 VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__dfrtp_1
X_4378_ _1404_ _1440_ VGND VGND VPWR VPWR _1441_ sky130_fd_sc_hd__nand2_1
XTAP_460 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3329_ _0403_ _0404_ cu.id.starting_int_service VGND VGND VPWR VPWR _0405_ sky130_fd_sc_hd__a21o_2
XTAP_471 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6048_ clknet_leaf_4_clk _0086_ net170 VGND VGND VPWR VPWR cu.reg_file.reg_l\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_95_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3430__A1 alu.Cin VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3430__B2 cu.reg_file.reg_a\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__2979__A net6 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6238__RESET_B net182 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4446__B1 _1296_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output120_A net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4997__A1 _1622_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4137__C _0773_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4749__A1 _1739_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5946__A0 _0373_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3421__A1 cu.reg_file.reg_d\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5964__S _2686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3680_ _0718_ _0755_ _0720_ VGND VGND VPWR VPWR _0756_ sky130_fd_sc_hd__a21oi_1
X_5350_ _1052_ net109 _2215_ VGND VGND VPWR VPWR _2217_ sky130_fd_sc_hd__mux2_1
X_5281_ net81 _1191_ _2170_ VGND VGND VPWR VPWR _2176_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4301_ cu.reg_file.reg_c\[2\] _1313_ _1363_ _1366_ VGND VGND VPWR VPWR _1367_ sky130_fd_sc_hd__a211o_1
XFILLER_0_10_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4232_ cu.id.state\[0\] VGND VGND VPWR VPWR _1300_ sky130_fd_sc_hd__buf_2
Xclkbuf_leaf_4_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_4_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__3488__A1 cu.reg_file.reg_a\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4163_ _2920_ VGND VGND VPWR VPWR _1233_ sky130_fd_sc_hd__buf_4
X_3114_ _2818_ _2819_ _2851_ VGND VGND VPWR VPWR _2852_ sky130_fd_sc_hd__or3_1
X_4094_ _1090_ _1164_ _1166_ _0611_ _1167_ VGND VGND VPWR VPWR _1168_ sky130_fd_sc_hd__o221a_1
X_3045_ ih.t.count\[24\] _2762_ _2782_ VGND VGND VPWR VPWR _2783_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4996_ _1982_ VGND VGND VPWR VPWR _0031_ sky130_fd_sc_hd__clkbuf_1
X_3947_ _1003_ _1011_ _1020_ _1022_ _2948_ VGND VGND VPWR VPWR _1023_ sky130_fd_sc_hd__o41a_2
XFILLER_0_45_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3878_ _0898_ _0953_ VGND VGND VPWR VPWR _0954_ sky130_fd_sc_hd__xnor2_1
X_5617_ net97 _2194_ _2431_ VGND VGND VPWR VPWR _2432_ sky130_fd_sc_hd__a21o_1
XFILLER_0_33_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5165__A1 _1260_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5548_ _2169_ _2358_ _2366_ _2136_ VGND VGND VPWR VPWR _2367_ sky130_fd_sc_hd__o211a_1
XANTENNA__3361__A_N _0308_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4510__C _1545_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5479_ _2301_ VGND VGND VPWR VPWR _0195_ sky130_fd_sc_hd__clkbuf_1
XTAP_290 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5625__C1 _1661_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5640__A2 _2147_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3651__B2 cu.reg_file.reg_a\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4254__A _1321_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5928__A0 _0359_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3333__A cu.id.starting_int_service VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output45_A net45 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5092__A0 _1191_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4850_ cu.pc.pc_o\[3\] _1848_ _1815_ VGND VGND VPWR VPWR _1849_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4164__A _1233_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_0_clk_A clknet_2_0__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3801_ _0875_ _0876_ VGND VGND VPWR VPWR _0877_ sky130_fd_sc_hd__or2_1
X_4781_ net199 _1785_ net201 VGND VGND VPWR VPWR _0003_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_82_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3732_ _0806_ _0807_ VGND VGND VPWR VPWR _0808_ sky130_fd_sc_hd__or2_1
X_3663_ _0738_ VGND VGND VPWR VPWR _0739_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_70_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5402_ _1369_ _2148_ VGND VGND VPWR VPWR _2246_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5333_ _1052_ net101 _2206_ VGND VGND VPWR VPWR _2208_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3594_ cu.reg_file.reg_l\[4\] _0422_ _0668_ _0669_ _0576_ VGND VGND VPWR VPWR _0670_
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_11_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5264_ ih.t.timer_max\[30\] _2165_ _2153_ VGND VGND VPWR VPWR _2166_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4215_ _1282_ VGND VGND VPWR VPWR _1283_ sky130_fd_sc_hd__buf_2
XANTENNA__4122__A2 _1186_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5195_ cu.reg_file.reg_sp\[0\] _2085_ _2116_ VGND VGND VPWR VPWR _2117_ sky130_fd_sc_hd__mux2_1
X_4146_ _0917_ _1215_ VGND VGND VPWR VPWR _1216_ sky130_fd_sc_hd__and2_1
XFILLER_0_92_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5083__A0 _1074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4077_ _0570_ _0684_ VGND VGND VPWR VPWR _1151_ sky130_fd_sc_hd__nor2_1
X_3028_ ih.t.timer_max\[30\] _2765_ VGND VGND VPWR VPWR _2766_ sky130_fd_sc_hd__nor2_1
XANTENNA__3633__A1 _2950_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5386__A1 net124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4979_ _1948_ _1956_ VGND VGND VPWR VPWR _1967_ sky130_fd_sc_hd__and2b_1
XANTENNA__3397__B1 _0293_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5138__A1 _1144_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5689__A2 _1650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3321__B1 cu.id.cb_opcode_x\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5074__A0 _0617_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4821__A0 _1050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3624__A1 cu.reg_file.reg_l\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5916__A3 _2666_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5808__A cu.reg_file.reg_sp\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5129__A1 _1073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5301__A1 net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4000_ _1073_ VGND VGND VPWR VPWR _1074_ sky130_fd_sc_hd__buf_4
XFILLER_0_1_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5951_ _2684_ VGND VGND VPWR VPWR _0284_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3615__A1 cu.reg_file.reg_sp\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4902_ _1894_ _1895_ VGND VGND VPWR VPWR _1896_ sky130_fd_sc_hd__nor2_1
XFILLER_0_62_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3615__B2 cu.reg_file.reg_d\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5882_ _1074_ ih.t.timer_max\[2\] _2645_ VGND VGND VPWR VPWR _2648_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4833_ _1831_ _1832_ VGND VGND VPWR VPWR _1833_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_7_313 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5718__A _2351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4764_ _1268_ _1747_ VGND VGND VPWR VPWR _1772_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5437__B _2225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3715_ _0566_ VGND VGND VPWR VPWR _0791_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_496 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_43_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4695_ _1714_ _1715_ _1672_ VGND VGND VPWR VPWR _1716_ sky130_fd_sc_hd__and3b_1
XFILLER_0_70_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3646_ _0652_ _0663_ _0685_ _0718_ _0721_ VGND VGND VPWR VPWR _0722_ sky130_fd_sc_hd__a221o_1
XFILLER_0_87_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5453__A _1374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3577_ _0507_ VGND VGND VPWR VPWR _0653_ sky130_fd_sc_hd__buf_6
X_5316_ _1075_ net94 _2195_ VGND VGND VPWR VPWR _2198_ sky130_fd_sc_hd__mux2_1
X_6296_ clknet_leaf_42_clk _0278_ net152 VGND VGND VPWR VPWR cu.id.cb_opcode_z\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__3551__B1 _0624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5247_ _2154_ VGND VGND VPWR VPWR _0110_ sky130_fd_sc_hd__clkbuf_1
Xhold37 ih.t.count\[21\] VGND VGND VPWR VPWR net233 sky130_fd_sc_hd__dlygate4sd3_1
Xhold26 ih.t.count\[10\] VGND VGND VPWR VPWR net222 sky130_fd_sc_hd__dlygate4sd3_1
Xhold15 _0097_ VGND VGND VPWR VPWR net211 sky130_fd_sc_hd__dlygate4sd3_1
X_5178_ _2104_ VGND VGND VPWR VPWR _0091_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5056__A0 cu.reg_file.reg_c\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4129_ _0959_ _1198_ VGND VGND VPWR VPWR _1199_ sky130_fd_sc_hd__or2_1
XFILLER_0_66_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4031__B2 _0566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5295__A0 _1075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4098__B2 _1032_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4098__A1 _0916_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5047__A0 cu.reg_file.reg_b\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4270__A1 cu.reg_file.reg_a\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4270__B2 cu.reg_file.reg_sp\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1083 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1072 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1061 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1050 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1094 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4558__C1 _1323_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4573__A2 _1052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3500_ _0440_ VGND VGND VPWR VPWR _0576_ sky130_fd_sc_hd__buf_4
XFILLER_0_40_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4480_ cu.reg_file.reg_d\[3\] _1282_ _1286_ cu.reg_file.reg_sp\[11\] VGND VGND VPWR
+ VPWR _1537_ sky130_fd_sc_hd__a22o_1
XANTENNA__3781__B1 _0741_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3431_ _0504_ VGND VGND VPWR VPWR _0507_ sky130_fd_sc_hd__inv_2
XANTENNA__4325__A2 _0993_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6150_ clknet_leaf_8_clk _0184_ net168 VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__dfrtp_4
XTAP_801 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3362_ _2880_ _0437_ _0323_ VGND VGND VPWR VPWR _0438_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_20_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_834 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5101_ _1791_ _0366_ _2037_ VGND VGND VPWR VPWR _2055_ sky130_fd_sc_hd__and3_1
X_6081_ clknet_leaf_14_clk _0115_ net180 VGND VGND VPWR VPWR ih.t.timer_max\[29\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_867 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_856 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3293_ _2951_ _0368_ VGND VGND VPWR VPWR _0369_ sky130_fd_sc_hd__and2_1
XTAP_889 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_878 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5032_ cu.reg_file.reg_b\[1\] _2008_ _2006_ VGND VGND VPWR VPWR _2009_ sky130_fd_sc_hd__mux2_1
XFILLER_0_32_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_73_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5038__A0 cu.reg_file.reg_b\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5934_ _2876_ _2486_ _2668_ VGND VGND VPWR VPWR _2676_ sky130_fd_sc_hd__mux2_1
X_5865_ _2157_ ih.t.timer_max\[10\] _2636_ VGND VGND VPWR VPWR _2639_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4816_ _1299_ cu.pc.pc_o\[1\] VGND VGND VPWR VPWR _1817_ sky130_fd_sc_hd__xor2_1
X_5796_ _1110_ _2580_ _2545_ VGND VGND VPWR VPWR _2581_ sky130_fd_sc_hd__mux2_1
XFILLER_0_71_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4747_ _1754_ _1747_ VGND VGND VPWR VPWR _1756_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4678_ _1704_ VGND VGND VPWR VPWR ih.t.next_count\[14\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_31_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5513__B2 net61 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3629_ cu.reg_file.reg_h\[2\] _0495_ _0499_ cu.reg_file.reg_a\[2\] VGND VGND VPWR
+ VPWR _0705_ sky130_fd_sc_hd__a22o_1
Xoutput38 net38 VGND VGND VPWR VPWR memory_address_out[12] sky130_fd_sc_hd__buf_2
XFILLER_0_3_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput49 net49 VGND VGND VPWR VPWR memory_address_out[8] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6279_ clknet_leaf_13_clk _0261_ net180 VGND VGND VPWR VPWR ih.t.timer_max\[19\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__5277__A0 net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5029__A0 cu.reg_file.reg_b\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4246__B _1311_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4961__S _1808_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3763__B1 _0748_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5504__A1 _1374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3818__A1 cu.reg_file.reg_b\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3818__B2 cu.reg_file.reg_d\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5032__S _2006_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3980_ _0395_ _1019_ VGND VGND VPWR VPWR _1055_ sky130_fd_sc_hd__nor2_1
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4243__A1 _2883_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3995__B _0824_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5650_ net74 _1648_ _2137_ _2274_ VGND VGND VPWR VPWR _2464_ sky130_fd_sc_hd__a31o_1
XFILLER_0_57_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_0_clk clk VGND VGND VPWR VPWR clknet_0_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_17_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4601_ _1364_ _1489_ _1644_ VGND VGND VPWR VPWR _1645_ sky130_fd_sc_hd__a21o_1
XFILLER_0_72_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5581_ net79 _1633_ _2394_ _2397_ VGND VGND VPWR VPWR _2398_ sky130_fd_sc_hd__o22a_1
XFILLER_0_53_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4532_ _1585_ _1586_ _1356_ VGND VGND VPWR VPWR _1587_ sky130_fd_sc_hd__a21oi_1
XANTENNA__4900__A cu.pc.pc_o\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3754__B1 _0748_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4463_ cu.pc.pc_o\[10\] VGND VGND VPWR VPWR _1521_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_13_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6202_ clknet_leaf_4_clk net15 net171 VGND VGND VPWR VPWR ih.ih.ih.prev_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_3414_ _0464_ _0487_ _0482_ cu.reg_file.reg_l\[0\] VGND VGND VPWR VPWR _0490_ sky130_fd_sc_hd__o211a_1
X_4394_ _1396_ _1455_ VGND VGND VPWR VPWR _1456_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_40_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6133_ clknet_leaf_9_clk _0167_ net175 VGND VGND VPWR VPWR net125 sky130_fd_sc_hd__dfrtp_1
X_3345_ _0409_ _0407_ VGND VGND VPWR VPWR _0421_ sky130_fd_sc_hd__nand2_4
XTAP_620 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6064_ clknet_leaf_23_clk _0098_ net192 VGND VGND VPWR VPWR mc.cc.count\[1\] sky130_fd_sc_hd__dfstp_1
XTAP_686 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3276_ _0348_ _0351_ VGND VGND VPWR VPWR _0352_ sky130_fd_sc_hd__nor2_2
XANTENNA__3809__A1 cu.reg_file.reg_mem\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_653 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5015_ cu.reg_file.reg_a\[5\] _1995_ _1985_ VGND VGND VPWR VPWR _1996_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout181_A net182 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4482__A1 cu.id.imm_i\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4482__B2 cu.pc.pc_o\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5917_ _1780_ _2532_ cu.id.can_be_interrupted VGND VGND VPWR VPWR _2667_ sky130_fd_sc_hd__o21ai_1
X_5848_ _2618_ _2621_ _2619_ VGND VGND VPWR VPWR _2626_ sky130_fd_sc_hd__a21boi_1
X_5779_ _2564_ _2565_ VGND VGND VPWR VPWR _2566_ sky130_fd_sc_hd__xnor2_1
XANTENNA__5991__RESET_B net161 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_550 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3161__A _2893_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6097__RESET_B net195 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_54_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3100__S ih.t.timer_max\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5816__A cu.reg_file.reg_sp\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5489__B1 _2247_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output75_A net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3130_ ih.t.count\[30\] _2866_ VGND VGND VPWR VPWR _2868_ sky130_fd_sc_hd__nand2_1
XFILLER_0_38_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3061_ _2758_ _2798_ ih.t.count\[18\] VGND VGND VPWR VPWR _2799_ sky130_fd_sc_hd__a21oi_1
XANTENNA__4464__B2 cu.reg_file.reg_sp\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4464__A1 cu.reg_file.reg_d\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4167__A _0617_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5413__A0 _1190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5964__A1 _2448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4767__A2 _1632_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3963_ _0918_ _1029_ _1034_ _1037_ VGND VGND VPWR VPWR _1038_ sky130_fd_sc_hd__o22a_1
X_5702_ ih.t.timer_max\[30\] _2151_ _2320_ ih.t.timer_max\[14\] VGND VGND VPWR VPWR
+ _2508_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_72_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3894_ _0967_ _0969_ _0328_ VGND VGND VPWR VPWR _0970_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_72_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5633_ _2444_ _2445_ _2447_ _1641_ VGND VGND VPWR VPWR _2448_ sky130_fd_sc_hd__o22a_4
XFILLER_0_45_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_33_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5564_ _1400_ _2381_ VGND VGND VPWR VPWR _2382_ sky130_fd_sc_hd__and2b_1
X_4515_ _1382_ _1564_ _1565_ _1570_ VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__a31o_1
XFILLER_0_79_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5495_ ih.t.enable _2257_ _2192_ ih.t.timer_max\[8\] VGND VGND VPWR VPWR _2315_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4446_ _1503_ _1504_ _1296_ VGND VGND VPWR VPWR _1505_ sky130_fd_sc_hd__o21a_1
X_4377_ _1415_ _1434_ VGND VGND VPWR VPWR _1440_ sky130_fd_sc_hd__nor2_1
XANTENNA__4152__B1 _0824_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6116_ clknet_leaf_24_clk _0150_ net190 VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__dfrtp_2
XFILLER_0_0_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3328_ _2925_ _2890_ _2932_ VGND VGND VPWR VPWR _0404_ sky130_fd_sc_hd__or3_1
XTAP_450 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_461 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6047_ clknet_leaf_4_clk _0085_ net170 VGND VGND VPWR VPWR cu.reg_file.reg_l\[5\]
+ sky130_fd_sc_hd__dfrtp_2
X_3259_ _0321_ _0322_ _0328_ _0334_ VGND VGND VPWR VPWR _0335_ sky130_fd_sc_hd__nor4_2
XFILLER_0_68_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5400__S _2237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3430__A2 _0498_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_output113_A net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5946__A1 _2448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3421__A2 _0492_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5280_ _2175_ VGND VGND VPWR VPWR _0122_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_49_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4300_ cu.pc.pc_o\[2\] _1322_ _1317_ cu.reg_file.reg_l\[2\] _1365_ VGND VGND VPWR
+ VPWR _1366_ sky130_fd_sc_hd__a221o_1
X_4231_ cu.pc.pc_o\[0\] VGND VGND VPWR VPWR _1299_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__5882__A0 _1074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3488__A2 _0499_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3893__C1 _0968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4162_ _1209_ _1213_ _1222_ _1231_ VGND VGND VPWR VPWR _1232_ sky130_fd_sc_hd__nor4_1
X_3113_ _2821_ _2823_ _2824_ _2850_ VGND VGND VPWR VPWR _2851_ sky130_fd_sc_hd__or4_1
X_4093_ _1090_ _1164_ VGND VGND VPWR VPWR _1167_ sky130_fd_sc_hd__nand2_1
X_3044_ ih.t.timer_max\[24\] _2761_ VGND VGND VPWR VPWR _2782_ sky130_fd_sc_hd__nand2_1
XANTENNA__4625__A _1666_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4995_ cu.pc.pc_o\[15\] _1981_ _1814_ VGND VGND VPWR VPWR _1982_ sky130_fd_sc_hd__mux2_1
X_3946_ _1012_ _0996_ _1016_ _1021_ VGND VGND VPWR VPWR _1022_ sky130_fd_sc_hd__or4_1
XFILLER_0_73_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3877_ _0737_ _0752_ _0899_ VGND VGND VPWR VPWR _0953_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_33_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5616_ net129 _2236_ _2247_ net137 VGND VGND VPWR VPWR _2431_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5547_ ih.gpio_interrupt_mask\[1\] _2326_ _2365_ _2125_ _2327_ VGND VGND VPWR VPWR
+ _2366_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5478_ net65 _0618_ _2300_ VGND VGND VPWR VPWR _2301_ sky130_fd_sc_hd__mux2_1
X_4429_ _1488_ VGND VGND VPWR VPWR _1489_ sky130_fd_sc_hd__buf_4
XANTENNA__5873__A0 _2165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_291 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_280 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6300__RESET_B net160 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5130__S _2069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4535__A cu.reg_file.reg_sp\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5928__A1 _2429_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_51_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5305__S _2182_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6041__RESET_B net162 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5616__B1 _2247_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5092__A1 _1209_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5040__S _2002_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4780_ _1768_ _1784_ _0350_ VGND VGND VPWR VPWR _1785_ sky130_fd_sc_hd__o21a_1
X_3800_ _0874_ _0871_ VGND VGND VPWR VPWR _0876_ sky130_fd_sc_hd__and2b_1
X_3731_ _0572_ _0510_ _0712_ VGND VGND VPWR VPWR _0807_ sky130_fd_sc_hd__or3b_1
XFILLER_0_27_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3662_ _2950_ _2913_ _0536_ VGND VGND VPWR VPWR _0738_ sky130_fd_sc_hd__and3_1
X_5401_ _2245_ VGND VGND VPWR VPWR _0173_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3593_ cu.reg_file.reg_mem\[4\] _0418_ _0433_ cu.reg_file.reg_a\[4\] VGND VGND VPWR
+ VPWR _0669_ sky130_fd_sc_hd__a22o_1
X_5332_ _2207_ VGND VGND VPWR VPWR _0142_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_2_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5263_ _1126_ _1624_ _1666_ VGND VGND VPWR VPWR _2165_ sky130_fd_sc_hd__mux2_1
XANTENNA__4339__B _1401_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5194_ _2115_ VGND VGND VPWR VPWR _2116_ sky130_fd_sc_hd__inv_2
X_4214_ _1279_ _1275_ VGND VGND VPWR VPWR _1282_ sky130_fd_sc_hd__nor2b_2
X_4145_ _1214_ _0779_ VGND VGND VPWR VPWR _1215_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5083__A1 _1226_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4076_ _0918_ _0766_ _1149_ _0517_ VGND VGND VPWR VPWR _1150_ sky130_fd_sc_hd__o211a_1
XFILLER_0_92_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3027_ ih.t.timer_max\[28\] ih.t.timer_max\[29\] _2764_ VGND VGND VPWR VPWR _2765_
+ sky130_fd_sc_hd__or3_1
XANTENNA__3633__A2 _0341_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4978_ _1233_ cu.pc.pc_o\[14\] VGND VGND VPWR VPWR _1966_ sky130_fd_sc_hd__xor2_1
XFILLER_0_80_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3929_ _0976_ _0980_ _1004_ VGND VGND VPWR VPWR _1005_ sky130_fd_sc_hd__or3_1
XFILLER_0_18_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5074__A1 _1622_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_504 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5824__A cu.reg_file.reg_sp\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5035__S _2006_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5837__A0 cu.reg_file.reg_sp\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5950_ _1233_ _2486_ _2666_ VGND VGND VPWR VPWR _2684_ sky130_fd_sc_hd__mux2_1
X_4901_ cu.pc.pc_o\[7\] _1872_ cu.pc.pc_o\[8\] VGND VGND VPWR VPWR _1895_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4812__A1 _2948_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4812__B2 _1484_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5881_ _2647_ VGND VGND VPWR VPWR _0251_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4832_ _0340_ cu.pc.pc_o\[1\] _1819_ VGND VGND VPWR VPWR _1832_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_62_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4763_ _1739_ _1770_ VGND VGND VPWR VPWR _1771_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_28_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4576__B1 _1213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4694_ ih.t.count\[18\] ih.t.count\[19\] _1708_ ih.t.count\[20\] VGND VGND VPWR VPWR
+ _1715_ sky130_fd_sc_hd__a31o_1
X_3714_ _0643_ _0632_ VGND VGND VPWR VPWR _0790_ sky130_fd_sc_hd__and2b_1
XFILLER_0_43_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5990__SET_B net188 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3645_ _0719_ _0720_ VGND VGND VPWR VPWR _0721_ sky130_fd_sc_hd__and2b_1
XFILLER_0_87_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3576_ _0576_ _0646_ _0648_ _0651_ VGND VGND VPWR VPWR _0652_ sky130_fd_sc_hd__o2bb2a_4
XFILLER_0_30_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5315_ _2197_ VGND VGND VPWR VPWR _0135_ sky130_fd_sc_hd__clkbuf_1
X_6295_ clknet_leaf_42_clk _0277_ net152 VGND VGND VPWR VPWR cu.id.cb_opcode_z\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__3551__B2 cu.reg_file.reg_sp\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3551__A1 cu.reg_file.reg_h\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5828__A0 _1222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5246_ ih.t.timer_max\[24\] _2144_ _2153_ VGND VGND VPWR VPWR _2154_ sky130_fd_sc_hd__mux2_1
XFILLER_0_53_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold27 ih.t.count\[13\] VGND VGND VPWR VPWR net223 sky130_fd_sc_hd__dlygate4sd3_1
Xhold16 ih.t.count\[19\] VGND VGND VPWR VPWR net212 sky130_fd_sc_hd__dlygate4sd3_1
Xhold38 ih.t.count\[15\] VGND VGND VPWR VPWR net234 sky130_fd_sc_hd__dlygate4sd3_1
X_5177_ _1647_ _2103_ VGND VGND VPWR VPWR _2104_ sky130_fd_sc_hd__and2_1
XANTENNA__5056__A1 _2022_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4128_ _0949_ _0958_ _0779_ VGND VGND VPWR VPWR _1198_ sky130_fd_sc_hd__a21o_1
X_4059_ _0917_ _0757_ _0804_ _0776_ VGND VGND VPWR VPWR _1133_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_93_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4813__A _1814_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5295__A1 net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1040 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1073 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1062 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1051 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1095 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1084 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_507 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4558__B1 _1343_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4161__C _1226_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3781__A1 cu.reg_file.reg_d\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3781__B2 cu.reg_file.reg_h\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3430_ alu.Cin _0498_ _0499_ cu.reg_file.reg_a\[0\] _0505_ VGND VGND VPWR VPWR _0506_
+ sky130_fd_sc_hd__a221o_1
X_3361_ _0308_ _0315_ _0435_ _0436_ VGND VGND VPWR VPWR _0437_ sky130_fd_sc_hd__and4bb_2
XANTENNA__4730__B1 _1644_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6080_ clknet_leaf_22_clk _0114_ net191 VGND VGND VPWR VPWR ih.t.timer_max\[28\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_835 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5100_ _2054_ VGND VGND VPWR VPWR _0063_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_57_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3717__A_N _0652_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_868 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_857 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5031_ _1051_ _1623_ _2002_ VGND VGND VPWR VPWR _2008_ sky130_fd_sc_hd__mux2_1
X_3292_ _2953_ _0339_ _0352_ _0367_ VGND VGND VPWR VPWR _0368_ sky130_fd_sc_hd__o211a_4
XTAP_879 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5933_ _2675_ VGND VGND VPWR VPWR _0275_ sky130_fd_sc_hd__clkbuf_1
X_5864_ _2638_ VGND VGND VPWR VPWR _0243_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4815_ _1816_ VGND VGND VPWR VPWR _0016_ sky130_fd_sc_hd__clkbuf_1
X_5795_ _2578_ _2579_ VGND VGND VPWR VPWR _2580_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3247__A_N _2878_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4746_ _1483_ _1748_ _1754_ VGND VGND VPWR VPWR _1755_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_16_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3772__A1 cu.pc.pc_o\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4677_ _1702_ _1703_ _1672_ VGND VGND VPWR VPWR _1704_ sky130_fd_sc_hd__and3b_1
XANTENNA__5464__A _2194_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3628_ cu.reg_file.reg_c\[2\] _0485_ _0489_ cu.reg_file.reg_e\[2\] _0703_ VGND VGND
+ VPWR VPWR _0704_ sky130_fd_sc_hd__a221o_1
Xoutput39 net39 VGND VGND VPWR VPWR memory_address_out[13] sky130_fd_sc_hd__buf_2
X_3559_ _0295_ _2921_ _0634_ VGND VGND VPWR VPWR _0635_ sky130_fd_sc_hd__or3_1
X_6278_ clknet_leaf_12_clk _0260_ net177 VGND VGND VPWR VPWR ih.t.timer_max\[18\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__5498__A1_N ih.t.timer_max\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5277__A1 _1187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5229_ _1306_ _2137_ VGND VGND VPWR VPWR _2138_ sky130_fd_sc_hd__and2_1
XFILLER_0_85_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_39_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_62_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3763__A1 cu.reg_file.reg_sp\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3763__B2 cu.reg_file.reg_h\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3515__A1 cu.reg_file.reg_sp\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3515__B2 cu.reg_file.reg_h\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_30_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3818__A2 _0426_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3341__B _0405_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_72_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4600_ _1632_ _1643_ VGND VGND VPWR VPWR _1644_ sky130_fd_sc_hd__nor2_4
XFILLER_0_57_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5580_ net111 _2147_ _2225_ net119 _2396_ VGND VGND VPWR VPWR _2397_ sky130_fd_sc_hd__a221o_1
XFILLER_0_25_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4531_ _1567_ _1579_ VGND VGND VPWR VPWR _1586_ sky130_fd_sc_hd__nand2_1
XANTENNA__4900__B cu.pc.pc_o\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3754__A1 cu.reg_file.reg_sp\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3754__B2 cu.reg_file.reg_h\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4462_ _1513_ _1514_ VGND VGND VPWR VPWR _1520_ sky130_fd_sc_hd__nand2_1
X_6201_ clknet_leaf_4_clk net14 net172 VGND VGND VPWR VPWR ih.ih.ih.prev_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_7_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3506__A1 _0341_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3413_ _0480_ _0487_ _0488_ VGND VGND VPWR VPWR _0489_ sky130_fd_sc_hd__a21o_2
X_4393_ _1449_ _1450_ _1454_ VGND VGND VPWR VPWR _1455_ sky130_fd_sc_hd__o21a_2
X_6132_ clknet_leaf_26_clk _0166_ net195 VGND VGND VPWR VPWR net124 sky130_fd_sc_hd__dfrtp_4
X_3344_ cu.reg_file.reg_mem\[0\] _0418_ _0419_ cu.reg_file.reg_h\[0\] VGND VGND VPWR
+ VPWR _0420_ sky130_fd_sc_hd__a22o_1
XTAP_610 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6063_ clknet_leaf_25_clk net211 net195 VGND VGND VPWR VPWR mc.cc.count\[0\] sky130_fd_sc_hd__dfrtp_1
XTAP_676 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3275_ _0299_ _2953_ _0349_ _2914_ _0350_ VGND VGND VPWR VPWR _0351_ sky130_fd_sc_hd__a221o_1
XTAP_654 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_687 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3809__A2 _0640_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5014_ _1191_ _1209_ _0368_ VGND VGND VPWR VPWR _1995_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5916_ _1484_ _2351_ _2666_ _2665_ cu.ir.idx\[1\] VGND VGND VPWR VPWR _0267_ sky130_fd_sc_hd__a32o_1
XFILLER_0_75_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5195__A0 cu.reg_file.reg_sp\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5847_ cu.reg_file.reg_sp\[14\] _1287_ VGND VGND VPWR VPWR _2625_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5778_ _2550_ _2551_ _2557_ _2556_ _2549_ VGND VGND VPWR VPWR _2565_ sky130_fd_sc_hd__a311o_1
X_4729_ _1738_ VGND VGND VPWR VPWR ih.t.next_count\[31\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_16_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5498__B2 _1400_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_180 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5133__S _2069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5670__A1 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4972__S _1808_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4704__C _1672_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__6066__RESET_B net195 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4933__A0 _1226_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5489__B2 net132 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5489__A1 net124 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5832__A cu.reg_file.reg_sp\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4448__A cu.reg_file.reg_h\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output68_A net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3060_ ih.t.timer_max\[18\] _2757_ VGND VGND VPWR VPWR _2798_ sky130_fd_sc_hd__nand2_1
XANTENNA__5043__S _2002_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5661__A1 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4464__A2 _1282_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4167__B _1050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5413__A1 net136 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5701_ net6 _1650_ _2488_ _2507_ VGND VGND VPWR VPWR _0211_ sky130_fd_sc_hd__a31o_1
XANTENNA__4767__A3 _1643_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3962_ _0572_ _0510_ _0401_ _1035_ _1036_ VGND VGND VPWR VPWR _1037_ sky130_fd_sc_hd__o311a_1
XFILLER_0_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3893_ _2893_ _0386_ _0308_ _0968_ VGND VGND VPWR VPWR _0969_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_45_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5632_ _1649_ _2446_ VGND VGND VPWR VPWR _2447_ sky130_fd_sc_hd__and2_1
XANTENNA__4630__B _1670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5563_ ih.t.timer_max\[10\] _2193_ _2314_ ih.t.timer_max\[2\] _2380_ VGND VGND VPWR
+ VPWR _2381_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4514_ _1402_ _1561_ _1569_ _1371_ VGND VGND VPWR VPWR _1570_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_79_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5494_ _1400_ _2287_ VGND VGND VPWR VPWR _2314_ sky130_fd_sc_hd__nor2_2
XFILLER_0_79_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4445_ cu.reg_file.reg_b\[1\] _1281_ _1283_ cu.reg_file.reg_d\[1\] VGND VGND VPWR
+ VPWR _1504_ sky130_fd_sc_hd__a22o_1
XANTENNA__5742__A _0296_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4376_ _1419_ _1423_ _1437_ VGND VGND VPWR VPWR _1439_ sky130_fd_sc_hd__nand3_1
XANTENNA__5461__B _2284_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6115_ clknet_leaf_27_clk _0149_ net186 VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__dfrtp_4
X_3327_ _2878_ _0402_ _2877_ VGND VGND VPWR VPWR _0403_ sky130_fd_sc_hd__a21o_1
XTAP_440 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_462 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3258_ _0329_ _0332_ _0333_ VGND VGND VPWR VPWR _0334_ sky130_fd_sc_hd__or3_2
XTAP_495 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6046_ clknet_leaf_3_clk _0084_ net156 VGND VGND VPWR VPWR cu.reg_file.reg_l\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_3189_ _2925_ _2901_ VGND VGND VPWR VPWR _2926_ sky130_fd_sc_hd__nor2_1
XFILLER_0_95_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4391__A1 cu.pc.pc_o\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5652__A _1649_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5643__A1 ih.t.timer_max\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_2_0__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_0__leaf_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA_output106_A net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_67_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_315 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5038__S _2006_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_23_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5331__A0 _0619_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4230_ _1297_ VGND VGND VPWR VPWR _1298_ sky130_fd_sc_hd__buf_2
XANTENNA__5882__A1 ih.t.timer_max\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4161_ _0516_ _0819_ _1226_ _1230_ VGND VGND VPWR VPWR _1231_ sky130_fd_sc_hd__or4b_1
XANTENNA__3082__A ih.t.timer_max\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3893__B1 _0308_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3112_ _2826_ _2827_ _2849_ VGND VGND VPWR VPWR _2850_ sky130_fd_sc_hd__or3_1
X_4092_ _0519_ _1165_ _0614_ _0551_ VGND VGND VPWR VPWR _1166_ sky130_fd_sc_hd__o211ai_1
XANTENNA__5634__A1 _2448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3043_ ih.t.count\[25\] _2780_ VGND VGND VPWR VPWR _2781_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_65_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5398__A0 _1194_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4994_ _1975_ _1980_ _1808_ VGND VGND VPWR VPWR _1981_ sky130_fd_sc_hd__mux2_1
X_3945_ _0982_ _0997_ _0986_ VGND VGND VPWR VPWR _1021_ sky130_fd_sc_hd__nor3b_2
XFILLER_0_85_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5615_ _2430_ VGND VGND VPWR VPWR _0202_ sky130_fd_sc_hd__clkbuf_1
X_3876_ _0887_ _0901_ VGND VGND VPWR VPWR _0952_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_33_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5546_ mc.cl.next_data\[1\] _2359_ _2324_ _2364_ VGND VGND VPWR VPWR _2365_ sky130_fd_sc_hd__a22o_1
X_5477_ _2299_ _2284_ VGND VGND VPWR VPWR _2300_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5472__A _2147_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4428_ _1269_ _1484_ VGND VGND VPWR VPWR _1488_ sky130_fd_sc_hd__nor2_1
XANTENNA__5322__A0 _1192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5873__A1 ih.t.timer_max\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4359_ _1397_ _1395_ _1421_ VGND VGND VPWR VPWR _1423_ sky130_fd_sc_hd__a21o_1
XANTENNA__4088__A _0617_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_292 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_270 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4816__A _1299_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6029_ clknet_leaf_1_clk _0067_ net153 VGND VGND VPWR VPWR cu.reg_file.reg_e\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_68_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5411__S _2248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4535__B _1286_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5366__B _2225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5696__A2_N _1643_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4116__B2 _1188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5616__A1 net129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5616__B2 net137 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3730_ _0759_ _0783_ VGND VGND VPWR VPWR _0806_ sky130_fd_sc_hd__xor2_1
XFILLER_0_27_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3661_ _0645_ _0722_ _0734_ _0736_ _0730_ VGND VGND VPWR VPWR _0737_ sky130_fd_sc_hd__a311o_1
XFILLER_0_70_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5400_ _1261_ net131 _2237_ VGND VGND VPWR VPWR _2245_ sky130_fd_sc_hd__mux2_1
X_3592_ cu.reg_file.reg_c\[4\] _0427_ _0430_ cu.reg_file.reg_e\[4\] VGND VGND VPWR
+ VPWR _0668_ sky130_fd_sc_hd__a22o_1
X_5331_ _0619_ net100 _2206_ VGND VGND VPWR VPWR _2207_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5262_ _2164_ VGND VGND VPWR VPWR _0115_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_55_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4213_ _1280_ VGND VGND VPWR VPWR _1281_ sky130_fd_sc_hd__buf_2
X_5193_ _2114_ VGND VGND VPWR VPWR _2115_ sky130_fd_sc_hd__buf_2
X_4144_ _0952_ _0955_ VGND VGND VPWR VPWR _1214_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4075_ _0767_ _0773_ _1145_ _1148_ VGND VGND VPWR VPWR _1149_ sky130_fd_sc_hd__a31o_1
X_3026_ ih.t.timer_max\[27\] _2763_ VGND VGND VPWR VPWR _2764_ sky130_fd_sc_hd__or2_2
XANTENNA__4355__B _1415_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4977_ _1963_ _1964_ VGND VGND VPWR VPWR _1965_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3928_ _0994_ _0989_ VGND VGND VPWR VPWR _1004_ sky130_fd_sc_hd__or2b_1
XFILLER_0_18_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3859_ _0898_ _0934_ VGND VGND VPWR VPWR _0935_ sky130_fd_sc_hd__xor2_1
XFILLER_0_33_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4346__A1 _0374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4346__B2 cu.pc.pc_o\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5529_ _1649_ _2347_ _2348_ _1641_ VGND VGND VPWR VPWR _2349_ sky130_fd_sc_hd__a31o_1
XANTENNA__3715__A _0566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3003__A_N net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5141__S _2066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_516 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5534__B1 _2247_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5316__S _2195_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5840__A cu.reg_file.reg_sp\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output50_A net50 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3360__A _2908_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5880_ _1051_ ih.t.timer_max\[1\] _2645_ VGND VGND VPWR VPWR _2647_ sky130_fd_sc_hd__mux2_1
X_4900_ cu.pc.pc_o\[7\] cu.pc.pc_o\[8\] _1872_ VGND VGND VPWR VPWR _1894_ sky130_fd_sc_hd__and3_1
XANTENNA__4812__A2 _1808_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5448__S0 _1354_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4831_ _1829_ _1830_ VGND VGND VPWR VPWR _1831_ sky130_fd_sc_hd__and2b_1
XFILLER_0_28_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4191__A _1110_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4762_ _1301_ _1300_ _1748_ _1268_ VGND VGND VPWR VPWR _1770_ sky130_fd_sc_hd__a31o_1
XANTENNA__5773__A0 cu.reg_file.reg_sp\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4576__A1 _2702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4576__B2 _2697_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4693_ ih.t.count\[19\] ih.t.count\[20\] _1711_ VGND VGND VPWR VPWR _1714_ sky130_fd_sc_hd__and3_1
X_3713_ _0664_ _0684_ _0787_ _0788_ VGND VGND VPWR VPWR _0789_ sky130_fd_sc_hd__nand4_1
X_3644_ _0671_ _0681_ VGND VGND VPWR VPWR _0720_ sky130_fd_sc_hd__and2_1
XFILLER_0_30_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3575_ cu.reg_file.reg_l\[5\] _0422_ _0649_ _0650_ _0576_ VGND VGND VPWR VPWR _0651_
+ sky130_fd_sc_hd__a2111o_1
X_5314_ _1052_ net93 _2195_ VGND VGND VPWR VPWR _2197_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_376 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6294_ clknet_leaf_41_clk _0276_ net151 VGND VGND VPWR VPWR cu.id.opcode\[7\] sky130_fd_sc_hd__dfrtp_2
XANTENNA__3551__A2 _0495_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5245_ _1667_ _2147_ _2152_ VGND VGND VPWR VPWR _2153_ sky130_fd_sc_hd__o21a_4
Xhold17 ih.t.next_count\[19\] VGND VGND VPWR VPWR net213 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__4500__A1 _1296_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold28 cu.ir.idx\[0\] VGND VGND VPWR VPWR net224 sky130_fd_sc_hd__dlygate4sd3_1
X_5176_ mc.cl.next_data\[11\] net21 mc.count VGND VGND VPWR VPWR _2103_ sky130_fd_sc_hd__mux2_1
Xhold39 cu.id.is_halted VGND VGND VPWR VPWR net235 sky130_fd_sc_hd__dlygate4sd3_1
X_4127_ _0916_ _0944_ _1196_ _1032_ _0918_ VGND VGND VPWR VPWR _1197_ sky130_fd_sc_hd__o221a_1
X_4058_ _0757_ _0767_ VGND VGND VPWR VPWR _1132_ sky130_fd_sc_hd__nand2_1
X_3009_ ih.t.timer_max\[3\] _2746_ VGND VGND VPWR VPWR _2747_ sky130_fd_sc_hd__or2_1
XFILLER_0_38_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_454 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5764__A0 _1089_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4319__B2 cu.reg_file.reg_sp\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4319__A1 cu.reg_file.reg_a\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3445__A _2936_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5136__S _2069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1030 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1074 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1063 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1052 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1041 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1096 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1085 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4558__A1 cu.reg_file.reg_sp\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3339__B _0405_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3781__A2 _0488_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output98_A net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5046__S _2002_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3360_ _2908_ _0342_ VGND VGND VPWR VPWR _0436_ sky130_fd_sc_hd__nor2_1
XANTENNA__4730__A1 _1364_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_825 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_858 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5030_ _2007_ VGND VGND VPWR VPWR _0040_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3291_ _0350_ _0358_ _0366_ VGND VGND VPWR VPWR _0367_ sky130_fd_sc_hd__o21a_1
XTAP_869 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5932_ _2875_ _2467_ _2668_ VGND VGND VPWR VPWR _2675_ sky130_fd_sc_hd__mux2_1
XFILLER_0_87_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4914__A cu.pc.pc_o\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5863_ _2155_ ih.t.timer_max\[9\] _2636_ VGND VGND VPWR VPWR _2638_ sky130_fd_sc_hd__mux2_1
X_4814_ _1299_ _1810_ _1815_ VGND VGND VPWR VPWR _1816_ sky130_fd_sc_hd__mux2_1
X_5794_ _2569_ _2572_ _2570_ VGND VGND VPWR VPWR _2579_ sky130_fd_sc_hd__a21bo_1
X_4745_ _0296_ _0320_ _1319_ _1753_ VGND VGND VPWR VPWR _1754_ sky130_fd_sc_hd__or4_1
XFILLER_0_28_295 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4676_ ih.t.count\[12\] ih.t.count\[13\] _1696_ ih.t.count\[14\] VGND VGND VPWR VPWR
+ _1703_ sky130_fd_sc_hd__a31o_1
XFILLER_0_31_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3772__A2 _0740_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3627_ _0464_ _0487_ _0482_ cu.reg_file.reg_l\[2\] VGND VGND VPWR VPWR _0703_ sky130_fd_sc_hd__o211a_1
X_3558_ _0322_ _0633_ _0443_ VGND VGND VPWR VPWR _0634_ sky130_fd_sc_hd__o21ba_1
XANTENNA__6184__RESET_B net162 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6277_ clknet_leaf_12_clk _0259_ net178 VGND VGND VPWR VPWR ih.t.timer_max\[17\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__5480__A _2236_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3489_ _0294_ _0372_ _0536_ VGND VGND VPWR VPWR _0565_ sky130_fd_sc_hd__o21ai_1
X_5228_ _1415_ _2136_ VGND VGND VPWR VPWR _2137_ sky130_fd_sc_hd__nor2_4
XANTENNA__4485__B1 _1343_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5159_ cu.reg_file.reg_l\[4\] _1189_ _2088_ VGND VGND VPWR VPWR _2093_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_36_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_36_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_78_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_168 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3515__A2 _0413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3279__A1 _0340_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output136_A net136 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_27_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_27_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__4453__B _1511_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4530_ _1567_ _1579_ VGND VGND VPWR VPWR _1585_ sky130_fd_sc_hd__or2_1
X_4461_ _1515_ _1516_ _1519_ VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__o21ai_4
XFILLER_0_13_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6200_ clknet_leaf_6_clk net13 net166 VGND VGND VPWR VPWR ih.ih.ih.prev_data\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_3412_ net146 _0473_ _0479_ _0486_ _0483_ VGND VGND VPWR VPWR _0488_ sky130_fd_sc_hd__o2111a_4
XFILLER_0_40_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6131_ clknet_leaf_19_clk _0165_ net190 VGND VGND VPWR VPWR net123 sky130_fd_sc_hd__dfrtp_2
X_4392_ cu.reg_file.reg_c\[6\] _1313_ _1451_ _1453_ VGND VGND VPWR VPWR _1454_ sky130_fd_sc_hd__a211o_1
XTAP_600 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_68_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3343_ _0412_ _0414_ _0405_ VGND VGND VPWR VPWR _0419_ sky130_fd_sc_hd__nor3b_4
XTAP_611 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4628__B _2869_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6062_ clknet_leaf_24_clk mc.rw.next_state\[2\] net195 VGND VGND VPWR VPWR mc.rw.state\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_677 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3274_ _0296_ VGND VGND VPWR VPWR _0350_ sky130_fd_sc_hd__clkbuf_4
XTAP_644 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_688 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5013_ _1994_ VGND VGND VPWR VPWR _0036_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_84_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_18_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_18_clk sky130_fd_sc_hd__clkbuf_16
X_5915_ _2663_ cu.ir.idx\[1\] VGND VGND VPWR VPWR _2666_ sky130_fd_sc_hd__nor2_4
X_5846_ _2624_ VGND VGND VPWR VPWR _0239_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_36_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_63_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2989_ net8 VGND VGND VPWR VPWR _2728_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5777_ _2562_ _2563_ VGND VGND VPWR VPWR _2564_ sky130_fd_sc_hd__nand2_1
XANTENNA__5195__A1 _2085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4728_ _1672_ _1736_ _1737_ VGND VGND VPWR VPWR _1738_ sky130_fd_sc_hd__and3_1
XFILLER_0_16_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4659_ net229 _1689_ _1687_ VGND VGND VPWR VPWR _1692_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_71_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5670__A2 _1648_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5958__A0 cu.id.imm_i\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3984__A2 _1052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_224 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5489__A2 _2236_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6035__RESET_B net161 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5324__S _2195_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4551__A2_N _1598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3352__B _0405_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5661__A2 _1633_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4167__C _1073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3961_ _0781_ _0712_ _0773_ VGND VGND VPWR VPWR _1036_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_70_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5700_ _2506_ _1643_ cu.reg_file.reg_mem\[13\] _1646_ VGND VGND VPWR VPWR _2507_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_18_508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3892_ _0379_ _0448_ VGND VGND VPWR VPWR _0968_ sky130_fd_sc_hd__or2_2
XFILLER_0_45_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5631_ net13 _2345_ _2369_ net6 VGND VGND VPWR VPWR _2446_ sky130_fd_sc_hd__a22o_1
XFILLER_0_57_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5562_ ih.t.timer_max\[26\] _2146_ _2204_ ih.t.timer_max\[18\] VGND VGND VPWR VPWR
+ _2380_ sky130_fd_sc_hd__a22o_1
XFILLER_0_26_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4513_ _1567_ _1568_ VGND VGND VPWR VPWR _1569_ sky130_fd_sc_hd__nand2_1
XFILLER_0_53_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5493_ mc.cl.cmp_o _1648_ _1631_ VGND VGND VPWR VPWR _2313_ sky130_fd_sc_hd__and3_2
Xclkbuf_leaf_7_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_7_clk sky130_fd_sc_hd__clkbuf_16
X_4444_ cu.reg_file.reg_sp\[9\] _1287_ _1285_ cu.reg_file.reg_h\[1\] VGND VGND VPWR
+ VPWR _1503_ sky130_fd_sc_hd__a22o_1
XANTENNA__3246__C _2935_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4639__A _1672_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4375_ _1419_ _1423_ _1437_ VGND VGND VPWR VPWR _1438_ sky130_fd_sc_hd__a21o_1
XANTENNA__5123__B1_N _2951_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3543__A _0618_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6114_ clknet_leaf_27_clk _0148_ net186 VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__dfrtp_4
X_3326_ _2899_ _2900_ _2894_ VGND VGND VPWR VPWR _0402_ sky130_fd_sc_hd__a21bo_1
XTAP_430 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6045_ clknet_leaf_4_clk _0083_ net170 VGND VGND VPWR VPWR cu.reg_file.reg_l\[3\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_452 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3257_ _2888_ _2927_ _2933_ _2934_ VGND VGND VPWR VPWR _0333_ sky130_fd_sc_hd__and4_1
XTAP_496 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3188_ _2892_ _2894_ VGND VGND VPWR VPWR _2925_ sky130_fd_sc_hd__nand2_4
XFILLER_0_95_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3415__B2 cu.reg_file.reg_e\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3415__A1 cu.reg_file.reg_c\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5829_ cu.reg_file.reg_sp\[11\] _2609_ _2538_ VGND VGND VPWR VPWR _2610_ sky130_fd_sc_hd__mux2_1
XANTENNA__5409__S _2248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5144__S _2066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3351__B1 _0426_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5643__A2 _2193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5159__A1 _1189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output80_A net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5331__A1 net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4160_ _1032_ _1227_ _1228_ _1229_ VGND VGND VPWR VPWR _1230_ sky130_fd_sc_hd__o211a_2
X_3111_ _2829_ _2831_ _2832_ _2848_ VGND VGND VPWR VPWR _2849_ sky130_fd_sc_hd__or4_1
XANTENNA__3893__A1 _2893_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4091_ _0820_ VGND VGND VPWR VPWR _1165_ sky130_fd_sc_hd__inv_2
XANTENNA__5095__A0 _1193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3042_ ih.t.timer_max\[25\] _2762_ VGND VGND VPWR VPWR _2780_ sky130_fd_sc_hd__xor2_1
XANTENNA__4194__A _0516_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5398__A1 net130 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4993_ _1978_ _1979_ _1798_ VGND VGND VPWR VPWR _1980_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3944_ _0531_ _1018_ _1019_ VGND VGND VPWR VPWR _1020_ sky130_fd_sc_hd__nand3_1
XFILLER_0_58_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3875_ _0877_ _0904_ VGND VGND VPWR VPWR _0951_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_45_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5614_ cu.reg_file.reg_mem\[4\] _2429_ _2351_ VGND VGND VPWR VPWR _2430_ sky130_fd_sc_hd__mux2_1
XFILLER_0_5_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5545_ _1666_ _2362_ _2363_ VGND VGND VPWR VPWR _2364_ sky130_fd_sc_hd__o21a_1
XANTENNA__5570__A1 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5476_ _2225_ VGND VGND VPWR VPWR _2299_ sky130_fd_sc_hd__inv_2
XANTENNA__5322__A1 net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4427_ cu.reg_file.reg_b\[0\] net143 _1284_ cu.reg_file.reg_h\[0\] _1486_ VGND VGND
+ VPWR VPWR _1487_ sky130_fd_sc_hd__a221o_1
X_4358_ _1397_ _1395_ _1421_ VGND VGND VPWR VPWR _1422_ sky130_fd_sc_hd__nand3_1
XTAP_260 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4088__B _1050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4289_ _1355_ VGND VGND VPWR VPWR _1356_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__5086__A0 _1187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3309_ _0359_ _2893_ VGND VGND VPWR VPWR _0385_ sky130_fd_sc_hd__nand2_1
XTAP_293 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6028_ clknet_leaf_1_clk _0066_ net164 VGND VGND VPWR VPWR cu.reg_file.reg_e\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__4816__B cu.pc.pc_o\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_68_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5139__S _2069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4116__A2 _1186_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4521__C1 _1323_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3183__A cu.id.cb_opcode_x\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5077__B1 _2951_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4824__A0 cu.pc.pc_o\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5616__A2 _2236_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5049__S _2002_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3660_ _0731_ _0735_ VGND VGND VPWR VPWR _0736_ sky130_fd_sc_hd__and2b_1
XFILLER_0_70_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3591_ cu.reg_file.reg_sp\[4\] _0413_ _0419_ cu.reg_file.reg_h\[4\] _0666_ VGND VGND
+ VPWR VPWR _0667_ sky130_fd_sc_hd__a221o_1
XFILLER_0_42_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5330_ _2205_ _2181_ VGND VGND VPWR VPWR _2206_ sky130_fd_sc_hd__nand2_8
XFILLER_0_2_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5261_ ih.t.timer_max\[29\] _2163_ _2153_ VGND VGND VPWR VPWR _2164_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4212_ _1272_ _1275_ _1276_ _1279_ VGND VGND VPWR VPWR _1280_ sky130_fd_sc_hd__nor4b_2
X_5192_ _1790_ _0352_ _2951_ VGND VGND VPWR VPWR _2114_ sky130_fd_sc_hd__or3b_1
XANTENNA__4917__A _2920_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5068__A0 cu.reg_file.reg_c\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4143_ _0516_ _1212_ VGND VGND VPWR VPWR _1213_ sky130_fd_sc_hd__nor2_4
X_4074_ _0776_ _0805_ _1147_ _0817_ _0777_ VGND VGND VPWR VPWR _1148_ sky130_fd_sc_hd__a221o_1
XANTENNA__3821__A _0895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3025_ ih.t.timer_max\[25\] ih.t.timer_max\[26\] _2762_ VGND VGND VPWR VPWR _2763_
+ sky130_fd_sc_hd__or3_1
XANTENNA__4291__B2 _1354_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4976_ cu.pc.pc_o\[13\] _1939_ cu.pc.pc_o\[14\] VGND VGND VPWR VPWR _1964_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_73_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3927_ _1001_ _1002_ VGND VGND VPWR VPWR _1003_ sky130_fd_sc_hd__nand2_1
XANTENNA__3268__A _0343_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3858_ _0920_ _0796_ VGND VGND VPWR VPWR _0934_ sky130_fd_sc_hd__nand2_1
XFILLER_0_61_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3789_ _0861_ _0864_ VGND VGND VPWR VPWR _0865_ sky130_fd_sc_hd__xnor2_2
X_5528_ net2 _2148_ _2344_ VGND VGND VPWR VPWR _2348_ sky130_fd_sc_hd__mux2_1
XANTENNA__3554__B1 _0499_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5459_ _2286_ VGND VGND VPWR VPWR _0190_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4546__B _1598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4806__B1 _1807_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5658__A net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3178__A _2908_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5534__A1 net125 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5534__B2 net133 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5470__A0 net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5448__S1 _1330_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4830_ _0341_ cu.pc.pc_o\[2\] VGND VGND VPWR VPWR _1830_ sky130_fd_sc_hd__nand2_1
XANTENNA__5287__B _1354_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4761_ _1769_ VGND VGND VPWR VPWR _0004_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4576__A2 _1190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4692_ net212 _1711_ _1713_ VGND VGND VPWR VPWR ih.t.next_count\[19\] sky130_fd_sc_hd__a21oi_1
XFILLER_0_15_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3712_ _0644_ _0733_ VGND VGND VPWR VPWR _0788_ sky130_fd_sc_hd__and2_1
XFILLER_0_28_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3643_ _0652_ _0663_ VGND VGND VPWR VPWR _0719_ sky130_fd_sc_hd__nor2_1
X_5313_ _2196_ VGND VGND VPWR VPWR _0134_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_23_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3574_ cu.reg_file.reg_mem\[5\] _0640_ _0433_ cu.reg_file.reg_a\[5\] VGND VGND VPWR
+ VPWR _0650_ sky130_fd_sc_hd__a22o_1
X_6293_ clknet_leaf_41_clk _0275_ net151 VGND VGND VPWR VPWR cu.id.opcode\[6\] sky130_fd_sc_hd__dfrtp_1
X_5244_ _1661_ _2151_ _2141_ VGND VGND VPWR VPWR _2152_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_11_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold29 ih.t.count\[9\] VGND VGND VPWR VPWR net225 sky130_fd_sc_hd__dlygate4sd3_1
Xhold18 ih.t.count\[22\] VGND VGND VPWR VPWR net214 sky130_fd_sc_hd__dlygate4sd3_1
X_5175_ _2102_ VGND VGND VPWR VPWR _0090_ sky130_fd_sc_hd__clkbuf_1
X_4126_ _0945_ _1195_ VGND VGND VPWR VPWR _1196_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5680__A2_N _1643_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4057_ _1121_ _1130_ _0817_ VGND VGND VPWR VPWR _1131_ sky130_fd_sc_hd__o21a_1
XFILLER_0_36_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3008_ ih.t.timer_max\[0\] ih.t.timer_max\[1\] ih.t.timer_max\[2\] VGND VGND VPWR
+ VPWR _2746_ sky130_fd_sc_hd__or3_1
XFILLER_0_38_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5213__A0 _1052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_411 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4959_ _1945_ _1947_ _1798_ VGND VGND VPWR VPWR _1949_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_46_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3775__B1 _0748_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5516__A1 _1369_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5417__S _2248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1031 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1020 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1064 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1053 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1042 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1097 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1086 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1075 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_458 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3636__A _0545_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4730__A2 _1489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_826 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3290_ _0359_ _2915_ _0316_ _0363_ _0365_ VGND VGND VPWR VPWR _0366_ sky130_fd_sc_hd__o2111a_1
XTAP_859 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5931_ _2674_ VGND VGND VPWR VPWR _0274_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5862_ _2637_ VGND VGND VPWR VPWR _0242_ sky130_fd_sc_hd__clkbuf_1
X_4813_ _1814_ VGND VGND VPWR VPWR _1815_ sky130_fd_sc_hd__buf_4
XFILLER_0_7_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5746__A1 _0986_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5793_ _2576_ _2577_ VGND VGND VPWR VPWR _2578_ sky130_fd_sc_hd__nand2_1
XFILLER_0_56_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4744_ _0338_ _1749_ _1750_ _1752_ VGND VGND VPWR VPWR _1753_ sky130_fd_sc_hd__o22a_1
XFILLER_0_22_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4675_ ih.t.count\[13\] ih.t.count\[14\] _1699_ VGND VGND VPWR VPWR _1702_ sky130_fd_sc_hd__and3_1
X_3626_ _0694_ _0701_ VGND VGND VPWR VPWR _0702_ sky130_fd_sc_hd__nor2_1
X_3557_ _0442_ _0437_ VGND VGND VPWR VPWR _0633_ sky130_fd_sc_hd__nand2_1
X_6276_ clknet_leaf_12_clk _0258_ net178 VGND VGND VPWR VPWR ih.t.timer_max\[16\]
+ sky130_fd_sc_hd__dfrtp_4
X_5227_ _1636_ VGND VGND VPWR VPWR _2136_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3488_ cu.reg_file.reg_a\[7\] _0499_ _0494_ cu.reg_file.reg_mem\[7\] _0563_ VGND
+ VGND VPWR VPWR _0564_ sky130_fd_sc_hd__a221o_1
XANTENNA__4377__A _1415_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4485__A1 cu.reg_file.reg_sp\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4485__B2 cu.id.imm_i\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5158_ _2092_ VGND VGND VPWR VPWR _0083_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5664__A_N _1400_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5089_ _1189_ _1213_ _2035_ VGND VGND VPWR VPWR _2047_ sky130_fd_sc_hd__mux2_1
X_4109_ _1168_ _1179_ _1180_ _1182_ _1023_ VGND VGND VPWR VPWR _1183_ sky130_fd_sc_hd__o221a_1
XFILLER_0_78_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_81_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4840__A cu.pc.pc_o\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4986__S _1814_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3576__A1_N _0576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4287__A _1348_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3279__B1_N _0343_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3279__A2 _0341_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output129_A net129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5520__S0 _1354_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5728__A1 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4460_ _1371_ _1517_ _1518_ _1511_ VGND VGND VPWR VPWR _1519_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__4896__S _1798_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3411_ _0483_ _0486_ VGND VGND VPWR VPWR _0487_ sky130_fd_sc_hd__nor2_2
X_4391_ cu.pc.pc_o\[6\] _1322_ _1315_ cu.reg_file.reg_e\[6\] _1452_ VGND VGND VPWR
+ VPWR _1453_ sky130_fd_sc_hd__a221o_1
X_6130_ clknet_leaf_4_clk _0164_ net171 VGND VGND VPWR VPWR net122 sky130_fd_sc_hd__dfrtp_4
X_3342_ _0407_ _0417_ _0409_ VGND VGND VPWR VPWR _0418_ sky130_fd_sc_hd__nor3b_4
XFILLER_0_0_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_601 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6061_ clknet_leaf_24_clk mc.rw.next_state\[1\] net193 VGND VGND VPWR VPWR mc.rw.state\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__4467__A1 _1296_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_667 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3273_ _2874_ _2927_ VGND VGND VPWR VPWR _0349_ sky130_fd_sc_hd__nor2_1
XTAP_645 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_689 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_678 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5012_ cu.reg_file.reg_a\[4\] _1993_ _1985_ VGND VGND VPWR VPWR _1994_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4925__A _1521_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5914_ _2351_ _2664_ _2665_ net224 VGND VGND VPWR VPWR _0266_ sky130_fd_sc_hd__a22o_1
XFILLER_0_75_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5845_ cu.reg_file.reg_sp\[13\] _2623_ _2538_ VGND VGND VPWR VPWR _2624_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2988_ net2 VGND VGND VPWR VPWR _2727_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5776_ cu.reg_file.reg_sp\[5\] _2535_ VGND VGND VPWR VPWR _2563_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4727_ ih.t.count\[30\] ih.t.count\[31\] _1732_ VGND VGND VPWR VPWR _1737_ sky130_fd_sc_hd__nand3_1
X_4658_ ih.t.count\[8\] _1689_ VGND VGND VPWR VPWR _1691_ sky130_fd_sc_hd__and2_1
XFILLER_0_31_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3609_ _0664_ _0684_ VGND VGND VPWR VPWR _0685_ sky130_fd_sc_hd__nor2_1
X_4589_ _1329_ _1401_ VGND VGND VPWR VPWR _1633_ sky130_fd_sc_hd__nand2_4
X_6259_ clknet_leaf_1_clk _0241_ net153 VGND VGND VPWR VPWR cu.reg_file.reg_sp\[15\]
+ sky130_fd_sc_hd__dfstp_2
XANTENNA__5407__A0 _1052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5958__A1 _2391_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4570__A _0824_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5385__B _2236_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4449__A1 cu.reg_file.reg_sp\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4449__B2 cu.id.imm_i\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4167__D _1089_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4745__A _0296_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3960_ _0781_ _0712_ VGND VGND VPWR VPWR _1035_ sky130_fd_sc_hd__or2_1
XFILLER_0_70_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3891_ _2883_ _0304_ _0966_ _2893_ _0301_ VGND VGND VPWR VPWR _0967_ sky130_fd_sc_hd__o221a_1
XFILLER_0_85_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5630_ net73 _1648_ _2137_ _2274_ VGND VGND VPWR VPWR _2445_ sky130_fd_sc_hd__a31o_1
XFILLER_0_5_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5561_ net78 _1633_ _2375_ _2378_ VGND VGND VPWR VPWR _2379_ sky130_fd_sc_hd__o22a_1
XFILLER_0_60_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4512_ _1566_ _1561_ VGND VGND VPWR VPWR _1568_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5492_ net76 _1633_ _2309_ _2311_ VGND VGND VPWR VPWR _2312_ sky130_fd_sc_hd__o22a_1
XFILLER_0_13_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4443_ _1382_ _1498_ _1499_ _1502_ VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__a31o_2
XFILLER_0_13_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4374_ _1435_ _1436_ VGND VGND VPWR VPWR _1437_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6113_ clknet_leaf_27_clk _0147_ net186 VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__dfrtp_1
X_3325_ _0395_ _0400_ VGND VGND VPWR VPWR _0401_ sky130_fd_sc_hd__or2_2
XTAP_420 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6044_ clknet_leaf_3_clk _0082_ net156 VGND VGND VPWR VPWR cu.reg_file.reg_l\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_3256_ _0330_ _0331_ _2932_ VGND VGND VPWR VPWR _0332_ sky130_fd_sc_hd__a21oi_1
XTAP_453 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_486 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3187_ _2901_ _2923_ _2874_ VGND VGND VPWR VPWR _2924_ sky130_fd_sc_hd__or3b_2
XFILLER_0_21_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_431 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5828_ _1222_ _2608_ _2545_ VGND VGND VPWR VPWR _2609_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5759_ cu.reg_file.reg_sp\[3\] _2534_ VGND VGND VPWR VPWR _2548_ sky130_fd_sc_hd__nor2_1
XANTENNA__4128__B1 _0779_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3453__B _0528_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_67_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3575__D1 _0576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3590__A1 cu.reg_file.reg_d\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5335__S _2206_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3590__B2 cu.reg_file.reg_b\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output73_A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3110_ _2834_ _2843_ _2844_ _2847_ VGND VGND VPWR VPWR _2848_ sky130_fd_sc_hd__or4_1
XFILLER_0_65_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4090_ _1129_ _1163_ VGND VGND VPWR VPWR _1164_ sky130_fd_sc_hd__xnor2_1
XANTENNA__5095__A1 _1624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3041_ _2763_ _2777_ ih.t.count\[26\] VGND VGND VPWR VPWR _2779_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_81_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4992_ _1263_ _1975_ _1794_ VGND VGND VPWR VPWR _1979_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3943_ _0971_ _0986_ VGND VGND VPWR VPWR _1019_ sky130_fd_sc_hd__or2_2
XFILLER_0_14_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3874_ _0856_ _0908_ VGND VGND VPWR VPWR _0950_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5613_ _2425_ _2426_ _2428_ _1641_ VGND VGND VPWR VPWR _2429_ sky130_fd_sc_hd__o22a_4
XFILLER_0_5_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_26_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3566__D1 _0576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5544_ ih.t.timer_max\[17\] _2151_ _2319_ ih.t.timer_max\[1\] _1661_ VGND VGND VPWR
+ VPWR _2363_ sky130_fd_sc_hd__a221o_1
XANTENNA__5570__A2 _1648_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5475_ _2298_ VGND VGND VPWR VPWR _0194_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3581__A1 cu.reg_file.reg_d\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4426_ cu.reg_file.reg_d\[0\] _1282_ _1286_ cu.reg_file.reg_sp\[8\] VGND VGND VPWR
+ VPWR _1486_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4357_ _1419_ _1420_ VGND VGND VPWR VPWR _1421_ sky130_fd_sc_hd__nand2_1
XTAP_250 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3704__D _0779_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4288_ _2698_ mc.rw.state\[1\] mc.rw.state\[0\] VGND VGND VPWR VPWR _1355_ sky130_fd_sc_hd__or3_1
XANTENNA__5086__A1 _1222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3308_ _0317_ _0379_ _0383_ VGND VGND VPWR VPWR _0384_ sky130_fd_sc_hd__or3_2
XTAP_283 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_261 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6027_ clknet_leaf_1_clk _0065_ net164 VGND VGND VPWR VPWR cu.reg_file.reg_e\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_294 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3239_ _0310_ _0311_ _0312_ _0314_ VGND VGND VPWR VPWR _0315_ sky130_fd_sc_hd__or4b_4
XFILLER_0_68_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5561__A2 _1633_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3572__B2 cu.reg_file.reg_h\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3572__A1 cu.reg_file.reg_sp\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3464__A cu.reg_file.reg_a\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6197__D net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4521__B1 _1343_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4994__S _1808_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5077__A1 _2035_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output111_A net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3639__A _0587_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_264 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_70_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3590_ cu.reg_file.reg_d\[4\] _0415_ _0432_ cu.reg_file.reg_b\[4\] VGND VGND VPWR
+ VPWR _0666_ sky130_fd_sc_hd__a22o_1
XFILLER_0_2_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3563__A1 cu.reg_file.reg_c\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5260_ _1144_ _1209_ _1666_ VGND VGND VPWR VPWR _2163_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3315__A1 _2936_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4211_ _2912_ _0583_ _1277_ _1278_ VGND VGND VPWR VPWR _1279_ sky130_fd_sc_hd__a31o_1
X_5191_ _2113_ VGND VGND VPWR VPWR _0095_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4917__B cu.pc.pc_o\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5068__A1 _1193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4142_ _0956_ _1205_ _1206_ _0957_ _1211_ VGND VGND VPWR VPWR _1212_ sky130_fd_sc_hd__o221a_1
X_4073_ _0811_ _1146_ VGND VGND VPWR VPWR _1147_ sky130_fd_sc_hd__nand2_1
X_3024_ ih.t.timer_max\[24\] _2761_ VGND VGND VPWR VPWR _2762_ sky130_fd_sc_hd__or2_2
XFILLER_0_93_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4975_ cu.pc.pc_o\[14\] cu.pc.pc_o\[13\] _1939_ VGND VGND VPWR VPWR _1963_ sky130_fd_sc_hd__and3_1
XANTENNA__4579__B1 _1624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3926_ _0981_ _0998_ VGND VGND VPWR VPWR _1002_ sky130_fd_sc_hd__nand2_1
XANTENNA__3549__A _0498_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6107__RESET_B net195 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3857_ _0865_ _0925_ VGND VGND VPWR VPWR _0933_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_41_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3788_ cu.reg_file.reg_mem\[12\] _0640_ _0862_ _0863_ VGND VGND VPWR VPWR _0864_
+ sky130_fd_sc_hd__a211oi_2
X_5527_ net2 _2345_ _2346_ VGND VGND VPWR VPWR _2347_ sky130_fd_sc_hd__a21o_1
XANTENNA__3554__A1 cu.reg_file.reg_b\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3554__B2 cu.reg_file.reg_a\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3284__A _0340_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5458_ net60 _2085_ _2285_ VGND VGND VPWR VPWR _2286_ sky130_fd_sc_hd__mux2_1
X_5389_ _2239_ VGND VGND VPWR VPWR _0167_ sky130_fd_sc_hd__clkbuf_1
X_4409_ cu.reg_file.reg_sp\[7\] _0993_ _1344_ cu.id.cb_opcode_x\[1\] _1324_ VGND VGND
+ VPWR VPWR _1470_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4806__A1 _2935_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4843__A cu.id.cb_opcode_y\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4562__B _1614_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3793__A1 cu.pc.pc_o\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5534__A2 _2236_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3922__A _0986_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output36_A net36 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5470__A1 _2085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_17 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4430__C1 _1489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4760_ net235 _1768_ VGND VGND VPWR VPWR _1769_ sky130_fd_sc_hd__or2_1
X_4691_ ih.t.count\[19\] _1711_ _1670_ VGND VGND VPWR VPWR _1713_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_15_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3711_ _0759_ _0763_ _0783_ _0785_ _0786_ VGND VGND VPWR VPWR _0787_ sky130_fd_sc_hd__a311o_2
XANTENNA__3784__B2 cu.reg_file.reg_mem\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3784__A1 cu.reg_file.reg_a\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3642_ _0702_ _0716_ _0717_ VGND VGND VPWR VPWR _0718_ sky130_fd_sc_hd__o21ai_2
X_5312_ _0619_ net92 _2195_ VGND VGND VPWR VPWR _2196_ sky130_fd_sc_hd__mux2_1
XFILLER_0_51_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3573_ cu.reg_file.reg_c\[5\] _0427_ _0430_ cu.reg_file.reg_e\[5\] VGND VGND VPWR
+ VPWR _0649_ sky130_fd_sc_hd__a22o_1
X_6292_ clknet_leaf_41_clk _0274_ net151 VGND VGND VPWR VPWR cu.id.alu_opcode\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_5243_ _2150_ VGND VGND VPWR VPWR _2151_ sky130_fd_sc_hd__buf_2
Xhold19 ih.t.count\[25\] VGND VGND VPWR VPWR net215 sky130_fd_sc_hd__dlygate4sd3_1
X_5174_ _1647_ _2101_ VGND VGND VPWR VPWR _2102_ sky130_fd_sc_hd__and2_1
X_4125_ _0942_ _0943_ _0944_ VGND VGND VPWR VPWR _1195_ sky130_fd_sc_hd__a21oi_1
X_4056_ _0804_ _0811_ VGND VGND VPWR VPWR _1130_ sky130_fd_sc_hd__and2_1
X_3007_ _2736_ _2737_ _2738_ _2744_ VGND VGND VPWR VPWR _2745_ sky130_fd_sc_hd__or4_4
XANTENNA__5759__A cu.reg_file.reg_sp\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4958_ _1945_ _1947_ VGND VGND VPWR VPWR _1948_ sky130_fd_sc_hd__or2_1
X_4889_ cu.pc.pc_o\[7\] _1872_ VGND VGND VPWR VPWR _1884_ sky130_fd_sc_hd__xor2_1
XFILLER_0_46_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3909_ _0310_ _0328_ _0740_ _0984_ VGND VGND VPWR VPWR _0985_ sky130_fd_sc_hd__nor4_1
XANTENNA__3775__A1 cu.reg_file.reg_sp\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3775__B2 cu.reg_file.reg_h\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5494__A _1400_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4724__B1 _1670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_394 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5452__A1 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5452__B2 net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1021 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1010 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1065 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1054 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1043 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1032 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1098 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1087 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1076 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3636__B _0598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3518__A1 _0340_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_40_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_816 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5343__S _2206_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_849 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5930_ _2936_ _2448_ _2668_ VGND VGND VPWR VPWR _2674_ sky130_fd_sc_hd__mux2_1
X_5861_ _2144_ ih.t.timer_max\[8\] _2636_ VGND VGND VPWR VPWR _2637_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4812_ _2948_ _1808_ _1813_ _1484_ VGND VGND VPWR VPWR _1814_ sky130_fd_sc_hd__a22o_4
X_5792_ cu.reg_file.reg_sp\[7\] _2535_ VGND VGND VPWR VPWR _2577_ sky130_fd_sc_hd__nand2_1
XANTENNA__5746__A2 _2532_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4743_ _2907_ _0311_ _0379_ _1751_ VGND VGND VPWR VPWR _1752_ sky130_fd_sc_hd__or4_1
XFILLER_0_7_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_22_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4674_ net223 _1699_ _1701_ VGND VGND VPWR VPWR ih.t.next_count\[13\] sky130_fd_sc_hd__a21oi_1
XANTENNA__5708__A2_N _1643_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3625_ _0576_ _0695_ _0697_ _0700_ VGND VGND VPWR VPWR _0701_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_31_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3556_ _0623_ _0627_ _0630_ _0631_ VGND VGND VPWR VPWR _0632_ sky130_fd_sc_hd__o31a_4
X_6275_ clknet_leaf_12_clk _0257_ net178 VGND VGND VPWR VPWR ih.t.timer_max\[7\] sky130_fd_sc_hd__dfrtp_4
X_5226_ _2135_ VGND VGND VPWR VPWR _0108_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3487_ cu.pc.pc_o\[7\] _0501_ _0498_ cu.alu_f\[7\] _0504_ VGND VGND VPWR VPWR _0563_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4377__B _1434_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5682__B2 ih.t.timer_max\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5157_ cu.reg_file.reg_l\[3\] _1187_ _2088_ VGND VGND VPWR VPWR _2092_ sky130_fd_sc_hd__mux2_1
X_5088_ _2046_ VGND VGND VPWR VPWR _0059_ sky130_fd_sc_hd__clkbuf_1
X_4108_ _0996_ _1003_ _1181_ _1010_ VGND VGND VPWR VPWR _1182_ sky130_fd_sc_hd__or4b_2
X_4039_ _1060_ _0599_ VGND VGND VPWR VPWR _1113_ sky130_fd_sc_hd__nand2_1
XPHY_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4173__A1 _0892_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5520__S1 _1330_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4936__A0 _1521_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3647__A _0293_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3410_ net148 _0460_ _0462_ VGND VGND VPWR VPWR _0486_ sky130_fd_sc_hd__a21oi_4
X_4390_ cu.reg_file.reg_sp\[6\] _0993_ _1344_ _0387_ _1324_ VGND VGND VPWR VPWR _1452_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_21_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3341_ _0412_ _0405_ VGND VGND VPWR VPWR _0417_ sky130_fd_sc_hd__or2_4
XANTENNA__5113__A0 cu.reg_file.reg_e\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_602 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6060_ clknet_leaf_23_clk mc.rw.next_state\[0\] net193 VGND VGND VPWR VPWR mc.rw.state\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_668 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3272_ _2942_ _0345_ _0347_ _0336_ VGND VGND VPWR VPWR _0348_ sky130_fd_sc_hd__o31a_1
XTAP_635 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_679 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5011_ _1189_ _1213_ _0368_ VGND VGND VPWR VPWR _1993_ sky130_fd_sc_hd__mux2_1
XFILLER_0_84_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3427__B1 _0293_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5913_ _2947_ _1482_ _2664_ VGND VGND VPWR VPWR _2665_ sky130_fd_sc_hd__a21o_1
XANTENNA__4941__A _2920_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5844_ _1209_ _2622_ _2115_ VGND VGND VPWR VPWR _2623_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5248__S _1667_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2987_ _2721_ ih.ih.ih.prev_data\[9\] _2722_ ih.ih.ih.prev_data\[14\] _2725_ VGND
+ VGND VPWR VPWR _2726_ sky130_fd_sc_hd__o221a_1
XFILLER_0_16_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5775_ cu.reg_file.reg_sp\[5\] _2535_ VGND VGND VPWR VPWR _2562_ sky130_fd_sc_hd__or2_1
XFILLER_0_44_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4726_ ih.t.count\[30\] _1732_ ih.t.count\[31\] VGND VGND VPWR VPWR _1736_ sky130_fd_sc_hd__a21o_1
X_4657_ _1689_ _1690_ VGND VGND VPWR VPWR ih.t.next_count\[7\] sky130_fd_sc_hd__nor2_1
XFILLER_0_16_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5352__A0 _1075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3608_ _0682_ _0683_ VGND VGND VPWR VPWR _0684_ sky130_fd_sc_hd__nor2_2
X_4588_ mc.cl.cmp_o _1631_ VGND VGND VPWR VPWR _1632_ sky130_fd_sc_hd__or2b_4
XFILLER_0_12_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3539_ _0572_ _0573_ _0608_ _0613_ _0614_ VGND VGND VPWR VPWR _0615_ sky130_fd_sc_hd__o2111a_1
XANTENNA__3902__B2 _0359_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6258_ clknet_leaf_3_clk _0240_ net156 VGND VGND VPWR VPWR cu.reg_file.reg_sp\[14\]
+ sky130_fd_sc_hd__dfstp_2
X_6189_ clknet_leaf_22_clk _0222_ net191 VGND VGND VPWR VPWR mc.cl.next_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_5209_ _1364_ _2125_ VGND VGND VPWR VPWR _2126_ sky130_fd_sc_hd__or2_1
XANTENNA__3666__B1 _0741_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5407__A1 net133 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4997__S _0368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5343__A0 _1194_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5894__A1 _1667_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5646__A1 _1665_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4449__A2 _0993_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4909__B1 _1798_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3890_ _2917_ _0965_ VGND VGND VPWR VPWR _0966_ sky130_fd_sc_hd__nand2_1
XFILLER_0_72_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5582__B1 _2204_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5560_ net110 _2147_ _2225_ net118 _2377_ VGND VGND VPWR VPWR _2378_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4385__B2 cu.reg_file.reg_l\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4511_ _1566_ _1561_ VGND VGND VPWR VPWR _1567_ sky130_fd_sc_hd__nand2_1
X_5491_ net100 _2205_ _2310_ _2257_ VGND VGND VPWR VPWR _2311_ sky130_fd_sc_hd__a211o_1
XFILLER_0_41_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4442_ _1496_ _1500_ _1501_ _1371_ VGND VGND VPWR VPWR _1502_ sky130_fd_sc_hd__a22o_1
XANTENNA__5592__A _1649_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4373_ _1396_ _1434_ VGND VGND VPWR VPWR _1436_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6112_ clknet_leaf_7_clk _0146_ net167 VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__dfrtp_1
XANTENNA__4001__A _1074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3324_ _2950_ _0399_ VGND VGND VPWR VPWR _0400_ sky130_fd_sc_hd__nand2_2
XFILLER_0_0_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_410 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5637__A1 net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6043_ clknet_leaf_4_clk _0081_ net170 VGND VGND VPWR VPWR cu.reg_file.reg_l\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_3255_ cu.id.opcode\[0\] cu.id.alu_opcode\[3\] cu.id.alu_opcode\[1\] _2892_ VGND
+ VGND VPWR VPWR _0331_ sky130_fd_sc_hd__or4bb_1
XTAP_443 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_487 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3186_ _2894_ VGND VGND VPWR VPWR _2923_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5767__A cu.reg_file.reg_sp\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5827_ _2606_ _2607_ VGND VGND VPWR VPWR _2608_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_36_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5758_ _2547_ VGND VGND VPWR VPWR _0228_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_44_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4709_ ih.t.count\[25\] _1723_ _1670_ VGND VGND VPWR VPWR _1725_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_32_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3584__C1 _0536_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5689_ net3 _1650_ _2488_ _2498_ VGND VGND VPWR VPWR _0208_ sky130_fd_sc_hd__a31o_1
XANTENNA__4300__A1 cu.pc.pc_o\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4565__B _1579_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5316__A0 _1075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4119__B2 _1190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3590__A2 _0415_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5619__A1 net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5619__B2 _1401_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output66_A net66 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3040_ ih.t.count\[26\] _2763_ _2777_ VGND VGND VPWR VPWR _2778_ sky130_fd_sc_hd__and3_1
XFILLER_0_58_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4991_ cu.pc.pc_o\[15\] _1977_ VGND VGND VPWR VPWR _1978_ sky130_fd_sc_hd__xor2_1
X_3942_ _1000_ _1008_ VGND VGND VPWR VPWR _1018_ sky130_fd_sc_hd__nand2_1
XFILLER_0_18_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3802__B1 _0741_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3873_ _0845_ _0910_ VGND VGND VPWR VPWR _0949_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5612_ _1649_ _2427_ VGND VGND VPWR VPWR _2428_ sky130_fd_sc_hd__and2_1
XFILLER_0_45_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5543_ _1400_ _2361_ VGND VGND VPWR VPWR _2362_ sky130_fd_sc_hd__and2b_1
XFILLER_0_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5474_ net64 _2085_ _2297_ VGND VGND VPWR VPWR _2298_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3581__A2 _0492_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4425_ _1269_ _1484_ VGND VGND VPWR VPWR _1485_ sky130_fd_sc_hd__or2_4
X_4356_ _1332_ _1417_ VGND VGND VPWR VPWR _1420_ sky130_fd_sc_hd__nand2_1
X_3307_ _2905_ _0380_ _0381_ _0382_ VGND VGND VPWR VPWR _0383_ sky130_fd_sc_hd__or4_1
XTAP_251 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4287_ _1348_ VGND VGND VPWR VPWR _1354_ sky130_fd_sc_hd__buf_4
XTAP_284 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_262 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6026_ clknet_leaf_1_clk _0064_ net153 VGND VGND VPWR VPWR cu.reg_file.reg_e\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_295 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3238_ _2910_ _0313_ _0305_ VGND VGND VPWR VPWR _0314_ sky130_fd_sc_hd__or3_1
X_3169_ _2887_ _2891_ _2905_ VGND VGND VPWR VPWR _2906_ sky130_fd_sc_hd__or3_1
XFILLER_0_49_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4349__A1 cu.pc.pc_o\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3464__B _0499_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4521__A1 cu.reg_file.reg_sp\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3911__C _0379_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_51_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3639__B _0710_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_27_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_82_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3655__A _0566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4210_ _2877_ _0336_ _0436_ _0293_ VGND VGND VPWR VPWR _1278_ sky130_fd_sc_hd__a31o_1
X_5190_ _2111_ _2112_ VGND VGND VPWR VPWR _2113_ sky130_fd_sc_hd__and2_1
XANTENNA__5081__S _2039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4141_ _0817_ _0942_ _1210_ _0933_ VGND VGND VPWR VPWR _1211_ sky130_fd_sc_hd__a22oi_1
XANTENNA__3079__A1 ih.t.timer_max\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4072_ _0808_ _0810_ _0805_ VGND VGND VPWR VPWR _1146_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_92_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3023_ ih.t.timer_max\[22\] ih.t.timer_max\[23\] _2760_ VGND VGND VPWR VPWR _2761_
+ sky130_fd_sc_hd__or3_2
XFILLER_0_78_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4974_ _1962_ VGND VGND VPWR VPWR _0029_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4579__A1 _2702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4579__B2 _2697_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3925_ _0998_ _1000_ VGND VGND VPWR VPWR _1001_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5528__A0 net2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3856_ _0829_ _0919_ _0931_ VGND VGND VPWR VPWR _0932_ sky130_fd_sc_hd__a21o_1
XFILLER_0_81_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3787_ cu.reg_file.reg_b\[4\] _0426_ _0429_ cu.reg_file.reg_d\[4\] VGND VGND VPWR
+ VPWR _0863_ sky130_fd_sc_hd__a22o_1
X_5526_ net16 _2179_ _2279_ ih.input_handler_enable VGND VGND VPWR VPWR _2346_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3554__A2 _0502_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5457_ _1633_ _2284_ VGND VGND VPWR VPWR _2285_ sky130_fd_sc_hd__nor2_1
XANTENNA__4503__A1 cu.pc.pc_o\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4408_ cu.reg_file.reg_l\[7\] _1317_ VGND VGND VPWR VPWR _1469_ sky130_fd_sc_hd__and2_1
X_5388_ _1052_ net125 _2237_ VGND VGND VPWR VPWR _2239_ sky130_fd_sc_hd__mux2_1
XANTENNA__5700__B1 cu.reg_file.reg_mem\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4503__B2 cu.reg_file.reg_d\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4339_ _1393_ _1401_ VGND VGND VPWR VPWR _1404_ sky130_fd_sc_hd__and2b_1
XFILLER_0_5_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6009_ clknet_leaf_31_clk _0047_ net185 VGND VGND VPWR VPWR cu.reg_file.reg_b\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__4806__A2 _1256_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4843__B cu.pc.pc_o\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_37_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4990__A1 _1233_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3793__A2 _0740_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3710_ _0701_ _0694_ VGND VGND VPWR VPWR _0786_ sky130_fd_sc_hd__and2b_1
XFILLER_0_28_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4690_ _1711_ _1712_ VGND VGND VPWR VPWR ih.t.next_count\[18\] sky130_fd_sc_hd__nor2_1
XFILLER_0_43_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3641_ _0694_ _0701_ VGND VGND VPWR VPWR _0717_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5930__A0 _2936_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3572_ cu.reg_file.reg_sp\[5\] _0636_ _0419_ cu.reg_file.reg_h\[5\] _0647_ VGND VGND
+ VPWR VPWR _0648_ sky130_fd_sc_hd__a221o_1
XANTENNA__6240__RESET_B net194 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5311_ _2181_ _2194_ VGND VGND VPWR VPWR _2195_ sky130_fd_sc_hd__nand2_8
XFILLER_0_51_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6291_ clknet_leaf_41_clk _0273_ net151 VGND VGND VPWR VPWR cu.id.alu_opcode\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_5242_ _2145_ _2149_ VGND VGND VPWR VPWR _2150_ sky130_fd_sc_hd__or2_2
XANTENNA__4497__B1 _1286_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5173_ mc.cl.next_data\[10\] net20 mc.count VGND VGND VPWR VPWR _2101_ sky130_fd_sc_hd__mux2_1
X_4124_ _1193_ VGND VGND VPWR VPWR _1194_ sky130_fd_sc_hd__buf_4
Xinput1 interrupt_gpio_in VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__dlymetal6s2s_1
X_4055_ _1127_ _1128_ VGND VGND VPWR VPWR _1129_ sky130_fd_sc_hd__nor2_1
XFILLER_0_78_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3006_ _2739_ net33 ih.gpio_interrupt_mask\[6\] _2742_ _2743_ VGND VGND VPWR VPWR
+ _2744_ sky130_fd_sc_hd__a311o_1
XANTENNA__5749__A0 cu.reg_file.reg_sp\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4957_ _1920_ _1922_ _1932_ _1946_ _1921_ VGND VGND VPWR VPWR _1947_ sky130_fd_sc_hd__o311a_1
XFILLER_0_19_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5775__A cu.reg_file.reg_sp\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4888_ _1883_ VGND VGND VPWR VPWR _0022_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_46_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3908_ _2918_ _0966_ VGND VGND VPWR VPWR _0984_ sky130_fd_sc_hd__nand2_1
XFILLER_0_19_479 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_61_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3839_ _0777_ _0914_ VGND VGND VPWR VPWR _0915_ sky130_fd_sc_hd__nand2_1
XANTENNA__3295__A _2950_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5509_ _2169_ _2312_ _2328_ _2136_ VGND VGND VPWR VPWR _2329_ sky130_fd_sc_hd__o211a_1
XFILLER_0_42_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4854__A _0374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1022 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1011 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1000 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1055 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1044 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1033 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1099 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1088 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1077 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1066 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_37_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5912__B1 _1484_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_817 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_57_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_839 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5860_ _1667_ _2194_ _2635_ VGND VGND VPWR VPWR _2636_ sky130_fd_sc_hd__o21ai_4
X_4811_ _1301_ _1775_ _1811_ _1812_ VGND VGND VPWR VPWR _1813_ sky130_fd_sc_hd__a211o_1
X_5791_ cu.reg_file.reg_sp\[7\] _2535_ VGND VGND VPWR VPWR _2576_ sky130_fd_sc_hd__or2_1
XFILLER_0_7_148 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4742_ _0314_ _1741_ VGND VGND VPWR VPWR _1751_ sky130_fd_sc_hd__nor2_1
X_4673_ ih.t.count\[13\] _1699_ _1670_ VGND VGND VPWR VPWR _1701_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_83_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3624_ cu.reg_file.reg_l\[3\] _0422_ _0698_ _0699_ _0440_ VGND VGND VPWR VPWR _0700_
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_43_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3555_ _0295_ _2921_ _0536_ VGND VGND VPWR VPWR _0631_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_24_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6274_ clknet_leaf_13_clk _0256_ net181 VGND VGND VPWR VPWR ih.t.timer_max\[6\] sky130_fd_sc_hd__dfstp_1
X_3486_ cu.reg_file.reg_h\[7\] _0495_ _0539_ cu.reg_file.reg_sp\[7\] _0561_ VGND VGND
+ VPWR VPWR _0562_ sky130_fd_sc_hd__a221o_1
X_5225_ _1261_ ih.gpio_interrupt_mask\[7\] _2127_ VGND VGND VPWR VPWR _2135_ sky130_fd_sc_hd__mux2_1
X_5156_ _2091_ VGND VGND VPWR VPWR _0082_ sky130_fd_sc_hd__clkbuf_1
X_5087_ cu.reg_file.reg_d\[3\] _2045_ _2039_ VGND VGND VPWR VPWR _2046_ sky130_fd_sc_hd__mux2_1
X_4107_ _1018_ _1019_ _0395_ VGND VGND VPWR VPWR _1181_ sky130_fd_sc_hd__a21oi_1
X_4038_ _0588_ _0610_ VGND VGND VPWR VPWR _1112_ sky130_fd_sc_hd__or2_1
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5989_ clknet_leaf_28_clk _0027_ net188 VGND VGND VPWR VPWR cu.pc.pc_o\[11\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_47_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4584__A _1511_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_84_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5189__A1 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5354__S _2215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output96_A net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3340_ cu.reg_file.reg_sp\[0\] _0413_ _0415_ cu.reg_file.reg_d\[0\] VGND VGND VPWR
+ VPWR _0416_ sky130_fd_sc_hd__a22o_1
XTAP_603 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5113__A1 _1191_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_625 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3271_ _0301_ _0346_ _0316_ VGND VGND VPWR VPWR _0347_ sky130_fd_sc_hd__o21ai_1
X_5010_ _1992_ VGND VGND VPWR VPWR _0035_ sky130_fd_sc_hd__clkbuf_1
XTAP_636 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_669 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3675__A1 cu.reg_file.reg_mem\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5912_ _2663_ _1644_ _1484_ VGND VGND VPWR VPWR _2664_ sky130_fd_sc_hd__o21a_1
XANTENNA__4941__B cu.pc.pc_o\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5843_ _2620_ _2621_ VGND VGND VPWR VPWR _2622_ sky130_fd_sc_hd__xnor2_1
X_2986_ _2723_ ih.ih.ih.prev_data\[5\] _2724_ ih.ih.ih.prev_data\[10\] VGND VGND VPWR
+ VPWR _2725_ sky130_fd_sc_hd__o22a_1
X_5774_ _2561_ VGND VGND VPWR VPWR _0230_ sky130_fd_sc_hd__clkbuf_1
X_4725_ net218 _1732_ _1735_ VGND VGND VPWR VPWR ih.t.next_count\[30\] sky130_fd_sc_hd__a21oi_1
XFILLER_0_44_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4656_ net226 _1686_ _1687_ VGND VGND VPWR VPWR _1690_ sky130_fd_sc_hd__o21ai_1
X_4587_ _1374_ _1625_ _1630_ _1417_ VGND VGND VPWR VPWR _1631_ sky130_fd_sc_hd__a211o_1
XANTENNA__5352__A1 net110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3607_ _0681_ _0671_ VGND VGND VPWR VPWR _0683_ sky130_fd_sc_hd__and2b_1
XFILLER_0_31_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3538_ _0549_ _0555_ VGND VGND VPWR VPWR _0614_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3469_ _0537_ _0538_ _0543_ _0544_ VGND VGND VPWR VPWR _0545_ sky130_fd_sc_hd__o31a_4
X_6257_ clknet_leaf_1_clk _0239_ net153 VGND VGND VPWR VPWR cu.reg_file.reg_sp\[13\]
+ sky130_fd_sc_hd__dfstp_2
X_6188_ clknet_leaf_21_clk _0221_ net191 VGND VGND VPWR VPWR mc.cl.next_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_5208_ _1634_ VGND VGND VPWR VPWR _2125_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__3666__A1 cu.reg_file.reg_d\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5139_ _2079_ cu.reg_file.reg_h\[5\] _2069_ VGND VGND VPWR VPWR _2080_ sky130_fd_sc_hd__mux2_1
XANTENNA__3666__B2 cu.reg_file.reg_h\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3748__A _0384_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5040__A0 _1189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5591__A1 net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5591__B2 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5343__A1 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5894__A2 _2205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_19_clk_A clknet_2_3__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output134_A net134 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5031__A0 _1051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4510_ _1517_ _1530_ _1545_ VGND VGND VPWR VPWR _1566_ sky130_fd_sc_hd__and3_1
XFILLER_0_79_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5490_ net108 _2146_ _2193_ net92 VGND VGND VPWR VPWR _2310_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4441_ _1478_ _1496_ VGND VGND VPWR VPWR _1501_ sky130_fd_sc_hd__nor2_1
XANTENNA__5084__S _2039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4372_ _1396_ _1434_ VGND VGND VPWR VPWR _1435_ sky130_fd_sc_hd__or2_1
X_6111_ clknet_leaf_30_clk _0145_ net187 VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__dfrtp_4
XTAP_400 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5098__A0 _1110_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3323_ _2893_ _0386_ _0324_ _0398_ VGND VGND VPWR VPWR _0399_ sky130_fd_sc_hd__a31o_2
XFILLER_0_0_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_411 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_95_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5637__A2 _2194_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3254_ _2894_ _2884_ VGND VGND VPWR VPWR _0330_ sky130_fd_sc_hd__or2b_1
XTAP_444 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3648__A1 cu.reg_file.reg_d\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6042_ clknet_leaf_3_clk _0080_ net156 VGND VGND VPWR VPWR cu.reg_file.reg_l\[0\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_477 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3185_ _2920_ _2921_ VGND VGND VPWR VPWR _2922_ sky130_fd_sc_hd__nor2_1
XFILLER_0_95_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5826_ _2597_ _2600_ _2598_ VGND VGND VPWR VPWR _2607_ sky130_fd_sc_hd__a21bo_1
X_2969_ _2708_ VGND VGND VPWR VPWR mc.cc.enable sky130_fd_sc_hd__inv_2
XFILLER_0_60_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5757_ cu.reg_file.reg_sp\[2\] _2546_ _2539_ VGND VGND VPWR VPWR _2547_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4708_ _1723_ _1724_ VGND VGND VPWR VPWR ih.t.next_count\[24\] sky130_fd_sc_hd__nor2_1
XANTENNA__5783__A cu.reg_file.reg_sp\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3584__B1 _0495_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5688_ _2497_ _1643_ cu.reg_file.reg_mem\[10\] _1646_ VGND VGND VPWR VPWR _2498_
+ sky130_fd_sc_hd__a2bb2o_1
X_4639_ _1672_ _1676_ _1677_ VGND VGND VPWR VPWR _1678_ sky130_fd_sc_hd__and3_1
XANTENNA__3336__B1 cu.id.starting_int_service VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6309_ clknet_leaf_18_clk _0291_ net184 VGND VGND VPWR VPWR cu.id.imm_i\[14\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__5089__A0 _1189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3909__C _0740_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5316__A1 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4119__A2 _1186_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3327__B1 _2877_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5619__A2 _2205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4827__B1 cu.pc.pc_o\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4990_ _1233_ _1969_ _1976_ VGND VGND VPWR VPWR _1977_ sky130_fd_sc_hd__o21ba_1
XFILLER_0_58_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3941_ _1013_ _1014_ VGND VGND VPWR VPWR _1017_ sky130_fd_sc_hd__and2b_1
XFILLER_0_14_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3802__A1 cu.reg_file.reg_d\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3802__B2 cu.reg_file.reg_h\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3872_ _0833_ _0912_ VGND VGND VPWR VPWR _0948_ sky130_fd_sc_hd__xor2_1
X_5611_ net12 _2345_ _2369_ net5 VGND VGND VPWR VPWR _2427_ sky130_fd_sc_hd__a22o_1
X_5542_ ih.t.timer_max\[9\] _2193_ _2314_ ih.t.timer_max\[1\] _2360_ VGND VGND VPWR
+ VPWR _2361_ sky130_fd_sc_hd__a221o_1
XFILLER_0_26_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5473_ _2296_ _2284_ VGND VGND VPWR VPWR _2297_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4424_ _1482_ _1483_ VGND VGND VPWR VPWR _1484_ sky130_fd_sc_hd__nand2_2
XFILLER_0_41_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4355_ _1396_ _1415_ VGND VGND VPWR VPWR _1419_ sky130_fd_sc_hd__nand2_1
XFILLER_0_39_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3306_ _2903_ _0313_ _0329_ VGND VGND VPWR VPWR _0382_ sky130_fd_sc_hd__o21bai_2
XTAP_241 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4286_ mc.rw.state\[1\] mc.rw.state\[0\] _2698_ VGND VGND VPWR VPWR _1353_ sky130_fd_sc_hd__o21a_2
XTAP_274 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_252 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6025_ clknet_leaf_30_clk _0063_ net183 VGND VGND VPWR VPWR cu.reg_file.reg_d\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_3237_ _2892_ cu.id.opcode\[0\] VGND VGND VPWR VPWR _0313_ sky130_fd_sc_hd__or2_2
XTAP_296 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3168_ _2893_ _2896_ _2904_ VGND VGND VPWR VPWR _2905_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_68_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3099_ ih.t.count\[0\] _2836_ VGND VGND VPWR VPWR _2837_ sky130_fd_sc_hd__nor2_1
XANTENNA__5988__RESET_B net188 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_211 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5809_ _2590_ _2591_ VGND VGND VPWR VPWR _2592_ sky130_fd_sc_hd__nand2_1
XFILLER_0_32_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4285__A1 _1335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5482__A0 net66 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4592__A _1434_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5644__A_N _1400_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3001__A net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3796__B1 _0748_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5537__A1 net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5537__B2 _1401_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3936__A _0296_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5362__S _2215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4140_ _0817_ _0941_ _0776_ VGND VGND VPWR VPWR _1210_ sky130_fd_sc_hd__a21o_1
X_4071_ _0765_ _0766_ VGND VGND VPWR VPWR _1145_ sky130_fd_sc_hd__or2_1
XFILLER_0_92_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3022_ ih.t.timer_max\[21\] _2759_ VGND VGND VPWR VPWR _2760_ sky130_fd_sc_hd__or2_2
XANTENNA__5598__A net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5225__A0 _1261_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_58_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4579__A2 _1194_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4973_ cu.pc.pc_o\[13\] _1961_ _1814_ VGND VGND VPWR VPWR _1962_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3924_ _0976_ _0999_ VGND VGND VPWR VPWR _1000_ sky130_fd_sc_hd__nor2_1
XANTENNA__3787__B1 _0429_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3855_ _0829_ _0919_ _0930_ VGND VGND VPWR VPWR _0931_ sky130_fd_sc_hd__o21a_1
X_3786_ cu.reg_file.reg_sp\[12\] _0636_ _0748_ cu.reg_file.reg_h\[4\] VGND VGND VPWR
+ VPWR _0862_ sky130_fd_sc_hd__a22o_1
X_5525_ _1625_ _2344_ VGND VGND VPWR VPWR _2345_ sky130_fd_sc_hd__nand2_4
XANTENNA__4751__A2 _1739_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5456_ _2283_ VGND VGND VPWR VPWR _2284_ sky130_fd_sc_hd__buf_2
X_4407_ cu.id.cb_opcode_x\[1\] _1295_ _1298_ cu.pc.pc_o\[7\] _1306_ VGND VGND VPWR
+ VPWR _1468_ sky130_fd_sc_hd__a221o_1
XANTENNA__4503__A2 _1321_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5387_ _2238_ VGND VGND VPWR VPWR _0166_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5700__B2 _1646_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4338_ _1356_ _1401_ _1402_ VGND VGND VPWR VPWR _1403_ sky130_fd_sc_hd__o21ai_1
X_4269_ _1330_ _1334_ _1336_ VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__a21oi_1
X_6008_ clknet_leaf_3_clk _0046_ net156 VGND VGND VPWR VPWR cu.reg_file.reg_b\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_96_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_77_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_49_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5519__A1 net31 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5519__B2 net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_24_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3491__A _0566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4258__A1 cu.reg_file.reg_sp\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4258__B2 _1299_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4753__C _0307_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4430__B2 cu.pc.pc_o\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3640_ _0711_ _0714_ _0715_ VGND VGND VPWR VPWR _0716_ sky130_fd_sc_hd__a21oi_2
XFILLER_0_36_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5930__A1 _2448_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3571_ cu.reg_file.reg_d\[5\] _0415_ _0432_ cu.reg_file.reg_b\[5\] VGND VGND VPWR
+ VPWR _0647_ sky130_fd_sc_hd__a22o_1
XFILLER_0_87_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5310_ _2193_ VGND VGND VPWR VPWR _2194_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_11_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_3_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6290_ clknet_leaf_41_clk _0272_ net151 VGND VGND VPWR VPWR cu.id.alu_opcode\[0\]
+ sky130_fd_sc_hd__dfrtp_2
X_5241_ _1374_ _2148_ VGND VGND VPWR VPWR _2149_ sky130_fd_sc_hd__nor2_1
XANTENNA__5092__S _2035_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4497__A1 cu.reg_file.reg_d\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4497__B2 cu.reg_file.reg_sp\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5172_ _2100_ VGND VGND VPWR VPWR _0089_ sky130_fd_sc_hd__clkbuf_1
X_4123_ _1126_ VGND VGND VPWR VPWR _1193_ sky130_fd_sc_hd__clkbuf_4
Xinput2 keypad_input[0] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__buf_2
X_4054_ _1110_ _1126_ VGND VGND VPWR VPWR _1128_ sky130_fd_sc_hd__and2_1
X_3005_ net75 net34 ih.gpio_interrupt_mask\[7\] VGND VGND VPWR VPWR _2743_ sky130_fd_sc_hd__and3b_1
XANTENNA__3457__C1 cu.reg_file.reg_l\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4956_ cu.pc.pc_o\[11\] _1521_ _1233_ VGND VGND VPWR VPWR _1946_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_52_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_19_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4887_ cu.pc.pc_o\[6\] _1882_ _1815_ VGND VGND VPWR VPWR _1883_ sky130_fd_sc_hd__mux2_1
X_3907_ _0982_ VGND VGND VPWR VPWR _0983_ sky130_fd_sc_hd__inv_2
XFILLER_0_34_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3838_ _0833_ _0912_ _0913_ VGND VGND VPWR VPWR _0914_ sky130_fd_sc_hd__o21a_1
XFILLER_0_61_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3295__B _0361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5508_ _2125_ _2325_ _2326_ ih.gpio_interrupt_mask\[0\] _2327_ VGND VGND VPWR VPWR
+ _2328_ sky130_fd_sc_hd__a221o_1
XFILLER_0_14_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5791__A cu.reg_file.reg_sp\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3769_ _0844_ VGND VGND VPWR VPWR _0845_ sky130_fd_sc_hd__inv_2
XFILLER_0_42_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5439_ _2269_ VGND VGND VPWR VPWR _0187_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4854__B cu.pc.pc_o\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3448__C1 _2918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1012 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1001 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1056 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1045 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1034 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1023 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_32_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1089 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1078 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1067 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_244 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4176__A0 _0566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6038__RESET_B net161 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_807 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_829 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4810_ _1300_ _1768_ VGND VGND VPWR VPWR _1812_ sky130_fd_sc_hd__xor2_1
XANTENNA__5600__B1 _2225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5790_ _2575_ VGND VGND VPWR VPWR _0232_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4403__A1 cu.reg_file.reg_a\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4403__B2 cu.reg_file.reg_sp\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5087__S _2039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4741_ _2922_ _0303_ VGND VGND VPWR VPWR _1750_ sky130_fd_sc_hd__and2b_1
XFILLER_0_22_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4672_ _1699_ _1700_ VGND VGND VPWR VPWR ih.t.next_count\[12\] sky130_fd_sc_hd__nor2_1
XFILLER_0_22_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5903__A1 _1189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3623_ cu.reg_file.reg_mem\[3\] _0418_ _0433_ cu.reg_file.reg_a\[3\] VGND VGND VPWR
+ VPWR _0699_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3554_ cu.reg_file.reg_b\[6\] _0502_ _0499_ cu.reg_file.reg_a\[6\] _0629_ VGND VGND
+ VPWR VPWR _0630_ sky130_fd_sc_hd__a221o_1
X_6273_ clknet_leaf_12_clk _0255_ net174 VGND VGND VPWR VPWR ih.t.timer_max\[5\] sky130_fd_sc_hd__dfrtp_4
X_3485_ cu.reg_file.reg_b\[7\] _0502_ _0492_ cu.reg_file.reg_d\[7\] VGND VGND VPWR
+ VPWR _0561_ sky130_fd_sc_hd__a22o_1
X_5224_ _2134_ VGND VGND VPWR VPWR _0107_ sky130_fd_sc_hd__clkbuf_1
XANTENNA_fanout195_A net196 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5419__A0 _1261_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5155_ cu.reg_file.reg_l\[2\] _1074_ _2088_ VGND VGND VPWR VPWR _2091_ sky130_fd_sc_hd__mux2_1
X_5086_ _1187_ _1222_ _2035_ VGND VGND VPWR VPWR _2045_ sky130_fd_sc_hd__mux2_1
X_4106_ cu.alu_f\[2\] _1013_ _1012_ VGND VGND VPWR VPWR _1180_ sky130_fd_sc_hd__o21a_1
X_4037_ _0611_ _0643_ VGND VGND VPWR VPWR _1111_ sky130_fd_sc_hd__nand2_1
XFILLER_0_78_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5988_ clknet_leaf_28_clk _0026_ net188 VGND VGND VPWR VPWR cu.pc.pc_o\[10\] sky130_fd_sc_hd__dfrtp_1
X_4939_ _1521_ _1907_ cu.pc.pc_o\[11\] VGND VGND VPWR VPWR _1930_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_47_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4584__B _1530_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_534 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output89_A net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3270_ _2874_ _2927_ VGND VGND VPWR VPWR _0346_ sky130_fd_sc_hd__or2_1
XTAP_604 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_626 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3675__A2 _0640_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4494__B _1545_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5911_ cu.ir.idx\[0\] VGND VGND VPWR VPWR _2663_ sky130_fd_sc_hd__inv_2
XANTENNA__5821__A0 cu.reg_file.reg_sp\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5842_ _2611_ _2614_ _2612_ VGND VGND VPWR VPWR _2621_ sky130_fd_sc_hd__a21bo_1
XANTENNA__5585__C1 _1661_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5773_ cu.reg_file.reg_sp\[4\] _2560_ _2539_ VGND VGND VPWR VPWR _2561_ sky130_fd_sc_hd__mux2_1
X_4724_ ih.t.count\[30\] _1732_ _1670_ VGND VGND VPWR VPWR _1735_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_90_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2985_ net3 VGND VGND VPWR VPWR _2724_ sky130_fd_sc_hd__inv_2
XFILLER_0_16_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4655_ ih.t.count\[6\] ih.t.count\[7\] _1683_ VGND VGND VPWR VPWR _1689_ sky130_fd_sc_hd__and3_1
XANTENNA__5888__A0 _1191_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_364 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_31_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4586_ _1434_ _1462_ _1473_ _1629_ VGND VGND VPWR VPWR _1630_ sky130_fd_sc_hd__or4_4
XFILLER_0_3_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3899__C1 _0296_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3606_ _0671_ _0681_ VGND VGND VPWR VPWR _0682_ sky130_fd_sc_hd__and2b_1
X_3537_ _0610_ _0612_ net142 _0601_ VGND VGND VPWR VPWR _0613_ sky130_fd_sc_hd__a211o_1
X_3468_ _0294_ _0360_ _0536_ VGND VGND VPWR VPWR _0544_ sky130_fd_sc_hd__o21ai_1
X_6256_ clknet_leaf_0_clk _0238_ net153 VGND VGND VPWR VPWR cu.reg_file.reg_sp\[12\]
+ sky130_fd_sc_hd__dfstp_2
X_5207_ _2124_ VGND VGND VPWR VPWR _0100_ sky130_fd_sc_hd__clkbuf_1
X_6187_ clknet_leaf_20_clk _0220_ net189 VGND VGND VPWR VPWR mc.cl.next_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_3399_ cu.id.cb_opcode_z\[1\] _2918_ _0364_ _0470_ _0474_ VGND VGND VPWR VPWR _0475_
+ sky130_fd_sc_hd__o221a_1
XANTENNA__3666__A2 _0488_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5138_ _1209_ _1144_ _2066_ VGND VGND VPWR VPWR _2079_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5069_ _2032_ VGND VGND VPWR VPWR _0054_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5812__A0 _1623_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_114 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5040__A1 _1213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output127_A net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5031__A1 _1623_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3593__B2 cu.reg_file.reg_a\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3593__A1 cu.reg_file.reg_mem\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4440_ _2701_ _1478_ _1353_ VGND VGND VPWR VPWR _1500_ sky130_fd_sc_hd__a21o_1
XFILLER_0_53_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4489__B _1545_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6110_ clknet_leaf_7_clk _0144_ net167 VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__dfrtp_1
XANTENNA__6200__D net13 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4371_ _1428_ _1429_ _1433_ VGND VGND VPWR VPWR _1434_ sky130_fd_sc_hd__o21a_2
XFILLER_0_95_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5098__A1 _1263_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3322_ _0361_ _0388_ _0397_ _2891_ _2887_ VGND VGND VPWR VPWR _0398_ sky130_fd_sc_hd__a311o_1
XTAP_401 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6041_ clknet_leaf_33_clk _0079_ net162 VGND VGND VPWR VPWR cu.reg_file.reg_h\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_3253_ _2925_ _2932_ VGND VGND VPWR VPWR _0329_ sky130_fd_sc_hd__nor2_1
XTAP_434 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3184_ cu.id.cb_opcode_x\[0\] VGND VGND VPWR VPWR _2921_ sky130_fd_sc_hd__inv_2
XTAP_478 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3648__A2 _0415_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout158_A net160 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5825_ _2604_ _2605_ VGND VGND VPWR VPWR _2606_ sky130_fd_sc_hd__nand2_1
XFILLER_0_36_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2968_ _2705_ _2707_ VGND VGND VPWR VPWR _2708_ sky130_fd_sc_hd__and2_1
X_5756_ _1073_ _2544_ _2545_ VGND VGND VPWR VPWR _2546_ sky130_fd_sc_hd__mux2_1
X_4707_ net230 _1720_ _1687_ VGND VGND VPWR VPWR _1724_ sky130_fd_sc_hd__o21ai_1
X_5687_ mc.cl.next_data\[10\] _2359_ _2490_ _2496_ VGND VGND VPWR VPWR _2497_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__5275__S _2170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3584__A1 cu.reg_file.reg_e\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3584__B2 cu.reg_file.reg_h\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4638_ ih.t.count\[0\] ih.t.count\[1\] ih.t.count\[2\] VGND VGND VPWR VPWR _1677_
+ sky130_fd_sc_hd__nand3_1
XFILLER_0_8_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4569_ _1382_ _1616_ _1617_ _1621_ VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__a31o_1
X_6308_ clknet_leaf_19_clk _0290_ net183 VGND VGND VPWR VPWR cu.id.imm_i\[13\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__5089__A1 _1213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6239_ clknet_leaf_22_clk ih.t.next_count\[27\] net191 VGND VGND VPWR VPWR ih.t.count\[27\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__4619__S _1661_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_990 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5261__A1 _2163_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_35_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3327__A1 _2878_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5721__C1 _2870_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4827__A1 _1299_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3940_ _0976_ _0981_ _1008_ VGND VGND VPWR VPWR _1016_ sky130_fd_sc_hd__and3_1
XFILLER_0_14_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3802__A2 _0488_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3871_ _0817_ _0945_ _0946_ VGND VGND VPWR VPWR _0947_ sky130_fd_sc_hd__and3_1
XFILLER_0_45_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5610_ net72 _1648_ _2137_ _2274_ VGND VGND VPWR VPWR _2426_ sky130_fd_sc_hd__a31o_1
XFILLER_0_26_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_90_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5541_ ih.t.timer_max\[25\] _2146_ _2204_ ih.t.timer_max\[17\] VGND VGND VPWR VPWR
+ _2360_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3566__A1 cu.reg_file.reg_l\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5095__S _2035_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5472_ _2147_ VGND VGND VPWR VPWR _2296_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4423_ _1268_ _2947_ VGND VGND VPWR VPWR _1483_ sky130_fd_sc_hd__or2_2
XFILLER_0_1_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4354_ _2701_ _1404_ _1417_ VGND VGND VPWR VPWR _1418_ sky130_fd_sc_hd__and3_1
X_3305_ _0361_ _0376_ _2926_ _2928_ VGND VGND VPWR VPWR _0381_ sky130_fd_sc_hd__a211o_1
XTAP_242 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4285_ _1335_ _1349_ _1351_ VGND VGND VPWR VPWR _1352_ sky130_fd_sc_hd__o21a_1
XTAP_275 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_253 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6024_ clknet_leaf_3_clk _0062_ net156 VGND VGND VPWR VPWR cu.reg_file.reg_d\[6\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__5491__A1 net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_297 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3236_ _2894_ _2916_ _2939_ VGND VGND VPWR VPWR _0312_ sky130_fd_sc_hd__a21oi_4
X_3167_ _2898_ _2903_ VGND VGND VPWR VPWR _2904_ sky130_fd_sc_hd__or2_2
X_3098_ ih.t.timer_max\[1\] ih.t.count\[1\] VGND VGND VPWR VPWR _2836_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_49_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_18_clk_A clknet_2_1__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5808_ cu.reg_file.reg_sp\[9\] _2536_ VGND VGND VPWR VPWR _2591_ sky130_fd_sc_hd__nand2_1
XANTENNA__4754__B1 _0350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5739_ cu.reg_file.reg_sp\[1\] VGND VGND VPWR VPWR _2530_ sky130_fd_sc_hd__inv_2
XFILLER_0_17_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_20_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5482__A1 _0618_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5234__A1 _2085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3796__A1 cu.reg_file.reg_sp\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3796__B2 cu.reg_file.reg_h\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5537__A2 _2205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3936__B _2918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5209__A _1364_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_50_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output71_A net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4070_ _1143_ VGND VGND VPWR VPWR _1144_ sky130_fd_sc_hd__buf_4
XFILLER_0_92_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3021_ ih.t.timer_max\[19\] ih.t.timer_max\[20\] _2758_ VGND VGND VPWR VPWR _2759_
+ sky130_fd_sc_hd__or3_1
XANTENNA__4783__A _0986_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5598__B _1330_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4433__C1 _1323_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4972_ _1953_ _1960_ _1808_ VGND VGND VPWR VPWR _1961_ sky130_fd_sc_hd__mux2_1
X_3923_ _0980_ VGND VGND VPWR VPWR _0999_ sky130_fd_sc_hd__inv_2
XANTENNA__3787__B2 cu.reg_file.reg_d\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3787__A1 cu.reg_file.reg_b\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3854_ _0842_ _0929_ _0843_ VGND VGND VPWR VPWR _0930_ sky130_fd_sc_hd__o21ai_2
XFILLER_0_6_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3785_ cu.id.imm_i\[12\] _0739_ _0860_ _0653_ VGND VGND VPWR VPWR _0861_ sky130_fd_sc_hd__a22oi_4
X_5524_ _1666_ _2191_ VGND VGND VPWR VPWR _2344_ sky130_fd_sc_hd__nand2_2
XANTENNA__4023__A _0918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5455_ _1364_ _2274_ _2275_ _2282_ VGND VGND VPWR VPWR _2283_ sky130_fd_sc_hd__or4_1
XFILLER_0_67_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4406_ _1271_ _1466_ VGND VGND VPWR VPWR _1467_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5386_ _0619_ net124 _2237_ VGND VGND VPWR VPWR _2238_ sky130_fd_sc_hd__mux2_1
X_4337_ mc.rw.state\[1\] mc.rw.state\[0\] _2698_ VGND VGND VPWR VPWR _1402_ sky130_fd_sc_hd__o21ai_4
XANTENNA__5692__A2_N _1643_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4268_ mc.rw.state\[2\] _2705_ _2707_ _1335_ VGND VGND VPWR VPWR _1336_ sky130_fd_sc_hd__o211a_1
X_6007_ clknet_leaf_18_clk _0045_ net185 VGND VGND VPWR VPWR cu.reg_file.reg_b\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_3219_ _0294_ VGND VGND VPWR VPWR _0295_ sky130_fd_sc_hd__clkbuf_4
X_4199_ _0323_ _1266_ _2912_ _2937_ VGND VGND VPWR VPWR _1267_ sky130_fd_sc_hd__o211a_1
XFILLER_0_69_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3491__B _0547_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4258__A2 _0993_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3466__B1 _0495_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4718__B1 _1670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_70_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3570_ _0295_ _0634_ _0373_ VGND VGND VPWR VPWR _0646_ sky130_fd_sc_hd__or3b_1
XFILLER_0_51_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5240_ _1329_ _1372_ VGND VGND VPWR VPWR _2148_ sky130_fd_sc_hd__or2_2
XANTENNA__5373__S _2226_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4497__A2 _1282_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5694__B2 ih.t.timer_max\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5171_ _1647_ _2099_ VGND VGND VPWR VPWR _2100_ sky130_fd_sc_hd__and2_1
X_4122_ net208 _1186_ _0370_ _1192_ VGND VGND VPWR VPWR _0012_ sky130_fd_sc_hd__a22o_1
X_4053_ _1110_ _1126_ VGND VGND VPWR VPWR _1127_ sky130_fd_sc_hd__nor2_1
XANTENNA__5402__A _1369_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3004_ _2740_ net32 ih.gpio_interrupt_mask\[5\] _2741_ VGND VGND VPWR VPWR _2742_
+ sky130_fd_sc_hd__a31o_1
Xinput3 keypad_input[10] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__buf_4
XFILLER_0_93_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4955_ _1943_ _1944_ VGND VGND VPWR VPWR _1945_ sky130_fd_sc_hd__or2_1
XFILLER_0_46_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3906_ _0976_ _0981_ VGND VGND VPWR VPWR _0982_ sky130_fd_sc_hd__nand2_1
X_4886_ _1874_ _1881_ _1809_ VGND VGND VPWR VPWR _1882_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4709__B1 _1670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3837_ _0829_ _0832_ VGND VGND VPWR VPWR _0913_ sky130_fd_sc_hd__or2_1
X_3768_ _0842_ _0843_ VGND VGND VPWR VPWR _0844_ sky130_fd_sc_hd__and2b_1
XFILLER_0_42_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5507_ _1415_ _1629_ _1637_ VGND VGND VPWR VPWR _2327_ sky130_fd_sc_hd__nor3_4
XFILLER_0_42_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5283__S _2170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3699_ _0620_ _0547_ VGND VGND VPWR VPWR _0775_ sky130_fd_sc_hd__nand2_1
X_5438_ _2022_ net73 _2268_ VGND VGND VPWR VPWR _2269_ sky130_fd_sc_hd__mux2_1
XANTENNA__5685__A1 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5369_ _1052_ net117 _2226_ VGND VGND VPWR VPWR _2228_ sky130_fd_sc_hd__mux2_1
XANTENNA__3448__B1 _0387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1013 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1002 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1046 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1035 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1024 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1079 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1068 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1057 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_407 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_37_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_37_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5373__A0 _1188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5912__A2 _1644_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4598__A _1415_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_808 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_819 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_73_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_145 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4939__B1 cu.pc.pc_o\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5600__B2 net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5600__A1 net112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_510 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4740_ _2908_ _0361_ _0968_ _0313_ _0326_ VGND VGND VPWR VPWR _1749_ sky130_fd_sc_hd__o32a_1
XFILLER_0_28_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4671_ ih.t.count\[12\] _1696_ _1687_ VGND VGND VPWR VPWR _1700_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_83_362 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__6203__D net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3622_ cu.reg_file.reg_c\[3\] _0427_ _0430_ cu.reg_file.reg_e\[3\] VGND VGND VPWR
+ VPWR _0698_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3914__A1 _2936_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3553_ cu.pc.pc_o\[6\] _0501_ _0628_ cu.reg_file.reg_mem\[6\] _0536_ VGND VGND VPWR
+ VPWR _0629_ sky130_fd_sc_hd__a221o_1
X_6272_ clknet_leaf_12_clk _0254_ net174 VGND VGND VPWR VPWR ih.t.timer_max\[4\] sky130_fd_sc_hd__dfstp_1
X_3484_ cu.reg_file.reg_c\[7\] _0485_ _0489_ cu.reg_file.reg_e\[7\] _0559_ VGND VGND
+ VPWR VPWR _0560_ sky130_fd_sc_hd__a221o_2
X_5223_ _1194_ ih.gpio_interrupt_mask\[6\] _2127_ VGND VGND VPWR VPWR _2134_ sky130_fd_sc_hd__mux2_1
X_5154_ _2090_ VGND VGND VPWR VPWR _0081_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5419__A1 net139 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4105_ _0395_ _1169_ _1170_ _1178_ VGND VGND VPWR VPWR _1179_ sky130_fd_sc_hd__o31ai_1
XANTENNA_fanout188_A net196 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5085_ _2044_ VGND VGND VPWR VPWR _0058_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4036_ _1109_ VGND VGND VPWR VPWR _1110_ sky130_fd_sc_hd__buf_4
XFILLER_0_78_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5987_ clknet_leaf_27_clk _0025_ net186 VGND VGND VPWR VPWR cu.pc.pc_o\[9\] sky130_fd_sc_hd__dfrtp_4
XPHY_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4938_ cu.pc.pc_o\[11\] _1521_ _1907_ VGND VGND VPWR VPWR _1929_ sky130_fd_sc_hd__and3_1
XFILLER_0_47_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3602__B1 _0499_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4869_ _1851_ _1854_ _1852_ VGND VGND VPWR VPWR _1866_ sky130_fd_sc_hd__o21a_1
XFILLER_0_62_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4158__B2 _0916_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4584__C _1545_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5594__A0 cu.reg_file.reg_mem\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5897__A1 _1051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4121__A _1191_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_605 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4321__A1 cu.reg_file.reg_c\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_627 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5910_ _2662_ VGND VGND VPWR VPWR _0265_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3427__A3 _0307_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_16_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4791__A _1186_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5098__S _2035_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5841_ _2618_ _2619_ VGND VGND VPWR VPWR _2620_ sky130_fd_sc_hd__nand2_1
X_2984_ net13 VGND VGND VPWR VPWR _2723_ sky130_fd_sc_hd__inv_2
XANTENNA__4388__B2 cu.pc.pc_o\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4388__A1 _0387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5772_ _1160_ _2559_ _2545_ VGND VGND VPWR VPWR _2560_ sky130_fd_sc_hd__mux2_1
X_4723_ _1734_ VGND VGND VPWR VPWR ih.t.next_count\[29\] sky130_fd_sc_hd__clkbuf_1
XANTENNA__3200__A _2936_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5337__A0 _1188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4654_ _1686_ _1688_ VGND VGND VPWR VPWR ih.t.next_count\[6\] sky130_fd_sc_hd__nor2_1
XFILLER_0_71_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4585_ _1393_ _1627_ _1628_ VGND VGND VPWR VPWR _1629_ sky130_fd_sc_hd__or3_4
XFILLER_0_12_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3605_ _0653_ _0673_ _0675_ _0680_ VGND VGND VPWR VPWR _0681_ sky130_fd_sc_hd__o22a_2
XANTENNA__4560__A1 cu.reg_file.reg_h\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3536_ _0447_ _0611_ VGND VGND VPWR VPWR _0612_ sky130_fd_sc_hd__nand2_1
X_6255_ clknet_leaf_42_clk _0237_ net155 VGND VGND VPWR VPWR cu.reg_file.reg_sp\[11\]
+ sky130_fd_sc_hd__dfstp_4
X_5206_ _2122_ mc.cc.count\[3\] _2120_ VGND VGND VPWR VPWR _2124_ sky130_fd_sc_hd__and3b_1
XANTENNA__4966__A _1233_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3467_ cu.reg_file.reg_sp\[1\] _0539_ _0540_ _0541_ _0542_ VGND VGND VPWR VPWR _0543_
+ sky130_fd_sc_hd__a2111o_1
X_6186_ clknet_leaf_24_clk _0219_ net190 VGND VGND VPWR VPWR mc.cl.next_data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_3398_ _2900_ _2878_ _0301_ VGND VGND VPWR VPWR _0474_ sky130_fd_sc_hd__a21o_1
X_5137_ _2078_ VGND VGND VPWR VPWR _0076_ sky130_fd_sc_hd__clkbuf_1
X_5068_ cu.reg_file.reg_c\[6\] _1193_ _2025_ VGND VGND VPWR VPWR _2032_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4019_ _0801_ _0812_ VGND VGND VPWR VPWR _1093_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5576__B1 _2247_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4876__A cu.pc.pc_o\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4595__B _1417_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4067__B1 _0663_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3290__A1 _0359_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4370_ cu.reg_file.reg_c\[5\] _1313_ _1430_ _1432_ VGND VGND VPWR VPWR _1433_ sky130_fd_sc_hd__a211o_1
XANTENNA__4542__B2 cu.reg_file.reg_d\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4542__A1 cu.pc.pc_o\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3321_ _0375_ _0396_ cu.id.cb_opcode_x\[1\] _0387_ VGND VGND VPWR VPWR _0397_ sky130_fd_sc_hd__a211o_1
XANTENNA__5381__S _2226_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4786__A _1299_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_402 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3252_ _2887_ _2891_ _0323_ _0327_ VGND VGND VPWR VPWR _0328_ sky130_fd_sc_hd__or4b_4
XTAP_435 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6040_ clknet_leaf_33_clk _0078_ net161 VGND VGND VPWR VPWR cu.reg_file.reg_h\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_3183_ cu.id.cb_opcode_x\[1\] VGND VGND VPWR VPWR _2920_ sky130_fd_sc_hd__buf_4
XTAP_468 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5824_ cu.reg_file.reg_sp\[11\] _2536_ VGND VGND VPWR VPWR _2605_ sky130_fd_sc_hd__nand2_1
XFILLER_0_29_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2967_ _2701_ _2706_ VGND VGND VPWR VPWR _2707_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5755_ _2115_ VGND VGND VPWR VPWR _2545_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_44_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4706_ ih.t.count\[24\] _1720_ VGND VGND VPWR VPWR _1723_ sky130_fd_sc_hd__and2_1
X_5686_ ih.t.timer_max\[26\] _2151_ _2320_ ih.t.timer_max\[10\] VGND VGND VPWR VPWR
+ _2496_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_17_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_44_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4637_ ih.t.count\[0\] ih.t.count\[1\] ih.t.count\[2\] VGND VGND VPWR VPWR _1676_
+ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_451 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4568_ _1618_ _1619_ _1620_ _1614_ VGND VGND VPWR VPWR _1621_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__5291__S _2182_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6307_ clknet_leaf_18_clk _0289_ net184 VGND VGND VPWR VPWR cu.id.imm_i\[12\] sky130_fd_sc_hd__dfrtp_4
X_4499_ cu.id.imm_i\[12\] _1294_ _1297_ cu.pc.pc_o\[12\] _1488_ VGND VGND VPWR VPWR
+ _1555_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3519_ cu.id.cb_opcode_y\[1\] _0361_ _0437_ _0340_ _0583_ VGND VGND VPWR VPWR _0595_
+ sky130_fd_sc_hd__a221o_1
X_6238_ clknet_leaf_15_clk ih.t.next_count\[26\] net182 VGND VGND VPWR VPWR ih.t.count\[26\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_980 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6169_ clknet_leaf_2_clk _0203_ net155 VGND VGND VPWR VPWR cu.reg_file.reg_mem\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_991 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5797__A0 cu.reg_file.reg_sp\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_20_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_20_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_35_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4524__A1 _1304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4827__A2 cu.pc.pc_o\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3015__A ih.t.timer_max\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5788__A0 _1126_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_85_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_58_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3870_ _0833_ _0930_ VGND VGND VPWR VPWR _0946_ sky130_fd_sc_hd__xor2_2
XFILLER_0_38_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_11_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_11_clk sky130_fd_sc_hd__clkbuf_16
X_5540_ _2313_ VGND VGND VPWR VPWR _2359_ sky130_fd_sc_hd__buf_2
XANTENNA__5960__A0 cu.id.imm_i\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5471_ _2295_ VGND VGND VPWR VPWR _0193_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_30_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4422_ _1301_ _1300_ VGND VGND VPWR VPWR _1482_ sky130_fd_sc_hd__or2_1
X_4353_ _1306_ _1410_ _1414_ VGND VGND VPWR VPWR _1417_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_1_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4284_ _2696_ _1333_ VGND VGND VPWR VPWR _1351_ sky130_fd_sc_hd__or2_2
X_3304_ _0296_ _2891_ _0318_ VGND VGND VPWR VPWR _0380_ sky130_fd_sc_hd__or3_1
XTAP_221 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_232 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6023_ clknet_leaf_18_clk _0061_ net185 VGND VGND VPWR VPWR cu.reg_file.reg_d\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_3235_ _2885_ _2927_ _0309_ VGND VGND VPWR VPWR _0311_ sky130_fd_sc_hd__and3_1
XTAP_265 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_254 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_243 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5491__A2 _2205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_298 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3166_ _2901_ _2902_ _2884_ VGND VGND VPWR VPWR _2903_ sky130_fd_sc_hd__or3b_1
X_3097_ ih.t.timer_max\[4\] _2747_ VGND VGND VPWR VPWR _2835_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_12_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_532 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3999_ _1063_ _1070_ _1072_ VGND VGND VPWR VPWR _1073_ sky130_fd_sc_hd__nand3b_4
X_5807_ cu.reg_file.reg_sp\[9\] _2535_ VGND VGND VPWR VPWR _2590_ sky130_fd_sc_hd__or2_1
XFILLER_0_91_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5738_ net25 _2519_ _2529_ VGND VGND VPWR VPWR _0226_ sky130_fd_sc_hd__a21o_1
XFILLER_0_32_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5669_ _2169_ _2474_ _2481_ _2136_ VGND VGND VPWR VPWR _2482_ sky130_fd_sc_hd__o211a_1
XFILLER_0_67_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5942__A0 cu.id.cb_opcode_y\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5924__S _2668_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5170__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output64_A net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3020_ ih.t.timer_max\[18\] _2757_ VGND VGND VPWR VPWR _2758_ sky130_fd_sc_hd__or2_2
Xclkbuf_leaf_0_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_0_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__3484__B2 cu.reg_file.reg_e\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_58_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6206__D net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4433__B1 _1343_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4971_ _1958_ _1959_ _1798_ VGND VGND VPWR VPWR _1960_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3922_ _0986_ _0997_ VGND VGND VPWR VPWR _0998_ sky130_fd_sc_hd__nor2_1
XANTENNA__3787__A2 _0426_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3853_ _0854_ _0927_ _0928_ VGND VGND VPWR VPWR _0929_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_6_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3784_ cu.reg_file.reg_a\[4\] _0625_ _0628_ cu.reg_file.reg_mem\[12\] _0859_ VGND
+ VGND VPWR VPWR _0860_ sky130_fd_sc_hd__a221o_1
X_5523_ _2275_ _2342_ _1648_ VGND VGND VPWR VPWR _2343_ sky130_fd_sc_hd__and3b_1
XFILLER_0_26_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5454_ _1369_ _2276_ _2281_ VGND VGND VPWR VPWR _2282_ sky130_fd_sc_hd__o21ai_1
X_5385_ _2181_ _2236_ VGND VGND VPWR VPWR _2237_ sky130_fd_sc_hd__nand2_8
XANTENNA__5161__A1 _1191_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4405_ cu.reg_file.reg_c\[7\] _1281_ _1465_ VGND VGND VPWR VPWR _1466_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_1_251 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4677__C _1672_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4336_ _1348_ _1373_ VGND VGND VPWR VPWR _1401_ sky130_fd_sc_hd__nor2_4
XFILLER_0_10_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4267_ _1329_ VGND VGND VPWR VPWR _1335_ sky130_fd_sc_hd__inv_2
XFILLER_0_66_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6006_ clknet_leaf_31_clk _0044_ net185 VGND VGND VPWR VPWR cu.reg_file.reg_b\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_4198_ _2877_ _0436_ _0469_ VGND VGND VPWR VPWR _1266_ sky130_fd_sc_hd__and3_1
X_3218_ _0293_ VGND VGND VPWR VPWR _0294_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_508 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3149_ cu.id.opcode\[6\] cu.id.opcode\[7\] cu.id.opcode\[2\] cu.id.opcode\[1\] VGND
+ VGND VPWR VPWR _2886_ sky130_fd_sc_hd__and4bb_1
XFILLER_0_49_243 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_20_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3702__A2 _0773_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3466__B2 cu.reg_file.reg_h\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_43_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4124__A _1193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5654__S _1739_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5170_ mc.cl.next_data\[9\] net19 mc.count VGND VGND VPWR VPWR _2099_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_17_clk_A clknet_2_2__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4121_ _1191_ VGND VGND VPWR VPWR _1192_ sky130_fd_sc_hd__buf_4
X_4052_ _1115_ _1116_ _1119_ _1125_ VGND VGND VPWR VPWR _1126_ sky130_fd_sc_hd__or4b_4
X_3003_ net72 net31 ih.gpio_interrupt_mask\[4\] VGND VGND VPWR VPWR _2741_ sky130_fd_sc_hd__and3b_1
Xinput4 keypad_input[11] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__buf_2
XFILLER_0_36_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_2_1__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_1__leaf_clk sky130_fd_sc_hd__clkbuf_16
X_4954_ _1233_ cu.pc.pc_o\[12\] VGND VGND VPWR VPWR _1944_ sky130_fd_sc_hd__nor2_1
X_3905_ _0350_ _0980_ VGND VGND VPWR VPWR _0981_ sky130_fd_sc_hd__nor2_1
X_4885_ _1879_ _1880_ _1799_ VGND VGND VPWR VPWR _1881_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_321 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3836_ _0845_ _0910_ _0911_ VGND VGND VPWR VPWR _0912_ sky130_fd_sc_hd__a21oi_1
X_3767_ _0841_ _0838_ VGND VGND VPWR VPWR _0843_ sky130_fd_sc_hd__or2b_1
X_5506_ _1489_ _2125_ VGND VGND VPWR VPWR _2326_ sky130_fd_sc_hd__nor2_2
X_3698_ _0514_ _0605_ VGND VGND VPWR VPWR _0774_ sky130_fd_sc_hd__or2_2
XFILLER_0_42_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5437_ _2139_ _2225_ VGND VGND VPWR VPWR _2268_ sky130_fd_sc_hd__nand2_1
X_5368_ _2227_ VGND VGND VPWR VPWR _0158_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5685__A2 _1650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5299_ _1190_ net88 _2182_ VGND VGND VPWR VPWR _2187_ sky130_fd_sc_hd__mux2_1
X_4319_ cu.reg_file.reg_a\[3\] _1276_ _1287_ cu.reg_file.reg_sp\[3\] VGND VGND VPWR
+ VPWR _1384_ sky130_fd_sc_hd__a22o_1
XANTENNA__4645__B1 _1670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4209__A _2883_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1003 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1047 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1036 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1025 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1014 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1069 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1058 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3620__B2 cu.reg_file.reg_b\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3620__A1 cu.reg_file.reg_d\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5373__A1 net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4879__A _0387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_809 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4884__A0 _1126_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4939__A1 _1521_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3958__A _1032_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5600__A2 _2147_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3611__A1 cu.reg_file.reg_c\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3611__B2 cu.reg_file.reg_e\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4670_ ih.t.count\[12\] _1696_ VGND VGND VPWR VPWR _1699_ sky130_fd_sc_hd__and2_1
XFILLER_0_83_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_16_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_430 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3621_ cu.reg_file.reg_sp\[3\] _0413_ _0419_ cu.reg_file.reg_h\[3\] _0696_ VGND VGND
+ VPWR VPWR _0697_ sky130_fd_sc_hd__a221o_1
XANTENNA__4789__A _0350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3552_ _0494_ VGND VGND VPWR VPWR _0628_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6271_ clknet_leaf_12_clk _0253_ net174 VGND VGND VPWR VPWR ih.t.timer_max\[3\] sky130_fd_sc_hd__dfrtp_2
XFILLER_0_51_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3483_ _0464_ _0487_ _0482_ cu.reg_file.reg_l\[7\] VGND VGND VPWR VPWR _0559_ sky130_fd_sc_hd__o211a_1
X_5222_ _2133_ VGND VGND VPWR VPWR _0106_ sky130_fd_sc_hd__clkbuf_1
X_5153_ cu.reg_file.reg_l\[1\] _1051_ _2088_ VGND VGND VPWR VPWR _2090_ sky130_fd_sc_hd__mux2_1
X_4104_ _0547_ _0833_ _1176_ _1177_ VGND VGND VPWR VPWR _1178_ sky130_fd_sc_hd__a211o_1
X_5084_ cu.reg_file.reg_d\[2\] _2043_ _2039_ VGND VGND VPWR VPWR _2044_ sky130_fd_sc_hd__mux2_1
X_4035_ _1099_ _1105_ _1108_ VGND VGND VPWR VPWR _1109_ sky130_fd_sc_hd__or3b_1
XFILLER_0_2_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5986_ clknet_leaf_27_clk _0024_ net186 VGND VGND VPWR VPWR cu.pc.pc_o\[8\] sky130_fd_sc_hd__dfrtp_4
XPHY_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4937_ _1928_ VGND VGND VPWR VPWR _0026_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3602__A1 cu.pc.pc_o\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3602__B2 cu.reg_file.reg_a\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4868_ _1863_ _1864_ VGND VGND VPWR VPWR _1865_ sky130_fd_sc_hd__and2b_1
XANTENNA_20 _1233_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3819_ cu.reg_file.reg_mem\[9\] _0640_ _0893_ _0894_ VGND VGND VPWR VPWR _0895_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_6_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4799_ _0310_ _0311_ VGND VGND VPWR VPWR _1801_ sky130_fd_sc_hd__nor2_1
XFILLER_0_42_282 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5307__B _1354_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5107__A1 _1074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3669__A1 cu.pc.pc_o\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5291__A0 _0619_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6140__RESET_B net195 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5043__A0 _1191_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_511 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5594__A1 _2410_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_53_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5932__S _2668_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3018__A ih.t.timer_max\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_606 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5379__S _2226_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5624__A_N _1400_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5034__A0 _1074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5840_ cu.reg_file.reg_sp\[13\] _2536_ VGND VGND VPWR VPWR _2619_ sky130_fd_sc_hd__nand2_1
X_2983_ net7 VGND VGND VPWR VPWR _2722_ sky130_fd_sc_hd__inv_2
X_5771_ _2557_ _2558_ VGND VGND VPWR VPWR _2559_ sky130_fd_sc_hd__xor2_1
XFILLER_0_33_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4722_ _1732_ _1733_ _1669_ VGND VGND VPWR VPWR _1734_ sky130_fd_sc_hd__and3b_1
XFILLER_0_56_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_56_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5337__A1 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4653_ net227 _1683_ _1687_ VGND VGND VPWR VPWR _1688_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_71_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3348__B1 _0293_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4584_ _1511_ _1530_ _1545_ _1496_ VGND VGND VPWR VPWR _1628_ sky130_fd_sc_hd__or4b_1
XANTENNA__3899__A1 _0359_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3604_ _0677_ _0679_ VGND VGND VPWR VPWR _0680_ sky130_fd_sc_hd__or2_1
X_3535_ _0377_ _0602_ VGND VGND VPWR VPWR _0611_ sky130_fd_sc_hd__nor2_2
XFILLER_0_12_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3466_ cu.reg_file.reg_mem\[1\] _0482_ _0493_ _0495_ cu.reg_file.reg_h\[1\] VGND
+ VGND VPWR VPWR _0542_ sky130_fd_sc_hd__a32o_1
X_6254_ clknet_leaf_0_clk _0236_ net154 VGND VGND VPWR VPWR cu.reg_file.reg_sp\[10\]
+ sky130_fd_sc_hd__dfstp_4
X_5205_ net220 mc.cc.enable_edge_detector.prev_data _2122_ _2123_ VGND VGND VPWR VPWR
+ _0099_ sky130_fd_sc_hd__a31o_1
XANTENNA__4966__B cu.pc.pc_o\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6185_ clknet_leaf_34_clk _0218_ net158 VGND VGND VPWR VPWR ih.interrupt_source\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_3397_ _0335_ _0469_ _0453_ _0472_ _0293_ VGND VGND VPWR VPWR _0473_ sky130_fd_sc_hd__a41o_4
XFILLER_0_42_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5136_ _2077_ cu.reg_file.reg_h\[4\] _2069_ VGND VGND VPWR VPWR _2078_ sky130_fd_sc_hd__mux2_1
X_5067_ _2031_ VGND VGND VPWR VPWR _0053_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4076__A1 _0918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4018_ _0776_ _0801_ _1091_ _0768_ VGND VGND VPWR VPWR _1092_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_66_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5025__A0 _0618_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4379__A2 _1417_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5576__A1 net127 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5576__B2 net135 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5969_ _2694_ VGND VGND VPWR VPWR _0292_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4921__S _1798_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_30_274 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5053__A _0350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3275__C1 _0350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3814__A1 cu.pc.pc_o\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_80_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5228__A _1415_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output94_A net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3320_ _0373_ _0374_ VGND VGND VPWR VPWR _0396_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3750__B1 _0624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_403 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3251_ _0324_ _0325_ _2897_ _2909_ _0326_ VGND VGND VPWR VPWR _0327_ sky130_fd_sc_hd__a2111o_1
XTAP_425 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6062__RESET_B net195 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3182_ cu.id.cb_opcode_z\[0\] cu.id.cb_opcode_z\[1\] cu.id.cb_opcode_z\[2\] VGND
+ VGND VPWR VPWR _2919_ sky130_fd_sc_hd__and3b_1
XTAP_469 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__6209__D net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3805__B2 cu.reg_file.reg_mem\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3805__A1 cu.reg_file.reg_a\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_44_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5823_ cu.reg_file.reg_sp\[11\] _2536_ VGND VGND VPWR VPWR _2604_ sky130_fd_sc_hd__or2_1
XFILLER_0_63_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_224 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2966_ _2698_ mc.rw.state\[1\] mc.rw.state\[0\] VGND VGND VPWR VPWR _2706_ sky130_fd_sc_hd__and3_1
XFILLER_0_8_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5754_ _2530_ _2543_ VGND VGND VPWR VPWR _2544_ sky130_fd_sc_hd__xnor2_1
X_4705_ _1722_ VGND VGND VPWR VPWR ih.t.next_count\[23\] sky130_fd_sc_hd__clkbuf_1
X_5685_ net17 _1650_ _2488_ _2495_ VGND VGND VPWR VPWR _0207_ sky130_fd_sc_hd__a31o_1
XFILLER_0_17_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4636_ _1675_ VGND VGND VPWR VPWR ih.t.next_count\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5730__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4533__A2 _1579_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4567_ _2701_ _1618_ _1353_ VGND VGND VPWR VPWR _1620_ sky130_fd_sc_hd__a21o_1
X_6306_ clknet_leaf_6_clk _0288_ net164 VGND VGND VPWR VPWR cu.id.imm_i\[11\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4498_ cu.reg_file.reg_b\[4\] net143 _1284_ cu.reg_file.reg_h\[4\] _1553_ VGND VGND
+ VPWR VPWR _1554_ sky130_fd_sc_hd__a221o_1
XFILLER_0_12_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3518_ _0340_ _0443_ _0336_ VGND VGND VPWR VPWR _0594_ sky130_fd_sc_hd__a21o_1
X_6237_ clknet_leaf_15_clk ih.t.next_count\[25\] net179 VGND VGND VPWR VPWR ih.t.count\[25\]
+ sky130_fd_sc_hd__dfrtp_1
X_3449_ _0359_ _0386_ _2887_ VGND VGND VPWR VPWR _0525_ sky130_fd_sc_hd__a21oi_1
XTAP_970 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6168_ clknet_leaf_2_clk _0202_ net157 VGND VGND VPWR VPWR cu.reg_file.reg_mem\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_85_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_992 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_981 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5119_ _2034_ _2023_ VGND VGND VPWR VPWR _2065_ sky130_fd_sc_hd__or2_1
X_6099_ clknet_leaf_4_clk _0133_ net164 VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__dfrtp_2
XANTENNA__4049__B2 _1032_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4217__A _1284_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5549__A1 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_54_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4221__A1 cu.reg_file.reg_e\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output132_A net132 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4460__B2 _1511_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5960__A1 _2410_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5470_ net63 _2085_ _2294_ VGND VGND VPWR VPWR _2295_ sky130_fd_sc_hd__mux2_1
XFILLER_0_26_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4421_ _1423_ _1437_ _1456_ _1474_ VGND VGND VPWR VPWR _1481_ sky130_fd_sc_hd__or4_1
XFILLER_0_41_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4797__A _1798_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5392__S _2237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4352_ _1356_ _1404_ _1402_ VGND VGND VPWR VPWR _1416_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_1_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4283_ _1335_ _1349_ VGND VGND VPWR VPWR _1350_ sky130_fd_sc_hd__nand2_1
XANTENNA__4279__A1 cu.pc.pc_o\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3303_ _0378_ _0309_ VGND VGND VPWR VPWR _0379_ sky130_fd_sc_hd__and2_2
XTAP_200 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_233 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6022_ clknet_leaf_30_clk _0060_ net183 VGND VGND VPWR VPWR cu.reg_file.reg_d\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__4279__B2 cu.reg_file.reg_e\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_266 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_255 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3234_ _2923_ _2874_ _0309_ VGND VGND VPWR VPWR _0310_ sky130_fd_sc_hd__and3_1
XTAP_244 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_277 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3165_ cu.id.alu_opcode\[1\] VGND VGND VPWR VPWR _2902_ sky130_fd_sc_hd__buf_4
X_3096_ ih.t.count\[5\] _2833_ VGND VGND VPWR VPWR _2834_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_fanout163_A net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4451__A1 cu.reg_file.reg_b\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3006__A2 net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5400__A0 _1261_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3998_ _0531_ _1071_ _1040_ VGND VGND VPWR VPWR _1072_ sky130_fd_sc_hd__mux2_1
XFILLER_0_29_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5806_ _2589_ VGND VGND VPWR VPWR _0234_ sky130_fd_sc_hd__clkbuf_1
X_5737_ _2518_ mc.cl.next_data\[7\] _2111_ VGND VGND VPWR VPWR _2529_ sky130_fd_sc_hd__and3_1
X_5668_ ih.gpio_interrupt_mask\[7\] _2326_ _2480_ _2125_ _2327_ VGND VGND VPWR VPWR
+ _2481_ sky130_fd_sc_hd__a221o_1
XFILLER_0_32_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4619_ _1650_ _1657_ _1661_ VGND VGND VPWR VPWR _1662_ sky130_fd_sc_hd__mux2_1
X_5599_ net104 _2205_ _2414_ _1401_ VGND VGND VPWR VPWR _2415_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_20_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5219__A0 _1190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_67_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3402__C1 _2935_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5942__A1 _2410_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5506__A _1489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5940__S _2666_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output57_A net57 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5241__A _1374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4433__A1 cu.reg_file.reg_sp\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4970_ _1209_ _1953_ _1794_ VGND VGND VPWR VPWR _1959_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_46_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3921_ _0989_ _0994_ VGND VGND VPWR VPWR _0997_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3852_ _0853_ _0850_ VGND VGND VPWR VPWR _0928_ sky130_fd_sc_hd__and2b_1
XFILLER_0_6_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5522_ _2336_ _2341_ _2282_ VGND VGND VPWR VPWR _2342_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3783_ cu.pc.pc_o\[12\] _0740_ _0857_ _0858_ VGND VGND VPWR VPWR _0859_ sky130_fd_sc_hd__a211o_1
XFILLER_0_81_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5453_ _1374_ _2278_ _2280_ VGND VGND VPWR VPWR _2281_ sky130_fd_sc_hd__or3_1
X_5384_ _2235_ VGND VGND VPWR VPWR _2236_ sky130_fd_sc_hd__clkbuf_8
X_4404_ cu.reg_file.reg_e\[7\] _1283_ _1285_ cu.reg_file.reg_l\[7\] _1464_ VGND VGND
+ VPWR VPWR _1465_ sky130_fd_sc_hd__a221o_1
X_4335_ _1393_ VGND VGND VPWR VPWR _1400_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4266_ _2697_ _1333_ VGND VGND VPWR VPWR _1334_ sky130_fd_sc_hd__nor2_1
XFILLER_0_66_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6005_ clknet_leaf_31_clk _0043_ net185 VGND VGND VPWR VPWR cu.reg_file.reg_b\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_3217_ cu.id.starting_int_service VGND VGND VPWR VPWR _0293_ sky130_fd_sc_hd__clkbuf_4
X_4197_ _0370_ _1261_ _1262_ _1264_ _1265_ VGND VGND VPWR VPWR _0014_ sky130_fd_sc_hd__a221o_1
X_3148_ cu.id.alu_opcode\[0\] cu.id.opcode\[0\] VGND VGND VPWR VPWR _2885_ sky130_fd_sc_hd__and2_2
XANTENNA__3337__A_N _0405_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3079_ ih.t.timer_max\[10\] _2752_ ih.t.timer_max\[11\] VGND VGND VPWR VPWR _2817_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_82_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_531 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5297__S _2182_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_92_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5924__A1 _2391_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4188__A0 cu.alu_f\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4514__A2_N _1561_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_60_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5688__B1 cu.reg_file.reg_mem\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_450 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3280__A1_N _2918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4120_ _1144_ VGND VGND VPWR VPWR _1191_ sky130_fd_sc_hd__clkbuf_4
X_4051_ _0570_ _0644_ _1124_ _1069_ VGND VGND VPWR VPWR _1125_ sky130_fd_sc_hd__o22a_1
XANTENNA__4103__B1 _0824_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput5 keypad_input[12] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_4
X_3002_ net73 VGND VGND VPWR VPWR _2740_ sky130_fd_sc_hd__inv_2
XANTENNA__5851__A0 cu.reg_file.reg_sp\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4953_ _2920_ cu.pc.pc_o\[12\] VGND VGND VPWR VPWR _1943_ sky130_fd_sc_hd__and2_1
XANTENNA__3614__C1 _0536_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3904_ _0449_ _0971_ _0979_ _2935_ VGND VGND VPWR VPWR _0980_ sky130_fd_sc_hd__and4b_2
XFILLER_0_74_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4884_ _1126_ _1874_ _1795_ VGND VGND VPWR VPWR _1880_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_333 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3835_ _0838_ _0841_ VGND VGND VPWR VPWR _0911_ sky130_fd_sc_hd__nor2_1
XFILLER_0_54_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3766_ _0838_ _0841_ VGND VGND VPWR VPWR _0842_ sky130_fd_sc_hd__and2b_1
X_5505_ mc.cl.next_data\[0\] _2313_ _2323_ _2324_ VGND VGND VPWR VPWR _2325_ sky130_fd_sc_hd__a22o_1
X_5436_ _2267_ VGND VGND VPWR VPWR _0186_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3697_ _0772_ VGND VGND VPWR VPWR _0773_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5367_ _0619_ net116 _2226_ VGND VGND VPWR VPWR _2227_ sky130_fd_sc_hd__mux2_1
X_4318_ _1377_ _1379_ _1378_ VGND VGND VPWR VPWR _1383_ sky130_fd_sc_hd__a21bo_1
X_5298_ _2186_ VGND VGND VPWR VPWR _0129_ sky130_fd_sc_hd__clkbuf_1
X_4249_ _1316_ VGND VGND VPWR VPWR _1317_ sky130_fd_sc_hd__buf_2
XFILLER_0_96_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1004 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_84_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_1037 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1026 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1015 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1059 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1048 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5070__A1 _1260_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4225__A _2950_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3620__A2 _0415_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4879__B cu.pc.pc_o\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3136__A1 _2745_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3304__A _0296_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3620_ cu.reg_file.reg_d\[3\] _0415_ _0432_ cu.reg_file.reg_b\[3\] VGND VGND VPWR
+ VPWR _0696_ sky130_fd_sc_hd__a22o_1
XFILLER_0_24_442 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3551_ cu.reg_file.reg_h\[6\] _0495_ _0624_ cu.reg_file.reg_sp\[6\] _0626_ VGND VGND
+ VPWR VPWR _0627_ sky130_fd_sc_hd__a221o_1
XFILLER_0_24_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6270_ clknet_leaf_9_clk _0252_ net174 VGND VGND VPWR VPWR ih.t.timer_max\[2\] sky130_fd_sc_hd__dfrtp_2
X_3482_ _0547_ _0549_ _0552_ _0554_ _0557_ VGND VGND VPWR VPWR _0558_ sky130_fd_sc_hd__a2111o_4
X_5221_ _1192_ ih.gpio_interrupt_mask\[5\] _2127_ VGND VGND VPWR VPWR _2133_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5152_ _2089_ VGND VGND VPWR VPWR _0080_ sky130_fd_sc_hd__clkbuf_1
X_4103_ _0547_ _0833_ _0824_ VGND VGND VPWR VPWR _1177_ sky130_fd_sc_hd__o21ai_1
X_5083_ _1074_ _1226_ _2035_ VGND VGND VPWR VPWR _2043_ sky130_fd_sc_hd__mux2_1
X_4034_ _0570_ _0733_ _1106_ _1107_ VGND VGND VPWR VPWR _1108_ sky130_fd_sc_hd__o211a_1
XFILLER_0_78_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5985_ clknet_leaf_27_clk _0023_ net186 VGND VGND VPWR VPWR cu.pc.pc_o\[7\] sky130_fd_sc_hd__dfrtp_4
XPHY_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4936_ _1521_ _1927_ _1814_ VGND VGND VPWR VPWR _1928_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3602__A2 _0501_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_21 mc.cl.next_data\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4867_ _0373_ cu.pc.pc_o\[5\] VGND VGND VPWR VPWR _1864_ sky130_fd_sc_hd__nand2_1
XANTENNA_10 keypad_input[5] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4158__A3 _0779_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3818_ cu.reg_file.reg_b\[1\] _0426_ _0429_ cu.reg_file.reg_d\[1\] VGND VGND VPWR
+ VPWR _0894_ sky130_fd_sc_hd__a22o_1
X_4798_ _1789_ _1796_ _1799_ VGND VGND VPWR VPWR _1800_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3749_ cu.reg_file.reg_d\[7\] _0488_ _0741_ cu.reg_file.reg_h\[7\] VGND VGND VPWR
+ VPWR _0825_ sky130_fd_sc_hd__a22o_1
X_5419_ _1261_ net139 _2248_ VGND VGND VPWR VPWR _2256_ sky130_fd_sc_hd__mux2_1
XANTENNA__3669__A2 _0740_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5291__A1 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5043__A1 _1209_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_2_0__f_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_16_clk_A clknet_2_2__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4554__B1 _1284_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5704__A2_N _1643_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_607 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_88_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5034__A1 _1226_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2982_ net17 VGND VGND VPWR VPWR _2721_ sky130_fd_sc_hd__inv_2
X_5770_ _2550_ _2551_ _2549_ VGND VGND VPWR VPWR _2558_ sky130_fd_sc_hd__a21o_1
XFILLER_0_29_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4721_ ih.t.count\[27\] ih.t.count\[28\] _1726_ ih.t.count\[29\] VGND VGND VPWR VPWR
+ _1733_ sky130_fd_sc_hd__a31o_1
XFILLER_0_90_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4652_ _1669_ VGND VGND VPWR VPWR _1687_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_56_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput30 programmable_gpio_in[3] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3603_ cu.reg_file.reg_sp\[4\] _0539_ _0492_ cu.reg_file.reg_d\[4\] _0678_ VGND VGND
+ VPWR VPWR _0679_ sky130_fd_sc_hd__a221o_1
XANTENNA__4312__B _1374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4583_ _1561_ _1626_ _1598_ _1614_ VGND VGND VPWR VPWR _1627_ sky130_fd_sc_hd__or4b_1
XFILLER_0_12_401 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3534_ _0609_ VGND VGND VPWR VPWR _0610_ sky130_fd_sc_hd__clkbuf_2
XFILLER_0_12_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3465_ cu.reg_file.reg_e\[1\] _0480_ _0487_ VGND VGND VPWR VPWR _0541_ sky130_fd_sc_hd__and3_1
X_6253_ clknet_leaf_0_clk _0235_ net154 VGND VGND VPWR VPWR cu.reg_file.reg_sp\[9\]
+ sky130_fd_sc_hd__dfstp_2
X_5204_ mc.cc.count\[1\] _2118_ _2120_ mc.cc.count\[2\] VGND VGND VPWR VPWR _2123_
+ sky130_fd_sc_hd__o211a_1
X_6184_ clknet_leaf_34_clk net198 net162 VGND VGND VPWR VPWR ih.interrupt_source\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_3396_ _2918_ _0355_ _0470_ _2902_ _0471_ VGND VGND VPWR VPWR _0472_ sky130_fd_sc_hd__o221a_1
XANTENNA_fanout193_A net194 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5135_ _1213_ _1160_ _2066_ VGND VGND VPWR VPWR _2077_ sky130_fd_sc_hd__mux2_1
X_5066_ cu.reg_file.reg_c\[5\] _1191_ _2025_ VGND VGND VPWR VPWR _2031_ sky130_fd_sc_hd__mux2_1
XANTENNA__5273__A1 _1051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4017_ _0770_ _0773_ VGND VGND VPWR VPWR _1091_ sky130_fd_sc_hd__nand2_1
XFILLER_0_79_478 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5025__A1 _1622_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5576__A2 _2236_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5968_ cu.id.imm_i\[15\] _2486_ _2686_ VGND VGND VPWR VPWR _2694_ sky130_fd_sc_hd__mux2_1
X_4919_ _1910_ _1911_ VGND VGND VPWR VPWR _1912_ sky130_fd_sc_hd__xor2_1
XFILLER_0_47_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5899_ ih.t.timer_max\[18\] _1074_ _2654_ VGND VGND VPWR VPWR _2657_ sky130_fd_sc_hd__mux2_1
XFILLER_0_7_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_35_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3511__A1 _0576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5264__A1 _2165_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3814__A2 _0740_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3750__B2 cu.reg_file.reg_sp\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_404 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3250_ _2899_ _2900_ VGND VGND VPWR VPWR _0326_ sky130_fd_sc_hd__nand2_1
XTAP_426 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3181_ _2916_ _2917_ VGND VGND VPWR VPWR _2918_ sky130_fd_sc_hd__nand2b_4
XTAP_459 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3502__A1 cu.reg_file.reg_b\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3502__B2 cu.reg_file.reg_a\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5822_ _2603_ VGND VGND VPWR VPWR _0236_ sky130_fd_sc_hd__clkbuf_1
X_5753_ _2541_ _2542_ VGND VGND VPWR VPWR _2543_ sky130_fd_sc_hd__and2_1
X_4704_ _1720_ _1721_ _1672_ VGND VGND VPWR VPWR _1722_ sky130_fd_sc_hd__and3b_1
X_2965_ _2704_ _2699_ VGND VGND VPWR VPWR _2705_ sky130_fd_sc_hd__nor2_1
XFILLER_0_60_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5684_ _2494_ _1643_ cu.reg_file.reg_mem\[9\] _1646_ VGND VGND VPWR VPWR _2495_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_60_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4635_ _1672_ _1673_ _1674_ VGND VGND VPWR VPWR _1675_ sky130_fd_sc_hd__and3_1
XFILLER_0_32_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4566_ _1356_ _1614_ VGND VGND VPWR VPWR _1619_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6305_ clknet_leaf_6_clk _0287_ net164 VGND VGND VPWR VPWR cu.id.imm_i\[10\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_12_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3517_ cu.reg_file.reg_l\[1\] _0422_ _0592_ VGND VGND VPWR VPWR _0593_ sky130_fd_sc_hd__a21o_1
X_4497_ cu.reg_file.reg_d\[4\] _1282_ _1286_ cu.reg_file.reg_sp\[12\] VGND VGND VPWR
+ VPWR _1553_ sky130_fd_sc_hd__a22o_1
X_6236_ clknet_leaf_15_clk ih.t.next_count\[24\] net179 VGND VGND VPWR VPWR ih.t.count\[24\]
+ sky130_fd_sc_hd__dfrtp_1
X_3448_ _0372_ _0522_ _0523_ _0387_ _2918_ VGND VGND VPWR VPWR _0524_ sky130_fd_sc_hd__a311o_1
XTAP_971 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_960 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3379_ _0298_ _2923_ _2901_ VGND VGND VPWR VPWR _0455_ sky130_fd_sc_hd__or3_1
X_6167_ clknet_leaf_2_clk _0201_ net155 VGND VGND VPWR VPWR cu.reg_file.reg_mem\[3\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_85_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_993 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_982 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5118_ _2064_ VGND VGND VPWR VPWR _0071_ sky130_fd_sc_hd__clkbuf_1
X_6098_ clknet_leaf_6_clk _0132_ net164 VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__dfrtp_4
X_5049_ _1260_ _1263_ _2002_ VGND VGND VPWR VPWR _2020_ sky130_fd_sc_hd__mux2_1
XFILLER_0_39_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5549__A2 _1649_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5329__A _2204_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_62_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_518 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_50_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output125_A net125 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3312__A cu.id.cb_opcode_x\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4408__A cu.reg_file.reg_l\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5938__S _2666_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3420__B1 _0495_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4143__A _0516_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4420_ _1440_ _1462_ _1473_ _1332_ VGND VGND VPWR VPWR _1480_ sky130_fd_sc_hd__a31o_1
XFILLER_0_1_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4920__A0 _1623_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4250__D_N _2936_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_540 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4351_ _1306_ _1410_ _1414_ VGND VGND VPWR VPWR _1415_ sky130_fd_sc_hd__o21a_4
X_4282_ _1332_ _1348_ VGND VGND VPWR VPWR _1349_ sky130_fd_sc_hd__xnor2_1
X_3302_ _2892_ _2894_ VGND VGND VPWR VPWR _0378_ sky130_fd_sc_hd__and2b_1
XTAP_201 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_212 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_223 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6021_ clknet_leaf_30_clk _0059_ net183 VGND VGND VPWR VPWR cu.reg_file.reg_d\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_3233_ cu.id.opcode\[1\] cu.id.opcode\[6\] cu.id.opcode\[7\] cu.id.opcode\[2\] VGND
+ VGND VPWR VPWR _0309_ sky130_fd_sc_hd__and4b_1
XTAP_256 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3487__B1 _0498_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3164_ _2899_ _2875_ _2876_ _2900_ VGND VGND VPWR VPWR _2901_ sky130_fd_sc_hd__or4b_4
X_3095_ ih.t.timer_max\[5\] _2749_ VGND VGND VPWR VPWR _2833_ sky130_fd_sc_hd__xor2_1
XFILLER_0_76_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5400__A1 net131 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3997_ _0588_ _1044_ _1061_ _0610_ _1045_ VGND VGND VPWR VPWR _1071_ sky130_fd_sc_hd__o221a_1
XANTENNA__5149__A _2951_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5805_ cu.reg_file.reg_sp\[8\] _2588_ _2539_ VGND VGND VPWR VPWR _2589_ sky130_fd_sc_hd__mux2_1
X_5736_ net24 _2519_ _2528_ VGND VGND VPWR VPWR _0225_ sky130_fd_sc_hd__a21o_1
XANTENNA__4053__A _1110_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5667_ mc.cl.next_data\[7\] _2313_ net141 _2479_ VGND VGND VPWR VPWR _2480_ sky130_fd_sc_hd__a22o_1
XFILLER_0_72_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4988__A cu.pc.pc_o\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4618_ _1660_ VGND VGND VPWR VPWR _1661_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__3892__A _0379_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5598_ net88 _1330_ VGND VGND VPWR VPWR _2414_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4549_ _1581_ _1601_ _1588_ VGND VGND VPWR VPWR _1603_ sky130_fd_sc_hd__nand3_1
XFILLER_0_96_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_6219_ clknet_leaf_11_clk ih.t.next_count\[7\] net176 VGND VGND VPWR VPWR ih.t.count\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__5612__A _1649_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_790 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2971__A net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3134__B_N _2869_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5458__A1 _2085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5630__A1 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3977__A _1051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3920_ _0995_ VGND VGND VPWR VPWR _0996_ sky130_fd_sc_hd__inv_2
XFILLER_0_25_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3696__B _0528_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3851_ _0866_ _0925_ _0926_ VGND VGND VPWR VPWR _0927_ sky130_fd_sc_hd__o21a_1
XANTENNA__5394__A0 _1190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3782_ cu.reg_file.reg_b\[4\] _0743_ _0624_ cu.reg_file.reg_sp\[12\] VGND VGND VPWR
+ VPWR _0858_ sky130_fd_sc_hd__a22o_1
X_5521_ _2337_ _2338_ _2339_ _2340_ _1369_ VGND VGND VPWR VPWR _2341_ sky130_fd_sc_hd__a32o_1
XFILLER_0_14_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_26_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5697__A1 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5452_ net71 _1638_ _2279_ net70 VGND VGND VPWR VPWR _2280_ sky130_fd_sc_hd__a22o_1
X_5383_ _1369_ _2191_ VGND VGND VPWR VPWR _2235_ sky130_fd_sc_hd__nor2_1
X_4403_ cu.reg_file.reg_a\[7\] _1276_ _1287_ cu.reg_file.reg_sp\[7\] VGND VGND VPWR
+ VPWR _1464_ sky130_fd_sc_hd__a22o_1
X_4334_ _1397_ _1394_ _1383_ VGND VGND VPWR VPWR _1399_ sky130_fd_sc_hd__a21o_1
XANTENNA__3217__A cu.id.starting_int_service VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4265_ _1332_ VGND VGND VPWR VPWR _1333_ sky130_fd_sc_hd__clkbuf_4
X_6004_ clknet_leaf_18_clk _0042_ net185 VGND VGND VPWR VPWR cu.reg_file.reg_b\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_3216_ _2896_ _2952_ VGND VGND VPWR VPWR _2953_ sky130_fd_sc_hd__nand2_2
X_4196_ cu.alu_f\[7\] _1027_ _1184_ VGND VGND VPWR VPWR _1265_ sky130_fd_sc_hd__and3_1
X_3147_ cu.id.alu_opcode\[3\] VGND VGND VPWR VPWR _2884_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3078_ _2754_ _2814_ ih.t.count\[12\] VGND VGND VPWR VPWR _2816_ sky130_fd_sc_hd__a21oi_1
XANTENNA__5621__A1 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5621__B2 _2435_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3887__A _0824_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3632__B1 _0492_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_49_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4188__A1 _1256_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3935__A1 _0986_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5719_ _2514_ _2519_ _2520_ _2518_ VGND VGND VPWR VPWR _0216_ sky130_fd_sc_hd__a22o_1
XFILLER_0_32_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5688__B2 _1646_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4112__A1 _1027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5860__A1 _1667_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4179__A1 _0545_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5517__A net32 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4050_ _1120_ _1096_ _1097_ _0754_ _1123_ VGND VGND VPWR VPWR _1124_ sky130_fd_sc_hd__o221a_1
XANTENNA__4103__A1 _0547_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3001_ net74 VGND VGND VPWR VPWR _2739_ sky130_fd_sc_hd__inv_2
Xinput6 keypad_input[13] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_4
XANTENNA__5603__A1 ih.t.timer_max\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5398__S _2237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4952_ _1213_ _1941_ _1795_ VGND VGND VPWR VPWR _1942_ sky130_fd_sc_hd__mux2_1
XANTENNA__3614__B1 _0502_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4883_ _1877_ _1878_ VGND VGND VPWR VPWR _1879_ sky130_fd_sc_hd__xor2_1
XFILLER_0_46_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3903_ _0308_ _0525_ _0977_ _0978_ VGND VGND VPWR VPWR _0979_ sky130_fd_sc_hd__and4b_1
XFILLER_0_19_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5367__A0 _0619_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3834_ _0856_ _0908_ _0909_ VGND VGND VPWR VPWR _0910_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_345 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3765_ cu.reg_file.reg_mem\[14\] _0640_ _0839_ _0840_ VGND VGND VPWR VPWR _0841_
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_42_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5504_ _1374_ _1625_ _1630_ _1489_ _1417_ VGND VGND VPWR VPWR _2324_ sky130_fd_sc_hd__a2111oi_4
X_3696_ _0512_ _0528_ VGND VGND VPWR VPWR _0772_ sky130_fd_sc_hd__and2_1
XFILLER_0_14_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5435_ _2022_ net72 _2266_ VGND VGND VPWR VPWR _2267_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4342__A1 cu.reg_file.reg_a\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5366_ _2181_ _2225_ VGND VGND VPWR VPWR _2226_ sky130_fd_sc_hd__nand2_4
XANTENNA__4342__B2 cu.reg_file.reg_sp\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4317_ _1370_ _1375_ _1381_ _1382_ VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__a22o_1
X_5297_ _1188_ net87 _2182_ VGND VGND VPWR VPWR _2186_ sky130_fd_sc_hd__mux2_1
X_4248_ _1309_ _1311_ VGND VGND VPWR VPWR _1316_ sky130_fd_sc_hd__nor2b_2
X_4179_ _0574_ _0545_ _0447_ VGND VGND VPWR VPWR _1249_ sky130_fd_sc_hd__mux2_1
XFILLER_0_96_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1038 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1027 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1016 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1005 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1049 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5358__A0 _1192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_33_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3136__A2 _2869_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5800__A cu.reg_file.reg_sp\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5011__S _0368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3320__A _0373_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5946__S _2666_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4135__B _0779_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_90 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_24_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3550_ cu.reg_file.reg_d\[6\] _0492_ _0625_ cu.alu_f\[6\] VGND VGND VPWR VPWR _0626_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_36_292 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5220_ _2132_ VGND VGND VPWR VPWR _0105_ sky130_fd_sc_hd__clkbuf_1
X_3481_ _0556_ VGND VGND VPWR VPWR _0557_ sky130_fd_sc_hd__inv_2
XFILLER_0_47_31 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5151_ cu.reg_file.reg_l\[0\] _2085_ _2088_ VGND VGND VPWR VPWR _2089_ sky130_fd_sc_hd__mux2_1
X_5082_ _2042_ VGND VGND VPWR VPWR _0057_ sky130_fd_sc_hd__clkbuf_1
X_4102_ _0829_ _1175_ VGND VGND VPWR VPWR _1176_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4033_ _0822_ _0632_ _0566_ _0531_ VGND VGND VPWR VPWR _1107_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5984_ clknet_leaf_28_clk _0022_ net188 VGND VGND VPWR VPWR cu.pc.pc_o\[6\] sky130_fd_sc_hd__dfrtp_4
X_4935_ _1917_ _1926_ _1808_ VGND VGND VPWR VPWR _1927_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_22 net61 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_11 memory_data_in[7] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4866_ _0373_ cu.pc.pc_o\[5\] VGND VGND VPWR VPWR _1863_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4797_ _1798_ VGND VGND VPWR VPWR _1799_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_6_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3817_ cu.reg_file.reg_sp\[9\] _0636_ _0748_ cu.reg_file.reg_h\[1\] VGND VGND VPWR
+ VPWR _0893_ sky130_fd_sc_hd__a22o_1
X_3748_ _0384_ _0392_ _0400_ VGND VGND VPWR VPWR _0824_ sky130_fd_sc_hd__and3_2
XFILLER_0_6_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3679_ _0684_ VGND VGND VPWR VPWR _0755_ sky130_fd_sc_hd__inv_2
X_5418_ _2255_ VGND VGND VPWR VPWR _0180_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5349_ _2216_ VGND VGND VPWR VPWR _0150_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4935__S _1808_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3287__D1 _0296_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4554__B2 cu.reg_file.reg_h\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_608 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3817__B1 _0748_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2981_ _2715_ ih.ih.ih.prev_data\[6\] _2716_ ih.ih.ih.prev_data\[12\] _2719_ VGND
+ VGND VPWR VPWR _2720_ sky130_fd_sc_hd__o221a_1
XFILLER_0_33_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4720_ ih.t.count\[28\] ih.t.count\[29\] _1729_ VGND VGND VPWR VPWR _1732_ sky130_fd_sc_hd__and3_1
Xclkbuf_leaf_41_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_41_clk sky130_fd_sc_hd__clkbuf_16
X_4651_ ih.t.count\[6\] _1683_ VGND VGND VPWR VPWR _1686_ sky130_fd_sc_hd__and2_1
XFILLER_0_83_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput20 memory_data_in[2] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_4
Xinput31 programmable_gpio_in[4] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__buf_2
X_3602_ cu.pc.pc_o\[4\] _0501_ _0499_ cu.reg_file.reg_a\[4\] _0504_ VGND VGND VPWR
+ VPWR _0678_ sky130_fd_sc_hd__a221o_1
X_4582_ _1579_ VGND VGND VPWR VPWR _1626_ sky130_fd_sc_hd__inv_2
XFILLER_0_12_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3533_ _0548_ _0393_ _0529_ VGND VGND VPWR VPWR _0609_ sky130_fd_sc_hd__or3_1
X_3464_ cu.reg_file.reg_a\[1\] _0499_ VGND VGND VPWR VPWR _0540_ sky130_fd_sc_hd__and2_1
X_6252_ clknet_leaf_0_clk _0234_ net154 VGND VGND VPWR VPWR cu.reg_file.reg_sp\[8\]
+ sky130_fd_sc_hd__dfstp_4
X_5203_ mc.cc.count\[2\] mc.cc.count\[1\] _2118_ VGND VGND VPWR VPWR _2122_ sky130_fd_sc_hd__nor3_1
X_6183_ clknet_leaf_23_clk _0216_ net193 VGND VGND VPWR VPWR mc.count sky130_fd_sc_hd__dfrtp_4
X_5134_ _2076_ VGND VGND VPWR VPWR _0075_ sky130_fd_sc_hd__clkbuf_1
X_3395_ _2878_ _0402_ _0301_ VGND VGND VPWR VPWR _0471_ sky130_fd_sc_hd__a21o_1
XANTENNA__5440__A _2139_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5065_ _2030_ VGND VGND VPWR VPWR _0052_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3808__B1 _0429_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4016_ _1073_ _1089_ VGND VGND VPWR VPWR _1090_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_28_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4481__B1 _1284_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5967_ _2693_ VGND VGND VPWR VPWR _0291_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4918_ _1899_ _1902_ VGND VGND VPWR VPWR _1911_ sky130_fd_sc_hd__or2b_1
XFILLER_0_35_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xclkbuf_leaf_32_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_32_clk sky130_fd_sc_hd__clkbuf_16
X_5898_ _2656_ VGND VGND VPWR VPWR _0259_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4849_ _1840_ _1847_ _1809_ VGND VGND VPWR VPWR _1848_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4536__A1 cu.reg_file.reg_d\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5543__A_N _1400_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_23_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_23_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_26_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_38_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3983__C1 _1027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4413__B _1473_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3750__A2 _0743_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_405 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_449 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3180_ _2899_ _2900_ _2875_ _2876_ VGND VGND VPWR VPWR _2917_ sky130_fd_sc_hd__and4b_2
XFILLER_0_28_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3699__B _0547_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5821_ cu.reg_file.reg_sp\[10\] _2602_ _2539_ VGND VGND VPWR VPWR _2603_ sky130_fd_sc_hd__mux2_1
X_2964_ _2695_ mc.rw.state\[0\] VGND VGND VPWR VPWR _2704_ sky130_fd_sc_hd__and2_1
XFILLER_0_60_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5752_ cu.reg_file.reg_sp\[2\] _2534_ VGND VGND VPWR VPWR _2542_ sky130_fd_sc_hd__or2_1
X_4703_ ih.t.count\[21\] ih.t.count\[22\] _1714_ ih.t.count\[23\] VGND VGND VPWR VPWR
+ _1721_ sky130_fd_sc_hd__a31o_1
Xclkbuf_leaf_14_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_14_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_17_538 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_29_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5683_ mc.cl.next_data\[9\] _2359_ _2490_ _2493_ VGND VGND VPWR VPWR _2494_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_17_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4634_ ih.t.count\[0\] ih.t.count\[1\] VGND VGND VPWR VPWR _1674_ sky130_fd_sc_hd__or2_1
XANTENNA__4518__B2 cu.pc.pc_o\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4565_ _1567_ _1579_ _1598_ VGND VGND VPWR VPWR _1618_ sky130_fd_sc_hd__or3b_1
X_6304_ clknet_leaf_6_clk _0286_ net164 VGND VGND VPWR VPWR cu.id.imm_i\[9\] sky130_fd_sc_hd__dfrtp_4
X_3516_ cu.reg_file.reg_b\[1\] _0432_ _0433_ cu.reg_file.reg_a\[1\] VGND VGND VPWR
+ VPWR _0592_ sky130_fd_sc_hd__a22o_1
X_4496_ _1351_ _1550_ _1551_ _1371_ _1552_ VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__a221o_1
X_6235_ clknet_leaf_15_clk ih.t.next_count\[23\] net179 VGND VGND VPWR VPWR ih.t.count\[23\]
+ sky130_fd_sc_hd__dfrtp_1
X_3447_ _0373_ cu.id.cb_opcode_y\[0\] VGND VGND VPWR VPWR _0523_ sky130_fd_sc_hd__or2_1
XANTENNA_clkbuf_leaf_15_clk_A clknet_2_2__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_961 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_950 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3378_ _0379_ _0450_ _0451_ _0453_ VGND VGND VPWR VPWR _0454_ sky130_fd_sc_hd__or4b_2
X_6166_ clknet_leaf_2_clk _0200_ net155 VGND VGND VPWR VPWR cu.reg_file.reg_mem\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_994 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_983 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_972 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6097_ clknet_leaf_26_clk _0131_ net195 VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__dfrtp_2
X_5117_ cu.reg_file.reg_e\[7\] _1260_ _2056_ VGND VGND VPWR VPWR _2064_ sky130_fd_sc_hd__mux2_1
X_5048_ _2019_ VGND VGND VPWR VPWR _0046_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4206__B1 _0293_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_62_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3312__B _0387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output118_A net118 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5954__S _2686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3420__A1 cu.reg_file.reg_sp\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3420__B2 cu.reg_file.reg_h\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5173__A1 net20 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4350_ cu.reg_file.reg_c\[4\] _1313_ _1411_ _1413_ VGND VGND VPWR VPWR _1414_ sky130_fd_sc_hd__a211o_2
X_3301_ _0371_ _0376_ VGND VGND VPWR VPWR _0377_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4281_ _1340_ _1341_ _1347_ VGND VGND VPWR VPWR _1348_ sky130_fd_sc_hd__o21a_2
XTAP_202 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_224 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6020_ clknet_leaf_18_clk _0058_ net184 VGND VGND VPWR VPWR cu.reg_file.reg_d\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_257 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3232_ _2902_ _0304_ _0307_ VGND VGND VPWR VPWR _0308_ sky130_fd_sc_hd__o21ai_2
XTAP_235 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3487__A1 cu.pc.pc_o\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_3_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_3_clk sky130_fd_sc_hd__clkbuf_16
X_3163_ cu.id.opcode\[1\] VGND VGND VPWR VPWR _2900_ sky130_fd_sc_hd__buf_2
XTAP_279 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3094_ _2750_ _2830_ ih.t.count\[6\] VGND VGND VPWR VPWR _2832_ sky130_fd_sc_hd__a21oi_1
XANTENNA__5421__C _1369_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5936__A0 _0343_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5804_ _1622_ _2587_ _2545_ VGND VGND VPWR VPWR _2588_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3996_ _0570_ _0759_ _1068_ _1069_ VGND VGND VPWR VPWR _1070_ sky130_fd_sc_hd__o22a_1
X_5735_ _2518_ mc.cl.next_data\[6\] _2111_ VGND VGND VPWR VPWR _2528_ sky130_fd_sc_hd__and3_1
XFILLER_0_17_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4053__B _1126_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5666_ _1665_ _2477_ _2478_ VGND VGND VPWR VPWR _2479_ sky130_fd_sc_hd__o21a_1
XFILLER_0_72_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4617_ _0315_ _1658_ _1659_ VGND VGND VPWR VPWR _1660_ sky130_fd_sc_hd__nor3b_4
X_5597_ net96 _2194_ _2412_ VGND VGND VPWR VPWR _2413_ sky130_fd_sc_hd__a21o_1
X_4548_ _1581_ _1588_ _1601_ VGND VGND VPWR VPWR _1602_ sky130_fd_sc_hd__a21o_1
Xmax_cap150 net238 VGND VGND VPWR VPWR net150 sky130_fd_sc_hd__clkbuf_2
X_4479_ _1382_ _1532_ _1533_ _1536_ VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__a31o_1
X_6218_ clknet_leaf_11_clk ih.t.next_count\[6\] net176 VGND VGND VPWR VPWR ih.t.count\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_6149_ clknet_leaf_8_clk _0183_ net168 VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__dfrtp_4
XTAP_791 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4427__B1 _1284_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3650__B2 cu.reg_file.reg_e\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5975__RESET_B net161 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_430 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3953__A2 _0619_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5155__A1 _1074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5014__S _0368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_500 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5630__A2 _1648_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3850_ _0861_ _0864_ VGND VGND VPWR VPWR _0926_ sky130_fd_sc_hd__or2b_1
XANTENNA__5394__A1 net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4197__A2 _1261_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3781_ cu.reg_file.reg_d\[4\] _0488_ _0741_ cu.reg_file.reg_h\[4\] VGND VGND VPWR
+ VPWR _0857_ sky130_fd_sc_hd__a22o_1
XFILLER_0_41_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5520_ net28 net30 net27 net29 _1354_ _1330_ VGND VGND VPWR VPWR _2340_ sky130_fd_sc_hd__mux4_1
XFILLER_0_54_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5451_ _1335_ _1372_ VGND VGND VPWR VPWR _2279_ sky130_fd_sc_hd__nor2_1
XFILLER_0_41_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5382_ _2234_ VGND VGND VPWR VPWR _0165_ sky130_fd_sc_hd__clkbuf_1
X_4402_ _1333_ _1462_ _1457_ VGND VGND VPWR VPWR _1463_ sky130_fd_sc_hd__o21a_1
XANTENNA__5697__A2 _1650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4333_ _1395_ _1397_ VGND VGND VPWR VPWR _1398_ sky130_fd_sc_hd__or2b_1
XFILLER_0_67_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4264_ _1331_ VGND VGND VPWR VPWR _1332_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_1_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6003_ clknet_leaf_4_clk _0041_ net170 VGND VGND VPWR VPWR cu.reg_file.reg_b\[1\]
+ sky130_fd_sc_hd__dfrtp_4
X_3215_ _2938_ _2932_ VGND VGND VPWR VPWR _2952_ sky130_fd_sc_hd__or2_2
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4195_ _0516_ _1260_ _1263_ _1027_ VGND VGND VPWR VPWR _1264_ sky130_fd_sc_hd__a22o_1
X_3146_ cu.id.alu_opcode\[1\] VGND VGND VPWR VPWR _2883_ sky130_fd_sc_hd__inv_2
X_3077_ ih.t.count\[12\] _2754_ _2814_ VGND VGND VPWR VPWR _2815_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5621__A2 _1633_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_77_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3632__A1 cu.reg_file.reg_sp\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3632__B2 cu.reg_file.reg_d\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5604__A_N _1400_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_92_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_227 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5718_ _2351_ _2514_ VGND VGND VPWR VPWR _2520_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3979_ _0372_ _0371_ _0774_ _1019_ _1053_ VGND VGND VPWR VPWR _1054_ sky130_fd_sc_hd__o2111a_1
XANTENNA__5594__S _2351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4511__B _1561_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5649_ _2169_ _2455_ _2462_ _2136_ VGND VGND VPWR VPWR _2463_ sky130_fd_sc_hd__o211a_1
XFILLER_0_32_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3143__A _2878_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4112__A2 _1075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5860__A2 _2194_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2982__A net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3623__A1 cu.reg_file.reg_mem\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3623__B2 cu.reg_file.reg_a\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_363 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_525 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5517__B _1330_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4887__A0 cu.pc.pc_o\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output62_A net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3000_ net71 net30 ih.gpio_interrupt_mask\[3\] VGND VGND VPWR VPWR _2738_ sky130_fd_sc_hd__and3b_1
Xinput7 keypad_input[14] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_4
XANTENNA__5603__A2 _2193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4951_ _1939_ _1940_ VGND VGND VPWR VPWR _1941_ sky130_fd_sc_hd__nor2_1
XANTENNA__3614__B2 cu.reg_file.reg_b\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3614__A1 cu.pc.pc_o\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4882_ _1863_ _1866_ _1864_ VGND VGND VPWR VPWR _1878_ sky130_fd_sc_hd__o21a_1
X_3902_ _2886_ _0965_ _0521_ _0359_ VGND VGND VPWR VPWR _0978_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_46_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3833_ _0850_ _0853_ VGND VGND VPWR VPWR _0909_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3764_ cu.reg_file.reg_b\[6\] _0426_ _0429_ cu.reg_file.reg_d\[6\] VGND VGND VPWR
+ VPWR _0840_ sky130_fd_sc_hd__a22o_1
X_5503_ _1661_ _2318_ _2322_ VGND VGND VPWR VPWR _2323_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_14_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3695_ _0768_ _0770_ _0753_ VGND VGND VPWR VPWR _0771_ sky130_fd_sc_hd__or3b_1
XFILLER_0_42_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5434_ _2139_ _2147_ VGND VGND VPWR VPWR _2266_ sky130_fd_sc_hd__nand2_1
XANTENNA__3228__A _2936_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5443__A _2139_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5365_ _2224_ VGND VGND VPWR VPWR _2225_ sky130_fd_sc_hd__buf_4
XFILLER_0_58_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4316_ _1351_ VGND VGND VPWR VPWR _1382_ sky130_fd_sc_hd__clkbuf_4
X_5296_ _2185_ VGND VGND VPWR VPWR _0128_ sky130_fd_sc_hd__clkbuf_1
X_4247_ _1314_ VGND VGND VPWR VPWR _1315_ sky130_fd_sc_hd__buf_2
X_4178_ _1246_ _1247_ _0600_ VGND VGND VPWR VPWR _1248_ sky130_fd_sc_hd__mux2_1
X_3129_ ih.t.count\[30\] _2866_ VGND VGND VPWR VPWR _2867_ sky130_fd_sc_hd__nor2_1
XANTENNA__5055__B1 _2951_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4506__B _1561_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1028 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1017 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1006 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1039 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5358__A1 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4225__C _1269_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5618__A net89 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2977__A net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5046__A0 _1193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5597__A1 net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output100_A net100 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3320__B _0374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5962__S _2686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3480_ _0550_ _0555_ VGND VGND VPWR VPWR _0556_ sky130_fd_sc_hd__nand2_1
XFILLER_0_24_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5521__B2 _1369_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5150_ _2087_ VGND VGND VPWR VPWR _2088_ sky130_fd_sc_hd__clkbuf_4
X_5081_ cu.reg_file.reg_d\[1\] _2041_ _2039_ VGND VGND VPWR VPWR _2042_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_43 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4101_ _0918_ _0948_ _1172_ _1174_ VGND VGND VPWR VPWR _1175_ sky130_fd_sc_hd__a2bb2o_2
XFILLER_0_44_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5285__A0 net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4032_ alu.Cin _0554_ _0556_ _0509_ VGND VGND VPWR VPWR _1106_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__5037__A0 _1187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5983_ clknet_leaf_28_clk _0021_ net188 VGND VGND VPWR VPWR cu.pc.pc_o\[5\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_59_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4934_ _1924_ _1925_ _1798_ VGND VGND VPWR VPWR _1926_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4260__A1 cu.reg_file.reg_c\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_12 programmable_gpio_in[0] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_23 net61 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4865_ _1860_ _1861_ VGND VGND VPWR VPWR _1862_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4796_ _2948_ _1797_ VGND VGND VPWR VPWR _1798_ sky130_fd_sc_hd__nand2_8
XFILLER_0_27_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3816_ cu.id.imm_i\[9\] _0739_ _0891_ _0653_ VGND VGND VPWR VPWR _0892_ sky130_fd_sc_hd__a22oi_4
X_3747_ _0574_ _0558_ _0822_ _0566_ VGND VGND VPWR VPWR _0823_ sky130_fd_sc_hd__a22o_1
XFILLER_0_15_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_70_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_15_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3771__B1 _0624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3678_ _0645_ _0722_ VGND VGND VPWR VPWR _0754_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5417_ _1194_ net138 _2248_ VGND VGND VPWR VPWR _2255_ sky130_fd_sc_hd__mux2_1
Xoutput130 net130 VGND VGND VPWR VPWR ss6[6] sky130_fd_sc_hd__buf_2
XANTENNA__5512__B2 net66 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5512__A1 net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5348_ _0619_ net108 _2215_ VGND VGND VPWR VPWR _2216_ sky130_fd_sc_hd__mux2_1
X_5279_ net80 _1189_ _2170_ VGND VGND VPWR VPWR _2175_ sky130_fd_sc_hd__mux2_1
XANTENNA__5028__B1 _2951_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5579__B2 _1401_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5579__A1 net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_61_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5503__A1 _1661_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3514__B1 _0415_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_609 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3817__B2 cu.reg_file.reg_h\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3817__A1 cu.reg_file.reg_sp\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_17_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_447 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2980_ _2717_ ih.ih.ih.prev_data\[4\] _2718_ ih.ih.ih.prev_data\[13\] VGND VGND VPWR
+ VPWR _2719_ sky130_fd_sc_hd__o22a_1
XFILLER_0_56_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4242__A1 _2908_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3450__C1 _2935_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4650_ _1685_ VGND VGND VPWR VPWR ih.t.next_count\[5\] sky130_fd_sc_hd__clkbuf_1
XANTENNA__4162__A _1209_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput21 memory_data_in[3] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_2
Xinput10 keypad_input[2] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_2
X_3601_ cu.reg_file.reg_b\[4\] _0502_ _0494_ cu.reg_file.reg_mem\[4\] _0676_ VGND
+ VGND VPWR VPWR _0677_ sky130_fd_sc_hd__a221o_1
Xinput32 programmable_gpio_in[5] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__buf_1
X_4581_ _1329_ _1372_ VGND VGND VPWR VPWR _1625_ sky130_fd_sc_hd__nand2_4
XFILLER_0_3_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3532_ _0574_ _0604_ _0607_ VGND VGND VPWR VPWR _0608_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3463_ _0480_ _0493_ VGND VGND VPWR VPWR _0539_ sky130_fd_sc_hd__and2_2
X_6251_ clknet_leaf_0_clk _0233_ net155 VGND VGND VPWR VPWR cu.reg_file.reg_sp\[7\]
+ sky130_fd_sc_hd__dfrtp_4
X_5202_ net228 _2118_ _2121_ VGND VGND VPWR VPWR _0098_ sky130_fd_sc_hd__a21o_1
X_6182_ clknet_leaf_18_clk _0215_ net173 VGND VGND VPWR VPWR ih.input_handler_enable
+ sky130_fd_sc_hd__dfrtp_1
X_5133_ _2075_ cu.reg_file.reg_h\[3\] _2069_ VGND VGND VPWR VPWR _2076_ sky130_fd_sc_hd__mux2_1
X_3394_ _0378_ _0309_ VGND VGND VPWR VPWR _0470_ sky130_fd_sc_hd__nand2_1
X_5064_ cu.reg_file.reg_c\[4\] _1189_ _2025_ VGND VGND VPWR VPWR _2030_ sky130_fd_sc_hd__mux2_1
XANTENNA__3808__A1 cu.reg_file.reg_b\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3808__B2 cu.reg_file.reg_d\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_403 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5440__B _2236_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4015_ _1081_ _1082_ _1085_ _1088_ VGND VGND VPWR VPWR _1089_ sky130_fd_sc_hd__or4_4
XFILLER_0_74_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4481__B2 cu.reg_file.reg_h\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4481__A1 cu.reg_file.reg_b\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5966_ cu.id.imm_i\[14\] _2467_ _2686_ VGND VGND VPWR VPWR _2693_ sky130_fd_sc_hd__mux2_1
X_5897_ ih.t.timer_max\[17\] _1051_ _2654_ VGND VGND VPWR VPWR _2656_ sky130_fd_sc_hd__mux2_1
X_4917_ _2920_ cu.pc.pc_o\[9\] VGND VGND VPWR VPWR _1910_ sky130_fd_sc_hd__xor2_1
X_4848_ _1845_ _1846_ _1799_ VGND VGND VPWR VPWR _1847_ sky130_fd_sc_hd__mux2_1
XFILLER_0_62_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_463 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4779_ _1775_ _1779_ VGND VGND VPWR VPWR _1784_ sky130_fd_sc_hd__nand2_1
XFILLER_0_43_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_30_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4946__S _1808_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2990__A net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4527__A2 _1561_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5724__A1 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_406 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5017__S _0368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_417 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_428 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5660__B1 _2225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5820_ _1226_ _2601_ _2545_ VGND VGND VPWR VPWR _2602_ sky130_fd_sc_hd__mux2_1
XFILLER_0_91_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_2963_ _2703_ VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__clkbuf_1
X_5751_ cu.reg_file.reg_sp\[2\] _2534_ VGND VGND VPWR VPWR _2541_ sky130_fd_sc_hd__nand2_1
X_4702_ ih.t.count\[22\] ih.t.count\[23\] _1717_ VGND VGND VPWR VPWR _1720_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5682_ ih.t.timer_max\[25\] _2151_ _2320_ ih.t.timer_max\[9\] VGND VGND VPWR VPWR
+ _2493_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_44_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4633_ ih.t.count\[0\] ih.t.count\[1\] VGND VGND VPWR VPWR _1673_ sky130_fd_sc_hd__nand2_1
XFILLER_0_44_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4564_ _1599_ _1602_ _1615_ VGND VGND VPWR VPWR _1617_ sky130_fd_sc_hd__nand3_1
XFILLER_0_69_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6040__RESET_B net161 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6303_ clknet_leaf_18_clk _0285_ net184 VGND VGND VPWR VPWR cu.id.imm_i\[8\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_52_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_12_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3515_ cu.reg_file.reg_sp\[1\] _0413_ _0419_ cu.reg_file.reg_h\[1\] _0590_ VGND VGND
+ VPWR VPWR _0591_ sky130_fd_sc_hd__a221o_1
XFILLER_0_40_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6234_ clknet_leaf_14_clk ih.t.next_count\[22\] net180 VGND VGND VPWR VPWR ih.t.count\[22\]
+ sky130_fd_sc_hd__dfrtp_1
X_4495_ _1402_ _1545_ VGND VGND VPWR VPWR _1552_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3446_ _0373_ cu.id.cb_opcode_y\[0\] VGND VGND VPWR VPWR _0522_ sky130_fd_sc_hd__nand2_1
XTAP_962 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_951 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_940 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5451__A _1335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3377_ _0452_ _0303_ VGND VGND VPWR VPWR _0453_ sky130_fd_sc_hd__nor2_1
X_6165_ clknet_leaf_2_clk _0199_ net155 VGND VGND VPWR VPWR cu.reg_file.reg_mem\[1\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_40_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_995 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_984 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_973 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6096_ clknet_leaf_7_clk _0130_ net165 VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__dfrtp_2
X_5116_ _2063_ VGND VGND VPWR VPWR _0070_ sky130_fd_sc_hd__clkbuf_1
X_5047_ cu.reg_file.reg_b\[6\] _2018_ _2006_ VGND VGND VPWR VPWR _2019_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5954__A1 _2350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5949_ _2683_ VGND VGND VPWR VPWR _0283_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5706__B2 ih.t.timer_max\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_7_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_328 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3193__A1 _2918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5890__A0 _1193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2985__A net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4445__A1 cu.reg_file.reg_b\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4445__B2 cu.reg_file.reg_d\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3956__B1 _0773_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output92_A net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3300_ _0372_ _2921_ _0375_ VGND VGND VPWR VPWR _0376_ sky130_fd_sc_hd__and3_1
X_4280_ cu.reg_file.reg_c\[1\] _1313_ _1342_ _1346_ VGND VGND VPWR VPWR _1347_ sky130_fd_sc_hd__a211o_1
XTAP_214 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_247 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3231_ _2897_ _2917_ _0305_ _0306_ VGND VGND VPWR VPWR _0307_ sky130_fd_sc_hd__o2bb2a_2
XANTENNA__4133__B1 _1032_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3162_ cu.id.opcode\[2\] VGND VGND VPWR VPWR _2899_ sky130_fd_sc_hd__buf_2
XTAP_269 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3487__A2 _0501_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3093_ ih.t.count\[6\] _2750_ _2830_ VGND VGND VPWR VPWR _2831_ sky130_fd_sc_hd__and3_1
XFILLER_0_89_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4615__A _0350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5803_ _2585_ _2586_ VGND VGND VPWR VPWR _2587_ sky130_fd_sc_hd__xnor2_1
X_3995_ _0620_ _0824_ VGND VGND VPWR VPWR _1069_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3947__B1 _2948_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5936__A1 _2350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5734_ net23 _2519_ _2527_ VGND VGND VPWR VPWR _0224_ sky130_fd_sc_hd__a21o_1
X_5665_ ih.t.timer_max\[23\] _2150_ _2319_ ih.t.timer_max\[7\] _1660_ VGND VGND VPWR
+ VPWR _2478_ sky130_fd_sc_hd__a221o_1
XFILLER_0_88_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4616_ _2923_ _2903_ VGND VGND VPWR VPWR _1659_ sky130_fd_sc_hd__or2_1
XFILLER_0_32_317 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5596_ net128 _2236_ _2247_ net136 VGND VGND VPWR VPWR _2412_ sky130_fd_sc_hd__a22o_1
X_4547_ _1599_ _1600_ VGND VGND VPWR VPWR _1601_ sky130_fd_sc_hd__nand2_1
Xmax_cap140 _2873_ VGND VGND VPWR VPWR net140 sky130_fd_sc_hd__buf_1
XFILLER_0_40_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4478_ _1530_ _1534_ _1535_ _1356_ VGND VGND VPWR VPWR _1536_ sky130_fd_sc_hd__o22ai_1
X_6217_ clknet_leaf_10_clk ih.t.next_count\[5\] net176 VGND VGND VPWR VPWR ih.t.count\[5\]
+ sky130_fd_sc_hd__dfrtp_1
X_3429_ cu.pc.pc_o\[0\] _0501_ _0502_ cu.reg_file.reg_b\[0\] _0504_ VGND VGND VPWR
+ VPWR _0505_ sky130_fd_sc_hd__a221o_1
X_6148_ clknet_leaf_18_clk _0182_ net184 VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__dfrtp_4
XTAP_770 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_792 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6079_ clknet_leaf_15_clk _0113_ net179 VGND VGND VPWR VPWR ih.t.timer_max\[27\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__4427__B2 cu.reg_file.reg_h\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4427__A1 cu.reg_file.reg_b\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4244__B _1309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4418__A1 _1473_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output130_A net130 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_512 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_46_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3780_ _0854_ _0855_ VGND VGND VPWR VPWR _0856_ sky130_fd_sc_hd__nand2_2
XANTENNA_clkbuf_leaf_14_clk_A clknet_2_2__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5450_ net68 _2277_ _2179_ net69 VGND VGND VPWR VPWR _2278_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4401_ _1455_ VGND VGND VPWR VPWR _1462_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5381_ _1261_ net123 _2226_ VGND VGND VPWR VPWR _2234_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_29_clk_A clknet_2_3__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4332_ _1396_ _1393_ VGND VGND VPWR VPWR _1397_ sky130_fd_sc_hd__nand2_1
X_4263_ mc.rw.state\[2\] _2699_ VGND VGND VPWR VPWR _1331_ sky130_fd_sc_hd__and2_1
XANTENNA__5713__B _1354_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_66_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6002_ clknet_leaf_31_clk _0040_ net185 VGND VGND VPWR VPWR cu.reg_file.reg_b\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_3214_ _2882_ _2906_ _2945_ _2948_ _2950_ VGND VGND VPWR VPWR _2951_ sky130_fd_sc_hd__o311a_4
XANTENNA__4329__B _1393_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4194_ _0516_ _1175_ VGND VGND VPWR VPWR _1263_ sky130_fd_sc_hd__nor2_4
X_3145_ _2874_ _2881_ VGND VGND VPWR VPWR _2882_ sky130_fd_sc_hd__nor2_1
XANTENNA__4409__A1 cu.reg_file.reg_sp\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4409__B2 cu.id.cb_opcode_x\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3076_ ih.t.timer_max\[12\] _2753_ VGND VGND VPWR VPWR _2814_ sky130_fd_sc_hd__nand2_1
XFILLER_0_49_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA_fanout161_A net162 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3632__A2 _0624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5909__A1 _1260_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3978_ _1021_ VGND VGND VPWR VPWR _1053_ sky130_fd_sc_hd__inv_2
X_5717_ _2518_ _2351_ VGND VGND VPWR VPWR _2519_ sky130_fd_sc_hd__nor2_4
XFILLER_0_17_144 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3396__A1 _2918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5648_ ih.gpio_interrupt_mask\[6\] _2326_ _2461_ _2125_ _2327_ VGND VGND VPWR VPWR
+ _2462_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_32_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5579_ net103 _2205_ _2395_ _1401_ VGND VGND VPWR VPWR _2396_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3424__A cu.id.starting_int_service VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5845__A0 cu.reg_file.reg_sp\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_556 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_83_537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_36_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5517__C _1354_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5025__S _2002_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5836__A0 _1213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output55_A net55 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput8 keypad_input[15] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_78_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5064__A1 _1189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4950_ cu.pc.pc_o\[12\] _1929_ VGND VGND VPWR VPWR _1940_ sky130_fd_sc_hd__nor2_1
XANTENNA__3614__A2 _0501_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4881_ _1875_ _1876_ VGND VGND VPWR VPWR _1877_ sky130_fd_sc_hd__or2b_1
X_3901_ _0361_ _0332_ VGND VGND VPWR VPWR _0977_ sky130_fd_sc_hd__nor2_1
X_3832_ _0866_ _0906_ _0907_ VGND VGND VPWR VPWR _0908_ sky130_fd_sc_hd__a21o_1
XANTENNA__4575__B1 _1222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5502_ ih.t.timer_max\[0\] _2320_ _2321_ VGND VGND VPWR VPWR _2322_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_54_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3763_ cu.reg_file.reg_sp\[14\] _0636_ _0748_ cu.reg_file.reg_h\[6\] VGND VGND VPWR
+ VPWR _0839_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3694_ _0769_ _0734_ VGND VGND VPWR VPWR _0770_ sky130_fd_sc_hd__xnor2_2
XFILLER_0_42_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5433_ _2265_ VGND VGND VPWR VPWR _0185_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5364_ _1374_ _2179_ VGND VGND VPWR VPWR _2224_ sky130_fd_sc_hd__and2_1
XFILLER_0_22_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4315_ _1377_ _1380_ VGND VGND VPWR VPWR _1381_ sky130_fd_sc_hd__xnor2_1
XANTENNA__5443__B _2247_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3550__A1 cu.reg_file.reg_d\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5295_ _1075_ net86 _2182_ VGND VGND VPWR VPWR _2185_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3550__B2 cu.alu_f\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4246_ _1309_ _1311_ VGND VGND VPWR VPWR _1314_ sky130_fd_sc_hd__nor2_2
X_4177_ _0663_ _0681_ _1060_ VGND VGND VPWR VPWR _1247_ sky130_fd_sc_hd__mux2_1
X_3128_ _2766_ _2865_ VGND VGND VPWR VPWR _2866_ sky130_fd_sc_hd__nor2_1
XFILLER_0_69_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5055__A1 _2002_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3059_ ih.t.count\[19\] _2796_ VGND VGND VPWR VPWR _2797_ sky130_fd_sc_hd__xnor2_1
XTAP_1029 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1018 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1007 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5618__B _1330_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3369__A1 cu.id.cb_opcode_y\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3369__B2 _0343_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5046__A1 _1624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5597__A2 _2194_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4309__B1 _1374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5080_ _1051_ _1623_ _2035_ VGND VGND VPWR VPWR _2041_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4100_ _0960_ _1173_ VGND VGND VPWR VPWR _1174_ sky130_fd_sc_hd__nand2_1
XANTENNA__5285__A1 _1260_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4031_ _1102_ _1103_ _1104_ _0566_ VGND VGND VPWR VPWR _1105_ sky130_fd_sc_hd__o22a_1
XFILLER_0_37_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5037__A1 _1222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5982_ clknet_leaf_27_clk _0020_ net186 VGND VGND VPWR VPWR cu.pc.pc_o\[4\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_59_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4933_ _1226_ _1917_ _1794_ VGND VGND VPWR VPWR _1925_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_74_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4864_ cu.pc.pc_o\[4\] _1838_ cu.pc.pc_o\[5\] VGND VGND VPWR VPWR _1861_ sky130_fd_sc_hd__a21oi_1
XANTENNA_13 programmable_gpio_in[4] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4795_ _0986_ _1005_ _1786_ _0983_ VGND VGND VPWR VPWR _1797_ sky130_fd_sc_hd__a2bb2o_2
XANTENNA_24 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3815_ cu.reg_file.reg_a\[1\] _0625_ _0628_ cu.reg_file.reg_mem\[9\] _0890_ VGND
+ VGND VPWR VPWR _0891_ sky130_fd_sc_hd__a221o_1
X_3746_ _0550_ _0820_ _0821_ VGND VGND VPWR VPWR _0822_ sky130_fd_sc_hd__a21o_2
XFILLER_0_15_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3771__A1 cu.reg_file.reg_b\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3771__B2 cu.reg_file.reg_sp\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5416_ _2254_ VGND VGND VPWR VPWR _0179_ sky130_fd_sc_hd__clkbuf_1
X_3677_ _0737_ _0752_ VGND VGND VPWR VPWR _0753_ sky130_fd_sc_hd__xor2_1
XFILLER_0_30_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput120 net120 VGND VGND VPWR VPWR ss5[4] sky130_fd_sc_hd__clkbuf_4
Xoutput131 net131 VGND VGND VPWR VPWR ss6[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5347_ _2147_ _2181_ VGND VGND VPWR VPWR _2215_ sky130_fd_sc_hd__nand2_4
XFILLER_0_10_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5278_ _2174_ VGND VGND VPWR VPWR _0121_ sky130_fd_sc_hd__clkbuf_1
X_4229_ _1296_ _1294_ VGND VGND VPWR VPWR _1297_ sky130_fd_sc_hd__nor2_2
XANTENNA__5028__A1 _2002_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5579__A2 _2205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_283 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5364__A _1374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2988__A net2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3514__B2 cu.reg_file.reg_d\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5303__S _2182_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_88_459 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4242__A2 _0361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4162__B _1213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput11 keypad_input[3] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__buf_2
XFILLER_0_71_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput22 memory_data_in[4] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_2
X_4580_ _2702_ _1261_ _1263_ _2697_ VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__a22o_1
X_3600_ cu.reg_file.reg_h\[4\] _0495_ _0498_ cu.alu_f\[4\] VGND VGND VPWR VPWR _0676_
+ sky130_fd_sc_hd__a22o_1
XFILLER_0_52_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3531_ _0603_ _0606_ VGND VGND VPWR VPWR _0607_ sky130_fd_sc_hd__or2_1
Xinput33 programmable_gpio_in[6] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_24_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3462_ cu.reg_file.reg_d\[1\] _0492_ _0498_ cu.alu_f\[1\] VGND VGND VPWR VPWR _0538_
+ sky130_fd_sc_hd__a22o_1
X_6250_ clknet_leaf_42_clk _0232_ net155 VGND VGND VPWR VPWR cu.reg_file.reg_sp\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_5201_ mc.cc.count\[1\] _2118_ _2120_ VGND VGND VPWR VPWR _2121_ sky130_fd_sc_hd__o21ai_1
X_6181_ clknet_leaf_23_clk _0214_ VGND VGND VPWR VPWR mc.cl.cmp_o sky130_fd_sc_hd__dfxtp_1
X_3393_ _0312_ _0449_ VGND VGND VPWR VPWR _0469_ sky130_fd_sc_hd__nor2_4
X_5132_ _1222_ _1089_ _2066_ VGND VGND VPWR VPWR _2075_ sky130_fd_sc_hd__mux2_1
XANTENNA__4618__A _1660_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5063_ _2029_ VGND VGND VPWR VPWR _0051_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4466__C1 _1489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3808__A2 _0426_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4014_ _0558_ _0681_ _0822_ _1040_ _1087_ VGND VGND VPWR VPWR _1088_ sky130_fd_sc_hd__a221o_1
XANTENNA__5449__A _1335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5965_ _2692_ VGND VGND VPWR VPWR _0290_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_90_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5896_ _2655_ VGND VGND VPWR VPWR _0258_ sky130_fd_sc_hd__clkbuf_1
X_4916_ _1907_ _1908_ VGND VGND VPWR VPWR _1909_ sky130_fd_sc_hd__nor2_1
XFILLER_0_47_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4847_ _1089_ _1840_ _1795_ VGND VGND VPWR VPWR _1846_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4778_ net140 _1783_ net205 VGND VGND VPWR VPWR _0015_ sky130_fd_sc_hd__a21boi_1
XFILLER_0_43_551 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3729_ _0755_ _0787_ VGND VGND VPWR VPWR _0805_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3135__C _2870_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4962__S _1814_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3983__A1 cu.alu_f\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5488__A1 net84 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_21_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_21_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_407 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4160__A1 _1032_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5660__B2 net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5660__A1 net115 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5968__S _2686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2962_ _2697_ _2702_ VGND VGND VPWR VPWR _2703_ sky130_fd_sc_hd__or2_1
XFILLER_0_8_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4066__A2_N _0663_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5750_ _2540_ VGND VGND VPWR VPWR _0227_ sky130_fd_sc_hd__clkbuf_1
X_4701_ net214 _1717_ _1719_ VGND VGND VPWR VPWR ih.t.next_count\[22\] sky130_fd_sc_hd__a21oi_1
X_5681_ net16 _1650_ _2488_ _2492_ VGND VGND VPWR VPWR _0206_ sky130_fd_sc_hd__a31o_1
XFILLER_0_60_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4632_ _1669_ VGND VGND VPWR VPWR _1672_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_60_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_56_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4923__A0 cu.pc.pc_o\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4563_ _1599_ _1602_ _1615_ VGND VGND VPWR VPWR _1616_ sky130_fd_sc_hd__a21o_1
XFILLER_0_71_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4494_ _1535_ _1545_ VGND VGND VPWR VPWR _1551_ sky130_fd_sc_hd__xor2_1
XFILLER_0_69_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6302_ clknet_leaf_35_clk _0284_ net160 VGND VGND VPWR VPWR cu.id.cb_opcode_x\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_4_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3514_ cu.reg_file.reg_mem\[1\] _0418_ _0415_ cu.reg_file.reg_d\[1\] VGND VGND VPWR
+ VPWR _0590_ sky130_fd_sc_hd__a22o_1
X_6233_ clknet_leaf_14_clk ih.t.next_count\[21\] net180 VGND VGND VPWR VPWR ih.t.count\[21\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_69_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3445_ _2936_ _0520_ VGND VGND VPWR VPWR _0521_ sky130_fd_sc_hd__nor2_1
XFILLER_0_40_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_952 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_941 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_930 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3376_ _2884_ _2885_ _2941_ VGND VGND VPWR VPWR _0452_ sky130_fd_sc_hd__and3_1
X_6164_ clknet_leaf_37_clk _0198_ net159 VGND VGND VPWR VPWR cu.reg_file.reg_mem\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA_fanout191_A net194 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_996 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_985 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_974 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_963 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6095_ clknet_leaf_7_clk _0129_ net165 VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__dfrtp_1
X_5115_ cu.reg_file.reg_e\[6\] _1193_ _2056_ VGND VGND VPWR VPWR _2063_ sky130_fd_sc_hd__mux2_1
X_5046_ _1193_ _1624_ _2002_ VGND VGND VPWR VPWR _2018_ sky130_fd_sc_hd__mux2_1
XFILLER_0_33_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5651__A1 net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5651__B2 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5948_ _0387_ _2467_ _2666_ VGND VGND VPWR VPWR _2683_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5879_ _2646_ VGND VGND VPWR VPWR _0250_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_250 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4530__B _1579_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4390__B2 _0387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4390__A1 cu.reg_file.reg_sp\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_93_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_38_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5536__B _1330_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5552__A _1649_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_215 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3230_ _2892_ _2899_ _2900_ _2923_ VGND VGND VPWR VPWR _0306_ sky130_fd_sc_hd__or4bb_1
XTAP_237 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3161_ _2893_ _2897_ VGND VGND VPWR VPWR _2898_ sky130_fd_sc_hd__nand2_1
XTAP_259 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4168__A _1144_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3092_ ih.t.timer_max\[5\] _2749_ ih.t.timer_max\[6\] VGND VGND VPWR VPWR _2830_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_89_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2998__A2 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5802_ _2576_ _2579_ _2577_ VGND VGND VPWR VPWR _2586_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_57_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3994_ _0918_ _0760_ _1065_ _1067_ VGND VGND VPWR VPWR _1068_ sky130_fd_sc_hd__a2bb2o_1
X_5733_ _2518_ mc.cl.next_data\[5\] _2111_ VGND VGND VPWR VPWR _2527_ sky130_fd_sc_hd__and3_1
XFILLER_0_72_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5664_ _1400_ _2476_ VGND VGND VPWR VPWR _2477_ sky130_fd_sc_hd__and2b_1
XFILLER_0_72_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_25_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4615_ _0350_ _2940_ _0379_ VGND VGND VPWR VPWR _1658_ sky130_fd_sc_hd__or3_2
X_5595_ _2411_ VGND VGND VPWR VPWR _0201_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_32_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4546_ _1333_ _1598_ VGND VGND VPWR VPWR _1600_ sky130_fd_sc_hd__nand2_1
XFILLER_0_4_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_96_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4477_ _1517_ _1530_ VGND VGND VPWR VPWR _1535_ sky130_fd_sc_hd__nand2_1
XFILLER_0_40_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6216_ clknet_leaf_10_clk ih.t.next_count\[4\] net176 VGND VGND VPWR VPWR ih.t.count\[4\]
+ sky130_fd_sc_hd__dfrtp_2
X_3428_ _2948_ _0501_ _0503_ VGND VGND VPWR VPWR _0504_ sky130_fd_sc_hd__a21bo_2
X_6147_ clknet_leaf_30_clk _0181_ net187 VGND VGND VPWR VPWR net139 sky130_fd_sc_hd__dfrtp_4
XTAP_760 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3359_ _2940_ _2942_ _0379_ VGND VGND VPWR VPWR _0435_ sky130_fd_sc_hd__nor3_1
XTAP_793 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6078_ clknet_leaf_15_clk _0112_ net179 VGND VGND VPWR VPWR ih.t.timer_max\[26\]
+ sky130_fd_sc_hd__dfrtp_2
X_5029_ cu.reg_file.reg_b\[0\] _2003_ _2006_ VGND VGND VPWR VPWR _2007_ sky130_fd_sc_hd__mux2_1
XANTENNA__4525__B _1579_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5388__A0 _1052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4244__C _1311_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3938__A1 alu.Cin VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4363__A1 cu.reg_file.reg_e\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5560__B1 _2225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2996__A net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5312__A0 _0619_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5984__RESET_B net188 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5863__A1 ih.t.timer_max\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output123_A net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_86_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5379__A0 _1194_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4400_ _1382_ _1457_ _1458_ _1461_ VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__a31o_2
X_5380_ _2233_ VGND VGND VPWR VPWR _0164_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3343__C_N _0405_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4331_ _1376_ VGND VGND VPWR VPWR _1396_ sky130_fd_sc_hd__clkbuf_4
X_4262_ _1329_ VGND VGND VPWR VPWR _1330_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__5303__A0 _1194_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3213_ _2949_ VGND VGND VPWR VPWR _2950_ sky130_fd_sc_hd__buf_4
X_6001_ clknet_leaf_2_clk _0039_ net157 VGND VGND VPWR VPWR cu.reg_file.reg_a\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_66_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4193_ _1184_ VGND VGND VPWR VPWR _1262_ sky130_fd_sc_hd__inv_2
XANTENNA__5606__A1 _1666_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3144_ _2877_ _2880_ VGND VGND VPWR VPWR _2881_ sky130_fd_sc_hd__and2_1
XANTENNA__4409__A2 _0993_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3075_ ih.t.count\[13\] _2812_ VGND VGND VPWR VPWR _2813_ sky130_fd_sc_hd__xnor2_1
XANTENNA__3617__B1 _0536_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_fanout154_A net163 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3977_ _1051_ VGND VGND VPWR VPWR _1052_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_45_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4042__B1 _0566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5716_ mc.count VGND VGND VPWR VPWR _2518_ sky130_fd_sc_hd__buf_2
XANTENNA__5457__A _1633_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_60_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5647_ mc.cl.next_data\[6\] _2313_ net141 _2460_ VGND VGND VPWR VPWR _2461_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5578_ net87 _1330_ VGND VGND VPWR VPWR _2395_ sky130_fd_sc_hd__or2_1
X_4529_ _1580_ _1581_ _1582_ _1334_ VGND VGND VPWR VPWR _1584_ sky130_fd_sc_hd__a31oi_1
XANTENNA__3553__C1 _0536_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_590 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2997__A_N net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_83_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_2_3__f_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4033__B1 _0566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5781__A0 cu.reg_file.reg_sp\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_51_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput9 keypad_input[1] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__buf_2
XANTENNA_output48_A net48 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5041__S _2006_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_332 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4880_ _0387_ cu.pc.pc_o\[6\] VGND VGND VPWR VPWR _1876_ sky130_fd_sc_hd__nand2_1
X_3900_ _0321_ _0970_ _0972_ _0975_ VGND VGND VPWR VPWR _0976_ sky130_fd_sc_hd__or4_4
XFILLER_0_52_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3831_ _0861_ _0864_ VGND VGND VPWR VPWR _0907_ sky130_fd_sc_hd__nor2_1
XANTENNA__5772__A0 _1160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4575__A1 _2702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3762_ cu.id.imm_i\[14\] _0739_ _0837_ _0653_ VGND VGND VPWR VPWR _0838_ sky130_fd_sc_hd__a22oi_4
X_5501_ ih.t.enable _2257_ _2150_ ih.t.timer_max\[16\] _1660_ VGND VGND VPWR VPWR
+ _2321_ sky130_fd_sc_hd__a221o_1
XANTENNA__4575__B2 _2697_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3693_ _0645_ _0722_ _0735_ VGND VGND VPWR VPWR _0769_ sky130_fd_sc_hd__a21o_1
X_5432_ _2022_ net71 _2264_ VGND VGND VPWR VPWR _2265_ sky130_fd_sc_hd__mux2_1
XANTENNA__4327__A1 cu.reg_file.reg_c\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5363_ _2223_ VGND VGND VPWR VPWR _0157_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4314_ _1378_ _1379_ VGND VGND VPWR VPWR _1380_ sky130_fd_sc_hd__nand2_1
XANTENNA__3550__A2 _0492_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5294_ _2184_ VGND VGND VPWR VPWR _0127_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4245_ _1312_ VGND VGND VPWR VPWR _1313_ sky130_fd_sc_hd__clkbuf_4
X_4176_ _0566_ _0632_ _1060_ VGND VGND VPWR VPWR _1246_ sky130_fd_sc_hd__mux2_1
X_3127_ ih.t.timer_max\[30\] _2765_ VGND VGND VPWR VPWR _2865_ sky130_fd_sc_hd__and2_1
X_3058_ ih.t.timer_max\[19\] _2758_ VGND VGND VPWR VPWR _2796_ sky130_fd_sc_hd__xor2_1
XTAP_1019 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1008 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_65_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3369__A2 _0361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5126__S _2066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3435__A alu.Cin VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_13_clk_A clknet_2_2__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4266__A _2697_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_28_clk_A clknet_2_3__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4557__A1 cu.pc.pc_o\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_47_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4030_ _0599_ _0603_ _1101_ _0729_ _0606_ VGND VGND VPWR VPWR _1104_ sky130_fd_sc_hd__a32o_1
X_5981_ clknet_leaf_27_clk _0019_ net187 VGND VGND VPWR VPWR cu.pc.pc_o\[3\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_59_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4904__A _2920_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4932_ _1920_ _1923_ VGND VGND VPWR VPWR _1924_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_86_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6034__RESET_B net188 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_14 net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4863_ cu.pc.pc_o\[5\] cu.pc.pc_o\[4\] _1838_ VGND VGND VPWR VPWR _1860_ sky130_fd_sc_hd__and3_1
XFILLER_0_6_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4794_ _0617_ _1788_ _1795_ VGND VGND VPWR VPWR _1796_ sky130_fd_sc_hd__mux2_1
X_3814_ cu.pc.pc_o\[9\] _0740_ _0889_ VGND VGND VPWR VPWR _0890_ sky130_fd_sc_hd__a21o_1
XFILLER_0_82_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3745_ _0614_ _0573_ VGND VGND VPWR VPWR _0821_ sky130_fd_sc_hd__nand2_1
XANTENNA__3771__A2 _0743_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5415_ _1192_ net137 _2248_ VGND VGND VPWR VPWR _2254_ sky130_fd_sc_hd__mux2_1
Xoutput110 net110 VGND VGND VPWR VPWR ss4[2] sky130_fd_sc_hd__clkbuf_4
X_3676_ _0747_ _0751_ VGND VGND VPWR VPWR _0752_ sky130_fd_sc_hd__xor2_2
Xoutput132 net132 VGND VGND VPWR VPWR ss7[0] sky130_fd_sc_hd__clkbuf_4
Xoutput121 net121 VGND VGND VPWR VPWR ss5[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_63_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5346_ _2214_ VGND VGND VPWR VPWR _0149_ sky130_fd_sc_hd__clkbuf_1
X_5277_ net79 _1187_ _2170_ VGND VGND VPWR VPWR _2174_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4228_ _1271_ VGND VGND VPWR VPWR _1296_ sky130_fd_sc_hd__inv_2
X_4159_ _0954_ _0778_ VGND VGND VPWR VPWR _1229_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_35_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_35_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_92_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4539__A1 _1296_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_560 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xclkbuf_leaf_26_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_26_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__4242__A3 _0968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_96_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_83_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4162__C _1222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput12 keypad_input[4] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__clkbuf_2
Xinput23 memory_data_in[5] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__buf_1
X_3530_ _0519_ _0605_ VGND VGND VPWR VPWR _0606_ sky130_fd_sc_hd__nor2_2
Xinput34 programmable_gpio_in[7] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_12_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3461_ cu.reg_file.reg_c\[1\] _0485_ _0533_ _0535_ _0536_ VGND VGND VPWR VPWR _0537_
+ sky130_fd_sc_hd__a2111o_1
X_5200_ mc.cc.enable_edge_detector.prev_data _2708_ VGND VGND VPWR VPWR _2120_ sky130_fd_sc_hd__or2_1
X_6180_ clknet_leaf_36_clk _0000_ net158 VGND VGND VPWR VPWR ih.interrupt_source\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_3392_ _0465_ net147 _0467_ VGND VGND VPWR VPWR _0468_ sky130_fd_sc_hd__nor3_1
XFILLER_0_58_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5131_ _2074_ VGND VGND VPWR VPWR _0074_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_20_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5290__A _2180_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5062_ cu.reg_file.reg_c\[3\] _1187_ _2025_ VGND VGND VPWR VPWR _2029_ sky130_fd_sc_hd__mux2_1
X_4013_ _0607_ _1086_ _0694_ VGND VGND VPWR VPWR _1087_ sky130_fd_sc_hd__o21a_1
XANTENNA__3269__A1 _0340_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_79_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_87_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xclkbuf_leaf_17_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_17_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__5449__B _1354_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5964_ cu.id.imm_i\[13\] _2448_ _2686_ VGND VGND VPWR VPWR _2692_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5895_ ih.t.timer_max\[16\] _0618_ _2654_ VGND VGND VPWR VPWR _2655_ sky130_fd_sc_hd__mux2_1
X_4915_ cu.pc.pc_o\[9\] _1894_ VGND VGND VPWR VPWR _1908_ sky130_fd_sc_hd__nor2_1
X_4846_ _1843_ _1844_ VGND VGND VPWR VPWR _1845_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_47_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4777_ net199 _1782_ VGND VGND VPWR VPWR _1783_ sky130_fd_sc_hd__nand2_1
X_3728_ _0664_ _0803_ VGND VGND VPWR VPWR _0804_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_15_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3659_ _0632_ _0643_ VGND VGND VPWR VPWR _0735_ sky130_fd_sc_hd__and2_1
X_5329_ _2204_ VGND VGND VPWR VPWR _2205_ sky130_fd_sc_hd__clkbuf_8
XANTENNA__4202__C_N _1269_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4339__A_N _1393_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3432__A1 _0343_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_34_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5488__A2 _2180_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_408 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5314__S _2195_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5645__C1 _1660_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5948__A0 _0387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2961_ _2698_ _2699_ _2701_ VGND VGND VPWR VPWR _2702_ sky130_fd_sc_hd__a21o_4
XFILLER_0_60_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3959__C1 _0918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1180 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4700_ ih.t.count\[22\] _1717_ _1670_ VGND VGND VPWR VPWR _1719_ sky130_fd_sc_hd__o21ai_1
X_5680_ _2491_ _1643_ cu.reg_file.reg_mem\[8\] _2111_ VGND VGND VPWR VPWR _2492_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_17_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5176__A1 net21 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4631_ _1671_ VGND VGND VPWR VPWR ih.t.next_count\[0\] sky130_fd_sc_hd__clkbuf_1
X_4562_ _1396_ _1614_ VGND VGND VPWR VPWR _1615_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_52_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4493_ _1548_ _1549_ VGND VGND VPWR VPWR _1550_ sky130_fd_sc_hd__xnor2_1
X_6301_ clknet_leaf_37_clk _0283_ net158 VGND VGND VPWR VPWR cu.id.cb_opcode_x\[0\]
+ sky130_fd_sc_hd__dfrtp_1
X_3513_ cu.reg_file.reg_c\[1\] _0427_ _0430_ cu.reg_file.reg_e\[1\] VGND VGND VPWR
+ VPWR _0589_ sky130_fd_sc_hd__a22o_1
XFILLER_0_40_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6232_ clknet_leaf_14_clk ih.t.next_count\[20\] net180 VGND VGND VPWR VPWR ih.t.count\[20\]
+ sky130_fd_sc_hd__dfrtp_1
Xclkbuf_leaf_6_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_6_clk sky130_fd_sc_hd__clkbuf_16
X_3444_ _2886_ _0378_ VGND VGND VPWR VPWR _0520_ sky130_fd_sc_hd__nand2_1
XFILLER_0_85_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_953 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_942 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_931 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_920 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6163_ clknet_leaf_6_clk _0197_ net166 VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__dfrtp_2
X_3375_ _2878_ _0301_ VGND VGND VPWR VPWR _0451_ sky130_fd_sc_hd__nor2_1
XTAP_986 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_975 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_964 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6094_ clknet_leaf_27_clk _0128_ net186 VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__dfrtp_4
X_5114_ _2062_ VGND VGND VPWR VPWR _0069_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_85_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_997 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5045_ _2017_ VGND VGND VPWR VPWR _0045_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5947_ _2682_ VGND VGND VPWR VPWR _0282_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_433 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5167__A1 net18 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5878_ _2022_ ih.t.timer_max\[0\] _2645_ VGND VGND VPWR VPWR _2646_ sky130_fd_sc_hd__mux2_1
XFILLER_0_35_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4829_ _0341_ cu.pc.pc_o\[2\] VGND VGND VPWR VPWR _1829_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4390__A2 _0993_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4127__C1 _0918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3443__A _0384_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4973__S _1814_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4850__A0 cu.pc.pc_o\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4381__A2 _1434_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_205 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5044__S _2006_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_238 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_39_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3160_ _2894_ VGND VGND VPWR VPWR _2897_ sky130_fd_sc_hd__inv_2
XTAP_249 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4168__B _1160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3091_ ih.t.count\[7\] _2828_ VGND VGND VPWR VPWR _2829_ sky130_fd_sc_hd__xnor2_1
Xhold1 ih.ip_ed.prev_data VGND VGND VPWR VPWR net197 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_49_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4615__C _0379_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5801_ _2583_ _2584_ VGND VGND VPWR VPWR _2585_ sky130_fd_sc_hd__nand2_1
X_5732_ net22 _2519_ _2526_ VGND VGND VPWR VPWR _0223_ sky130_fd_sc_hd__a21o_1
XFILLER_0_71_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3993_ _1033_ _1066_ _0806_ VGND VGND VPWR VPWR _1067_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_549 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5663_ ih.t.timer_max\[23\] _2204_ _2314_ ih.t.timer_max\[7\] _2475_ VGND VGND VPWR
+ VPWR _2476_ sky130_fd_sc_hd__a221o_1
XFILLER_0_29_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4614_ _1656_ VGND VGND VPWR VPWR _1657_ sky130_fd_sc_hd__inv_2
XFILLER_0_72_488 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5594_ cu.reg_file.reg_mem\[3\] _2410_ _2351_ VGND VGND VPWR VPWR _2411_ sky130_fd_sc_hd__mux2_1
X_4545_ _1333_ _1598_ VGND VGND VPWR VPWR _1599_ sky130_fd_sc_hd__or2_1
XFILLER_0_25_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xmax_cap142 _0509_ VGND VGND VPWR VPWR net142 sky130_fd_sc_hd__buf_2
X_4476_ _1356_ _1517_ _1402_ VGND VGND VPWR VPWR _1534_ sky130_fd_sc_hd__o21a_1
X_6215_ clknet_leaf_10_clk ih.t.next_count\[3\] net176 VGND VGND VPWR VPWR ih.t.count\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3427_ _2913_ _2952_ _0307_ _0293_ VGND VGND VPWR VPWR _0503_ sky130_fd_sc_hd__a31o_1
XANTENNA__3263__A _0296_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6146_ clknet_leaf_7_clk _0180_ net167 VGND VGND VPWR VPWR net138 sky130_fd_sc_hd__dfrtp_2
XTAP_761 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3358_ cu.reg_file.reg_b\[0\] _0432_ _0433_ cu.reg_file.reg_a\[0\] VGND VGND VPWR
+ VPWR _0434_ sky130_fd_sc_hd__a22o_1
XTAP_794 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6077_ clknet_leaf_15_clk _0111_ net179 VGND VGND VPWR VPWR ih.t.timer_max\[25\]
+ sky130_fd_sc_hd__dfrtp_4
X_3289_ _2940_ _2953_ _0364_ VGND VGND VPWR VPWR _0365_ sky130_fd_sc_hd__o21bai_1
X_5028_ _2002_ _2005_ _2951_ VGND VGND VPWR VPWR _2006_ sky130_fd_sc_hd__o21a_4
XANTENNA__5388__A1 net125 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5129__S _2066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3438__A _0384_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4348__C1 _1364_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5560__A1 net110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5560__B2 net118 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5312__A1 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3901__A _0361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5379__A1 net122 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4587__C1 _1417_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_179 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5000__A0 cu.reg_file.reg_a\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5551__B2 net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5551__A1 net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4330_ _1383_ _1394_ VGND VGND VPWR VPWR _1395_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5303__A1 net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4261_ _1291_ _1307_ _1328_ VGND VGND VPWR VPWR _1329_ sky130_fd_sc_hd__o21bai_4
XFILLER_0_5_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3314__B1 _2918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3212_ cu.id.starting_int_service VGND VGND VPWR VPWR _2949_ sky130_fd_sc_hd__inv_2
X_6000_ clknet_leaf_3_clk _0038_ net156 VGND VGND VPWR VPWR cu.reg_file.reg_a\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_4192_ _1260_ VGND VGND VPWR VPWR _1261_ sky130_fd_sc_hd__buf_4
X_3143_ _2878_ _2879_ VGND VGND VPWR VPWR _2880_ sky130_fd_sc_hd__or2_2
X_3074_ ih.t.timer_max\[13\] _2754_ VGND VGND VPWR VPWR _2812_ sky130_fd_sc_hd__xor2_1
XANTENNA__4814__A0 _1299_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_82_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3976_ _1050_ VGND VGND VPWR VPWR _1051_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_45_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5457__B _2284_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5715_ _2517_ VGND VGND VPWR VPWR _0215_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_93_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5646_ _1665_ _2458_ _2459_ VGND VGND VPWR VPWR _2460_ sky130_fd_sc_hd__o21a_1
XFILLER_0_5_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5542__B2 ih.t.timer_max\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5542__A1 ih.t.timer_max\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5577_ net95 _2194_ _2393_ VGND VGND VPWR VPWR _2394_ sky130_fd_sc_hd__a21o_1
XFILLER_0_60_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4528_ _1580_ _1581_ _1582_ VGND VGND VPWR VPWR _1583_ sky130_fd_sc_hd__a21o_1
X_4459_ _1356_ _1501_ _1402_ VGND VGND VPWR VPWR _1518_ sky130_fd_sc_hd__o21a_1
XANTENNA__4502__C1 _1323_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6129_ clknet_leaf_19_clk _0163_ net184 VGND VGND VPWR VPWR net121 sky130_fd_sc_hd__dfrtp_1
XANTENNA__4817__A _0340_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5058__A0 cu.reg_file.reg_c\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_580 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_591 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_55_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3792__B1 _0741_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5383__A _1369_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5297__A0 _1188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5322__S _2195_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5049__A0 _1260_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4272__A1 cu.reg_file.reg_c\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5558__A net86 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5221__A0 _1192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4024__A1 _1032_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3830_ _0877_ _0904_ _0905_ VGND VGND VPWR VPWR _0906_ sky130_fd_sc_hd__a21o_1
XFILLER_0_6_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4575__A2 _1188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3761_ cu.reg_file.reg_a\[6\] _0625_ _0628_ cu.reg_file.reg_mem\[14\] _0836_ VGND
+ VGND VPWR VPWR _0837_ sky130_fd_sc_hd__a221o_1
XFILLER_0_82_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5500_ _2319_ VGND VGND VPWR VPWR _2320_ sky130_fd_sc_hd__buf_2
X_3692_ _0754_ _0757_ _0767_ VGND VGND VPWR VPWR _0768_ sky130_fd_sc_hd__or3_2
XFILLER_0_42_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5431_ _2139_ _2205_ VGND VGND VPWR VPWR _2264_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5362_ _1261_ net115 _2215_ VGND VGND VPWR VPWR _2223_ sky130_fd_sc_hd__mux2_1
XFILLER_0_72_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4313_ _1332_ _1368_ VGND VGND VPWR VPWR _1379_ sky130_fd_sc_hd__nand2_1
XFILLER_0_65_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5293_ _1052_ net85 _2182_ VGND VGND VPWR VPWR _2184_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4244_ _0992_ _1309_ _1311_ VGND VGND VPWR VPWR _1312_ sky130_fd_sc_hd__and3b_2
X_4175_ _1241_ _1244_ _0588_ VGND VGND VPWR VPWR _1245_ sky130_fd_sc_hd__mux2_1
X_3126_ _2770_ _2771_ _2863_ VGND VGND VPWR VPWR _2864_ sky130_fd_sc_hd__or3_1
XANTENNA__4356__B _1417_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3057_ ih.t.count\[20\] _2759_ _2793_ VGND VGND VPWR VPWR _2795_ sky130_fd_sc_hd__and3_1
XTAP_1009 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5468__A _2205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_18_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_73_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3959_ _0758_ _1031_ _1033_ _0918_ VGND VGND VPWR VPWR _1034_ sky130_fd_sc_hd__o211ai_1
XFILLER_0_9_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_241 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5629_ _2169_ _2436_ _2443_ _2136_ VGND VGND VPWR VPWR _2444_ sky130_fd_sc_hd__o211a_1
XANTENNA__5407__S _2248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5279__A0 net80 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5142__S _2069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XPHY_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3214__C1 _2950_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_47_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5980_ clknet_leaf_30_clk _0018_ net187 VGND VGND VPWR VPWR cu.pc.pc_o\[2\] sky130_fd_sc_hd__dfrtp_4
XFILLER_0_59_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4931_ _1921_ _1922_ VGND VGND VPWR VPWR _1923_ sky130_fd_sc_hd__nand2_1
XANTENNA__4904__B cu.pc.pc_o\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5288__A _1369_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4192__A _1260_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4862_ _1859_ VGND VGND VPWR VPWR _0020_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3813_ cu.reg_file.reg_d\[1\] _0488_ _0741_ cu.reg_file.reg_h\[1\] _0888_ VGND VGND
+ VPWR VPWR _0889_ sky130_fd_sc_hd__a221o_1
XANTENNA_15 net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4793_ _1794_ VGND VGND VPWR VPWR _1795_ sky130_fd_sc_hd__buf_4
XFILLER_0_55_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_157 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3744_ _0605_ _0553_ VGND VGND VPWR VPWR _0820_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3675_ cu.reg_file.reg_mem\[8\] _0640_ _0749_ _0750_ VGND VGND VPWR VPWR _0751_ sky130_fd_sc_hd__a211oi_4
XFILLER_0_42_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5414_ _2253_ VGND VGND VPWR VPWR _0178_ sky130_fd_sc_hd__clkbuf_1
Xoutput100 net100 VGND VGND VPWR VPWR ss3[0] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_30_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput133 net133 VGND VGND VPWR VPWR ss7[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput122 net122 VGND VGND VPWR VPWR ss5[6] sky130_fd_sc_hd__clkbuf_4
Xoutput111 net111 VGND VGND VPWR VPWR ss4[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_42_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5345_ _1261_ net107 _2206_ VGND VGND VPWR VPWR _2214_ sky130_fd_sc_hd__mux2_1
XANTENNA__5751__A cu.reg_file.reg_sp\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5276_ _2173_ VGND VGND VPWR VPWR _0120_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4227_ _1294_ VGND VGND VPWR VPWR _1295_ sky130_fd_sc_hd__buf_2
XANTENNA__4484__A1 cu.pc.pc_o\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3287__A2 _0361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4158_ _0771_ _0954_ _0779_ _0935_ _0916_ VGND VGND VPWR VPWR _1228_ sky130_fd_sc_hd__o32a_1
X_3109_ ih.t.count\[3\] _2846_ VGND VGND VPWR VPWR _2847_ sky130_fd_sc_hd__xor2_1
X_4089_ _1161_ _1162_ VGND VGND VPWR VPWR _1163_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_77_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4830__A _0341_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3446__A _0373_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4277__A _1343_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput13 keypad_input[5] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__buf_2
Xinput24 memory_data_in[6] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__buf_1
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5047__S _2006_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3460_ _0504_ VGND VGND VPWR VPWR _0536_ sky130_fd_sc_hd__clkbuf_4
X_3391_ _2923_ _0354_ net150 _0382_ _0466_ VGND VGND VPWR VPWR _0467_ sky130_fd_sc_hd__a311o_1
X_5130_ _2073_ cu.reg_file.reg_h\[2\] _2069_ VGND VGND VPWR VPWR _2074_ sky130_fd_sc_hd__mux2_1
XFILLER_0_20_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5061_ _2028_ VGND VGND VPWR VPWR _0050_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4466__A1 cu.id.imm_i\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4466__B2 _1521_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4012_ _0610_ _1083_ _0701_ _0611_ VGND VGND VPWR VPWR _1086_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__3269__A2 _0341_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4915__A cu.pc.pc_o\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5415__A0 _1192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5963_ _2691_ VGND VGND VPWR VPWR _0289_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5966__A1 _2467_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4769__A2 _1644_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4914_ cu.pc.pc_o\[9\] _1894_ VGND VGND VPWR VPWR _1907_ sky130_fd_sc_hd__and2_1
XFILLER_0_59_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5894_ _1667_ _2205_ _2152_ VGND VGND VPWR VPWR _2654_ sky130_fd_sc_hd__o21a_4
X_4845_ _1829_ _1832_ _1830_ VGND VGND VPWR VPWR _1844_ sky130_fd_sc_hd__o21a_1
XFILLER_0_35_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4776_ _0980_ _1781_ VGND VGND VPWR VPWR _1782_ sky130_fd_sc_hd__or2_1
XFILLER_0_15_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_12_clk_A clknet_2_2__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5465__B _2284_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3727_ _0684_ _0787_ _0682_ VGND VGND VPWR VPWR _0803_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_43_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3658_ _0733_ VGND VGND VPWR VPWR _0734_ sky130_fd_sc_hd__inv_2
XFILLER_0_30_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3589_ _0294_ _0634_ _0374_ VGND VGND VPWR VPWR _0665_ sky130_fd_sc_hd__or3b_1
X_5328_ _2149_ VGND VGND VPWR VPWR _2204_ sky130_fd_sc_hd__clkbuf_4
XANTENNA_clkbuf_leaf_27_clk_A clknet_2_3__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5700__A2_N _1643_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5259_ _2162_ VGND VGND VPWR VPWR _0114_ sky130_fd_sc_hd__clkbuf_1
Xclkbuf_2_2__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_2__leaf_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_65_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_65_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5709__A1 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_19_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_93_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5978__RESET_B net188 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2999__B net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_409 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_28_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout190 net194 VGND VGND VPWR VPWR net190 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_44_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4454__B _1511_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5948__A1 _2467_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2960_ _2700_ VGND VGND VPWR VPWR _2701_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_29_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1181 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1170 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4630_ ih.t.count\[0\] _1670_ VGND VGND VPWR VPWR _1671_ sky130_fd_sc_hd__and2b_1
XFILLER_0_84_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4561_ _1305_ _1610_ _1613_ VGND VGND VPWR VPWR _1614_ sky130_fd_sc_hd__o21a_1
X_6300_ clknet_leaf_38_clk _0282_ net160 VGND VGND VPWR VPWR cu.id.cb_opcode_y\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_4492_ _1332_ _1530_ _1532_ VGND VGND VPWR VPWR _1549_ sky130_fd_sc_hd__o21a_1
XFILLER_0_52_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3512_ _0587_ VGND VGND VPWR VPWR _0588_ sky130_fd_sc_hd__buf_2
X_6231_ clknet_leaf_14_clk net213 net180 VGND VGND VPWR VPWR ih.t.count\[19\] sky130_fd_sc_hd__dfrtp_1
X_3443_ _0384_ _0392_ VGND VGND VPWR VPWR _0519_ sky130_fd_sc_hd__or2_1
XANTENNA__5884__A0 _1187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_910 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6162_ clknet_leaf_6_clk _0196_ net165 VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_85_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_943 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_932 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_921 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3374_ _0312_ _0448_ _0449_ VGND VGND VPWR VPWR _0450_ sky130_fd_sc_hd__or3_1
XANTENNA__4151__A3 _0773_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5113_ cu.reg_file.reg_e\[5\] _1191_ _2056_ VGND VGND VPWR VPWR _2062_ sky130_fd_sc_hd__mux2_1
XFILLER_0_85_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_987 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_976 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_965 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_954 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6093_ clknet_leaf_10_clk _0127_ net175 VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__dfrtp_1
XANTENNA__5636__B1 _2247_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_998 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5044_ cu.reg_file.reg_b\[5\] _2016_ _2006_ VGND VGND VPWR VPWR _2017_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4611__A1 _1650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5946_ _0373_ _2448_ _2666_ VGND VGND VPWR VPWR _2682_ sky130_fd_sc_hd__mux2_1
X_5877_ _1667_ _2180_ _2635_ VGND VGND VPWR VPWR _2645_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_75_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4828_ _1826_ _1827_ VGND VGND VPWR VPWR _1828_ sky130_fd_sc_hd__nor2_1
XANTENNA__5476__A _2225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_445 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3708__B _0587_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_50_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4759_ _1760_ _1766_ _1767_ VGND VGND VPWR VPWR _1768_ sky130_fd_sc_hd__or3_2
XFILLER_0_7_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_43_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5415__S _2248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_423 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_206 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_239 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3090_ ih.t.timer_max\[7\] _2750_ VGND VGND VPWR VPWR _2828_ sky130_fd_sc_hd__xor2_1
Xhold2 _0217_ VGND VGND VPWR VPWR net198 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_55_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3992_ _0816_ _0807_ _0776_ VGND VGND VPWR VPWR _1066_ sky130_fd_sc_hd__a21oi_1
X_5800_ cu.reg_file.reg_sp\[8\] _2535_ VGND VGND VPWR VPWR _2584_ sky130_fd_sc_hd__nand2_1
X_5731_ _2518_ mc.cl.next_data\[4\] _2111_ VGND VGND VPWR VPWR _2526_ sky130_fd_sc_hd__and3_1
XFILLER_0_9_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_261 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5662_ ih.t.timer_max\[31\] _2145_ _2192_ ih.t.timer_max\[15\] VGND VGND VPWR VPWR
+ _2475_ sky130_fd_sc_hd__a22o_1
X_4613_ mc.cl.cmp_o _1364_ _1613_ VGND VGND VPWR VPWR _1656_ sky130_fd_sc_hd__or3b_1
X_5593_ _2406_ _2407_ _2409_ _1641_ VGND VGND VPWR VPWR _2410_ sky130_fd_sc_hd__o22a_2
XFILLER_0_4_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4544_ _1305_ _1594_ _1597_ VGND VGND VPWR VPWR _1598_ sky130_fd_sc_hd__o21ai_4
XANTENNA__3247__C _2908_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4475_ _1512_ _1531_ _1520_ VGND VGND VPWR VPWR _1533_ sky130_fd_sc_hd__nand3_1
X_6214_ clknet_leaf_10_clk ih.t.next_count\[2\] net175 VGND VGND VPWR VPWR ih.t.count\[2\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__5857__A0 cu.reg_file.reg_sp\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3426_ net146 _0473_ _0479_ _0486_ _0458_ VGND VGND VPWR VPWR _0502_ sky130_fd_sc_hd__o2111a_4
XTAP_751 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6145_ clknet_leaf_6_clk _0179_ net165 VGND VGND VPWR VPWR net137 sky130_fd_sc_hd__dfrtp_2
XTAP_740 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3332__A1 _2877_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3357_ _0412_ _0405_ _0424_ VGND VGND VPWR VPWR _0433_ sky130_fd_sc_hd__and3_2
X_6076_ clknet_leaf_21_clk _0110_ net189 VGND VGND VPWR VPWR ih.t.timer_max\[24\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_795 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_762 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3288_ _2902_ _2884_ VGND VGND VPWR VPWR _0364_ sky130_fd_sc_hd__xnor2_4
X_5027_ _1792_ _2004_ VGND VGND VPWR VPWR _2005_ sky130_fd_sc_hd__nor2_1
XANTENNA__4832__A1 _0340_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4060__A2 _0773_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5929_ _2673_ VGND VGND VPWR VPWR _0273_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_35_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5560__A2 _2147_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3571__A1 cu.reg_file.reg_d\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3571__B2 cu.reg_file.reg_b\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5145__S _2069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3323__A1 _2893_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3087__B1 ih.t.timer_max\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5993__RESET_B net161 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_81_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_14_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_26_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output90_A net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3562__A1 cu.reg_file.reg_sp\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3364__A _0293_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3562__B2 cu.reg_file.reg_h\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4260_ cu.reg_file.reg_c\[0\] _1313_ _1327_ VGND VGND VPWR VPWR _1328_ sky130_fd_sc_hd__a21oi_1
X_4191_ _1110_ VGND VGND VPWR VPWR _1260_ sky130_fd_sc_hd__buf_4
X_3211_ _2946_ _2947_ VGND VGND VPWR VPWR _2948_ sky130_fd_sc_hd__nor2_8
XFILLER_0_5_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3142_ _2875_ _2876_ VGND VGND VPWR VPWR _2879_ sky130_fd_sc_hd__nand2_1
XFILLER_0_89_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3073_ _2755_ _2809_ ih.t.count\[14\] VGND VGND VPWR VPWR _2811_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_49_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3975_ _0517_ _1038_ _1039_ _1049_ VGND VGND VPWR VPWR _1050_ sky130_fd_sc_hd__a211o_4
X_5714_ ih.input_handler_enable _0618_ _2516_ VGND VGND VPWR VPWR _2517_ sky130_fd_sc_hd__mux2_1
XFILLER_0_9_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_17_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5645_ ih.t.timer_max\[22\] _2150_ _2319_ ih.t.timer_max\[6\] _1660_ VGND VGND VPWR
+ VPWR _2459_ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5542__A2 _2193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5576_ net127 _2236_ _2247_ net135 VGND VGND VPWR VPWR _2393_ sky130_fd_sc_hd__a22o_1
XANTENNA__5473__B _2284_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3553__A1 cu.pc.pc_o\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4527_ _1333_ _1561_ _1565_ VGND VGND VPWR VPWR _1582_ sky130_fd_sc_hd__o21ai_2
XANTENNA__3274__A _0296_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4458_ _1501_ _1511_ VGND VGND VPWR VPWR _1517_ sky130_fd_sc_hd__and2_1
XANTENNA__3305__A1 _0361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3409_ _0464_ _0480_ _0482_ _0484_ VGND VGND VPWR VPWR _0485_ sky130_fd_sc_hd__a22o_2
XANTENNA__4502__B1 _1343_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6128_ clknet_leaf_20_clk _0162_ net189 VGND VGND VPWR VPWR net120 sky130_fd_sc_hd__dfrtp_4
X_4389_ cu.reg_file.reg_l\[6\] _1317_ VGND VGND VPWR VPWR _1451_ sky130_fd_sc_hd__and2_1
XTAP_570 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4817__B cu.pc.pc_o\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5058__A1 _1051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_581 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4805__A1 _0359_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6059_ clknet_2_0__leaf_clk _0096_ net157 VGND VGND VPWR VPWR cu.reg_file.reg_sp\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_63_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3792__B2 cu.reg_file.reg_h\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3792__A1 cu.reg_file.reg_d\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_31_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5049__A1 _1263_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5839__A cu.reg_file.reg_sp\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5558__B _1330_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3232__B1 _0307_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3760_ cu.pc.pc_o\[14\] _0740_ _0834_ _0835_ VGND VGND VPWR VPWR _0836_ sky130_fd_sc_hd__a211o_1
XFILLER_0_54_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3783__A1 cu.pc.pc_o\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5430_ _2263_ VGND VGND VPWR VPWR _0184_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3691_ _0765_ _0766_ VGND VGND VPWR VPWR _0767_ sky130_fd_sc_hd__nand2_1
XFILLER_0_2_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5361_ _2222_ VGND VGND VPWR VPWR _0156_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4732__A0 cu.alu_f\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5292_ _2183_ VGND VGND VPWR VPWR _0126_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_77_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4312_ _1376_ _1374_ VGND VGND VPWR VPWR _1378_ sky130_fd_sc_hd__nand2_1
XFILLER_0_10_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4243_ _2883_ _0320_ _1310_ _0295_ _2914_ VGND VGND VPWR VPWR _1311_ sky130_fd_sc_hd__a2111o_2
X_4174_ _1242_ _1243_ _0600_ VGND VGND VPWR VPWR _1244_ sky130_fd_sc_hd__mux2_1
X_3125_ _2773_ _2775_ _2776_ _2862_ VGND VGND VPWR VPWR _2863_ sky130_fd_sc_hd__or4_1
X_3056_ _2759_ _2793_ ih.t.count\[20\] VGND VGND VPWR VPWR _2794_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4372__B _1434_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_45_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3958_ _1032_ _0807_ VGND VGND VPWR VPWR _1033_ sky130_fd_sc_hd__or2_1
XFILLER_0_18_456 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5484__A _2247_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3889_ _2897_ _0324_ VGND VGND VPWR VPWR _0965_ sky130_fd_sc_hd__nor2_1
XFILLER_0_18_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5628_ ih.gpio_interrupt_mask\[5\] _2326_ _2442_ _2125_ _2327_ VGND VGND VPWR VPWR
+ _2443_ sky130_fd_sc_hd__a221o_1
X_5559_ net102 _2205_ _2376_ _1401_ VGND VGND VPWR VPWR _2377_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5279__A1 _1189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3462__B1 _0498_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4282__B _1348_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3214__B1 _2948_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4962__A0 cu.pc.pc_o\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_36_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3517__A1 cu.reg_file.reg_l\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6302__RESET_B net160 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5333__S _2206_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4930_ _1902_ _1910_ VGND VGND VPWR VPWR _1922_ sky130_fd_sc_hd__or2b_1
XFILLER_0_59_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4861_ cu.pc.pc_o\[4\] _1858_ _1815_ VGND VGND VPWR VPWR _1859_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_59_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3812_ cu.reg_file.reg_b\[1\] _0743_ _0624_ cu.reg_file.reg_sp\[9\] VGND VGND VPWR
+ VPWR _0888_ sky130_fd_sc_hd__a22o_1
XFILLER_0_27_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_16 net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3756__A1 cu.reg_file.reg_mem\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4792_ _1793_ VGND VGND VPWR VPWR _1794_ sky130_fd_sc_hd__buf_2
XFILLER_0_27_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3743_ _0753_ _0778_ _0780_ _0818_ VGND VGND VPWR VPWR _0819_ sky130_fd_sc_hd__a211o_1
XFILLER_0_88_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3674_ cu.reg_file.reg_b\[0\] _0426_ _0429_ cu.reg_file.reg_d\[0\] VGND VGND VPWR
+ VPWR _0750_ sky130_fd_sc_hd__a22o_1
XFILLER_0_70_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5413_ _1190_ net136 _2248_ VGND VGND VPWR VPWR _2253_ sky130_fd_sc_hd__mux2_1
Xoutput101 net101 VGND VGND VPWR VPWR ss3[1] sky130_fd_sc_hd__clkbuf_4
XANTENNA__3508__B2 _0341_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput123 net123 VGND VGND VPWR VPWR ss5[7] sky130_fd_sc_hd__buf_2
Xoutput134 net134 VGND VGND VPWR VPWR ss7[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5344_ _2213_ VGND VGND VPWR VPWR _0148_ sky130_fd_sc_hd__clkbuf_1
Xoutput112 net112 VGND VGND VPWR VPWR ss4[4] sky130_fd_sc_hd__clkbuf_4
X_5275_ net78 _1074_ _2170_ VGND VGND VPWR VPWR _2173_ sky130_fd_sc_hd__mux2_1
X_4226_ _1293_ VGND VGND VPWR VPWR _1294_ sky130_fd_sc_hd__buf_2
XFILLER_0_49_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5681__A1 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4157_ _0935_ _0813_ VGND VGND VPWR VPWR _1227_ sky130_fd_sc_hd__xnor2_1
X_3108_ _2747_ _2845_ VGND VGND VPWR VPWR _2846_ sky130_fd_sc_hd__nand2_1
X_4088_ _0617_ _1050_ VGND VGND VPWR VPWR _1162_ sky130_fd_sc_hd__xor2_1
X_3039_ ih.t.timer_max\[25\] _2762_ ih.t.timer_max\[26\] VGND VGND VPWR VPWR _2777_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_77_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4944__A0 _1222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4830__B cu.pc.pc_o\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3747__B2 _0566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3446__B cu.id.cb_opcode_y\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5121__A0 _1622_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6195__D net2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_56_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput14 keypad_input[6] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_2
Xinput25 memory_data_in[7] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_64_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_543 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3356__B _0405_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5360__A0 _1194_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3390_ _0300_ _0353_ _2912_ VGND VGND VPWR VPWR _0466_ sky130_fd_sc_hd__a21oi_1
X_5060_ cu.reg_file.reg_c\[2\] _1074_ _2025_ VGND VGND VPWR VPWR _2028_ sky130_fd_sc_hd__mux2_1
X_4011_ _0606_ _0701_ _1083_ _0603_ _1084_ VGND VGND VPWR VPWR _1085_ sky130_fd_sc_hd__a221o_1
XANTENNA__3674__B1 _0429_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5415__A1 net137 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5962_ cu.id.imm_i\[12\] _2429_ _2686_ VGND VGND VPWR VPWR _2691_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4913_ _1906_ VGND VGND VPWR VPWR _0024_ sky130_fd_sc_hd__clkbuf_1
X_5893_ _2653_ VGND VGND VPWR VPWR _0257_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_62_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4844_ _1841_ _1842_ VGND VGND VPWR VPWR _1843_ sky130_fd_sc_hd__and2b_1
XFILLER_0_7_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4775_ _0976_ _0989_ _1780_ _0994_ VGND VGND VPWR VPWR _1781_ sky130_fd_sc_hd__or4b_1
X_3726_ _0645_ _0799_ VGND VGND VPWR VPWR _0802_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_43_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_70_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4982__B1_N _1798_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3657_ _0732_ VGND VGND VPWR VPWR _0733_ sky130_fd_sc_hd__buf_2
X_3588_ _0652_ _0663_ VGND VGND VPWR VPWR _0664_ sky130_fd_sc_hd__xnor2_4
X_5327_ _2203_ VGND VGND VPWR VPWR _0141_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5481__B _2284_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5103__A0 cu.reg_file.reg_e\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5258_ ih.t.timer_max\[28\] _2161_ _2153_ VGND VGND VPWR VPWR _2162_ sky130_fd_sc_hd__mux2_1
XANTENNA__5654__A1 _2467_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5189_ mc.cl.next_data\[15\] net25 mc.count VGND VGND VPWR VPWR _2112_ sky130_fd_sc_hd__mux2_1
X_4209_ _2883_ _2937_ VGND VGND VPWR VPWR _1277_ sky130_fd_sc_hd__or2_1
XFILLER_0_3_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5709__A2 _1650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_80_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3176__B _2878_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5672__A _1649_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout180 net182 VGND VGND VPWR VPWR net180 sky130_fd_sc_hd__clkbuf_4
Xfanout191 net194 VGND VGND VPWR VPWR net191 sky130_fd_sc_hd__clkbuf_4
XANTENNA_output139_A net139 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5847__A cu.reg_file.reg_sp\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1182 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1171 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1160 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4560_ cu.reg_file.reg_h\[7\] _1316_ _1312_ cu.reg_file.reg_b\[7\] _1612_ VGND VGND
+ VPWR VPWR _1613_ sky130_fd_sc_hd__a221o_1
XFILLER_0_37_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4384__A1 cu.reg_file.reg_a\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4384__B2 cu.reg_file.reg_sp\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4491_ _1546_ _1547_ VGND VGND VPWR VPWR _1548_ sky130_fd_sc_hd__and2_1
XFILLER_0_52_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3511_ _0576_ _0581_ _0586_ VGND VGND VPWR VPWR _0587_ sky130_fd_sc_hd__o21ai_4
X_6230_ clknet_leaf_14_clk ih.t.next_count\[18\] net180 VGND VGND VPWR VPWR ih.t.count\[18\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__5333__A0 _1052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3442_ _0401_ _0511_ _0513_ _0517_ VGND VGND VPWR VPWR _0518_ sky130_fd_sc_hd__o211a_1
XFILLER_0_40_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_900 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6161_ clknet_leaf_8_clk _0195_ net167 VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__dfrtp_2
X_3373_ _2894_ _2874_ _0309_ _2941_ _0378_ VGND VGND VPWR VPWR _0449_ sky130_fd_sc_hd__a32o_2
XANTENNA__4198__A _2877_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_944 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_933 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_922 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_911 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5112_ _2061_ VGND VGND VPWR VPWR _0068_ sky130_fd_sc_hd__clkbuf_1
X_6092_ clknet_leaf_23_clk _0126_ net192 VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__dfrtp_1
XTAP_977 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_966 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_955 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5636__A1 net130 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_999 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_988 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5636__B2 net138 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5043_ _1191_ _1209_ _2002_ VGND VGND VPWR VPWR _2016_ sky130_fd_sc_hd__mux2_1
XANTENNA__4926__A _2920_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4611__A2 _1644_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5945_ _2681_ VGND VGND VPWR VPWR _0281_ sky130_fd_sc_hd__clkbuf_1
X_5876_ _2644_ VGND VGND VPWR VPWR _0249_ sky130_fd_sc_hd__clkbuf_1
X_4827_ _1299_ cu.pc.pc_o\[1\] cu.pc.pc_o\[2\] VGND VGND VPWR VPWR _1827_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_7_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_457 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4758_ _1268_ _1300_ _1756_ _1301_ VGND VGND VPWR VPWR _1767_ sky130_fd_sc_hd__and4bb_1
X_4689_ net231 _1708_ _1687_ VGND VGND VPWR VPWR _1712_ sky130_fd_sc_hd__o21ai_1
X_3709_ _0762_ _0784_ VGND VGND VPWR VPWR _0785_ sky130_fd_sc_hd__and2b_1
XANTENNA__5324__A0 _1194_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4127__B2 _1032_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4127__A1 _0916_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5875__A1 ih.t.timer_max\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5627__A1 mc.cl.next_data\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3638__B1 _0545_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_14_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_435 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4290__B _1354_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4366__A1 _0373_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4366__B2 cu.pc.pc_o\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_218 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_229 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3005__A_N net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5341__S _2206_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold3 cu.id.interrupt_requested VGND VGND VPWR VPWR net199 sky130_fd_sc_hd__buf_1
XANTENNA__3629__B1 _0499_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_11_clk_A clknet_2_2__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3991_ _0758_ _0760_ _1064_ VGND VGND VPWR VPWR _1065_ sky130_fd_sc_hd__o21bai_1
X_5730_ net21 _2519_ _2525_ VGND VGND VPWR VPWR _0222_ sky130_fd_sc_hd__a21o_1
XANTENNA_clkbuf_leaf_26_clk_A clknet_2_3__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_71_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5661_ net83 _1633_ _2470_ _2473_ VGND VGND VPWR VPWR _2474_ sky130_fd_sc_hd__o22a_1
X_4612_ _2704_ _1647_ _1655_ VGND VGND VPWR VPWR mc.rw.next_state\[0\] sky130_fd_sc_hd__a21o_1
XFILLER_0_72_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5592_ _1649_ _2408_ VGND VGND VPWR VPWR _2409_ sky130_fd_sc_hd__and2_1
XFILLER_0_88_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4543_ cu.reg_file.reg_h\[6\] _1317_ _1313_ cu.reg_file.reg_b\[6\] _1596_ VGND VGND
+ VPWR VPWR _1597_ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4474_ _1512_ _1520_ _1531_ VGND VGND VPWR VPWR _1532_ sky130_fd_sc_hd__a21o_1
X_6213_ clknet_leaf_10_clk ih.t.next_count\[1\] net175 VGND VGND VPWR VPWR ih.t.count\[1\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_0_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3425_ _0500_ VGND VGND VPWR VPWR _0501_ sky130_fd_sc_hd__clkbuf_4
XTAP_752 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6144_ clknet_leaf_6_clk _0178_ net166 VGND VGND VPWR VPWR net136 sky130_fd_sc_hd__dfrtp_4
XANTENNA__3332__A2 _2878_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3356_ _0412_ _0405_ _0424_ VGND VGND VPWR VPWR _0432_ sky130_fd_sc_hd__and3b_2
X_6075_ clknet_leaf_21_clk _0109_ net189 VGND VGND VPWR VPWR ih.t.enable sky130_fd_sc_hd__dfrtp_1
XTAP_785 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3287_ _0360_ _0361_ _0362_ _0297_ _0296_ VGND VGND VPWR VPWR _0363_ sky130_fd_sc_hd__a2111oi_1
XFILLER_0_29_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5251__S _1667_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_796 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3560__A _0413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5026_ _1790_ _0352_ VGND VGND VPWR VPWR _2004_ sky130_fd_sc_hd__nand2_1
XANTENNA__4832__A2 cu.pc.pc_o\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4045__B1 _0663_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5928_ _0359_ _2429_ _2668_ VGND VGND VPWR VPWR _2673_ sky130_fd_sc_hd__mux2_1
XANTENNA__3399__A2 _2918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5859_ _2141_ _2320_ VGND VGND VPWR VPWR _2635_ sky130_fd_sc_hd__and2b_2
XFILLER_0_90_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4348__A1 cu.reg_file.reg_sp\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4348__B2 _0374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3571__A2 _0415_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4520__A1 cu.pc.pc_o\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3470__A _0296_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_58_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4587__A1 _1374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_62_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_output83_A net83 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3210_ cu.id.state\[1\] cu.id.state\[0\] VGND VGND VPWR VPWR _2947_ sky130_fd_sc_hd__nand2_2
XFILLER_0_5_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4190_ _1259_ VGND VGND VPWR VPWR _0013_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_66_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3141_ cu.id.opcode\[0\] cu.id.opcode\[2\] cu.id.opcode\[1\] VGND VGND VPWR VPWR
+ _2878_ sky130_fd_sc_hd__nand3b_4
X_3072_ ih.t.count\[14\] _2755_ _2809_ VGND VGND VPWR VPWR _2810_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3974_ _0558_ _1040_ _1043_ _1048_ VGND VGND VPWR VPWR _1049_ sky130_fd_sc_hd__a211o_1
X_5713_ _1328_ _1354_ _2274_ VGND VGND VPWR VPWR _2516_ sky130_fd_sc_hd__and3_1
X_5644_ _1400_ _2457_ VGND VGND VPWR VPWR _2458_ sky130_fd_sc_hd__and2b_1
XFILLER_0_60_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5575_ _2392_ VGND VGND VPWR VPWR _0200_ sky130_fd_sc_hd__clkbuf_1
X_4526_ _1396_ _1579_ VGND VGND VPWR VPWR _1581_ sky130_fd_sc_hd__nand2_1
XANTENNA__4750__B2 _1269_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3553__A2 _0501_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4457_ _1512_ _1513_ _1514_ _1334_ VGND VGND VPWR VPWR _1516_ sky130_fd_sc_hd__a31o_1
XANTENNA__4502__B2 cu.id.imm_i\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3408_ _0483_ _0463_ VGND VGND VPWR VPWR _0484_ sky130_fd_sc_hd__nor2_1
XANTENNA__4502__A1 cu.reg_file.reg_sp\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6127_ clknet_leaf_7_clk _0161_ net165 VGND VGND VPWR VPWR net119 sky130_fd_sc_hd__dfrtp_4
X_4388_ _0387_ _1295_ _1298_ cu.pc.pc_o\[6\] _1306_ VGND VGND VPWR VPWR _1450_ sky130_fd_sc_hd__a221o_1
XTAP_560 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3339_ _0414_ _0405_ _0412_ VGND VGND VPWR VPWR _0415_ sky130_fd_sc_hd__and3b_4
XTAP_571 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6058_ clknet_leaf_23_clk mc.cc.enable net192 VGND VGND VPWR VPWR mc.cc.enable_edge_detector.prev_data
+ sky130_fd_sc_hd__dfrtp_1
X_5009_ cu.reg_file.reg_a\[3\] _1991_ _1985_ VGND VGND VPWR VPWR _1992_ sky130_fd_sc_hd__mux2_1
XFILLER_0_36_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5518__B1 _1374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3792__A2 _0488_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3465__A cu.reg_file.reg_e\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6198__D net11 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4995__S _1814_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5757__A0 cu.reg_file.reg_sp\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3783__A2 _0740_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5855__A cu.reg_file.reg_sp\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3690_ _0718_ _0684_ VGND VGND VPWR VPWR _0766_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_42_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3375__A _2878_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5360_ _1194_ net114 _2215_ VGND VGND VPWR VPWR _2222_ sky130_fd_sc_hd__mux2_1
XANTENNA__4732__A1 alu.Cin VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5291_ _0619_ net84 _2182_ VGND VGND VPWR VPWR _2183_ sky130_fd_sc_hd__mux2_1
X_4311_ _1376_ _1348_ _1349_ _1335_ VGND VGND VPWR VPWR _1377_ sky130_fd_sc_hd__a22o_1
XFILLER_0_22_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4242_ _2908_ _0361_ _0968_ _0336_ VGND VGND VPWR VPWR _1310_ sky130_fd_sc_hd__o31a_1
X_4173_ _0747_ _0892_ _0447_ VGND VGND VPWR VPWR _1243_ sky130_fd_sc_hd__mux2_1
X_3124_ _2778_ _2779_ _2861_ VGND VGND VPWR VPWR _2862_ sky130_fd_sc_hd__or3_1
X_3055_ ih.t.timer_max\[19\] _2758_ ih.t.timer_max\[20\] VGND VGND VPWR VPWR _2793_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_26_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_fanout152_A net163 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_92_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3957_ _0401_ _0528_ VGND VGND VPWR VPWR _1032_ sky130_fd_sc_hd__or2_4
XFILLER_0_18_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_18_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3888_ _0620_ _0819_ _0823_ _0963_ VGND VGND VPWR VPWR _0964_ sky130_fd_sc_hd__a211o_1
X_5627_ mc.cl.next_data\[5\] _2313_ net141 _2441_ VGND VGND VPWR VPWR _2442_ sky130_fd_sc_hd__a22o_1
XFILLER_0_33_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5558_ net86 _1330_ VGND VGND VPWR VPWR _2376_ sky130_fd_sc_hd__or2_1
XFILLER_0_60_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5920__A0 _2923_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4509_ _1546_ _1563_ _1562_ VGND VGND VPWR VPWR _1565_ sky130_fd_sc_hd__a21o_1
X_5489_ net124 _2236_ _2247_ net132 _2308_ VGND VGND VPWR VPWR _2309_ sky130_fd_sc_hd__a221o_1
XTAP_390 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_38_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_38_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_95_132 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_30 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3462__A1 cu.reg_file.reg_d\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3462__B2 cu.alu_f\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_22_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3765__A2 _0640_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5614__S _2351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output46_A net46 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_29_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_29_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__4473__B _1530_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4860_ _1850_ _1857_ _1809_ VGND VGND VPWR VPWR _1858_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3811_ _0886_ VGND VGND VPWR VPWR _0887_ sky130_fd_sc_hd__inv_2
XFILLER_0_55_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4791_ _1186_ _1790_ _0352_ _1792_ VGND VGND VPWR VPWR _1793_ sky130_fd_sc_hd__or4_2
XANTENNA_17 net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3742_ _0776_ _0798_ _0815_ _0817_ VGND VGND VPWR VPWR _0818_ sky130_fd_sc_hd__a22o_1
XANTENNA__3756__A2 _0640_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3673_ cu.reg_file.reg_sp\[8\] _0636_ _0748_ cu.reg_file.reg_h\[0\] VGND VGND VPWR
+ VPWR _0749_ sky130_fd_sc_hd__a22o_1
XFILLER_0_88_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5412_ _2252_ VGND VGND VPWR VPWR _0177_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3508__A2 _0361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5343_ _1194_ net106 _2206_ VGND VGND VPWR VPWR _2213_ sky130_fd_sc_hd__mux2_1
Xoutput102 net102 VGND VGND VPWR VPWR ss3[2] sky130_fd_sc_hd__clkbuf_4
Xoutput113 net113 VGND VGND VPWR VPWR ss4[5] sky130_fd_sc_hd__clkbuf_4
Xoutput124 net124 VGND VGND VPWR VPWR ss6[0] sky130_fd_sc_hd__buf_2
Xoutput135 net135 VGND VGND VPWR VPWR ss7[3] sky130_fd_sc_hd__clkbuf_4
X_5274_ _2172_ VGND VGND VPWR VPWR _0119_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5130__A1 cu.reg_file.reg_h\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4225_ _2950_ _1292_ _1269_ VGND VGND VPWR VPWR _1293_ sky130_fd_sc_hd__and3_2
XANTENNA__5681__A2 _1650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4156_ _0516_ _1225_ VGND VGND VPWR VPWR _1226_ sky130_fd_sc_hd__nor2_4
X_3107_ ih.t.timer_max\[3\] _2746_ VGND VGND VPWR VPWR _2845_ sky130_fd_sc_hd__nand2_1
X_4087_ _1144_ _1160_ VGND VGND VPWR VPWR _1161_ sky130_fd_sc_hd__xor2_1
X_3038_ ih.t.count\[27\] _2764_ _2774_ VGND VGND VPWR VPWR _2776_ sky130_fd_sc_hd__and3_1
X_4989_ cu.pc.pc_o\[14\] _1968_ _1233_ VGND VGND VPWR VPWR _1976_ sky130_fd_sc_hd__o21a_1
XFILLER_0_73_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4839__A cu.pc.pc_o\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5121__A1 _0617_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput26 nrst VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_52_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput15 keypad_input[7] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5360__A1 net114 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5663__A2 _2204_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4010_ _0531_ _0694_ VGND VGND VPWR VPWR _1084_ sky130_fd_sc_hd__nor2_1
XFILLER_0_74_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4871__A0 _1144_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3674__B2 cu.reg_file.reg_d\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3674__A1 cu.reg_file.reg_b\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5961_ _2690_ VGND VGND VPWR VPWR _0288_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_87_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4912_ cu.pc.pc_o\[8\] _1905_ _1815_ VGND VGND VPWR VPWR _1906_ sky130_fd_sc_hd__mux2_1
XANTENNA__5179__A1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5892_ _1260_ ih.t.timer_max\[7\] _2645_ VGND VGND VPWR VPWR _2653_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4843_ cu.id.cb_opcode_y\[0\] cu.pc.pc_o\[3\] VGND VGND VPWR VPWR _1842_ sky130_fd_sc_hd__nand2_1
X_4774_ _2948_ _0986_ VGND VGND VPWR VPWR _1780_ sky130_fd_sc_hd__nand2_1
X_3725_ _0733_ _0800_ VGND VGND VPWR VPWR _0801_ sky130_fd_sc_hd__xnor2_2
Xclkbuf_leaf_9_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_9_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_70_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3656_ _0730_ _0731_ VGND VGND VPWR VPWR _0732_ sky130_fd_sc_hd__or2_1
XANTENNA__5254__S _1667_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_173 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3587_ _0653_ _0655_ _0657_ _0662_ VGND VGND VPWR VPWR _0663_ sky130_fd_sc_hd__o22a_4
X_5326_ _1261_ net99 _2195_ VGND VGND VPWR VPWR _2203_ sky130_fd_sc_hd__mux2_1
X_5257_ _1160_ _1213_ _1667_ VGND VGND VPWR VPWR _2161_ sky130_fd_sc_hd__mux2_1
XANTENNA__5103__A1 _2022_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4208_ _2912_ _2937_ _0583_ _1274_ VGND VGND VPWR VPWR _1276_ sky130_fd_sc_hd__a31o_4
X_5188_ _1646_ VGND VGND VPWR VPWR _2111_ sky130_fd_sc_hd__clkbuf_2
X_4139_ _1203_ _1208_ _0516_ VGND VGND VPWR VPWR _1209_ sky130_fd_sc_hd__a21oi_4
XFILLER_0_3_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_93_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_530 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5590__A1 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5953__A _2685_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout192 net193 VGND VGND VPWR VPWR net192 sky130_fd_sc_hd__clkbuf_4
Xfanout181 net182 VGND VGND VPWR VPWR net181 sky130_fd_sc_hd__clkbuf_4
Xfanout170 net173 VGND VGND VPWR VPWR net170 sky130_fd_sc_hd__clkbuf_4
XTAP_1150 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1183 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1172 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1161 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5339__S _2206_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5581__A1 net79 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_427 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3510_ _0294_ _0585_ _0576_ VGND VGND VPWR VPWR _0586_ sky130_fd_sc_hd__o21ai_2
X_4490_ _1333_ _1545_ VGND VGND VPWR VPWR _1547_ sky130_fd_sc_hd__nand2_1
XANTENNA__5333__A1 net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5074__S _2035_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3441_ _0395_ _0516_ VGND VGND VPWR VPWR _0517_ sky130_fd_sc_hd__nand2_2
XTAP_901 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6160_ clknet_leaf_18_clk _0194_ net173 VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__dfrtp_4
X_3372_ _2925_ _0313_ _0325_ _2910_ _2879_ VGND VGND VPWR VPWR _0448_ sky130_fd_sc_hd__a2111oi_2
XTAP_934 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_923 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_912 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3895__B2 _2923_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3895__A1 _2893_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5111_ cu.reg_file.reg_e\[4\] _1189_ _2056_ VGND VGND VPWR VPWR _2061_ sky130_fd_sc_hd__mux2_1
XTAP_978 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_967 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_956 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_945 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6091_ clknet_leaf_19_clk _0125_ net190 VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__dfrtp_4
XANTENNA__5636__A2 _2236_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_989 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4926__B _1521_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5042_ _2015_ VGND VGND VPWR VPWR _0044_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_18_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5944_ _0374_ _2429_ _2666_ VGND VGND VPWR VPWR _2681_ sky130_fd_sc_hd__mux2_1
X_5875_ _2167_ ih.t.timer_max\[15\] _2636_ VGND VGND VPWR VPWR _2644_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_75_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4826_ _1299_ cu.pc.pc_o\[1\] cu.pc.pc_o\[2\] VGND VGND VPWR VPWR _1826_ sky130_fd_sc_hd__and3_1
XANTENNA__5021__A0 cu.reg_file.reg_a\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_90_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4757_ _1761_ _1764_ _1765_ VGND VGND VPWR VPWR _1766_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_31_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4688_ ih.t.count\[18\] _1708_ VGND VGND VPWR VPWR _1711_ sky130_fd_sc_hd__and2_1
X_3708_ _0710_ _0587_ VGND VGND VPWR VPWR _0784_ sky130_fd_sc_hd__and2b_1
XANTENNA__5324__A1 net98 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4389__A cu.reg_file.reg_l\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3639_ _0587_ _0710_ VGND VGND VPWR VPWR _0715_ sky130_fd_sc_hd__nor2_1
XFILLER_0_31_558 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3335__B1 _2877_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3293__A _2951_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5309_ _2192_ VGND VGND VPWR VPWR _2193_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__3886__A1 _0918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6289_ clknet_leaf_41_clk _0271_ net151 VGND VGND VPWR VPWR cu.id.opcode\[2\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__3740__B _0528_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4852__A cu.pc.pc_o\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5260__A0 _1144_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5012__A0 cu.reg_file.reg_a\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3187__B _2923_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5563__A1 ih.t.timer_max\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5563__B2 ih.t.timer_max\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_34_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3915__B _0968_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_219 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_208 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xhold4 _0001_ VGND VGND VPWR VPWR net200 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3629__A1 cu.reg_file.reg_h\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3629__B2 cu.reg_file.reg_a\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5251__A0 _1073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3990_ _0761_ _0772_ _0777_ VGND VGND VPWR VPWR _1064_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_69_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5660_ net115 _2146_ _2225_ net123 _2472_ VGND VGND VPWR VPWR _2473_ sky130_fd_sc_hd__a221o_1
XFILLER_0_57_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5003__A0 cu.reg_file.reg_a\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3378__A _0379_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4611_ _1650_ _1644_ _1651_ _1654_ VGND VGND VPWR VPWR _1655_ sky130_fd_sc_hd__a31o_1
XFILLER_0_72_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5591_ net11 _2345_ _2369_ net4 VGND VGND VPWR VPWR _2408_ sky130_fd_sc_hd__a22o_1
XANTENNA__5554__A1 _2372_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4542_ cu.pc.pc_o\[14\] _1322_ _1315_ cu.reg_file.reg_d\[6\] _1595_ VGND VGND VPWR
+ VPWR _1596_ sky130_fd_sc_hd__a221o_1
X_4473_ _1332_ _1530_ VGND VGND VPWR VPWR _1531_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_4_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_536 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_13_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6212_ clknet_leaf_10_clk ih.t.next_count\[0\] net176 VGND VGND VPWR VPWR ih.t.count\[0\]
+ sky130_fd_sc_hd__dfrtp_4
X_3424_ cu.id.starting_int_service net149 VGND VGND VPWR VPWR _0500_ sky130_fd_sc_hd__or2_1
Xmax_cap145 net236 VGND VGND VPWR VPWR net145 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_40_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6143_ clknet_leaf_8_clk _0177_ net168 VGND VGND VPWR VPWR net135 sky130_fd_sc_hd__dfrtp_1
XTAP_742 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5532__S _2351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3355_ cu.reg_file.reg_c\[0\] _0427_ _0430_ cu.reg_file.reg_e\[0\] VGND VGND VPWR
+ VPWR _0431_ sky130_fd_sc_hd__a22o_1
X_6074_ clknet_leaf_16_clk _0108_ net181 VGND VGND VPWR VPWR ih.gpio_interrupt_mask\[7\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_786 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3286_ _2888_ _2890_ _2933_ _2934_ VGND VGND VPWR VPWR _0362_ sky130_fd_sc_hd__and4_1
XTAP_797 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5025_ _0618_ _1622_ _2002_ VGND VGND VPWR VPWR _2003_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout182_A net196 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5490__B1 _2193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5768__A cu.reg_file.reg_sp\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_48_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5927_ _2672_ VGND VGND VPWR VPWR _0272_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5858_ _2634_ VGND VGND VPWR VPWR _0241_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5545__A1 _1666_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4809_ _1301_ _1775_ _1779_ _1268_ VGND VGND VPWR VPWR _1811_ sky130_fd_sc_hd__o22ai_1
XFILLER_0_16_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5789_ cu.reg_file.reg_sp\[6\] _2574_ _2539_ VGND VGND VPWR VPWR _2575_ sky130_fd_sc_hd__mux2_1
XANTENNA__4348__A2 _0993_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4566__B _1614_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3470__B _0528_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5678__A _1489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4582__A _1579_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_54_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_255 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_22_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_22_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output76_A net76 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5352__S _2215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3140_ _2875_ _2876_ VGND VGND VPWR VPWR _2877_ sky130_fd_sc_hd__nand2b_4
X_3071_ ih.t.timer_max\[13\] _2754_ ih.t.timer_max\[14\] VGND VGND VPWR VPWR _2809_
+ sky130_fd_sc_hd__o21ai_1
XANTENNA__3483__C1 cu.reg_file.reg_l\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_15_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5712_ net193 _2707_ _2514_ _2515_ VGND VGND VPWR VPWR _0214_ sky130_fd_sc_hd__a31o_1
XFILLER_0_85_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3973_ _0574_ _0822_ _1046_ _0545_ _1047_ VGND VGND VPWR VPWR _1048_ sky130_fd_sc_hd__a221o_1
XANTENNA__3786__B1 _0748_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6037__RESET_B net188 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5643_ ih.t.timer_max\[14\] _2193_ _2314_ ih.t.timer_max\[6\] _2456_ VGND VGND VPWR
+ VPWR _2457_ sky130_fd_sc_hd__a221o_1
XFILLER_0_72_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5527__A1 net2 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5574_ cu.reg_file.reg_mem\[2\] _2391_ _2351_ VGND VGND VPWR VPWR _2392_ sky130_fd_sc_hd__mux2_1
XFILLER_0_31_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4525_ _1396_ _1579_ VGND VGND VPWR VPWR _1580_ sky130_fd_sc_hd__or2_1
XFILLER_0_13_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4456_ _1512_ _1513_ _1514_ VGND VGND VPWR VPWR _1515_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_13_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4387_ _1271_ _1448_ VGND VGND VPWR VPWR _1449_ sky130_fd_sc_hd__nor2_1
X_3407_ net147 _0454_ _0457_ VGND VGND VPWR VPWR _0483_ sky130_fd_sc_hd__a21o_1
X_6126_ clknet_leaf_7_clk _0160_ net165 VGND VGND VPWR VPWR net118 sky130_fd_sc_hd__dfrtp_4
X_3338_ _0293_ _0407_ _0408_ VGND VGND VPWR VPWR _0414_ sky130_fd_sc_hd__or3b_4
XTAP_550 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6057_ clknet_leaf_24_clk _0095_ net190 VGND VGND VPWR VPWR mc.cl.next_data\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3269_ _0340_ _0341_ _0342_ _0344_ VGND VGND VPWR VPWR _0345_ sky130_fd_sc_hd__o211a_1
X_5008_ _1187_ _1222_ _0368_ VGND VGND VPWR VPWR _1991_ sky130_fd_sc_hd__mux2_1
XANTENNA__5215__A0 _1075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_48_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_36_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5518__A1 net33 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_10_clk_A clknet_2_2__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_25_clk_A clknet_2_3__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4257__A1 _0343_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output114_A net114 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4743__C _0379_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3359__C _0379_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_42_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4310_ mc.rw.state\[2\] _2699_ VGND VGND VPWR VPWR _1376_ sky130_fd_sc_hd__nand2_1
X_5290_ _2180_ _2181_ VGND VGND VPWR VPWR _2182_ sky130_fd_sc_hd__nand2_8
XFILLER_0_50_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4241_ _0336_ _0436_ _1308_ _0295_ VGND VGND VPWR VPWR _1309_ sky130_fd_sc_hd__a211o_2
X_4172_ _0871_ _0902_ _1060_ VGND VGND VPWR VPWR _1242_ sky130_fd_sc_hd__mux2_1
X_3123_ _2781_ _2783_ _2784_ _2860_ VGND VGND VPWR VPWR _2861_ sky130_fd_sc_hd__or4_1
X_3054_ _2760_ _2790_ ih.t.count\[21\] VGND VGND VPWR VPWR _2792_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_89_174 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_65_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_9_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4950__A cu.pc.pc_o\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3956_ _1030_ _1029_ _0773_ VGND VGND VPWR VPWR _1031_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_9_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3759__B1 _0624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5626_ _1666_ _2439_ _2440_ VGND VGND VPWR VPWR _2441_ sky130_fd_sc_hd__o21a_1
XANTENNA__5257__S _1667_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3887_ _0824_ _0915_ _0962_ VGND VGND VPWR VPWR _0963_ sky130_fd_sc_hd__and3_1
X_5557_ net94 _2194_ _2374_ VGND VGND VPWR VPWR _2375_ sky130_fd_sc_hd__a21o_1
XANTENNA__5920__A1 _2350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4508_ _1546_ _1562_ _1563_ VGND VGND VPWR VPWR _1564_ sky130_fd_sc_hd__nand3_1
X_5488_ net84 _2180_ _2224_ net116 VGND VGND VPWR VPWR _2308_ sky130_fd_sc_hd__a22o_1
X_4439_ _1497_ _1480_ _1481_ VGND VGND VPWR VPWR _1499_ sky130_fd_sc_hd__nand3_1
Xwire2 _0481_ VGND VGND VPWR VPWR net237 sky130_fd_sc_hd__buf_1
XANTENNA__5684__B1 cu.reg_file.reg_mem\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4487__B2 cu.reg_file.reg_b\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4487__A1 cu.reg_file.reg_h\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6109_ clknet_leaf_27_clk _0143_ net186 VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__dfrtp_4
XANTENNA__4239__A1 _0343_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_380 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4239__B2 _1299_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3462__A2 _0492_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_42 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_36_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3476__A _0528_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_288 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4478__A1 _1530_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_86_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3810_ _0882_ _0885_ VGND VGND VPWR VPWR _0886_ sky130_fd_sc_hd__xor2_1
X_4790_ _1791_ _0366_ VGND VGND VPWR VPWR _1792_ sky130_fd_sc_hd__or2_2
XFILLER_0_6_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3741_ _0816_ VGND VGND VPWR VPWR _0817_ sky130_fd_sc_hd__buf_2
XANTENNA_18 net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3610__C1 cu.reg_file.reg_l\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3672_ _0417_ _0421_ VGND VGND VPWR VPWR _0748_ sky130_fd_sc_hd__nor2_4
X_5411_ _1188_ net135 _2248_ VGND VGND VPWR VPWR _2252_ sky130_fd_sc_hd__mux2_1
Xoutput114 net114 VGND VGND VPWR VPWR ss4[6] sky130_fd_sc_hd__clkbuf_4
Xoutput125 net125 VGND VGND VPWR VPWR ss6[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_88_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5342_ _2212_ VGND VGND VPWR VPWR _0147_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3913__B1 _0296_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput103 net103 VGND VGND VPWR VPWR ss3[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_23_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput136 net136 VGND VGND VPWR VPWR ss7[4] sky130_fd_sc_hd__clkbuf_4
X_5273_ net77 _1051_ _2170_ VGND VGND VPWR VPWR _2172_ sky130_fd_sc_hd__mux2_1
XANTENNA__4469__A1 cu.reg_file.reg_sp\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4469__B2 cu.id.imm_i\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4224_ _2904_ _2924_ VGND VGND VPWR VPWR _1292_ sky130_fd_sc_hd__nand2_1
X_4155_ _0955_ _1215_ _1216_ _0952_ _1224_ VGND VGND VPWR VPWR _1225_ sky130_fd_sc_hd__o221a_1
X_3106_ _2749_ _2835_ ih.t.count\[4\] VGND VGND VPWR VPWR _2844_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_37_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4086_ _1159_ VGND VGND VPWR VPWR _1160_ sky130_fd_sc_hd__buf_4
X_3037_ _2764_ _2774_ ih.t.count\[27\] VGND VGND VPWR VPWR _2775_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_77_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5776__A cu.reg_file.reg_sp\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4988_ cu.pc.pc_o\[15\] _1963_ VGND VGND VPWR VPWR _1975_ sky130_fd_sc_hd__xor2_1
XFILLER_0_18_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3939_ _0983_ _0996_ _1003_ _1011_ _1014_ VGND VGND VPWR VPWR _1015_ sky130_fd_sc_hd__a2111o_1
XANTENNA__3296__A cu.id.cb_opcode_x\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5609_ _2169_ _2417_ _2424_ _2136_ VGND VGND VPWR VPWR _2425_ sky130_fd_sc_hd__o211a_1
XANTENNA__5409__A0 _1075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4590__A _1415_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3821__B_N _0892_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput27 programmable_gpio_in[0] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_64_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xinput16 keypad_input[8] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__buf_2
XFILLER_0_52_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5360__S _2215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3674__A2 _0426_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5960_ cu.id.imm_i\[11\] _2410_ _2686_ VGND VGND VPWR VPWR _2690_ sky130_fd_sc_hd__mux2_1
XANTENNA__3595__A1_N _0576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5820__A0 _1226_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5891_ _2652_ VGND VGND VPWR VPWR _0256_ sky130_fd_sc_hd__clkbuf_1
X_4911_ _1896_ _1904_ _1809_ VGND VGND VPWR VPWR _1905_ sky130_fd_sc_hd__mux2_1
XFILLER_0_47_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4842_ cu.id.cb_opcode_y\[0\] cu.pc.pc_o\[3\] VGND VGND VPWR VPWR _1841_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_28_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4773_ net206 _1779_ VGND VGND VPWR VPWR _0006_ sky130_fd_sc_hd__nor2_1
XFILLER_0_23_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_553 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_15_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3724_ _0644_ _0799_ _0790_ VGND VGND VPWR VPWR _0800_ sky130_fd_sc_hd__a21oi_1
X_3655_ _0566_ _0729_ VGND VGND VPWR VPWR _0731_ sky130_fd_sc_hd__nor2_1
XANTENNA__4139__B1 _0516_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_2_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3586_ _0659_ _0660_ _0661_ VGND VGND VPWR VPWR _0662_ sky130_fd_sc_hd__or3_2
X_5325_ _2202_ VGND VGND VPWR VPWR _0140_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5256_ _2160_ VGND VGND VPWR VPWR _0113_ sky130_fd_sc_hd__clkbuf_1
X_4207_ _2912_ _0583_ _1273_ _1274_ VGND VGND VPWR VPWR _1275_ sky130_fd_sc_hd__a31o_2
X_5187_ _2110_ VGND VGND VPWR VPWR _0094_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4394__B _1455_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4138_ _0916_ _0943_ _1206_ _0950_ _1207_ VGND VGND VPWR VPWR _1208_ sky130_fd_sc_hd__o221a_1
XFILLER_0_64_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4069_ _1135_ _1138_ _1141_ _1142_ VGND VGND VPWR VPWR _1143_ sky130_fd_sc_hd__or4_1
XFILLER_0_19_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_80_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5590__A2 _1648_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5878__A0 _2022_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3904__D _2935_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xfanout182 net196 VGND VGND VPWR VPWR net182 sky130_fd_sc_hd__buf_2
XANTENNA__4585__A _1393_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout171 net173 VGND VGND VPWR VPWR net171 sky130_fd_sc_hd__buf_2
Xfanout160 net162 VGND VGND VPWR VPWR net160 sky130_fd_sc_hd__buf_2
Xfanout193 net194 VGND VGND VPWR VPWR net193 sky130_fd_sc_hd__buf_2
XFILLER_0_69_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1140 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1173 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1162 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1151 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_60_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5581__A2 _1633_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_439 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_52_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3664__A _0501_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3440_ _0515_ VGND VGND VPWR VPWR _0516_ sky130_fd_sc_hd__buf_8
XFILLER_0_20_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3344__B2 cu.reg_file.reg_h\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3371_ _0416_ _0420_ _0441_ _0446_ VGND VGND VPWR VPWR _0447_ sky130_fd_sc_hd__o31a_4
XTAP_935 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_924 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_913 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_902 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6090_ clknet_leaf_4_clk _0124_ net172 VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__dfrtp_4
X_5110_ _2060_ VGND VGND VPWR VPWR _0067_ sky130_fd_sc_hd__clkbuf_1
XTAP_968 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_957 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_946 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5041_ cu.reg_file.reg_b\[4\] _2014_ _2006_ VGND VGND VPWR VPWR _2015_ sky130_fd_sc_hd__mux2_1
XTAP_979 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5090__S _2039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5943_ _2680_ VGND VGND VPWR VPWR _0280_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_34_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5874_ _2643_ VGND VGND VPWR VPWR _0248_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3280__B1 _2883_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4825_ _1825_ VGND VGND VPWR VPWR _0017_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_47_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_16_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_394 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4756_ _1268_ _1301_ _1300_ VGND VGND VPWR VPWR _1765_ sky130_fd_sc_hd__or3b_1
XFILLER_0_7_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3583__A1 cu.reg_file.reg_sp\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4687_ _1710_ VGND VGND VPWR VPWR ih.t.next_count\[17\] sky130_fd_sc_hd__clkbuf_1
X_3707_ _0781_ _0712_ _0782_ VGND VGND VPWR VPWR _0783_ sky130_fd_sc_hd__a21bo_1
XANTENNA__4780__B1 _0350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3638_ _0712_ _0713_ _0545_ _0599_ VGND VGND VPWR VPWR _0714_ sky130_fd_sc_hd__a2bb2o_1
X_3569_ _0644_ VGND VGND VPWR VPWR _0645_ sky130_fd_sc_hd__inv_2
XANTENNA__3293__B _0368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5308_ _1374_ _2191_ VGND VGND VPWR VPWR _2192_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3886__A2 _0779_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6288_ clknet_leaf_41_clk _0270_ net151 VGND VGND VPWR VPWR cu.id.opcode\[1\] sky130_fd_sc_hd__dfrtp_4
X_5239_ _2146_ VGND VGND VPWR VPWR _2147_ sky130_fd_sc_hd__buf_4
XANTENNA__5260__A1 _1209_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5563__A2 _2193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_46_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3574__B2 cu.reg_file.reg_a\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_209 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3629__A2 _0495_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xhold5 cu.id.is_interrupted VGND VGND VPWR VPWR net201 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5251__A1 _1226_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_423 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_84_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4610_ _2701_ _2706_ _1653_ VGND VGND VPWR VPWR _1654_ sky130_fd_sc_hd__mux2_1
X_5590_ net71 _1648_ _2137_ _2274_ VGND VGND VPWR VPWR _2407_ sky130_fd_sc_hd__a31o_1
XFILLER_0_4_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_515 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_20_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3565__B2 cu.reg_file.reg_a\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4541_ cu.reg_file.reg_sp\[14\] _0992_ _1344_ cu.id.imm_i\[14\] _1324_ VGND VGND
+ VPWR VPWR _1595_ sky130_fd_sc_hd__a221o_1
X_4472_ _1305_ _1526_ _1529_ VGND VGND VPWR VPWR _1530_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_20_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6211_ clknet_leaf_4_clk ih.ih.int_f.data_in net172 VGND VGND VPWR VPWR ih.ih.int_f.prev_data
+ sky130_fd_sc_hd__dfrtp_1
X_3423_ net146 _0473_ net145 _0486_ _0458_ VGND VGND VPWR VPWR _0499_ sky130_fd_sc_hd__o2111a_4
Xmax_cap146 _0468_ VGND VGND VPWR VPWR net146 sky130_fd_sc_hd__clkbuf_4
X_6142_ clknet_leaf_9_clk _0176_ net175 VGND VGND VPWR VPWR net134 sky130_fd_sc_hd__dfrtp_1
XTAP_710 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3354_ _0425_ _0414_ _0429_ VGND VGND VPWR VPWR _0430_ sky130_fd_sc_hd__o21bai_4
X_6073_ clknet_leaf_17_clk _0107_ net172 VGND VGND VPWR VPWR ih.gpio_interrupt_mask\[6\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_776 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3841__B _0916_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3285_ _0342_ VGND VGND VPWR VPWR _0361_ sky130_fd_sc_hd__clkbuf_4
XTAP_798 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5024_ _2001_ VGND VGND VPWR VPWR _2002_ sky130_fd_sc_hd__buf_4
XANTENNA__5490__A1 net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5490__B2 net92 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4953__A _2920_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5926_ _2893_ _2410_ _2668_ VGND VGND VPWR VPWR _2672_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_264 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_467 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_90_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_426 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5784__A cu.reg_file.reg_sp\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5857_ cu.reg_file.reg_sp\[15\] _2633_ _2538_ VGND VGND VPWR VPWR _2634_ sky130_fd_sc_hd__mux2_1
X_4808_ _1788_ _1800_ _1809_ VGND VGND VPWR VPWR _1810_ sky130_fd_sc_hd__mux2_1
X_5788_ _1126_ _2573_ _2545_ VGND VGND VPWR VPWR _2574_ sky130_fd_sc_hd__mux2_1
X_4739_ _1012_ _1747_ VGND VGND VPWR VPWR _1748_ sky130_fd_sc_hd__or2_1
XFILLER_0_31_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6170__CLK clknet_2_1__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4863__A cu.pc.pc_o\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3492__B1 _0545_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3994__A1_N _0918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3795__A1 cu.id.imm_i\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4992__A0 _1263_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3547__A1 cu.reg_file.reg_c\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_239 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_66_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output69_A net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3070_ ih.t.count\[15\] _2756_ _2806_ VGND VGND VPWR VPWR _2808_ sky130_fd_sc_hd__and3_1
XANTENNA_wire143_A _1280_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5711_ net193 mc.cl.cmp_o VGND VGND VPWR VPWR _2515_ sky130_fd_sc_hd__and2b_1
XFILLER_0_57_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4983__A0 _1624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3972_ _0531_ _0545_ VGND VGND VPWR VPWR _1047_ sky130_fd_sc_hd__nor2_1
XANTENNA__3786__A1 cu.reg_file.reg_sp\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_426 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3786__B2 cu.reg_file.reg_h\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5642_ ih.t.timer_max\[30\] _2146_ _2149_ ih.t.timer_max\[22\] VGND VGND VPWR VPWR
+ _2456_ sky130_fd_sc_hd__a22o_1
XFILLER_0_31_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5573_ _2387_ _2388_ _2390_ _1641_ VGND VGND VPWR VPWR _2391_ sky130_fd_sc_hd__o22a_2
X_4524_ _1304_ _1575_ _1578_ VGND VGND VPWR VPWR _1579_ sky130_fd_sc_hd__o21a_2
XFILLER_0_13_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_40_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4455_ _1396_ _1496_ _1498_ VGND VGND VPWR VPWR _1514_ sky130_fd_sc_hd__a21bo_1
X_4386_ cu.reg_file.reg_c\[6\] _1281_ _1447_ VGND VGND VPWR VPWR _1448_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_0_261 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3406_ net146 _0473_ net145 VGND VGND VPWR VPWR _0482_ sky130_fd_sc_hd__nor3_4
X_6125_ clknet_leaf_9_clk _0159_ net175 VGND VGND VPWR VPWR net117 sky130_fd_sc_hd__dfrtp_1
X_3337_ _0405_ _0407_ _0409_ _0412_ VGND VGND VPWR VPWR _0413_ sky130_fd_sc_hd__and4bb_4
XTAP_540 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_562 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6056_ clknet_leaf_22_clk _0094_ net191 VGND VGND VPWR VPWR mc.cl.next_data\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_3268_ _0343_ cu.id.cb_opcode_z\[1\] cu.id.cb_opcode_z\[2\] VGND VGND VPWR VPWR _0344_
+ sky130_fd_sc_hd__nand3_1
XTAP_595 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5007_ _1990_ VGND VGND VPWR VPWR _0034_ sky130_fd_sc_hd__clkbuf_1
X_3199_ _2884_ VGND VGND VPWR VPWR _2936_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_95_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_95_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3299__A _0373_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3777__A1 cu.reg_file.reg_mem\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5909_ ih.t.timer_max\[23\] _1260_ _2654_ VGND VGND VPWR VPWR _2662_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4032__A1_N alu.Cin VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5454__A1 _1369_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4257__A2 _2950_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4593__A _1434_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_86_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3002__A net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output107_A net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6170__RESET_B net161 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5390__A0 _1075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_120 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_77_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4240_ _0359_ _0320_ _0336_ _2914_ VGND VGND VPWR VPWR _1308_ sky130_fd_sc_hd__a211oi_1
XFILLER_0_22_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5693__A1 net4 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4171_ _1239_ _1240_ _0600_ VGND VGND VPWR VPWR _1241_ sky130_fd_sc_hd__mux2_1
X_3122_ _2786_ _2787_ _2859_ VGND VGND VPWR VPWR _2860_ sky130_fd_sc_hd__or3_1
XFILLER_0_93_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3053_ ih.t.count\[21\] _2760_ _2790_ VGND VGND VPWR VPWR _2791_ sky130_fd_sc_hd__and3_1
XFILLER_0_89_186 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3824__A1_N _0892_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_370 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4956__B1 _1233_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3955_ _0511_ VGND VGND VPWR VPWR _1030_ sky130_fd_sc_hd__inv_2
XFILLER_0_18_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3759__B2 cu.reg_file.reg_sp\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3759__A1 cu.reg_file.reg_b\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5625_ ih.t.timer_max\[21\] _2150_ _2319_ ih.t.timer_max\[5\] _1661_ VGND VGND VPWR
+ VPWR _2440_ sky130_fd_sc_hd__a221o_1
X_3886_ _0918_ _0779_ _0932_ _0947_ _0961_ VGND VGND VPWR VPWR _0962_ sky130_fd_sc_hd__a311o_1
XANTENNA__5381__A0 _1261_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5556_ net126 _2236_ _2247_ net134 VGND VGND VPWR VPWR _2374_ sky130_fd_sc_hd__a22o_1
XFILLER_0_13_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4507_ _1333_ _1545_ _1549_ VGND VGND VPWR VPWR _1563_ sky130_fd_sc_hd__a21o_1
XANTENNA__5273__S _2170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5487_ _2307_ VGND VGND VPWR VPWR _0197_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4438_ _1480_ _1481_ _1497_ VGND VGND VPWR VPWR _1498_ sky130_fd_sc_hd__a21o_1
XANTENNA__5684__B2 _1646_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xwire3 _2895_ VGND VGND VPWR VPWR net238 sky130_fd_sc_hd__buf_1
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4369_ cu.pc.pc_o\[5\] _1322_ _1315_ cu.reg_file.reg_e\[5\] _1431_ VGND VGND VPWR
+ VPWR _1432_ sky130_fd_sc_hd__a221o_1
X_6108_ clknet_leaf_26_clk _0142_ net195 VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__dfrtp_4
XTAP_370 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6039_ clknet_leaf_33_clk _0077_ net161 VGND VGND VPWR VPWR cu.reg_file.reg_h\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_68_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4947__A0 cu.pc.pc_o\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_87 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_470 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_259 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_59_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3989__B2 _0545_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5358__S _2215_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3740_ _0401_ _0528_ VGND VGND VPWR VPWR _0816_ sky130_fd_sc_hd__nor2_1
XANTENNA_19 net49 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_395 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3671_ cu.id.imm_i\[8\] _0739_ _0746_ _0653_ VGND VGND VPWR VPWR _0747_ sky130_fd_sc_hd__a22oi_4
X_5410_ _2251_ VGND VGND VPWR VPWR _0176_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_42_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput115 net115 VGND VGND VPWR VPWR ss4[7] sky130_fd_sc_hd__buf_2
XFILLER_0_88_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput104 net104 VGND VGND VPWR VPWR ss3[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_70_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5341_ _1192_ net105 _2206_ VGND VGND VPWR VPWR _2212_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5093__S _2039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput137 net137 VGND VGND VPWR VPWR ss7[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_23_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput126 net126 VGND VGND VPWR VPWR ss6[2] sky130_fd_sc_hd__clkbuf_4
XANTENNA__5666__A1 _1665_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5272_ _2171_ VGND VGND VPWR VPWR _0118_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_56_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4223_ _1271_ _1290_ VGND VGND VPWR VPWR _1291_ sky130_fd_sc_hd__nor2_1
X_4154_ _0817_ _0939_ _1223_ _0938_ VGND VGND VPWR VPWR _1224_ sky130_fd_sc_hd__o2bb2a_1
X_3105_ ih.t.count\[4\] _2749_ _2835_ _2842_ VGND VGND VPWR VPWR _2843_ sky130_fd_sc_hd__a31o_1
X_4085_ _1150_ _1151_ _1152_ _1158_ VGND VGND VPWR VPWR _1159_ sky130_fd_sc_hd__or4b_1
XANTENNA__3429__B1 _0502_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3036_ ih.t.timer_max\[27\] _2763_ VGND VGND VPWR VPWR _2774_ sky130_fd_sc_hd__nand2_1
XFILLER_0_77_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4929__B1 _1233_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_24_clk_A clknet_2_3__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4987_ _1974_ VGND VGND VPWR VPWR _0030_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_46_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3938_ alu.Cin _1013_ _1012_ VGND VGND VPWR VPWR _1014_ sky130_fd_sc_hd__o21a_1
XFILLER_0_18_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5792__A cu.reg_file.reg_sp\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3869_ _0942_ _0943_ _0944_ VGND VGND VPWR VPWR _0945_ sky130_fd_sc_hd__and3_1
X_5608_ ih.gpio_interrupt_mask\[4\] _2326_ _2423_ _2125_ _2327_ VGND VGND VPWR VPWR
+ _2424_ sky130_fd_sc_hd__a221o_1
XFILLER_0_61_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5354__A0 _1188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5539_ net77 _1633_ _2354_ _2357_ VGND VGND VPWR VPWR _2358_ sky130_fd_sc_hd__o22a_1
XFILLER_0_14_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5657__A1 net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3668__B1 _0624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5409__A1 net134 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput17 keypad_input[9] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_4
Xinput28 programmable_gpio_in[1] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__buf_1
XFILLER_0_64_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5345__A0 _1261_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_32_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4320__A1 cu.reg_file.reg_e\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4320__B2 cu.reg_file.reg_l\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_90_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5890_ _1193_ ih.t.timer_max\[6\] _2645_ VGND VGND VPWR VPWR _2652_ sky130_fd_sc_hd__mux2_1
X_4910_ _1799_ _1897_ _1902_ _1903_ VGND VGND VPWR VPWR _1904_ sky130_fd_sc_hd__a22o_1
XFILLER_0_59_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_90_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_87_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4841_ _1838_ _1839_ VGND VGND VPWR VPWR _1840_ sky130_fd_sc_hd__nor2_1
XFILLER_0_7_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4772_ _1301_ _1777_ _1778_ _1303_ VGND VGND VPWR VPWR _1779_ sky130_fd_sc_hd__o211a_1
XFILLER_0_28_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_43_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3723_ _0664_ _0684_ _0787_ _0794_ VGND VGND VPWR VPWR _0799_ sky130_fd_sc_hd__a31o_1
XFILLER_0_43_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3654_ _0566_ _0729_ VGND VGND VPWR VPWR _0730_ sky130_fd_sc_hd__and2_1
XFILLER_0_11_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3585_ cu.reg_file.reg_c\[5\] _0485_ _0621_ cu.reg_file.reg_l\[5\] VGND VGND VPWR
+ VPWR _0661_ sky130_fd_sc_hd__a22o_1
XANTENNA__5639__A1 net106 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5324_ _1194_ net98 _2195_ VGND VGND VPWR VPWR _2202_ sky130_fd_sc_hd__mux2_1
XFILLER_0_2_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5255_ ih.t.timer_max\[27\] _2159_ _2153_ VGND VGND VPWR VPWR _2160_ sky130_fd_sc_hd__mux2_1
XANTENNA__5639__B2 _1401_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4311__B2 _1335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4206_ _0336_ _1266_ _0293_ VGND VGND VPWR VPWR _1274_ sky130_fd_sc_hd__a21o_1
X_5186_ _1647_ _2109_ VGND VGND VPWR VPWR _2110_ sky130_fd_sc_hd__and2_1
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4137_ _0950_ _1204_ _0773_ VGND VGND VPWR VPWR _1207_ sky130_fd_sc_hd__nand3_1
XFILLER_0_78_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4068_ _0570_ _0664_ VGND VGND VPWR VPWR _1142_ sky130_fd_sc_hd__nor2_1
X_3019_ ih.t.timer_max\[16\] ih.t.timer_max\[17\] _2756_ VGND VGND VPWR VPWR _2757_
+ sky130_fd_sc_hd__or3_1
XFILLER_0_78_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_395 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5878__A1 ih.t.timer_max\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4866__A _0373_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout183 net196 VGND VGND VPWR VPWR net183 sky130_fd_sc_hd__clkbuf_4
Xfanout172 net173 VGND VGND VPWR VPWR net172 sky130_fd_sc_hd__buf_4
Xfanout161 net162 VGND VGND VPWR VPWR net161 sky130_fd_sc_hd__buf_4
Xfanout194 net195 VGND VGND VPWR VPWR net194 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_44_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_69_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1141 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1130 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3813__B1 _0741_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1174 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1163 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1152 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4369__B2 cu.reg_file.reg_e\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4369__A1 cu.pc.pc_o\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5318__A0 _1188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5869__A1 ih.t.timer_max\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output99_A net99 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3370_ _2949_ _0445_ _0440_ VGND VGND VPWR VPWR _0446_ sky130_fd_sc_hd__a21bo_1
XANTENNA__4541__A1 cu.reg_file.reg_sp\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_925 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_914 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_903 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_85_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_958 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_947 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_936 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5371__S _2226_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5040_ _1189_ _1213_ _2002_ VGND VGND VPWR VPWR _2014_ sky130_fd_sc_hd__mux2_1
XANTENNA__4495__B _1545_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_969 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_18_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5942_ cu.id.cb_opcode_y\[0\] _2410_ _2666_ VGND VGND VPWR VPWR _2680_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5873_ _2165_ ih.t.timer_max\[14\] _2636_ VGND VGND VPWR VPWR _2643_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_75_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4824_ cu.pc.pc_o\[1\] _1824_ _1815_ VGND VGND VPWR VPWR _1825_ sky130_fd_sc_hd__mux2_1
XANTENNA__4016__A _1073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_351 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4755_ _1756_ _1763_ VGND VGND VPWR VPWR _1764_ sky130_fd_sc_hd__nand2_1
XFILLER_0_28_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3706_ _0545_ _0600_ VGND VGND VPWR VPWR _0782_ sky130_fd_sc_hd__nand2_1
XFILLER_0_7_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4686_ _1708_ _1709_ _1672_ VGND VGND VPWR VPWR _1710_ sky130_fd_sc_hd__and3b_1
XFILLER_0_31_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3637_ _0575_ net142 VGND VGND VPWR VPWR _0713_ sky130_fd_sc_hd__or2_1
XFILLER_0_11_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3335__A2 _2878_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3568_ _0632_ _0643_ VGND VGND VPWR VPWR _0644_ sky130_fd_sc_hd__xnor2_2
X_5307_ _1329_ _1354_ VGND VGND VPWR VPWR _2191_ sky130_fd_sc_hd__nand2_2
XFILLER_0_11_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5281__S _2170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6287_ clknet_leaf_41_clk _0269_ net151 VGND VGND VPWR VPWR cu.id.opcode\[0\] sky130_fd_sc_hd__dfrtp_4
X_3499_ _0416_ _0420_ _0441_ _0446_ VGND VGND VPWR VPWR _0575_ sky130_fd_sc_hd__o31ai_2
X_5238_ _2145_ VGND VGND VPWR VPWR _2146_ sky130_fd_sc_hd__clkbuf_4
X_5169_ _2098_ VGND VGND VPWR VPWR _0088_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4048__B1 _0916_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5796__A0 _1110_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5310__A _2193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3574__A2 _0640_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4523__A1 cu.reg_file.reg_h\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4523__B2 cu.reg_file.reg_b\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xhold6 _0268_ VGND VGND VPWR VPWR net202 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA_output137_A net137 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_84_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_37_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xclkbuf_leaf_10_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_10_clk sky130_fd_sc_hd__clkbuf_16
X_4540_ cu.pc.pc_o\[14\] _1485_ _1593_ VGND VGND VPWR VPWR _1594_ sky130_fd_sc_hd__o21a_1
XFILLER_0_4_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_13_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3565__A2 _0640_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4471_ cu.reg_file.reg_h\[2\] _1317_ _1312_ cu.reg_file.reg_b\[2\] _1528_ VGND VGND
+ VPWR VPWR _1529_ sky130_fd_sc_hd__a221o_1
XFILLER_0_13_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_20_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_96_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_96_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6201__D net14 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6210_ clknet_leaf_4_clk net8 net171 VGND VGND VPWR VPWR ih.ih.ih.prev_data\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_0_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3422_ _0468_ _0473_ net237 _0486_ _0483_ VGND VGND VPWR VPWR _0498_ sky130_fd_sc_hd__o2111a_2
Xmax_cap147 net148 VGND VGND VPWR VPWR net147 sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_0_40_357 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6141_ clknet_leaf_23_clk _0175_ net192 VGND VGND VPWR VPWR net133 sky130_fd_sc_hd__dfrtp_4
XTAP_700 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_733 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3353_ _0428_ VGND VGND VPWR VPWR _0429_ sky130_fd_sc_hd__clkbuf_4
X_6072_ clknet_leaf_13_clk _0106_ net181 VGND VGND VPWR VPWR ih.gpio_interrupt_mask\[5\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_777 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3284_ _0340_ VGND VGND VPWR VPWR _0360_ sky130_fd_sc_hd__inv_2
XTAP_799 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5023_ _1790_ _0352_ _1791_ _0366_ VGND VGND VPWR VPWR _2001_ sky130_fd_sc_hd__and4b_1
XANTENNA__4953__B cu.pc.pc_o\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5925_ _2671_ VGND VGND VPWR VPWR _0271_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5856_ _1263_ _2632_ _2115_ VGND VGND VPWR VPWR _2633_ sky130_fd_sc_hd__mux2_1
X_4807_ _1808_ VGND VGND VPWR VPWR _1809_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_8_543 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2999_ net70 net29 ih.gpio_interrupt_mask\[2\] VGND VGND VPWR VPWR _2737_ sky130_fd_sc_hd__and3b_1
X_5787_ _2571_ _2572_ VGND VGND VPWR VPWR _2573_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_71_471 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5950__A0 _1233_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4738_ _0456_ _1746_ _2950_ VGND VGND VPWR VPWR _1747_ sky130_fd_sc_hd__o21ai_2
X_4669_ _1698_ VGND VGND VPWR VPWR ih.t.next_count\[11\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4863__B cu.pc.pc_o\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5678__C _1661_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_1_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_89_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4680__B1 _1687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3971_ _0600_ _1044_ _1042_ _0610_ _1045_ VGND VGND VPWR VPWR _1046_ sky130_fd_sc_hd__o221ai_1
X_5710_ _2708_ _1653_ VGND VGND VPWR VPWR _2514_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5641_ net82 _1633_ _2451_ _2454_ VGND VGND VPWR VPWR _2455_ sky130_fd_sc_hd__o22a_1
XFILLER_0_45_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5096__S _2039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_279 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5572_ _1649_ _2389_ VGND VGND VPWR VPWR _2390_ sky130_fd_sc_hd__and2_1
X_4523_ cu.reg_file.reg_h\[5\] _1316_ _1312_ cu.reg_file.reg_b\[5\] _1577_ VGND VGND
+ VPWR VPWR _1578_ sky130_fd_sc_hd__a221o_1
XFILLER_0_13_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4454_ _1332_ _1511_ VGND VGND VPWR VPWR _1513_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3405_ net148 _0476_ _0478_ _0382_ _0465_ VGND VGND VPWR VPWR _0481_ sky130_fd_sc_hd__a2111oi_1
X_4385_ cu.reg_file.reg_e\[6\] _1283_ _1285_ cu.reg_file.reg_l\[6\] _1446_ VGND VGND
+ VPWR VPWR _1447_ sky130_fd_sc_hd__a221o_1
X_6124_ clknet_leaf_20_clk _0158_ net189 VGND VGND VPWR VPWR net116 sky130_fd_sc_hd__dfrtp_1
X_3336_ _0410_ _0411_ cu.id.starting_int_service VGND VGND VPWR VPWR _0412_ sky130_fd_sc_hd__a21o_2
XTAP_530 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6055_ clknet_leaf_23_clk _0093_ net192 VGND VGND VPWR VPWR mc.cl.next_data\[13\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__4964__A cu.pc.pc_o\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_563 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3267_ cu.id.cb_opcode_z\[0\] VGND VGND VPWR VPWR _0343_ sky130_fd_sc_hd__buf_4
XTAP_596 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5006_ cu.reg_file.reg_a\[2\] _1989_ _1985_ VGND VGND VPWR VPWR _1990_ sky130_fd_sc_hd__mux2_1
XANTENNA__4671__B1 _1687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3198_ _2888_ _2890_ _2933_ _2934_ VGND VGND VPWR VPWR _2935_ sky130_fd_sc_hd__nand4_4
XFILLER_0_95_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3299__B _0374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5908_ _2661_ VGND VGND VPWR VPWR _0264_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3777__A2 _0640_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5839_ cu.reg_file.reg_sp\[13\] _2536_ VGND VGND VPWR VPWR _2618_ sky130_fd_sc_hd__or2_1
XFILLER_0_36_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_151 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_31_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_16_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5151__A1 _2085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4662__B1 _1687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4114__A _1089_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5390__A1 net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output81_A net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5142__A1 cu.reg_file.reg_h\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5693__A2 _1650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4170_ _0850_ _0861_ _1060_ VGND VGND VPWR VPWR _1240_ sky130_fd_sc_hd__mux2_1
X_3121_ _2789_ _2791_ _2792_ _2858_ VGND VGND VPWR VPWR _2859_ sky130_fd_sc_hd__or4_1
XANTENNA__4653__B1 _1687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3052_ ih.t.timer_max\[21\] _2759_ VGND VGND VPWR VPWR _2790_ sky130_fd_sc_hd__nand2_1
XFILLER_0_26_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_89_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_89_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_89_198 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_77_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4956__A1 cu.pc.pc_o\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3954_ _0712_ _0713_ VGND VGND VPWR VPWR _1029_ sky130_fd_sc_hd__xor2_1
XANTENNA__3759__A2 _0743_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4420__A3 _1473_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_73_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3885_ _0914_ _0960_ _0773_ _0777_ VGND VGND VPWR VPWR _0961_ sky130_fd_sc_hd__o2bb2a_1
X_5624_ _1400_ _2438_ VGND VGND VPWR VPWR _2439_ sky130_fd_sc_hd__and2b_1
XFILLER_0_5_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_268 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_60_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5381__A1 net123 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5555_ _2373_ VGND VGND VPWR VPWR _0199_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5554__S _2351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4506_ _1333_ _1561_ VGND VGND VPWR VPWR _1562_ sky130_fd_sc_hd__xnor2_1
X_5486_ net67 _0618_ _2306_ VGND VGND VPWR VPWR _2307_ sky130_fd_sc_hd__mux2_1
X_4437_ _1396_ _1496_ VGND VGND VPWR VPWR _1497_ sky130_fd_sc_hd__xnor2_1
XANTENNA__5133__A1 cu.reg_file.reg_h\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6107_ clknet_leaf_26_clk _0141_ net195 VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__dfrtp_2
XTAP_360 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4368_ cu.reg_file.reg_sp\[5\] _0993_ _1344_ _0373_ _1364_ VGND VGND VPWR VPWR _1431_
+ sky130_fd_sc_hd__a221o_1
X_4299_ cu.reg_file.reg_sp\[2\] _0993_ _1344_ _0341_ _1364_ VGND VGND VPWR VPWR _1365_
+ sky130_fd_sc_hd__a221o_1
X_3319_ _0394_ VGND VGND VPWR VPWR _0395_ sky130_fd_sc_hd__buf_2
XTAP_371 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6038_ clknet_leaf_33_clk _0076_ net161 VGND VGND VPWR VPWR cu.reg_file.reg_h\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_68_316 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_555 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_32_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5124__A1 cu.reg_file.reg_h\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3570__C_N _0373_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_27_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_352 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3670_ cu.reg_file.reg_a\[0\] _0625_ _0628_ cu.reg_file.reg_mem\[8\] _0745_ VGND
+ VGND VPWR VPWR _0746_ sky130_fd_sc_hd__a221o_1
XFILLER_0_88_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput116 net116 VGND VGND VPWR VPWR ss5[0] sky130_fd_sc_hd__buf_2
XFILLER_0_88_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5340_ _2211_ VGND VGND VPWR VPWR _0146_ sky130_fd_sc_hd__clkbuf_1
Xoutput105 net105 VGND VGND VPWR VPWR ss3[5] sky130_fd_sc_hd__buf_2
Xoutput138 net138 VGND VGND VPWR VPWR ss7[6] sky130_fd_sc_hd__clkbuf_4
X_5271_ net76 _2085_ _2170_ VGND VGND VPWR VPWR _2171_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput127 net127 VGND VGND VPWR VPWR ss6[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_368 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5115__A1 _1193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4222_ cu.reg_file.reg_c\[0\] _1281_ _1289_ VGND VGND VPWR VPWR _1290_ sky130_fd_sc_hd__a21oi_1
XANTENNA__4874__A0 cu.pc.pc_o\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4153_ _0816_ _0936_ _0776_ VGND VGND VPWR VPWR _1223_ sky130_fd_sc_hd__a21oi_1
X_3104_ _2837_ _2838_ _2840_ _2841_ VGND VGND VPWR VPWR _2842_ sky130_fd_sc_hd__or4_1
X_4084_ _1045_ _0681_ _1155_ _1157_ _0531_ VGND VGND VPWR VPWR _1158_ sky130_fd_sc_hd__a32o_1
XANTENNA__3429__A1 cu.pc.pc_o\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3035_ ih.t.count\[28\] _2772_ VGND VGND VPWR VPWR _2773_ sky130_fd_sc_hd__xnor2_1
XANTENNA__3429__B2 cu.reg_file.reg_b\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_61 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4929__A1 cu.pc.pc_o\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4986_ cu.pc.pc_o\[14\] _1973_ _1814_ VGND VGND VPWR VPWR _1974_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_149 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3937_ _0372_ _2921_ _1012_ VGND VGND VPWR VPWR _1013_ sky130_fd_sc_hd__and3_1
XFILLER_0_73_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3601__A1 cu.reg_file.reg_b\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3601__B2 cu.reg_file.reg_mem\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_33_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3868_ _0844_ _0929_ VGND VGND VPWR VPWR _0944_ sky130_fd_sc_hd__xnor2_1
X_5607_ mc.cl.next_data\[4\] _2313_ net141 _2422_ VGND VGND VPWR VPWR _2423_ sky130_fd_sc_hd__a22o_1
XANTENNA__5354__A1 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3799_ _0871_ _0874_ VGND VGND VPWR VPWR _0875_ sky130_fd_sc_hd__and2b_1
XANTENNA__4379__B1_N _1434_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5538_ net109 _2147_ _2225_ net117 _2356_ VGND VGND VPWR VPWR _2357_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5657__A2 _2193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5469_ _2293_ _2284_ VGND VGND VPWR VPWR _2294_ sky130_fd_sc_hd__nor2_1
XANTENNA__3668__B2 cu.reg_file.reg_sp\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3668__A1 cu.reg_file.reg_b\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4590__C _1633_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3918__D _0993_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_566 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput18 memory_data_in[0] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_2
XANTENNA__5345__A1 net107 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xinput29 programmable_gpio_in[2] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_2
XANTENNA__3008__A ih.t.timer_max\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5922__S _2668_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output44_A net44 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5281__A0 net81 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_87_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5369__S _2226_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4840_ cu.pc.pc_o\[3\] _1826_ VGND VGND VPWR VPWR _1839_ sky130_fd_sc_hd__nor2_1
XFILLER_0_28_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__6204__D net17 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4771_ _1268_ _1012_ _1646_ _1301_ VGND VGND VPWR VPWR _1778_ sky130_fd_sc_hd__or4b_1
XFILLER_0_7_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3722_ _0796_ _0797_ VGND VGND VPWR VPWR _0798_ sky130_fd_sc_hd__and2_1
XFILLER_0_82_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3653_ _0576_ _0723_ _0725_ _0728_ VGND VGND VPWR VPWR _0729_ sky130_fd_sc_hd__o2bb2a_2
XFILLER_0_43_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5323_ _2201_ VGND VGND VPWR VPWR _0139_ sky130_fd_sc_hd__clkbuf_1
X_3584_ cu.reg_file.reg_e\[5\] _0489_ _0495_ cu.reg_file.reg_h\[5\] _0536_ VGND VGND
+ VPWR VPWR _0660_ sky130_fd_sc_hd__a221o_1
XFILLER_0_11_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5639__A2 _2204_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5254_ _1089_ _1222_ _1667_ VGND VGND VPWR VPWR _2159_ sky130_fd_sc_hd__mux2_1
XANTENNA__4847__A0 _1089_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5185_ mc.cl.next_data\[14\] net24 mc.count VGND VGND VPWR VPWR _2109_ sky130_fd_sc_hd__mux2_1
XANTENNA__4311__A2 _1348_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_72 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4205_ _0359_ _2937_ VGND VGND VPWR VPWR _1273_ sky130_fd_sc_hd__or2_1
X_4136_ _0918_ _1205_ VGND VGND VPWR VPWR _1206_ sky130_fd_sc_hd__and2_1
XFILLER_0_78_411 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4067_ _0558_ _0632_ _0663_ _1139_ _1140_ VGND VGND VPWR VPWR _1141_ sky130_fd_sc_hd__a221o_1
X_3018_ ih.t.timer_max\[15\] _2755_ VGND VGND VPWR VPWR _2756_ sky130_fd_sc_hd__or2_2
XFILLER_0_78_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5279__S _2170_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3588__A _0652_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4969_ _1956_ _1957_ VGND VGND VPWR VPWR _1958_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5308__A _1374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4866__B cu.pc.pc_o\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout173 net182 VGND VGND VPWR VPWR net173 sky130_fd_sc_hd__clkbuf_2
Xfanout162 net163 VGND VGND VPWR VPWR net162 sky130_fd_sc_hd__buf_2
XANTENNA__3510__B1 _0576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout151 net152 VGND VGND VPWR VPWR net151 sky130_fd_sc_hd__clkbuf_4
Xfanout195 net196 VGND VGND VPWR VPWR net195 sky130_fd_sc_hd__buf_4
Xfanout184 net185 VGND VGND VPWR VPWR net184 sky130_fd_sc_hd__clkbuf_4
XANTENNA__5263__A0 _1126_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3813__A1 cu.reg_file.reg_d\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1131 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1120 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3813__B2 cu.reg_file.reg_h\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1164 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1153 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1142 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5015__A0 cu.reg_file.reg_a\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1175 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5566__A1 _1666_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_60_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_71_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5318__A1 net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3329__B1 cu.id.starting_int_service VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_926 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_915 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_904 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_959 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_948 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_937 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_23_clk_A clknet_2_3__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5254__A0 _1089_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4792__A _1793_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_38_clk_A clknet_2_1__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5941_ _2679_ VGND VGND VPWR VPWR _0279_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5099__S _2039_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_34_63 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5872_ _2642_ VGND VGND VPWR VPWR _0247_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5006__A0 cu.reg_file.reg_a\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5557__A1 net94 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4823_ _1817_ _1823_ _1809_ VGND VGND VPWR VPWR _1824_ sky130_fd_sc_hd__mux2_1
XANTENNA__4016__B _1089_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4754_ _2904_ _2924_ _1318_ _1762_ _0350_ VGND VGND VPWR VPWR _1763_ sky130_fd_sc_hd__a41o_1
XFILLER_0_28_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3705_ _0447_ net142 VGND VGND VPWR VPWR _0781_ sky130_fd_sc_hd__nand2_1
X_4685_ ih.t.count\[15\] ih.t.count\[16\] _1702_ ih.t.count\[17\] VGND VGND VPWR VPWR
+ _1709_ sky130_fd_sc_hd__a31o_1
XFILLER_0_70_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3636_ _0545_ _0598_ VGND VGND VPWR VPWR _0712_ sky130_fd_sc_hd__xnor2_4
X_3567_ _0576_ _0635_ _0638_ _0642_ VGND VGND VPWR VPWR _0643_ sky130_fd_sc_hd__o2bb2a_2
X_5306_ _2190_ VGND VGND VPWR VPWR _0133_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6286_ clknet_leaf_36_clk net202 net158 VGND VGND VPWR VPWR cu.id.can_be_interrupted
+ sky130_fd_sc_hd__dfrtp_1
X_5237_ _1369_ _1625_ VGND VGND VPWR VPWR _2145_ sky130_fd_sc_hd__nor2_1
XFILLER_0_11_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3498_ net142 VGND VGND VPWR VPWR _0574_ sky130_fd_sc_hd__inv_2
XANTENNA__4296__B2 cu.pc.pc_o\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4296__A1 _0341_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5168_ _1647_ _2097_ VGND VGND VPWR VPWR _2098_ sky130_fd_sc_hd__and2_1
X_5099_ cu.reg_file.reg_d\[7\] _2053_ _2039_ VGND VGND VPWR VPWR _2054_ sky130_fd_sc_hd__mux2_1
XANTENNA__4048__A1 _1032_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4119_ net209 _1186_ _0370_ _1190_ VGND VGND VPWR VPWR _0011_ sky130_fd_sc_hd__a22o_1
XFILLER_0_66_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_108 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4220__A1 cu.reg_file.reg_a\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4220__B2 cu.reg_file.reg_sp\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_528 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4877__A cu.pc.pc_o\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xhold7 ih.interrupt_source\[1\] VGND VGND VPWR VPWR net203 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5236__A0 _0617_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3005__B net34 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4117__A _1160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4470_ _1521_ _1321_ _1314_ cu.reg_file.reg_d\[2\] _1527_ VGND VGND VPWR VPWR _1528_
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_20_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_40_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4787__A _0343_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmax_cap148 _0335_ VGND VGND VPWR VPWR net148 sky130_fd_sc_hd__clkbuf_2
X_3421_ cu.reg_file.reg_d\[0\] _0492_ _0494_ cu.reg_file.reg_mem\[0\] _0496_ VGND
+ VGND VPWR VPWR _0497_ sky130_fd_sc_hd__a221o_1
XFILLER_0_40_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6140_ clknet_leaf_24_clk _0174_ net195 VGND VGND VPWR VPWR net132 sky130_fd_sc_hd__dfrtp_2
XTAP_701 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3352_ _0412_ _0405_ _0409_ _0407_ VGND VGND VPWR VPWR _0428_ sky130_fd_sc_hd__and4b_1
XFILLER_0_21_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_734 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6071_ clknet_leaf_17_clk _0105_ net172 VGND VGND VPWR VPWR ih.gpio_interrupt_mask\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_767 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4278__A1 cu.reg_file.reg_sp\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4278__B2 _0340_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3283_ _2902_ VGND VGND VPWR VPWR _0359_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_29_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_29_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_789 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5022_ _2000_ VGND VGND VPWR VPWR _0039_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_45_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_48_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4450__A1 cu.pc.pc_o\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5924_ _2899_ _2391_ _2668_ VGND VGND VPWR VPWR _2671_ sky130_fd_sc_hd__mux2_1
XANTENNA__4450__B2 cu.reg_file.reg_d\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5855_ cu.reg_file.reg_sp\[15\] _2631_ VGND VGND VPWR VPWR _2632_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_90_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_555 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4806_ _2935_ _1256_ _1807_ VGND VGND VPWR VPWR _1808_ sky130_fd_sc_hd__o21ai_4
X_2998_ _2734_ net28 ih.gpio_interrupt_mask\[1\] _2735_ VGND VGND VPWR VPWR _2736_
+ sky130_fd_sc_hd__a31o_1
X_5786_ _2562_ _2565_ _2563_ VGND VGND VPWR VPWR _2572_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_9_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5950__A1 _2486_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4737_ _0302_ _1266_ _1745_ VGND VGND VPWR VPWR _1746_ sky130_fd_sc_hd__nor3b_1
X_4668_ _1696_ _1697_ _1672_ VGND VGND VPWR VPWR _1698_ sky130_fd_sc_hd__and3b_1
XFILLER_0_71_483 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3961__B1 _0773_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3619_ _0294_ _0692_ _0634_ VGND VGND VPWR VPWR _0695_ sky130_fd_sc_hd__or3_1
XANTENNA__5702__B2 ih.t.timer_max\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4599_ _1634_ _1636_ _1641_ _1642_ VGND VGND VPWR VPWR _1643_ sky130_fd_sc_hd__nand4_4
XANTENNA__4269__A1 _1330_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6269_ clknet_leaf_9_clk _0251_ net174 VGND VGND VPWR VPWR ih.t.timer_max\[1\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__5466__A0 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_94_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_81_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3952__B1 _1027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5930__S _2668_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3016__A ih.t.timer_max\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4432__A1 cu.pc.pc_o\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3970_ _0603_ _0606_ VGND VGND VPWR VPWR _1045_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5377__S _2226_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5640_ net114 _2147_ _2225_ net122 _2453_ VGND VGND VPWR VPWR _2454_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5571_ net10 _2345_ _2369_ net3 VGND VGND VPWR VPWR _2389_ sky130_fd_sc_hd__a22o_1
XFILLER_0_60_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5932__A1 _2467_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_483 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4522_ cu.pc.pc_o\[13\] _1321_ _1314_ cu.reg_file.reg_d\[5\] _1576_ VGND VGND VPWR
+ VPWR _1577_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4453_ _1332_ _1511_ VGND VGND VPWR VPWR _1512_ sky130_fd_sc_hd__or2_1
XFILLER_0_40_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5696__B1 cu.reg_file.reg_mem\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4499__A1 cu.id.imm_i\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4499__B2 cu.pc.pc_o\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_13_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3404_ net146 _0473_ _0479_ VGND VGND VPWR VPWR _0480_ sky130_fd_sc_hd__nor3_2
XFILLER_0_40_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4384_ cu.reg_file.reg_a\[6\] _1276_ _1287_ cu.reg_file.reg_sp\[6\] VGND VGND VPWR
+ VPWR _1446_ sky130_fd_sc_hd__a22o_1
X_6123_ clknet_leaf_13_clk _0157_ net174 VGND VGND VPWR VPWR net115 sky130_fd_sc_hd__dfrtp_2
XANTENNA__5448__A0 net73 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3335_ _2900_ _2878_ _2877_ VGND VGND VPWR VPWR _0411_ sky130_fd_sc_hd__a21o_1
XTAP_520 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6054_ clknet_leaf_20_clk _0092_ net189 VGND VGND VPWR VPWR mc.cl.next_data\[12\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_56_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3266_ _2885_ _2927_ _2917_ VGND VGND VPWR VPWR _0342_ sky130_fd_sc_hd__and3_1
XTAP_553 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5005_ _1074_ _1226_ _0368_ VGND VGND VPWR VPWR _1989_ sky130_fd_sc_hd__mux2_1
XTAP_586 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_fanout180_A net182 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3197_ cu.id.alu_opcode\[0\] cu.id.opcode\[0\] VGND VGND VPWR VPWR _2934_ sky130_fd_sc_hd__nor2_2
XFILLER_0_88_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5907_ ih.t.timer_max\[22\] _1193_ _2654_ VGND VGND VPWR VPWR _2661_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5620__B1 _2225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3631__C1 _0536_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5838_ _2617_ VGND VGND VPWR VPWR _0238_ sky130_fd_sc_hd__clkbuf_1
X_5769_ _2555_ _2556_ VGND VGND VPWR VPWR _2557_ sky130_fd_sc_hd__nor2_1
XFILLER_0_16_163 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_71_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_122 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_31_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4890__A _2920_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_82_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5914__A1 _2351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_42_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_62_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output74_A net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3120_ _2794_ _2795_ _2857_ VGND VGND VPWR VPWR _2858_ sky130_fd_sc_hd__or3_1
XFILLER_0_93_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3051_ ih.t.count\[22\] _2788_ VGND VGND VPWR VPWR _2789_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_89_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5850__A0 _1624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6207__D net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5602__B1 _2204_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__4956__A2 _1521_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3953_ _0370_ _0619_ _1026_ _1028_ VGND VGND VPWR VPWR _0007_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_45_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3884_ _0948_ _0959_ VGND VGND VPWR VPWR _0960_ sky130_fd_sc_hd__nand2_1
XANTENNA__5905__A1 _1191_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5623_ ih.t.timer_max\[13\] _2193_ _2314_ ih.t.timer_max\[5\] _2437_ VGND VGND VPWR
+ VPWR _2438_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5554_ cu.reg_file.reg_mem\[1\] _2372_ _2351_ VGND VGND VPWR VPWR _2373_ sky130_fd_sc_hd__mux2_1
XFILLER_0_41_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5485_ _2305_ _2284_ VGND VGND VPWR VPWR _2306_ sky130_fd_sc_hd__nor2_1
X_4505_ _1305_ _1557_ _1560_ VGND VGND VPWR VPWR _1561_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_5_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_453 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4436_ _1305_ _1492_ _1495_ VGND VGND VPWR VPWR _1496_ sky130_fd_sc_hd__o21a_2
XFILLER_0_6_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4367_ cu.reg_file.reg_l\[5\] _1317_ VGND VGND VPWR VPWR _1430_ sky130_fd_sc_hd__and2_1
XANTENNA__4975__A cu.pc.pc_o\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6106_ clknet_leaf_27_clk _0140_ net186 VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__dfrtp_4
X_3318_ _0377_ _0393_ VGND VGND VPWR VPWR _0394_ sky130_fd_sc_hd__or2_1
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_350 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4298_ _1324_ VGND VGND VPWR VPWR _1364_ sky130_fd_sc_hd__clkbuf_8
XTAP_361 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6037_ clknet_leaf_28_clk _0075_ net188 VGND VGND VPWR VPWR cu.reg_file.reg_h\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_3249_ cu.id.alu_opcode\[1\] cu.id.alu_opcode\[3\] VGND VGND VPWR VPWR _0325_ sky130_fd_sc_hd__or2_1
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_34 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_56 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_95_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_545 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_64_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4215__A _1282_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_397 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4580__B1 _1263_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_19 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3013__B ih.t.timer_max\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_328 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output112_A net112 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_74_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5060__A1 _1074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3071__B1 ih.t.timer_max\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_27_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_27_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_70_537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_88_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput106 net106 VGND VGND VPWR VPWR ss3[6] sky130_fd_sc_hd__buf_2
XANTENNA__4571__B1 _1622_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput117 net117 VGND VGND VPWR VPWR ss5[1] sky130_fd_sc_hd__clkbuf_4
X_5270_ _2169_ _2140_ VGND VGND VPWR VPWR _2170_ sky130_fd_sc_hd__nor2_4
Xoutput139 net139 VGND VGND VPWR VPWR ss7[7] sky130_fd_sc_hd__buf_2
Xoutput128 net128 VGND VGND VPWR VPWR ss6[4] sky130_fd_sc_hd__clkbuf_4
X_4221_ cu.reg_file.reg_e\[0\] _1283_ _1285_ cu.reg_file.reg_l\[0\] _1288_ VGND VGND
+ VPWR VPWR _1289_ sky130_fd_sc_hd__a221o_1
XANTENNA__5390__S _2237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4152_ _1217_ _1221_ _0824_ VGND VGND VPWR VPWR _1222_ sky130_fd_sc_hd__o21a_4
X_3103_ _2746_ _2839_ ih.t.count\[2\] VGND VGND VPWR VPWR _2841_ sky130_fd_sc_hd__a21oi_1
X_4083_ _0606_ _0671_ _0681_ _1156_ VGND VGND VPWR VPWR _1157_ sky130_fd_sc_hd__a211oi_1
XANTENNA__3429__A2 _0501_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3034_ ih.t.timer_max\[28\] _2764_ VGND VGND VPWR VPWR _2772_ sky130_fd_sc_hd__xor2_1
XFILLER_0_77_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4929__A2 cu.pc.pc_o\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4985_ _1965_ _1972_ _1808_ VGND VGND VPWR VPWR _1973_ sky130_fd_sc_hd__mux2_1
X_3936_ _0296_ _2918_ VGND VGND VPWR VPWR _1012_ sky130_fd_sc_hd__nor2_2
XFILLER_0_46_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3601__A2 _0502_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3867_ _0856_ _0927_ VGND VGND VPWR VPWR _0943_ sky130_fd_sc_hd__xnor2_2
X_5606_ _1666_ _2420_ _2421_ VGND VGND VPWR VPWR _2422_ sky130_fd_sc_hd__o21a_1
XFILLER_0_5_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3798_ cu.reg_file.reg_mem\[11\] _0640_ _0872_ _0873_ VGND VGND VPWR VPWR _0874_
+ sky130_fd_sc_hd__a211oi_2
X_5537_ net101 _2205_ _2355_ _1401_ VGND VGND VPWR VPWR _2356_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5468_ _2205_ VGND VGND VPWR VPWR _2293_ sky130_fd_sc_hd__inv_2
XFILLER_0_1_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4419_ _1382_ _1475_ _1476_ _1479_ VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__a31o_1
X_5399_ _2244_ VGND VGND VPWR VPWR _0172_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3668__A2 _0743_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput19 memory_data_in[1] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_52_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_52_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_24_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4553__B1 _1286_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3008__B ih.t.timer_max\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5805__A0 cu.reg_file.reg_sp\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output37_A net37 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5281__A1 _1191_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_87_456 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_74_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_523 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_342 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4770_ _1300_ _1761_ _1776_ VGND VGND VPWR VPWR _1777_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_23_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_386 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3595__B2 _0670_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3721_ _0752_ _0789_ _0792_ _0795_ VGND VGND VPWR VPWR _0797_ sky130_fd_sc_hd__nand4_1
X_3652_ cu.reg_file.reg_l\[7\] _0422_ _0726_ _0727_ _0440_ VGND VGND VPWR VPWR _0728_
+ sky130_fd_sc_hd__a2111o_1
XFILLER_0_43_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3583_ cu.reg_file.reg_sp\[5\] _0539_ _0494_ cu.reg_file.reg_mem\[5\] _0658_ VGND
+ VGND VPWR VPWR _0659_ sky130_fd_sc_hd__a221o_1
X_5322_ _1192_ net97 _2195_ VGND VGND VPWR VPWR _2201_ sky130_fd_sc_hd__mux2_1
XFILLER_0_11_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5253_ _2158_ VGND VGND VPWR VPWR _0112_ sky130_fd_sc_hd__clkbuf_1
X_5184_ _2108_ VGND VGND VPWR VPWR _0093_ sky130_fd_sc_hd__clkbuf_1
X_4204_ _0469_ VGND VGND VPWR VPWR _1272_ sky130_fd_sc_hd__inv_2
X_4135_ _1204_ _0779_ VGND VGND VPWR VPWR _1205_ sky130_fd_sc_hd__or2_1
XANTENNA__4075__A2 _0773_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4066_ _0531_ _0663_ _0681_ _0822_ VGND VGND VPWR VPWR _1140_ sky130_fd_sc_hd__a2bb2o_1
X_3017_ ih.t.timer_max\[13\] ih.t.timer_max\[14\] _2754_ VGND VGND VPWR VPWR _2755_
+ sky130_fd_sc_hd__or3_1
XANTENNA__3588__B _0663_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_117 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4968_ _1943_ _1948_ VGND VGND VPWR VPWR _1957_ sky130_fd_sc_hd__and2b_1
XFILLER_0_73_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5295__S _2182_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4899_ _1893_ VGND VGND VPWR VPWR _0023_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_375 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3919_ _0986_ _0989_ _0994_ VGND VGND VPWR VPWR _0995_ sky130_fd_sc_hd__nand3b_1
XFILLER_0_34_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_548 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_14_294 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4299__C1 _1364_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout174 net175 VGND VGND VPWR VPWR net174 sky130_fd_sc_hd__clkbuf_4
Xfanout163 net26 VGND VGND VPWR VPWR net163 sky130_fd_sc_hd__buf_2
Xfanout152 net163 VGND VGND VPWR VPWR net152 sky130_fd_sc_hd__clkbuf_2
Xfanout196 net26 VGND VGND VPWR VPWR net196 sky130_fd_sc_hd__buf_2
Xfanout185 net196 VGND VGND VPWR VPWR net185 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5263__A1 _1624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1132 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1121 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1110 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3813__A2 _0488_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_286 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1165 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1154 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1143 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1176 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_64_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_52_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_916 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_905 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_20_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_949 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_938 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_927 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5254__A1 _1222_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5940_ _0341_ _2391_ _2666_ VGND VGND VPWR VPWR _2679_ sky130_fd_sc_hd__mux2_1
XANTENNA__3804__A2 _0740_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5871_ _2163_ ih.t.timer_max\[13\] _2636_ VGND VGND VPWR VPWR _2642_ sky130_fd_sc_hd__mux2_1
XANTENNA__5557__A2 _2194_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4822_ _1821_ _1822_ _1799_ VGND VGND VPWR VPWR _1823_ sky130_fd_sc_hd__mux2_1
XFILLER_0_50_41 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4753_ net149 _2952_ _0307_ VGND VGND VPWR VPWR _1762_ sky130_fd_sc_hd__and3b_1
XFILLER_0_7_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_50_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_269 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3704_ _0768_ _0770_ _0753_ _0779_ VGND VGND VPWR VPWR _0780_ sky130_fd_sc_hd__nor4_1
XFILLER_0_43_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4684_ ih.t.count\[16\] ih.t.count\[17\] _1705_ VGND VGND VPWR VPWR _1708_ sky130_fd_sc_hd__and3_1
XANTENNA__4517__B1 _1284_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_453 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3635_ _0587_ _0710_ VGND VGND VPWR VPWR _0711_ sky130_fd_sc_hd__nand2_1
XFILLER_0_31_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3566_ cu.reg_file.reg_l\[6\] _0422_ _0639_ _0641_ _0576_ VGND VGND VPWR VPWR _0642_
+ sky130_fd_sc_hd__a2111o_1
X_5305_ _1261_ net91 _2182_ VGND VGND VPWR VPWR _2190_ sky130_fd_sc_hd__mux2_1
X_3497_ _0514_ _0529_ VGND VGND VPWR VPWR _0573_ sky130_fd_sc_hd__or2_1
X_6285_ clknet_leaf_37_clk _0267_ net160 VGND VGND VPWR VPWR cu.ir.idx\[1\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__4686__C _1672_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5236_ _0617_ _1622_ _1667_ VGND VGND VPWR VPWR _2144_ sky130_fd_sc_hd__mux2_1
XFILLER_0_52_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5167_ mc.cl.next_data\[8\] net18 mc.count VGND VGND VPWR VPWR _2097_ sky130_fd_sc_hd__mux2_1
XANTENNA__5245__A1 _1667_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4118_ _1189_ VGND VGND VPWR VPWR _1190_ sky130_fd_sc_hd__buf_4
X_5098_ _1110_ _1263_ _2035_ VGND VGND VPWR VPWR _2053_ sky130_fd_sc_hd__mux2_1
X_4049_ _0802_ _1122_ _0812_ _1032_ VGND VGND VPWR VPWR _1123_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_93_289 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_356 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xhold8 ih.interrupt_source\[2\] VGND VGND VPWR VPWR net204 sky130_fd_sc_hd__dlygate4sd3_1
XFILLER_0_89_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5236__A1 _1622_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_69_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3798__A1 cu.reg_file.reg_mem\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4995__A0 cu.pc.pc_o\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_415 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5928__S _2668_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5539__A2 _1633_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_25_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4787__B _1299_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xmax_cap149 _0448_ VGND VGND VPWR VPWR net149 sky130_fd_sc_hd__buf_1
XFILLER_0_0_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3420_ cu.reg_file.reg_sp\[0\] _0480_ _0493_ _0495_ cu.reg_file.reg_h\[0\] VGND VGND
+ VPWR VPWR _0496_ sky130_fd_sc_hd__a32o_1
X_3351_ _0423_ _0424_ _0426_ VGND VGND VPWR VPWR _0427_ sky130_fd_sc_hd__a21o_2
XTAP_724 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_702 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_489 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6070_ clknet_leaf_5_clk _0104_ net172 VGND VGND VPWR VPWR ih.gpio_interrupt_mask\[3\]
+ sky130_fd_sc_hd__dfrtp_1
XTAP_768 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4278__A2 _0993_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3282_ _2915_ _0353_ _0357_ VGND VGND VPWR VPWR _0358_ sky130_fd_sc_hd__o21ba_1
XTAP_779 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5021_ cu.reg_file.reg_a\[7\] _1999_ _1985_ VGND VGND VPWR VPWR _2000_ sky130_fd_sc_hd__mux2_1
XANTENNA__4986__A0 cu.pc.pc_o\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3212__A cu.id.starting_int_service VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5923_ _2670_ VGND VGND VPWR VPWR _0270_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_512 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5854_ _1589_ _2630_ _2626_ VGND VGND VPWR VPWR _2631_ sky130_fd_sc_hd__mux2_1
XFILLER_0_63_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_84 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4805_ _0359_ _0304_ _1801_ _1804_ _1806_ VGND VGND VPWR VPWR _1807_ sky130_fd_sc_hd__o2111a_2
XANTENNA__4738__B1 _2950_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_2997_ net68 net27 ih.gpio_interrupt_mask\[0\] VGND VGND VPWR VPWR _2735_ sky130_fd_sc_hd__and3b_1
XFILLER_0_8_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_28_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5785_ _2569_ _2570_ VGND VGND VPWR VPWR _2571_ sky130_fd_sc_hd__nand2_1
X_4736_ _2897_ _2941_ _1742_ _1744_ VGND VGND VPWR VPWR _1745_ sky130_fd_sc_hd__a31o_1
X_4667_ ih.t.count\[10\] _1693_ ih.t.count\[11\] VGND VGND VPWR VPWR _1697_ sky130_fd_sc_hd__a21o_1
XFILLER_0_71_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4978__A _1233_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5163__A0 cu.reg_file.reg_l\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3618_ _0687_ _0689_ _0691_ _0693_ VGND VGND VPWR VPWR _0694_ sky130_fd_sc_hd__o31a_4
XFILLER_0_31_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4598_ _1415_ _1629_ _1637_ VGND VGND VPWR VPWR _1642_ sky130_fd_sc_hd__or3_2
XFILLER_0_12_551 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4189__S _1027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3549_ _0498_ VGND VGND VPWR VPWR _0625_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__5466__A1 _2085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6268_ clknet_leaf_9_clk _0250_ net175 VGND VGND VPWR VPWR ih.t.timer_max\[0\] sky130_fd_sc_hd__dfrtp_4
X_5219_ _1190_ ih.gpio_interrupt_mask\[4\] _2127_ VGND VGND VPWR VPWR _2132_ sky130_fd_sc_hd__mux2_1
X_6199_ clknet_leaf_5_clk net12 net169 VGND VGND VPWR VPWR ih.ih.ih.prev_data\[4\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_66_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_22_clk_A clknet_2_3__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3952__A1 alu.Cin VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4901__B1 cu.pc.pc_o\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_37_clk_A clknet_2_1__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_66_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3468__B1 _0536_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_2_3__f_clk clknet_0_clk VGND VGND VPWR VPWR clknet_2_3__leaf_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__6314__RESET_B net160 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_234 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_57_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5570_ net70 _1648_ _2137_ _2274_ VGND VGND VPWR VPWR _2388_ sky130_fd_sc_hd__a31o_1
XFILLER_0_25_131 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_462 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4521_ cu.reg_file.reg_sp\[13\] _0992_ _1343_ cu.id.imm_i\[13\] _1323_ VGND VGND
+ VPWR VPWR _1576_ sky130_fd_sc_hd__a221o_1
XFILLER_0_5_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4452_ _1505_ _1506_ _1510_ VGND VGND VPWR VPWR _1511_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_13_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_112 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5696__B2 _1646_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3403_ net148 _0476_ _0478_ _0382_ _0465_ VGND VGND VPWR VPWR _0479_ sky130_fd_sc_hd__a2111o_2
X_4383_ _1423_ _1437_ VGND VGND VPWR VPWR _1445_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6122_ clknet_leaf_7_clk _0156_ net167 VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__dfrtp_2
XANTENNA__5448__A1 net75 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3334_ _2925_ _2932_ _0364_ VGND VGND VPWR VPWR _0410_ sky130_fd_sc_hd__or3_1
XTAP_510 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_521 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6053_ clknet_leaf_22_clk _0091_ net192 VGND VGND VPWR VPWR mc.cl.next_data\[11\]
+ sky130_fd_sc_hd__dfrtp_1
X_3265_ cu.id.cb_opcode_z\[2\] VGND VGND VPWR VPWR _0341_ sky130_fd_sc_hd__buf_4
XANTENNA__3459__B1 _0502_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_554 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_56_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5004_ _1988_ VGND VGND VPWR VPWR _0033_ sky130_fd_sc_hd__clkbuf_1
XTAP_587 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3196_ _2899_ _2900_ VGND VGND VPWR VPWR _2933_ sky130_fd_sc_hd__nor2_2
XANTENNA_fanout173_A net182 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4959__B1 _1798_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5906_ _2660_ VGND VGND VPWR VPWR _0263_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5620__A1 net113 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3631__B1 _0502_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5837_ cu.reg_file.reg_sp\[12\] _2616_ _2538_ VGND VGND VPWR VPWR _2617_ sky130_fd_sc_hd__mux2_1
XFILLER_0_8_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_16_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5768_ cu.reg_file.reg_sp\[4\] _2534_ VGND VGND VPWR VPWR _2556_ sky130_fd_sc_hd__and2_1
X_4719_ net216 _1729_ _1731_ VGND VGND VPWR VPWR ih.t.next_count\[28\] sky130_fd_sc_hd__a21oi_1
XFILLER_0_16_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5699_ mc.cl.next_data\[13\] _2359_ _2490_ _2505_ VGND VGND VPWR VPWR _2506_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_16_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4890__B cu.pc.pc_o\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5611__B2 net5 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5611__A1 net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5375__A0 _1190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_473 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5507__A _1415_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3653__A1_N _0576_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output67_A net67 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3050_ ih.t.timer_max\[22\] _2760_ VGND VGND VPWR VPWR _2788_ sky130_fd_sc_hd__xor2_1
XANTENNA__5388__S _2237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3952_ alu.Cin _1023_ _1027_ VGND VGND VPWR VPWR _1028_ sky130_fd_sc_hd__o21a_1
XFILLER_0_18_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_535 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3883_ _0949_ _0958_ VGND VGND VPWR VPWR _0959_ sky130_fd_sc_hd__nor2_1
XFILLER_0_45_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5622_ ih.t.timer_max\[29\] _2146_ _2204_ ih.t.timer_max\[21\] VGND VGND VPWR VPWR
+ _2437_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5553_ _2367_ _2368_ _2371_ _1641_ VGND VGND VPWR VPWR _2372_ sky130_fd_sc_hd__o22a_2
XFILLER_0_26_451 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4504_ cu.reg_file.reg_h\[4\] _1316_ _1312_ cu.reg_file.reg_b\[4\] _1559_ VGND VGND
+ VPWR VPWR _1560_ sky130_fd_sc_hd__a221o_1
XFILLER_0_41_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5484_ _2247_ VGND VGND VPWR VPWR _2305_ sky130_fd_sc_hd__inv_2
XFILLER_0_13_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4435_ cu.reg_file.reg_h\[0\] _1316_ _1312_ cu.reg_file.reg_b\[0\] _1494_ VGND VGND
+ VPWR VPWR _1495_ sky130_fd_sc_hd__a221o_1
X_4366_ _0373_ _1295_ _1298_ cu.pc.pc_o\[5\] _1306_ VGND VGND VPWR VPWR _1429_ sky130_fd_sc_hd__a221o_1
XFILLER_0_6_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6105_ clknet_leaf_6_clk _0139_ net164 VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__dfrtp_4
X_3317_ _0384_ _0392_ VGND VGND VPWR VPWR _0393_ sky130_fd_sc_hd__or2b_1
XTAP_340 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4975__B cu.pc.pc_o\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4297_ cu.reg_file.reg_e\[2\] _1315_ VGND VGND VPWR VPWR _1363_ sky130_fd_sc_hd__and2_1
XTAP_362 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6036_ clknet_leaf_29_clk _0074_ net188 VGND VGND VPWR VPWR cu.reg_file.reg_h\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_3248_ cu.id.alu_opcode\[1\] cu.id.alu_opcode\[3\] VGND VGND VPWR VPWR _0324_ sky130_fd_sc_hd__nand2_2
XTAP_395 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4991__A cu.pc.pc_o\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3179_ cu.id.alu_opcode\[1\] cu.id.alu_opcode\[3\] cu.id.opcode\[0\] cu.id.alu_opcode\[0\]
+ VGND VGND VPWR VPWR _2916_ sky130_fd_sc_hd__or4bb_4
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5109__A0 cu.reg_file.reg_e\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4580__A1 _2702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4580__B2 _2697_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4231__A cu.pc.pc_o\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_59_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_86_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4399__A1 _1455_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output105_A net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5596__B1 _2247_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3310__A _2877_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5348__A0 _0619_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5936__S _2666_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5899__A1 _1074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5237__A _1369_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_70_549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_421 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4571__B2 _2697_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4571__A1 _2702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput107 net107 VGND VGND VPWR VPWR ss3[7] sky130_fd_sc_hd__clkbuf_4
Xoutput129 net129 VGND VGND VPWR VPWR ss6[5] sky130_fd_sc_hd__clkbuf_4
Xoutput118 net118 VGND VGND VPWR VPWR ss5[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_23_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5520__A0 net28 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4323__B2 cu.pc.pc_o\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4323__A1 cu.id.cb_opcode_y\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4220_ cu.reg_file.reg_a\[0\] _1276_ _1287_ cu.reg_file.reg_sp\[0\] VGND VGND VPWR
+ VPWR _1288_ sky130_fd_sc_hd__a22o_1
X_4151_ _0951_ _1214_ _0773_ _1220_ VGND VGND VPWR VPWR _1221_ sky130_fd_sc_hd__a31o_1
X_3102_ ih.t.count\[2\] _2746_ _2839_ VGND VGND VPWR VPWR _2840_ sky130_fd_sc_hd__and3_1
X_4082_ _1153_ _1117_ VGND VGND VPWR VPWR _1156_ sky130_fd_sc_hd__nor2_1
X_3033_ _2765_ _2769_ ih.t.count\[29\] VGND VGND VPWR VPWR _2771_ sky130_fd_sc_hd__a21oi_1
XANTENNA__4626__A2 _1667_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4984_ _1969_ _1970_ _1971_ _1799_ VGND VGND VPWR VPWR _1972_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_58_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3935_ _0986_ _1006_ _1010_ VGND VGND VPWR VPWR _1011_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_18_226 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5339__A0 _1190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5605_ ih.t.timer_max\[20\] _2150_ _2319_ ih.t.timer_max\[4\] _1661_ VGND VGND VPWR
+ VPWR _2421_ sky130_fd_sc_hd__a221o_1
XFILLER_0_33_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3866_ _0933_ _0941_ VGND VGND VPWR VPWR _0942_ sky130_fd_sc_hd__nor2_1
XFILLER_0_82_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5147__A _0618_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_14_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3797_ cu.reg_file.reg_b\[3\] _0426_ _0429_ cu.reg_file.reg_d\[3\] VGND VGND VPWR
+ VPWR _0873_ sky130_fd_sc_hd__a22o_1
X_5536_ net85 _1330_ VGND VGND VPWR VPWR _2355_ sky130_fd_sc_hd__or2_1
XFILLER_0_41_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5467_ _2292_ VGND VGND VPWR VPWR _0192_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_14_487 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4418_ _1473_ _1477_ _1478_ _1356_ VGND VGND VPWR VPWR _1479_ sky130_fd_sc_hd__o22ai_1
X_5398_ _1194_ net130 _2237_ VGND VGND VPWR VPWR _2244_ sky130_fd_sc_hd__mux2_1
X_4349_ cu.pc.pc_o\[4\] _1322_ _1315_ cu.reg_file.reg_e\[4\] _1412_ VGND VGND VPWR
+ VPWR _1413_ sky130_fd_sc_hd__a221o_1
X_6019_ clknet_leaf_3_clk _0057_ net170 VGND VGND VPWR VPWR cu.reg_file.reg_d\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_68_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4226__A _1293_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_492 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4553__B2 cu.reg_file.reg_sp\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4553__A1 cu.reg_file.reg_d\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_32_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_20_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3008__C ih.t.timer_max\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4136__A _0918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3720_ _0789_ _0792_ _0795_ _0752_ VGND VGND VPWR VPWR _0796_ sky130_fd_sc_hd__a31o_1
XFILLER_0_28_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_43_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3651_ cu.reg_file.reg_mem\[7\] _0418_ _0433_ cu.reg_file.reg_a\[7\] VGND VGND VPWR
+ VPWR _0727_ sky130_fd_sc_hd__a22o_1
X_3582_ cu.reg_file.reg_b\[5\] _0502_ _0499_ cu.reg_file.reg_a\[5\] VGND VGND VPWR
+ VPWR _0658_ sky130_fd_sc_hd__a22o_1
X_5321_ _2200_ VGND VGND VPWR VPWR _0138_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_262 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5252_ ih.t.timer_max\[26\] _2157_ _2153_ VGND VGND VPWR VPWR _2158_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5183_ _1647_ _2107_ VGND VGND VPWR VPWR _2108_ sky130_fd_sc_hd__and2_1
X_4203_ _1270_ VGND VGND VPWR VPWR _1271_ sky130_fd_sc_hd__buf_2
X_4134_ _0956_ _0957_ VGND VGND VPWR VPWR _1204_ sky130_fd_sc_hd__nor2_1
XFILLER_0_64_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4065_ _0610_ _1136_ _0652_ _0611_ VGND VGND VPWR VPWR _1139_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__3807__B1 _0748_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3016_ ih.t.timer_max\[12\] _2753_ VGND VGND VPWR VPWR _2754_ sky130_fd_sc_hd__or2_2
XANTENNA__4480__B1 _1286_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_502 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_449 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4967_ _1954_ _1955_ VGND VGND VPWR VPWR _1956_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3230__D_N _2923_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_546 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_73_151 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4898_ cu.pc.pc_o\[7\] _1892_ _1815_ VGND VGND VPWR VPWR _1893_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_31_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_31_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_46_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3918_ _0449_ _0972_ _0990_ _0993_ VGND VGND VPWR VPWR _0994_ sky130_fd_sc_hd__or4_2
XFILLER_0_61_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3849_ _0876_ _0924_ _0875_ VGND VGND VPWR VPWR _0925_ sky130_fd_sc_hd__o21ba_1
X_5519_ net31 _1625_ _2148_ net34 VGND VGND VPWR VPWR _2339_ sky130_fd_sc_hd__o22a_1
XFILLER_0_14_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xfanout164 net166 VGND VGND VPWR VPWR net164 sky130_fd_sc_hd__clkbuf_4
Xfanout153 net154 VGND VGND VPWR VPWR net153 sky130_fd_sc_hd__clkbuf_4
Xfanout175 net178 VGND VGND VPWR VPWR net175 sky130_fd_sc_hd__clkbuf_4
Xfanout186 net187 VGND VGND VPWR VPWR net186 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_69_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1122 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1111 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1100 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_457 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1155 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1144 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1133 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1177 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1166 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xclkbuf_leaf_22_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_22_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_25_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_64_184 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_346 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_379 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5515__A _1374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_917 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_906 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_939 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_928 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_18_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5974__RESET_B net161 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5870_ _2641_ VGND VGND VPWR VPWR _0246_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_75_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4821_ _1050_ _1817_ _1795_ VGND VGND VPWR VPWR _1822_ sky130_fd_sc_hd__mux2_1
XFILLER_0_34_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_75_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5396__S _2237_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_13_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_13_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__5962__A0 cu.id.imm_i\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4752_ _2880_ _2913_ _2935_ _0977_ _0350_ VGND VGND VPWR VPWR _1761_ sky130_fd_sc_hd__a41o_1
X_4683_ net217 _1705_ _1707_ VGND VGND VPWR VPWR ih.t.next_count\[16\] sky130_fd_sc_hd__a21oi_1
XFILLER_0_55_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3703_ _0512_ _0528_ VGND VGND VPWR VPWR _0779_ sky130_fd_sc_hd__nand2_2
XANTENNA__4517__B2 cu.reg_file.reg_h\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4517__A1 cu.reg_file.reg_b\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3634_ _0704_ _0706_ _0708_ _0709_ VGND VGND VPWR VPWR _0710_ sky130_fd_sc_hd__o31ai_4
XANTENNA__5425__A _2139_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_11_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_465 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3565_ cu.reg_file.reg_mem\[6\] _0640_ _0433_ cu.reg_file.reg_a\[6\] VGND VGND VPWR
+ VPWR _0641_ sky130_fd_sc_hd__a22o_1
X_5304_ _2189_ VGND VGND VPWR VPWR _0132_ sky130_fd_sc_hd__clkbuf_1
X_3496_ alu.Cin VGND VGND VPWR VPWR _0572_ sky130_fd_sc_hd__inv_2
X_6284_ clknet_leaf_35_clk _0266_ net159 VGND VGND VPWR VPWR cu.ir.idx\[0\] sky130_fd_sc_hd__dfrtp_2
X_5235_ _2143_ VGND VGND VPWR VPWR _0109_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5166_ _2096_ VGND VGND VPWR VPWR _0087_ sky130_fd_sc_hd__clkbuf_1
X_4117_ _1160_ VGND VGND VPWR VPWR _1189_ sky130_fd_sc_hd__buf_4
X_5097_ _2052_ VGND VGND VPWR VPWR _0062_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5245__A2 _2147_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4048_ _1032_ _1121_ _0916_ VGND VGND VPWR VPWR _1122_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_91_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_490 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5999_ clknet_leaf_1_clk _0037_ net153 VGND VGND VPWR VPWR cu.reg_file.reg_a\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_74_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xhold9 cu.id.can_be_interrupted VGND VGND VPWR VPWR net205 sky130_fd_sc_hd__dlygate4sd3_1
XANTENNA__3798__A2 _0640_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_57_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_57_438 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5944__A0 _0374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_110 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5944__S _2666_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output97_A net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3972__B _0545_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_40_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3350_ _0425_ _0421_ VGND VGND VPWR VPWR _0426_ sky130_fd_sc_hd__nor2_4
XTAP_725 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_703 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_758 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3281_ _0354_ _2953_ _0297_ _0356_ _2942_ VGND VGND VPWR VPWR _0357_ sky130_fd_sc_hd__a2111o_1
X_5020_ _1260_ _1263_ _0368_ VGND VGND VPWR VPWR _1999_ sky130_fd_sc_hd__mux2_1
XTAP_769 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3486__B2 cu.reg_file.reg_sp\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3486__A1 cu.reg_file.reg_h\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_2_clk clknet_2_0__leaf_clk VGND VGND VPWR VPWR clknet_leaf_2_clk sky130_fd_sc_hd__clkbuf_16
X_5922_ _2900_ _2372_ _2668_ VGND VGND VPWR VPWR _2670_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5853_ cu.reg_file.reg_sp\[14\] _1287_ VGND VGND VPWR VPWR _2630_ sky130_fd_sc_hd__or2_1
XANTENNA__4324__A cu.reg_file.reg_l\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_524 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4804_ _0306_ _0305_ _1805_ _2950_ VGND VGND VPWR VPWR _1806_ sky130_fd_sc_hd__o211a_1
X_5784_ cu.reg_file.reg_sp\[6\] _2535_ VGND VGND VPWR VPWR _2570_ sky130_fd_sc_hd__nand2_1
X_2996_ net69 VGND VGND VPWR VPWR _2734_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4735_ _0303_ _0449_ _1743_ VGND VGND VPWR VPWR _1744_ sky130_fd_sc_hd__or3_1
XFILLER_0_71_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4666_ ih.t.count\[10\] ih.t.count\[11\] _1693_ VGND VGND VPWR VPWR _1696_ sky130_fd_sc_hd__and3_1
XANTENNA__4978__B cu.pc.pc_o\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4597_ _1640_ VGND VGND VPWR VPWR _1641_ sky130_fd_sc_hd__clkinv_4
XANTENNA__5163__A1 _1193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_97 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3617_ _0294_ _0692_ _0536_ VGND VGND VPWR VPWR _0693_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_12_563 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3548_ _0539_ VGND VGND VPWR VPWR _0624_ sky130_fd_sc_hd__clkbuf_4
X_6267_ clknet_leaf_21_clk _0249_ net181 VGND VGND VPWR VPWR ih.t.timer_max\[15\]
+ sky130_fd_sc_hd__dfstp_2
X_3479_ _0400_ _0546_ VGND VGND VPWR VPWR _0555_ sky130_fd_sc_hd__and2_1
X_5218_ _2131_ VGND VGND VPWR VPWR _0104_ sky130_fd_sc_hd__clkbuf_1
X_6198_ clknet_leaf_7_clk net11 net168 VGND VGND VPWR VPWR ih.ih.ih.prev_data\[3\]
+ sky130_fd_sc_hd__dfrtp_1
X_5149_ _2951_ _2004_ _2086_ VGND VGND VPWR VPWR _2087_ sky130_fd_sc_hd__and3_1
XANTENNA__4426__B1 _1286_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_39_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_94_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_54_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5926__A0 _2893_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4901__A1 cu.pc.pc_o\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output135_A net135 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5231__C _2139_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3313__A _0374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5090__A0 cu.reg_file.reg_d\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_202 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_57_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5674__S _1739_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4520_ cu.pc.pc_o\[13\] _1485_ _1574_ VGND VGND VPWR VPWR _1575_ sky130_fd_sc_hd__o21a_1
XFILLER_0_25_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4451_ cu.reg_file.reg_b\[1\] _1313_ _1507_ _1509_ VGND VGND VPWR VPWR _1510_ sky130_fd_sc_hd__a211o_1
XANTENNA__5145__A1 cu.reg_file.reg_h\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3402_ _2896_ _0364_ _0477_ _2935_ _2949_ VGND VGND VPWR VPWR _0478_ sky130_fd_sc_hd__o2111ai_2
X_4382_ _1382_ _1438_ _1439_ _1444_ VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__a31o_2
X_6121_ clknet_leaf_30_clk _0155_ net183 VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__dfrtp_4
XTAP_500 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3333_ cu.id.starting_int_service _0408_ VGND VGND VPWR VPWR _0409_ sky130_fd_sc_hd__nor2_2
XTAP_511 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6052_ clknet_leaf_23_clk _0090_ net193 VGND VGND VPWR VPWR mc.cl.next_data\[10\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__5448__A2 net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3264_ cu.id.cb_opcode_z\[1\] VGND VGND VPWR VPWR _0340_ sky130_fd_sc_hd__buf_4
XANTENNA__3459__A1 cu.reg_file.reg_e\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_544 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4656__B1 _1687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5003_ cu.reg_file.reg_a\[1\] _1987_ _1985_ VGND VGND VPWR VPWR _1988_ sky130_fd_sc_hd__mux2_1
XANTENNA__3459__B2 cu.reg_file.reg_b\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_577 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_588 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3195_ _2931_ VGND VGND VPWR VPWR _2932_ sky130_fd_sc_hd__buf_2
XANTENNA__5605__C1 _1661_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5081__A0 cu.reg_file.reg_d\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5905_ ih.t.timer_max\[21\] _1191_ _2654_ VGND VGND VPWR VPWR _2660_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_73 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5620__A2 _2147_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3631__A1 cu.pc.pc_o\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_48_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4054__A _1110_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3631__B2 cu.reg_file.reg_b\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5836_ _1213_ _2615_ _2115_ VGND VGND VPWR VPWR _2616_ sky130_fd_sc_hd__mux2_1
X_2979_ net6 VGND VGND VPWR VPWR _2718_ sky130_fd_sc_hd__inv_2
XFILLER_0_8_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5767_ cu.reg_file.reg_sp\[4\] _2534_ VGND VGND VPWR VPWR _2555_ sky130_fd_sc_hd__nor2_1
XFILLER_0_29_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4718_ ih.t.count\[28\] _1729_ _1670_ VGND VGND VPWR VPWR _1731_ sky130_fd_sc_hd__o21ai_1
X_5698_ ih.t.timer_max\[29\] _2151_ _2320_ ih.t.timer_max\[13\] VGND VGND VPWR VPWR
+ _2505_ sky130_fd_sc_hd__a22oi_1
X_4649_ _1683_ _1684_ _1672_ VGND VGND VPWR VPWR _1685_ sky130_fd_sc_hd__and3b_1
XFILLER_0_16_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5136__A1 cu.reg_file.reg_h\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4895__A0 _1110_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6059__CLK clknet_2_0__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4229__A _1296_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3133__A _2870_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2972__A net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_94_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3622__B2 cu.reg_file.reg_e\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3622__A1 cu.reg_file.reg_c\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_27_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5375__A1 net120 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_35_485 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5127__A1 cu.reg_file.reg_h\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_77_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_500 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3951_ _2951_ _0368_ VGND VGND VPWR VPWR _1027_ sky130_fd_sc_hd__nand2_4
XANTENNA__3613__B2 cu.reg_file.reg_mem\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_374 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3882_ _0950_ _0956_ _0957_ VGND VGND VPWR VPWR _0958_ sky130_fd_sc_hd__or3_1
XFILLER_0_42_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_45_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5621_ net81 _1633_ _2432_ _2435_ VGND VGND VPWR VPWR _2436_ sky130_fd_sc_hd__o22a_1
X_5552_ _1649_ _2370_ VGND VGND VPWR VPWR _2371_ sky130_fd_sc_hd__and2_1
XFILLER_0_5_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4503_ cu.pc.pc_o\[12\] _1321_ _1314_ cu.reg_file.reg_d\[4\] _1558_ VGND VGND VPWR
+ VPWR _1559_ sky130_fd_sc_hd__a221o_1
XFILLER_0_13_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5483_ _2304_ VGND VGND VPWR VPWR _0196_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_13_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3218__A _0293_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4434_ cu.pc.pc_o\[8\] _1321_ _1314_ cu.reg_file.reg_d\[0\] _1493_ VGND VGND VPWR
+ VPWR _1494_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4365_ _1271_ _1427_ VGND VGND VPWR VPWR _1428_ sky130_fd_sc_hd__nor2_1
XFILLER_0_6_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_21_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_6104_ clknet_leaf_6_clk _0138_ net165 VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__dfrtp_2
XTAP_330 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3316_ _2887_ _0391_ _2950_ VGND VGND VPWR VPWR _0392_ sky130_fd_sc_hd__o21ai_2
XTAP_341 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_4296_ _0341_ _1295_ _1298_ cu.pc.pc_o\[2\] _1361_ VGND VGND VPWR VPWR _1362_ sky130_fd_sc_hd__a221o_1
X_6035_ clknet_leaf_33_clk _0073_ net161 VGND VGND VPWR VPWR cu.reg_file.reg_h\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_352 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_clkbuf_leaf_21_clk_A clknet_2_3__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3247_ _2878_ _2907_ _2908_ VGND VGND VPWR VPWR _0323_ sky130_fd_sc_hd__and3b_1
XTAP_396 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3178_ _2908_ _2914_ VGND VGND VPWR VPWR _2915_ sky130_fd_sc_hd__nor2_1
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_47 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_36_clk_A clknet_2_1__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_29_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5819_ _2599_ _2600_ VGND VGND VPWR VPWR _2601_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_17_496 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5109__A1 _1187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4580__A2 _1261_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_444 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5293__A0 _1052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_330 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5596__A1 net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5596__B2 net136 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_55_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5348__A1 net108 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4571__A2 _0619_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput108 net108 VGND VGND VPWR VPWR ss4[0] sky130_fd_sc_hd__buf_2
Xoutput119 net119 VGND VGND VPWR VPWR ss5[3] sky130_fd_sc_hd__clkbuf_4
XANTENNA__5520__A1 net30 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4150_ _0916_ _0940_ _1219_ _0817_ VGND VGND VPWR VPWR _1220_ sky130_fd_sc_hd__a2bb2o_1
X_3101_ ih.t.timer_max\[0\] ih.t.timer_max\[1\] ih.t.timer_max\[2\] VGND VGND VPWR
+ VPWR _2839_ sky130_fd_sc_hd__o21ai_1
Xoutput90 net90 VGND VGND VPWR VPWR ss1[6] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4081_ _1153_ _1112_ _1154_ _0610_ VGND VGND VPWR VPWR _1155_ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_37_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3032_ ih.t.count\[29\] _2765_ _2769_ VGND VGND VPWR VPWR _2770_ sky130_fd_sc_hd__and3_1
XFILLER_0_77_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4983_ _1624_ _1965_ _1795_ VGND VGND VPWR VPWR _1971_ sky130_fd_sc_hd__mux2_1
XFILLER_0_58_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3934_ _1007_ _0981_ _1009_ VGND VGND VPWR VPWR _1010_ sky130_fd_sc_hd__or3_1
XFILLER_0_85_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_58_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_18_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3865_ _0939_ _0940_ VGND VGND VPWR VPWR _0941_ sky130_fd_sc_hd__nand2_1
X_5604_ _1400_ _2419_ VGND VGND VPWR VPWR _2420_ sky130_fd_sc_hd__and2b_1
XFILLER_0_73_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5428__A _2139_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3796_ cu.reg_file.reg_sp\[11\] _0636_ _0748_ cu.reg_file.reg_h\[3\] VGND VGND VPWR
+ VPWR _0872_ sky130_fd_sc_hd__a22o_1
X_5535_ net93 _2194_ _2353_ VGND VGND VPWR VPWR _2354_ sky130_fd_sc_hd__a21o_1
XFILLER_0_5_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5466_ net62 _2085_ _2291_ VGND VGND VPWR VPWR _2292_ sky130_fd_sc_hd__mux2_1
XFILLER_0_14_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3770__B1 _0741_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4417_ _1460_ _1473_ VGND VGND VPWR VPWR _1478_ sky130_fd_sc_hd__nand2_1
XANTENNA__5511__A1 net64 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5511__B2 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5397_ _2243_ VGND VGND VPWR VPWR _0171_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5192__C_N _2951_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4348_ cu.reg_file.reg_sp\[4\] _0993_ _1344_ _0374_ _1364_ VGND VGND VPWR VPWR _1412_
+ sky130_fd_sc_hd__a221o_1
X_4279_ cu.pc.pc_o\[1\] _1322_ _1315_ cu.reg_file.reg_e\[1\] _1345_ VGND VGND VPWR
+ VPWR _1346_ sky130_fd_sc_hd__a221o_1
X_6018_ clknet_leaf_30_clk _0056_ net183 VGND VGND VPWR VPWR cu.reg_file.reg_d\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_96_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_49_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_300 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_49_363 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_37_514 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4538__C1 _1489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_64_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4553__A2 _1282_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_230 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5502__A1 ih.t.timer_max\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5266__A0 _1110_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3816__A1 cu.id.imm_i\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5018__A0 cu.reg_file.reg_a\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_87_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_15_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_28_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_43_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3650_ cu.reg_file.reg_c\[7\] _0427_ _0430_ cu.reg_file.reg_e\[7\] VGND VGND VPWR
+ VPWR _0726_ sky130_fd_sc_hd__a22o_1
XFILLER_0_43_539 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3581_ cu.reg_file.reg_d\[5\] _0492_ _0625_ cu.alu_f\[5\] _0656_ VGND VGND VPWR VPWR
+ _0657_ sky130_fd_sc_hd__a221o_1
X_5320_ _1190_ net96 _2195_ VGND VGND VPWR VPWR _2200_ sky130_fd_sc_hd__mux2_1
XFILLER_0_23_252 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5251_ _1073_ _1226_ _1667_ VGND VGND VPWR VPWR _2157_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4202_ _0294_ _1267_ _1269_ VGND VGND VPWR VPWR _1270_ sky130_fd_sc_hd__or3b_1
X_5182_ mc.cl.next_data\[13\] net23 mc.count VGND VGND VPWR VPWR _2107_ sky130_fd_sc_hd__mux2_1
XFILLER_0_48_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5257__A0 _1160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_7 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4133_ _1201_ _1202_ _1032_ VGND VGND VPWR VPWR _1203_ sky130_fd_sc_hd__a21o_1
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4064_ _0719_ _1137_ _1045_ VGND VGND VPWR VPWR _1138_ sky130_fd_sc_hd__a21oi_1
X_3015_ ih.t.timer_max\[10\] ih.t.timer_max\[11\] _2752_ VGND VGND VPWR VPWR _2753_
+ sky130_fd_sc_hd__or3_1
XANTENNA__3807__A1 cu.reg_file.reg_sp\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3807__B2 cu.reg_file.reg_h\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_436 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_78_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4480__B2 cu.reg_file.reg_sp\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4480__A1 cu.reg_file.reg_d\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5009__A0 cu.reg_file.reg_a\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4966_ _1233_ cu.pc.pc_o\[13\] VGND VGND VPWR VPWR _1955_ sky130_fd_sc_hd__and2_1
X_4897_ _1884_ _1891_ _1809_ VGND VGND VPWR VPWR _1892_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3917_ _0992_ VGND VGND VPWR VPWR _0993_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_46_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_452 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3848_ _0882_ _0885_ _0923_ VGND VGND VPWR VPWR _0924_ sky130_fd_sc_hd__a21boi_1
XANTENNA__5732__A1 net22 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3779_ _0853_ _0850_ VGND VGND VPWR VPWR _0855_ sky130_fd_sc_hd__or2b_1
XFILLER_0_89_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5518_ net33 _2191_ _1374_ VGND VGND VPWR VPWR _2338_ sky130_fd_sc_hd__o21a_1
XFILLER_0_14_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5496__B1 _2204_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5449_ _1335_ _1354_ VGND VGND VPWR VPWR _2277_ sky130_fd_sc_hd__nor2_1
XANTENNA__4299__A1 cu.reg_file.reg_sp\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4299__B2 _0341_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5248__A0 _1050_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4936__S _1814_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout165 net169 VGND VGND VPWR VPWR net165 sky130_fd_sc_hd__clkbuf_4
Xfanout154 net163 VGND VGND VPWR VPWR net154 sky130_fd_sc_hd__clkbuf_4
Xfanout176 net178 VGND VGND VPWR VPWR net176 sky130_fd_sc_hd__clkbuf_4
Xfanout187 net188 VGND VGND VPWR VPWR net187 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4237__A _1304_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4471__A1 cu.reg_file.reg_h\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1123 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1112 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1101 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4471__B2 cu.reg_file.reg_b\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1156 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1145 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1134 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1178 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1167 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_174 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_52_358 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_907 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_929 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_918 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5531__A _1739_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output42_A net42 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_200 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4820_ _1819_ _1820_ VGND VGND VPWR VPWR _1821_ sky130_fd_sc_hd__nor2_1
XANTENNA__5411__A0 _1188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_322 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_90_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_83_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5962__A1 _2429_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_152 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4751_ _1300_ _1739_ _1740_ _1759_ VGND VGND VPWR VPWR _1760_ sky130_fd_sc_hd__o22a_1
XFILLER_0_7_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4682_ ih.t.count\[16\] _1705_ _1670_ VGND VGND VPWR VPWR _1707_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_83_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3702_ _0771_ _0773_ _0777_ VGND VGND VPWR VPWR _0778_ sky130_fd_sc_hd__a21o_1
XANTENNA__5714__A1 _0618_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_196 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3633_ _2950_ _0341_ _0507_ VGND VGND VPWR VPWR _0709_ sky130_fd_sc_hd__a21o_1
XFILLER_0_24_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_51_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3564_ _0418_ VGND VGND VPWR VPWR _0640_ sky130_fd_sc_hd__clkbuf_8
X_6283_ clknet_leaf_13_clk _0265_ net181 VGND VGND VPWR VPWR ih.t.timer_max\[23\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__5425__B _2180_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5478__A0 net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5303_ _1194_ net90 _2182_ VGND VGND VPWR VPWR _2189_ sky130_fd_sc_hd__mux2_1
X_3495_ _0570_ _0510_ VGND VGND VPWR VPWR _0571_ sky130_fd_sc_hd__and2b_1
X_5234_ ih.t.enable _2085_ _2142_ VGND VGND VPWR VPWR _2143_ sky130_fd_sc_hd__mux2_1
X_5165_ cu.reg_file.reg_l\[7\] _1260_ _2088_ VGND VGND VPWR VPWR _2096_ sky130_fd_sc_hd__mux2_1
XANTENNA_fanout196_A net26 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4116_ net207 _1186_ _0370_ _1188_ VGND VGND VPWR VPWR _0010_ sky130_fd_sc_hd__a22o_1
XFILLER_0_38_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5096_ cu.reg_file.reg_d\[6\] _2051_ _2039_ VGND VGND VPWR VPWR _2052_ sky130_fd_sc_hd__mux2_1
X_4047_ _0804_ _0811_ VGND VGND VPWR VPWR _1121_ sky130_fd_sc_hd__nor2_1
XFILLER_0_93_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_66_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3896__A _2935_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5998_ clknet_leaf_0_clk _0036_ net153 VGND VGND VPWR VPWR cu.reg_file.reg_a\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_81_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4949_ cu.pc.pc_o\[12\] _1929_ VGND VGND VPWR VPWR _1939_ sky130_fd_sc_hd__and2_1
XFILLER_0_19_366 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_399 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5705__A1 net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_61_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_61_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_282 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_30_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4444__A1 cu.reg_file.reg_sp\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4444__B2 cu.reg_file.reg_h\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5944__A1 _2429_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_163 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_80_431 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5960__S _2686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_715 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_704 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3280_ _2918_ _0355_ _2883_ _2940_ VGND VGND VPWR VPWR _0356_ sky130_fd_sc_hd__a2bb2o_1
XTAP_759 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5880__A0 _1051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3486__A2 _0495_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4435__A1 cu.reg_file.reg_h\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4435__B2 cu.reg_file.reg_b\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5921_ _2669_ VGND VGND VPWR VPWR _0269_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4605__A _1648_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5852_ _2629_ VGND VGND VPWR VPWR _0240_ sky130_fd_sc_hd__clkbuf_1
X_4803_ _2939_ _2916_ _2932_ _0331_ VGND VGND VPWR VPWR _1805_ sky130_fd_sc_hd__o22a_1
X_5783_ cu.reg_file.reg_sp\[6\] _2535_ VGND VGND VPWR VPWR _2569_ sky130_fd_sc_hd__or2_1
X_2995_ _2714_ _2733_ VGND VGND VPWR VPWR ih.ih.int_f.data_in sky130_fd_sc_hd__nand2_1
X_4734_ _2939_ _2916_ _2878_ VGND VGND VPWR VPWR _1743_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_71_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4665_ net222 _1693_ _1695_ VGND VGND VPWR VPWR ih.t.next_count\[10\] sky130_fd_sc_hd__a21oi_1
X_4596_ _1629_ _1639_ VGND VGND VPWR VPWR _1640_ sky130_fd_sc_hd__nor2_1
X_3616_ cu.id.cb_opcode_y\[0\] VGND VGND VPWR VPWR _0692_ sky130_fd_sc_hd__inv_2
X_3547_ cu.reg_file.reg_c\[6\] _0485_ _0622_ VGND VGND VPWR VPWR _0623_ sky130_fd_sc_hd__a21o_1
X_6266_ clknet_leaf_22_clk _0248_ net191 VGND VGND VPWR VPWR ih.t.timer_max\[14\]
+ sky130_fd_sc_hd__dfstp_1
XFILLER_0_86_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_86_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3478_ _0514_ _0553_ VGND VGND VPWR VPWR _0554_ sky130_fd_sc_hd__nor2_1
XANTENNA__5871__A0 _2163_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_6197_ clknet_leaf_7_clk net10 net168 VGND VGND VPWR VPWR ih.ih.ih.prev_data\[2\]
+ sky130_fd_sc_hd__dfrtp_1
X_5217_ _1188_ ih.gpio_interrupt_mask\[3\] _2127_ VGND VGND VPWR VPWR _2131_ sky130_fd_sc_hd__mux2_1
X_5148_ _2023_ VGND VGND VPWR VPWR _2086_ sky130_fd_sc_hd__inv_2
X_5079_ _2040_ VGND VGND VPWR VPWR _0056_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4426__A1 cu.reg_file.reg_d\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4426__B2 cu.reg_file.reg_sp\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_94_567 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_66_258 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5926__A1 _2410_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4250__A _2893_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_339 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3313__B cu.id.cb_opcode_x\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output128_A net128 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5614__A0 cu.reg_file.reg_mem\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4425__A _1269_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5020__S _0368_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_25_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_25_155 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_25_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4450_ cu.pc.pc_o\[9\] _1322_ _1315_ cu.reg_file.reg_d\[1\] _1508_ VGND VGND VPWR
+ VPWR _1509_ sky130_fd_sc_hd__a221o_1
XFILLER_0_25_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4381_ _1353_ _1434_ _1443_ _1371_ VGND VGND VPWR VPWR _1444_ sky130_fd_sc_hd__a22o_1
X_3401_ _2902_ _0300_ _2912_ VGND VGND VPWR VPWR _0477_ sky130_fd_sc_hd__a21o_1
XFILLER_0_40_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6120_ clknet_leaf_7_clk _0154_ net167 VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_0_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3332_ _2877_ _2878_ _2932_ _2925_ VGND VGND VPWR VPWR _0408_ sky130_fd_sc_hd__o22a_1
XFILLER_0_0_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_501 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6051_ clknet_leaf_22_clk _0089_ net191 VGND VGND VPWR VPWR mc.cl.next_data\[9\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__5448__A3 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_56_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4105__B1 _1178_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3263_ _0296_ _0297_ _0337_ _0338_ VGND VGND VPWR VPWR _0339_ sky130_fd_sc_hd__or4_2
XANTENNA__3459__A2 _0488_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_545 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5002_ _1051_ _1623_ _0368_ VGND VGND VPWR VPWR _1987_ sky130_fd_sc_hd__mux2_1
X_3194_ cu.id.opcode\[2\] cu.id.opcode\[1\] cu.id.opcode\[6\] cu.id.opcode\[7\] VGND
+ VGND VPWR VPWR _2931_ sky130_fd_sc_hd__or4_1
XTAP_578 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_589 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_72_52 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5904_ _2659_ VGND VGND VPWR VPWR _0262_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4335__A _1393_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout159_A net160 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3631__A2 _0501_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5835_ _2613_ _2614_ VGND VGND VPWR VPWR _2615_ sky130_fd_sc_hd__xnor2_1
XANTENNA__4054__B _1126_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_239 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2978_ net12 VGND VGND VPWR VPWR _2717_ sky130_fd_sc_hd__inv_2
X_5766_ _2554_ VGND VGND VPWR VPWR _0229_ sky130_fd_sc_hd__clkbuf_1
X_4717_ _1729_ _1730_ VGND VGND VPWR VPWR ih.t.next_count\[27\] sky130_fd_sc_hd__nor2_1
X_5697_ net5 _1650_ _2488_ _2504_ VGND VGND VPWR VPWR _0210_ sky130_fd_sc_hd__a31o_1
XANTENNA__3395__A1 _2878_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4648_ ih.t.count\[4\] _1679_ ih.t.count\[5\] VGND VGND VPWR VPWR _1684_ sky130_fd_sc_hd__a21o_1
XFILLER_0_4_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_103 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_486 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4579_ _2702_ _1194_ _1624_ _2697_ VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__a22o_1
X_6249_ clknet_leaf_42_clk _0231_ net155 VGND VGND VPWR VPWR cu.reg_file.reg_sp\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__5844__A0 _1209_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_309 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_79_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_272 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3308__B _0379_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3324__A _2950_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_136 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3950_ _0964_ _1015_ _1016_ _1017_ _1025_ VGND VGND VPWR VPWR _1026_ sky130_fd_sc_hd__a2111o_1
XANTENNA__3613__A2 _0498_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3881_ _0866_ _0906_ VGND VGND VPWR VPWR _0957_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_73_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5620_ net113 _2147_ _2225_ net121 _2434_ VGND VGND VPWR VPWR _2435_ sky130_fd_sc_hd__a221o_1
X_5551_ net9 _2345_ _2369_ net17 VGND VGND VPWR VPWR _2370_ sky130_fd_sc_hd__a22o_1
XFILLER_0_5_314 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4574__B1 _1226_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4502_ cu.reg_file.reg_sp\[12\] _0992_ _1343_ cu.id.imm_i\[12\] _1323_ VGND VGND
+ VPWR VPWR _1558_ sky130_fd_sc_hd__a221o_1
XFILLER_0_41_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5482_ net66 _0618_ _2303_ VGND VGND VPWR VPWR _2304_ sky130_fd_sc_hd__mux2_1
X_4433_ cu.reg_file.reg_sp\[8\] _0992_ _1343_ cu.id.imm_i\[8\] _1323_ VGND VGND VPWR
+ VPWR _1493_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4364_ cu.reg_file.reg_c\[5\] _1281_ _1426_ VGND VGND VPWR VPWR _1427_ sky130_fd_sc_hd__a21oi_1
X_6103_ clknet_leaf_30_clk _0137_ net187 VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__dfrtp_4
X_4295_ _1271_ _1360_ VGND VGND VPWR VPWR _1361_ sky130_fd_sc_hd__nor2_1
XTAP_320 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3315_ _2936_ _0385_ _0386_ _2928_ _0390_ VGND VGND VPWR VPWR _0391_ sky130_fd_sc_hd__a311o_1
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_331 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6034_ clknet_leaf_28_clk _0072_ net188 VGND VGND VPWR VPWR cu.reg_file.reg_h\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__3234__A _2923_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_353 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3246_ _2896_ _2911_ _2935_ VGND VGND VPWR VPWR _0322_ sky130_fd_sc_hd__nand3_2
XTAP_364 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3177_ _2912_ _2913_ VGND VGND VPWR VPWR _2914_ sky130_fd_sc_hd__nand2_2
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4801__A1 _2923_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_59 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_91_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_76_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5818_ _2590_ _2593_ _2591_ VGND VGND VPWR VPWR _2600_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_91_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4512__B _1561_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_17_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5749_ cu.reg_file.reg_sp\[1\] _2531_ _2539_ VGND VGND VPWR VPWR _2540_ sky130_fd_sc_hd__mux2_1
XFILLER_0_12_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3144__A _2877_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2983__A net7 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5596__A2 _2236_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xoutput109 net109 VGND VGND VPWR VPWR ss4[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_50_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5520__A2 net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output72_A net72 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput80 net80 VGND VGND VPWR VPWR ss0[4] sky130_fd_sc_hd__clkbuf_4
X_3100_ _2836_ ih.t.count\[0\] ih.t.timer_max\[0\] VGND VGND VPWR VPWR _2838_ sky130_fd_sc_hd__mux2_1
Xoutput91 net91 VGND VGND VPWR VPWR ss1[7] sky130_fd_sc_hd__clkbuf_4
X_4080_ _0611_ _0671_ VGND VGND VPWR VPWR _1154_ sky130_fd_sc_hd__nand2_1
X_3031_ ih.t.timer_max\[28\] _2764_ ih.t.timer_max\[29\] VGND VGND VPWR VPWR _2769_
+ sky130_fd_sc_hd__o21ai_1
XFILLER_0_53_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4982_ _1966_ _1968_ _1798_ VGND VGND VPWR VPWR _1970_ sky130_fd_sc_hd__o21bai_1
XFILLER_0_46_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3933_ _0998_ _1008_ VGND VGND VPWR VPWR _1009_ sky130_fd_sc_hd__nor2_1
XFILLER_0_85_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_73_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_312 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_537 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3864_ _0877_ _0924_ VGND VGND VPWR VPWR _0940_ sky130_fd_sc_hd__xnor2_1
X_5603_ ih.t.timer_max\[12\] _2193_ _2314_ ih.t.timer_max\[4\] _2418_ VGND VGND VPWR
+ VPWR _2419_ sky130_fd_sc_hd__a221o_1
XANTENNA__5428__B _2194_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4332__B _1393_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3795_ cu.id.imm_i\[11\] _0739_ _0870_ _0653_ VGND VGND VPWR VPWR _0871_ sky130_fd_sc_hd__a22oi_4
X_5534_ net125 _2236_ _2247_ net133 VGND VGND VPWR VPWR _2353_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5465_ _2290_ _2284_ VGND VGND VPWR VPWR _2291_ sky130_fd_sc_hd__nor2_1
XANTENNA__3770__B2 cu.reg_file.reg_h\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3770__A1 cu.reg_file.reg_d\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4416_ _1356_ _1460_ _1402_ VGND VGND VPWR VPWR _1477_ sky130_fd_sc_hd__o21a_1
XFILLER_0_78_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5396_ _1192_ net129 _2237_ VGND VGND VPWR VPWR _2243_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_372 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4347_ cu.reg_file.reg_l\[4\] _1317_ VGND VGND VPWR VPWR _1411_ sky130_fd_sc_hd__and2_1
XANTENNA__5275__A1 _1074_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4278_ cu.reg_file.reg_sp\[1\] _0993_ _1344_ _0340_ _1324_ VGND VGND VPWR VPWR _1345_
+ sky130_fd_sc_hd__a221o_1
XANTENNA__4078__A2 _0663_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_94_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_6017_ clknet_leaf_3_clk _0055_ net156 VGND VGND VPWR VPWR cu.reg_file.reg_c\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_194 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3229_ _2902_ _2884_ _2875_ _2876_ VGND VGND VPWR VPWR _0305_ sky130_fd_sc_hd__or4bb_1
XFILLER_0_49_331 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_32_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__2978__A net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_404 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3761__A1 cu.reg_file.reg_a\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3513__A1 cu.reg_file.reg_c\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3513__B2 cu.reg_file.reg_e\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5266__A1 _1263_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4417__B _1473_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output110_A net110 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_481 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_55_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA_clkbuf_leaf_20_clk_A clknet_2_3__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3580_ cu.pc.pc_o\[5\] _0501_ VGND VGND VPWR VPWR _0656_ sky130_fd_sc_hd__and2_1
XANTENNA__3752__A1 cu.reg_file.reg_a\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3752__B2 cu.reg_file.reg_mem\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5250_ _2156_ VGND VGND VPWR VPWR _0111_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_54_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4201_ cu.id.state\[1\] cu.id.state\[0\] _1268_ VGND VGND VPWR VPWR _1269_ sky130_fd_sc_hd__and3b_4
XANTENNA_clkbuf_leaf_35_clk_A clknet_2_1__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3504__A1 cu.reg_file.reg_mem\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5181_ _2106_ VGND VGND VPWR VPWR _0092_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_48_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3504__B2 cu.reg_file.reg_h\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4132_ _0942_ _0943_ VGND VGND VPWR VPWR _1202_ sky130_fd_sc_hd__or2_1
XANTENNA__5257__A1 _1213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4063_ _0603_ _1136_ VGND VGND VPWR VPWR _1137_ sky130_fd_sc_hd__nand2_1
X_3014_ ih.t.timer_max\[9\] _2751_ VGND VGND VPWR VPWR _2752_ sky130_fd_sc_hd__or2_2
XANTENNA__3512__A _0587_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4480__A2 _1282_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4965_ _1233_ cu.pc.pc_o\[13\] VGND VGND VPWR VPWR _1954_ sky130_fd_sc_hd__nor2_1
XFILLER_0_19_515 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3916_ _0991_ VGND VGND VPWR VPWR _0992_ sky130_fd_sc_hd__buf_2
X_4896_ _1889_ _1890_ _1798_ VGND VGND VPWR VPWR _1891_ sky130_fd_sc_hd__mux2_1
XFILLER_0_73_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3847_ _0887_ _0922_ VGND VGND VPWR VPWR _0923_ sky130_fd_sc_hd__or2_1
XFILLER_0_34_518 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_464 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_231 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3778_ _0850_ _0853_ VGND VGND VPWR VPWR _0854_ sky130_fd_sc_hd__or2b_1
X_5517_ net32 _1330_ _1354_ VGND VGND VPWR VPWR _2337_ sky130_fd_sc_hd__or3_1
XFILLER_0_14_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5448_ net73 net75 net72 net74 _1354_ _1330_ VGND VGND VPWR VPWR _2276_ sky130_fd_sc_hd__mux4_1
XANTENNA__4299__A2 _0993_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5379_ _1194_ net122 _2226_ VGND VGND VPWR VPWR _2233_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_481 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xfanout155 net163 VGND VGND VPWR VPWR net155 sky130_fd_sc_hd__clkbuf_4
Xfanout177 net178 VGND VGND VPWR VPWR net177 sky130_fd_sc_hd__buf_2
Xfanout188 net196 VGND VGND VPWR VPWR net188 sky130_fd_sc_hd__clkbuf_4
XANTENNA__5248__A1 _1623_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xfanout166 net169 VGND VGND VPWR VPWR net166 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_96_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_1113 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1102 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_96_278 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1146 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1135 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1124 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1179 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1168 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1157 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3982__A1 _0298_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_64_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_908 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_919 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4428__A _1269_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5958__S _2686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5411__A1 net135 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4750_ _1645_ _1755_ _1758_ _1269_ VGND VGND VPWR VPWR _1759_ sky130_fd_sc_hd__o22a_1
XANTENNA__4163__A _2920_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4681_ _1705_ _1706_ VGND VGND VPWR VPWR ih.t.next_count\[15\] sky130_fd_sc_hd__nor2_1
XANTENNA__5983__RESET_B net188 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3701_ _0512_ _0776_ VGND VGND VPWR VPWR _0777_ sky130_fd_sc_hd__nor2_2
XANTENNA__3973__B2 _0545_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_28_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_50_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3632_ cu.reg_file.reg_sp\[2\] _0624_ _0492_ cu.reg_file.reg_d\[2\] _0707_ VGND VGND
+ VPWR VPWR _0708_ sky130_fd_sc_hd__a221o_1
X_5302_ _2188_ VGND VGND VPWR VPWR _0131_ sky130_fd_sc_hd__clkbuf_1
X_3563_ cu.reg_file.reg_c\[6\] _0427_ _0430_ cu.reg_file.reg_e\[6\] VGND VGND VPWR
+ VPWR _0639_ sky130_fd_sc_hd__a22o_1
X_6282_ clknet_leaf_13_clk _0264_ net181 VGND VGND VPWR VPWR ih.t.timer_max\[22\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__5478__A1 _0618_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3494_ _0569_ VGND VGND VPWR VPWR _0570_ sky130_fd_sc_hd__buf_2
XFILLER_0_3_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5233_ _2140_ _2141_ VGND VGND VPWR VPWR _2142_ sky130_fd_sc_hd__nor2_1
XANTENNA__3489__B1 _0536_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5164_ _2095_ VGND VGND VPWR VPWR _0086_ sky130_fd_sc_hd__clkbuf_1
X_4115_ _1187_ VGND VGND VPWR VPWR _1188_ sky130_fd_sc_hd__buf_4
X_5095_ _1193_ _1624_ _2035_ VGND VGND VPWR VPWR _2051_ sky130_fd_sc_hd__mux2_1
XANTENNA__4989__B1 _1233_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4046_ _0757_ _0767_ VGND VGND VPWR VPWR _1120_ sky130_fd_sc_hd__or2_1
XANTENNA__3354__B1_N _0429_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5650__A1 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5997_ clknet_leaf_1_clk _0035_ net153 VGND VGND VPWR VPWR cu.reg_file.reg_a\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_4948_ _1938_ VGND VGND VPWR VPWR _0027_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3413__B1 _0488_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4879_ _0387_ cu.pc.pc_o\[6\] VGND VGND VPWR VPWR _1875_ sky130_fd_sc_hd__nor2_1
XFILLER_0_46_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_348 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5705__A2 _1650_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4947__S _1814_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5632__A _1649_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4248__A _1309_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5641__A1 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2991__A net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3903__A_N _0308_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_495 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5157__A0 cu.reg_file.reg_l\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5807__A cu.reg_file.reg_sp\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_716 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_705 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_0_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_749 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5880__A1 ih.t.timer_max\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_2_2__f_clk_A clknet_0_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5920_ _2923_ _2350_ _2668_ VGND VGND VPWR VPWR _2669_ sky130_fd_sc_hd__mux2_1
X_5851_ cu.reg_file.reg_sp\[14\] _2628_ _2538_ VGND VGND VPWR VPWR _2629_ sky130_fd_sc_hd__mux2_1
X_2994_ _2720_ _2726_ _2732_ VGND VGND VPWR VPWR _2733_ sky130_fd_sc_hd__and3_1
XFILLER_0_61_65 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5396__A0 _1192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4802_ _1803_ _1742_ VGND VGND VPWR VPWR _1804_ sky130_fd_sc_hd__or2b_1
XFILLER_0_0_79 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5782_ _2568_ VGND VGND VPWR VPWR _0231_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_28_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_270 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4733_ _2893_ _1741_ VGND VGND VPWR VPWR _1742_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_16_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_28_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4664_ ih.t.count\[10\] _1693_ _1670_ VGND VGND VPWR VPWR _1695_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_71_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4595_ _1373_ _1417_ _1637_ _1638_ VGND VGND VPWR VPWR _1639_ sky130_fd_sc_hd__or4_1
X_3615_ cu.reg_file.reg_sp\[3\] _0539_ _0492_ cu.reg_file.reg_d\[3\] _0690_ VGND VGND
+ VPWR VPWR _0691_ sky130_fd_sc_hd__a221o_1
X_3546_ cu.reg_file.reg_e\[6\] _0489_ _0621_ cu.reg_file.reg_l\[6\] VGND VGND VPWR
+ VPWR _0622_ sky130_fd_sc_hd__a22o_1
X_6265_ clknet_leaf_15_clk _0247_ net179 VGND VGND VPWR VPWR ih.t.timer_max\[13\]
+ sky130_fd_sc_hd__dfrtp_4
X_5216_ _2130_ VGND VGND VPWR VPWR _0103_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5320__A0 _1190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3477_ _0400_ _0528_ VGND VGND VPWR VPWR _0553_ sky130_fd_sc_hd__or2b_1
X_6196_ clknet_leaf_7_clk net9 net167 VGND VGND VPWR VPWR ih.ih.ih.prev_data\[1\]
+ sky130_fd_sc_hd__dfrtp_1
X_5147_ _0618_ VGND VGND VPWR VPWR _2085_ sky130_fd_sc_hd__clkbuf_4
X_5078_ cu.reg_file.reg_d\[0\] _2036_ _2039_ VGND VGND VPWR VPWR _2040_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_521 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4426__A2 _1282_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4029_ _0611_ _0729_ _0607_ _0552_ VGND VGND VPWR VPWR _1103_ sky130_fd_sc_hd__a211o_1
XFILLER_0_94_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_39_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_94_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_47_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_19_164 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4362__A1 cu.reg_file.reg_a\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4362__B2 cu.reg_file.reg_sp\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_373 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5614__A1 _2429_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5301__S _2182_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4425__B _1484_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_57_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5917__A2 _2532_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_65_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_80_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_13_329 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4380_ _1441_ _1442_ VGND VGND VPWR VPWR _1443_ sky130_fd_sc_hd__nand2_1
XFILLER_0_0_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3400_ _0452_ _0303_ _0450_ _0475_ VGND VGND VPWR VPWR _0476_ sky130_fd_sc_hd__or4b_1
X_3331_ _0299_ _0329_ _0406_ _2877_ VGND VGND VPWR VPWR _0407_ sky130_fd_sc_hd__o2bb2a_4
XTAP_502 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6050_ clknet_leaf_24_clk _0088_ net190 VGND VGND VPWR VPWR mc.cl.next_data\[8\]
+ sky130_fd_sc_hd__dfrtp_1
X_3262_ _2907_ _2914_ VGND VGND VPWR VPWR _0338_ sky130_fd_sc_hd__and2_1
XTAP_535 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3193_ _2918_ _2919_ _2922_ _2924_ _2929_ VGND VGND VPWR VPWR _2930_ sky130_fd_sc_hd__o311a_1
XTAP_568 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5001_ _1986_ VGND VGND VPWR VPWR _0032_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4616__A _2923_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5903_ ih.t.timer_max\[20\] _1189_ _2654_ VGND VGND VPWR VPWR _2659_ sky130_fd_sc_hd__mux2_1
XFILLER_0_76_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5369__A0 _1052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5834_ _2604_ _2607_ _2605_ VGND VGND VPWR VPWR _2614_ sky130_fd_sc_hd__a21bo_1
XFILLER_0_91_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_229 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_462 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5447__A _1417_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2977_ net5 VGND VGND VPWR VPWR _2716_ sky130_fd_sc_hd__inv_2
X_5765_ cu.reg_file.reg_sp\[3\] _2553_ _2539_ VGND VGND VPWR VPWR _2554_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4716_ net232 _1726_ _1687_ VGND VGND VPWR VPWR _1730_ sky130_fd_sc_hd__o21ai_1
X_5696_ _2503_ _1643_ cu.reg_file.reg_mem\[12\] _1646_ VGND VGND VPWR VPWR _2504_
+ sky130_fd_sc_hd__a2bb2o_1
X_4647_ ih.t.count\[4\] ih.t.count\[5\] _1679_ VGND VGND VPWR VPWR _1683_ sky130_fd_sc_hd__and3_1
XFILLER_0_71_295 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_71_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5541__B1 _2204_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_340 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_159 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4578_ _0516_ _1200_ VGND VGND VPWR VPWR _1624_ sky130_fd_sc_hd__nor2_4
X_3529_ _0399_ _0546_ VGND VGND VPWR VPWR _0605_ sky130_fd_sc_hd__or2_1
X_6248_ clknet_leaf_41_clk _0230_ net151 VGND VGND VPWR VPWR cu.reg_file.reg_sp\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_6179_ clknet_leaf_19_clk _0213_ net183 VGND VGND VPWR VPWR cu.reg_file.reg_mem\[15\]
+ sky130_fd_sc_hd__dfrtp_2
XANTENNA__5121__S _2066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4804__C1 _2950_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_35_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5780__A0 _1144_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5523__C _1648_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4099__B1 _0773_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5031__S _2002_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5966__S _2686_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3880_ _0951_ _0952_ _0955_ VGND VGND VPWR VPWR _0956_ sky130_fd_sc_hd__or3_1
XFILLER_0_26_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5550_ _1335_ _1372_ _1661_ VGND VGND VPWR VPWR _2369_ sky130_fd_sc_hd__and3_2
XFILLER_0_53_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_337 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4574__B2 _2697_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4574__A1 _2702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_84_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5481_ _2302_ _2284_ VGND VGND VPWR VPWR _2303_ sky130_fd_sc_hd__nor2_1
X_4501_ cu.pc.pc_o\[12\] _1485_ _1556_ VGND VGND VPWR VPWR _1557_ sky130_fd_sc_hd__o21a_1
XFILLER_0_41_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4432_ cu.pc.pc_o\[8\] _1485_ _1491_ VGND VGND VPWR VPWR _1492_ sky130_fd_sc_hd__o21a_1
XANTENNA__4326__A1 cu.pc.pc_o\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4326__B2 cu.reg_file.reg_e\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4363_ cu.reg_file.reg_e\[5\] _1283_ _1285_ cu.reg_file.reg_l\[5\] _1425_ VGND VGND
+ VPWR VPWR _1426_ sky130_fd_sc_hd__a221o_1
X_6102_ clknet_leaf_9_clk _0136_ net174 VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__dfrtp_2
X_4294_ cu.reg_file.reg_c\[2\] _1281_ _1359_ VGND VGND VPWR VPWR _1360_ sky130_fd_sc_hd__a21oi_1
XTAP_321 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_310 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3314_ _0388_ _0389_ _2918_ VGND VGND VPWR VPWR _0390_ sky130_fd_sc_hd__a21oi_1
XTAP_332 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3245_ _0318_ _0319_ _0320_ _2913_ VGND VGND VPWR VPWR _0321_ sky130_fd_sc_hd__or4b_4
XTAP_343 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6033_ clknet_leaf_1_clk _0071_ net153 VGND VGND VPWR VPWR cu.reg_file.reg_e\[7\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_387 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3176_ _2909_ _2878_ VGND VGND VPWR VPWR _2913_ sky130_fd_sc_hd__or2_2
XFILLER_0_13_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_95_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_49_513 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_38 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_76_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_321 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_527 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_36_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_324 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_131 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5817_ _2597_ _2598_ VGND VGND VPWR VPWR _2599_ sky130_fd_sc_hd__nand2_1
XFILLER_0_8_175 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_17_454 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5748_ _2538_ VGND VGND VPWR VPWR _2539_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_44_240 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_273 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_44_284 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5679_ mc.cl.next_data\[8\] _2359_ _2489_ _2490_ VGND VGND VPWR VPWR _2491_ sky130_fd_sc_hd__o2bb2a_1
XANTENNA__6285__RESET_B net160 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_170 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4150__A1_N _0916_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4256__A _1323_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_310 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4795__A1_N _0986_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3461__D1 _0536_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4556__A1 _1296_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5815__A cu.reg_file.reg_sp\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_265 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput70 net70 VGND VGND VPWR VPWR programmable_gpio_wr[2] sky130_fd_sc_hd__buf_2
XANTENNA__5520__A3 net29 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output65_A net65 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput81 net81 VGND VGND VPWR VPWR ss0[5] sky130_fd_sc_hd__clkbuf_4
Xoutput92 net92 VGND VGND VPWR VPWR ss2[0] sky130_fd_sc_hd__clkbuf_4
XANTENNA__5550__A _1335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3030_ ih.t.timer_max\[31\] _2767_ VGND VGND VPWR VPWR _2768_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_37_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4981_ _1966_ _1968_ VGND VGND VPWR VPWR _1969_ sky130_fd_sc_hd__and2_1
XFILLER_0_58_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3932_ _1004_ _0986_ VGND VGND VPWR VPWR _1008_ sky130_fd_sc_hd__and2b_1
XANTENNA_clkbuf_leaf_9_clk_A clknet_2_2__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4613__B _1364_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3863_ _0936_ _0938_ VGND VGND VPWR VPWR _0939_ sky130_fd_sc_hd__and2b_1
X_5602_ ih.t.timer_max\[28\] _2146_ _2204_ ih.t.timer_max\[20\] VGND VGND VPWR VPWR
+ _2418_ sky130_fd_sc_hd__a22o_1
X_5533_ _2352_ VGND VGND VPWR VPWR _0198_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_26_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3794_ cu.reg_file.reg_a\[3\] _0625_ _0628_ cu.reg_file.reg_mem\[11\] _0869_ VGND
+ VGND VPWR VPWR _0870_ sky130_fd_sc_hd__a221o_1
XFILLER_0_41_232 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5464_ _2194_ VGND VGND VPWR VPWR _2290_ sky130_fd_sc_hd__inv_2
XFILLER_0_41_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3770__A2 _0488_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4415_ _1463_ _1474_ VGND VGND VPWR VPWR _1476_ sky130_fd_sc_hd__nand2_1
X_5395_ _2242_ VGND VGND VPWR VPWR _0170_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_4346_ _0374_ _1295_ _1298_ cu.pc.pc_o\[4\] _1409_ VGND VGND VPWR VPWR _1410_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_384 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5460__A _1369_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4277_ _1343_ VGND VGND VPWR VPWR _1344_ sky130_fd_sc_hd__clkbuf_4
X_6016_ clknet_leaf_4_clk _0054_ net170 VGND VGND VPWR VPWR cu.reg_file.reg_c\[6\]
+ sky130_fd_sc_hd__dfrtp_4
X_3228_ _2936_ _2885_ _2941_ VGND VGND VPWR VPWR _0304_ sky130_fd_sc_hd__nand3_2
XTAP_195 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3159_ _2894_ net238 VGND VGND VPWR VPWR _2896_ sky130_fd_sc_hd__nand2_4
XFILLER_0_68_129 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_96_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_34_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_34_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_76_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_91_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4538__B2 cu.pc.pc_o\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_484 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_25_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_25_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA_output103_A net103 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_493 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_55_302 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_51_552 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_2_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_23_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_427 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_2_148 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4200_ cu.id.state\[2\] VGND VGND VPWR VPWR _1268_ sky130_fd_sc_hd__buf_2
X_5180_ _1647_ _2105_ VGND VGND VPWR VPWR _2106_ sky130_fd_sc_hd__and2_1
X_4131_ _0942_ _0943_ VGND VGND VPWR VPWR _1201_ sky130_fd_sc_hd__nand2_1
X_4062_ _0599_ _1100_ VGND VGND VPWR VPWR _1136_ sky130_fd_sc_hd__nor2_1
X_3013_ ih.t.timer_max\[7\] ih.t.timer_max\[8\] _2750_ VGND VGND VPWR VPWR _2751_
+ sky130_fd_sc_hd__or3_1
XANTENNA__4465__B1 _1284_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4624__A _1665_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xclkbuf_leaf_16_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_16_clk sky130_fd_sc_hd__clkbuf_16
X_4964_ cu.pc.pc_o\[13\] _1939_ VGND VGND VPWR VPWR _1953_ sky130_fd_sc_hd__xor2_1
XFILLER_0_80_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3915_ _0295_ _0968_ VGND VGND VPWR VPWR _0991_ sky130_fd_sc_hd__or2_1
X_4895_ _1110_ _1884_ _1794_ VGND VGND VPWR VPWR _1890_ sky130_fd_sc_hd__mux2_1
XFILLER_0_6_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3846_ _0920_ _0896_ _0796_ _0921_ VGND VGND VPWR VPWR _0922_ sky130_fd_sc_hd__a31o_1
XFILLER_0_80_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3777_ cu.reg_file.reg_mem\[13\] _0640_ _0851_ _0852_ VGND VGND VPWR VPWR _0853_
+ sky130_fd_sc_hd__a211oi_2
XFILLER_0_42_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_62 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5455__A _1364_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5516_ _1369_ _2331_ _2332_ _2335_ VGND VGND VPWR VPWR _2336_ sky130_fd_sc_hd__o31a_1
XFILLER_0_14_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_89_95 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5447_ _1417_ _2136_ VGND VGND VPWR VPWR _2275_ sky130_fd_sc_hd__or2_1
XFILLER_0_14_298 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5378_ _2232_ VGND VGND VPWR VPWR _0163_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4329_ _1376_ _1393_ VGND VGND VPWR VPWR _1394_ sky130_fd_sc_hd__or2_1
Xfanout156 net157 VGND VGND VPWR VPWR net156 sky130_fd_sc_hd__clkbuf_4
Xfanout178 net182 VGND VGND VPWR VPWR net178 sky130_fd_sc_hd__clkbuf_2
Xfanout189 net190 VGND VGND VPWR VPWR net189 sky130_fd_sc_hd__clkbuf_4
Xfanout167 net168 VGND VGND VPWR VPWR net167 sky130_fd_sc_hd__clkbuf_4
XFILLER_0_69_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1114 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1103 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_69_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_1147 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1136 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1125 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_84_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5956__A0 cu.id.imm_i\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1169 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1158 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_92_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5708__B1 cu.reg_file.reg_mem\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__2989__A net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_20_257 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_909 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4428__B _1484_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3670__A1 cu.reg_file.reg_a\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_34_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3670__B2 cu.reg_file.reg_mem\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_68_471 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_68_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3700_ _0774_ _0775_ VGND VGND VPWR VPWR _0776_ sky130_fd_sc_hd__nand2_4
X_4680_ net234 _1702_ _1687_ VGND VGND VPWR VPWR _1706_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_55_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3631_ cu.pc.pc_o\[2\] _0501_ _0502_ cu.reg_file.reg_b\[2\] _0536_ VGND VGND VPWR
+ VPWR _0707_ sky130_fd_sc_hd__a221o_1
XFILLER_0_36_390 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3562_ cu.reg_file.reg_sp\[6\] _0636_ _0419_ cu.reg_file.reg_h\[6\] _0637_ VGND VGND
+ VPWR VPWR _0638_ sky130_fd_sc_hd__a221o_1
X_5301_ _1192_ net89 _2182_ VGND VGND VPWR VPWR _2188_ sky130_fd_sc_hd__mux2_1
XFILLER_0_59_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_51_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6281_ clknet_leaf_13_clk _0263_ net180 VGND VGND VPWR VPWR ih.t.timer_max\[21\]
+ sky130_fd_sc_hd__dfrtp_1
X_3493_ _0519_ _0553_ VGND VGND VPWR VPWR _0569_ sky130_fd_sc_hd__or2_1
X_5232_ _1364_ _1631_ VGND VGND VPWR VPWR _2141_ sky130_fd_sc_hd__or2_1
Xclkbuf_leaf_5_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_5_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_11_268 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5163_ cu.reg_file.reg_l\[6\] _1193_ _2088_ VGND VGND VPWR VPWR _2095_ sky130_fd_sc_hd__mux2_1
XFILLER_0_75_31 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4114_ _1089_ VGND VGND VPWR VPWR _1187_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__3523__A _0598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5094_ _2050_ VGND VGND VPWR VPWR _0061_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4989__A1 cu.pc.pc_o\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4045_ _0606_ _0643_ _0663_ _0822_ _1118_ VGND VGND VPWR VPWR _1119_ sky130_fd_sc_hd__a221o_1
XANTENNA__5650__A2 _1648_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5938__A0 _0340_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_482 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5996_ clknet_leaf_0_clk _0034_ net154 VGND VGND VPWR VPWR cu.reg_file.reg_a\[2\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_19_313 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4947_ cu.pc.pc_o\[11\] _1937_ _1814_ VGND VGND VPWR VPWR _1938_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_485 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_74_463 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4878_ _1872_ _1873_ VGND VGND VPWR VPWR _1874_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_46_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3829_ _0871_ _0874_ VGND VGND VPWR VPWR _0905_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5124__S _2069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3101__B1 ih.t.timer_max\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_213 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5641__A2 _1633_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3652__A1 cu.reg_file.reg_l\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_57_419 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_84_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_clkbuf_leaf_34_clk_A clknet_2_1__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4601__B1 _1644_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_143 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5157__A1 _1187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_25_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_80_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_706 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_13 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5823__A cu.reg_file.reg_sp\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_739 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5034__S _2002_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3340__B1 _0415_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3891__B2 _2893_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3891__A1 _2883_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5093__A0 cu.reg_file.reg_d\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xmax_cap1 net237 VGND VGND VPWR VPWR net236 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_61_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5850_ _1624_ _2627_ _2115_ VGND VGND VPWR VPWR _2628_ sky130_fd_sc_hd__mux2_1
XFILLER_0_61_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2993_ _2727_ ih.ih.ih.prev_data\[0\] _2728_ ih.ih.ih.prev_data\[15\] _2731_ VGND
+ VGND VPWR VPWR _2732_ sky130_fd_sc_hd__o221a_1
XANTENNA__5396__A1 net129 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_8_516 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4801_ _2923_ _2899_ _2879_ _0314_ _1802_ VGND VGND VPWR VPWR _1803_ sky130_fd_sc_hd__o311a_1
X_5781_ cu.reg_file.reg_sp\[5\] _2567_ _2539_ VGND VGND VPWR VPWR _2568_ sky130_fd_sc_hd__mux2_1
XFILLER_0_90_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_61_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4732_ cu.alu_f\[6\] alu.Cin _0359_ VGND VGND VPWR VPWR _1741_ sky130_fd_sc_hd__mux2_1
X_4663_ _1693_ _1694_ VGND VGND VPWR VPWR ih.t.next_count\[9\] sky130_fd_sc_hd__nor2_1
XANTENNA__5717__B _2351_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3614_ cu.pc.pc_o\[3\] _0501_ _0502_ cu.reg_file.reg_b\[3\] _0536_ VGND VGND VPWR
+ VPWR _0690_ sky130_fd_sc_hd__a221o_1
X_4594_ _1329_ _1372_ VGND VGND VPWR VPWR _1638_ sky130_fd_sc_hd__nor2_1
XFILLER_0_9_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_3_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3545_ _0464_ _0487_ _0482_ VGND VGND VPWR VPWR _0621_ sky130_fd_sc_hd__o21a_1
X_6264_ clknet_leaf_22_clk _0246_ net191 VGND VGND VPWR VPWR ih.t.timer_max\[12\]
+ sky130_fd_sc_hd__dfrtp_4
X_3476_ _0528_ _0551_ VGND VGND VPWR VPWR _0552_ sky130_fd_sc_hd__nor2_1
XANTENNA__4659__B1 _1687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5215_ _1075_ ih.gpio_interrupt_mask\[2\] _2127_ VGND VGND VPWR VPWR _2130_ sky130_fd_sc_hd__mux2_1
XANTENNA__5320__A1 net96 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6195_ clknet_leaf_4_clk net2 net171 VGND VGND VPWR VPWR ih.ih.ih.prev_data\[0\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_43_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5146_ _2084_ VGND VGND VPWR VPWR _0079_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5084__A0 cu.reg_file.reg_d\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5077_ _2035_ _2038_ _2951_ VGND VGND VPWR VPWR _2039_ sky130_fd_sc_hd__o21a_4
XANTENNA__5623__A2 _2193_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4028_ _0599_ _1101_ _0610_ VGND VGND VPWR VPWR _1102_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_94_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5979_ clknet_leaf_30_clk _0017_ net187 VGND VGND VPWR VPWR cu.pc.pc_o\[1\] sky130_fd_sc_hd__dfrtp_4
XANTENNA__5139__A1 cu.reg_file.reg_h\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4531__B _1579_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4898__A0 cu.pc.pc_o\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4250__C _2923_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_308 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_85_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_15_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_422 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5029__S _2006_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_466 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3338__A _0293_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_263 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output95_A net95 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3330_ _2889_ _2933_ VGND VGND VPWR VPWR _0406_ sky130_fd_sc_hd__or2_1
XFILLER_0_21_396 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_503 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3261_ _0302_ _0303_ _0317_ _0336_ VGND VGND VPWR VPWR _0337_ sky130_fd_sc_hd__o31a_1
XTAP_536 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5000_ cu.reg_file.reg_a\[0\] _1983_ _1985_ VGND VGND VPWR VPWR _1986_ sky130_fd_sc_hd__mux2_1
X_3192_ _2926_ _2928_ VGND VGND VPWR VPWR _2929_ sky130_fd_sc_hd__nor2_1
XTAP_569 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_341 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_88_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5902_ _2658_ VGND VGND VPWR VPWR _0261_ sky130_fd_sc_hd__clkbuf_1
X_5833_ _2611_ _2612_ VGND VGND VPWR VPWR _2613_ sky130_fd_sc_hd__nand2_1
XFILLER_0_91_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_63_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_29_474 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_2976_ net14 VGND VGND VPWR VPWR _2715_ sky130_fd_sc_hd__inv_2
XFILLER_0_56_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5764_ _1089_ _2552_ _2545_ VGND VGND VPWR VPWR _2553_ sky130_fd_sc_hd__mux2_1
XFILLER_0_44_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4715_ ih.t.count\[27\] _1726_ VGND VGND VPWR VPWR _1729_ sky130_fd_sc_hd__and2_1
X_5695_ mc.cl.next_data\[12\] _2359_ _2490_ _2502_ VGND VGND VPWR VPWR _2503_ sky130_fd_sc_hd__o2bb2a_1
XFILLER_0_16_135 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4646_ net219 _1679_ _1682_ VGND VGND VPWR VPWR ih.t.next_count\[4\] sky130_fd_sc_hd__a21oi_1
X_4577_ _2702_ _1192_ _1209_ _2697_ VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__a22o_1
X_6316_ clknet_leaf_36_clk _0002_ net158 VGND VGND VPWR VPWR cu.id.is_interrupted
+ sky130_fd_sc_hd__dfrtp_1
X_3528_ _0447_ _0601_ _0603_ VGND VGND VPWR VPWR _0604_ sky130_fd_sc_hd__mux2_1
X_6247_ clknet_leaf_42_clk _0229_ net151 VGND VGND VPWR VPWR cu.reg_file.reg_sp\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_3459_ cu.reg_file.reg_e\[1\] _0488_ _0502_ cu.reg_file.reg_b\[1\] _0534_ VGND VGND
+ VPWR VPWR _0535_ sky130_fd_sc_hd__a221o_1
X_6178_ clknet_leaf_19_clk _0212_ net184 VGND VGND VPWR VPWR cu.reg_file.reg_mem\[14\]
+ sky130_fd_sc_hd__dfrtp_1
X_5129_ _1226_ _1073_ _2066_ VGND VGND VPWR VPWR _2073_ sky130_fd_sc_hd__mux2_1
XANTENNA__4807__A _1808_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4526__B _1579_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4280__A1 cu.reg_file.reg_c\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_39_238 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_82_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5638__A net90 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_433 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3791__B1 _0624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5532__A1 _2350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_127 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_22_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA_output133_A net133 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5312__S _2195_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5599__B2 _1401_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4271__A1 cu.reg_file.reg_e\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4271__B2 cu.reg_file.reg_l\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_208 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_73_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3068__A ih.t.timer_max\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4574__A2 _1075_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_5480_ _2236_ VGND VGND VPWR VPWR _2302_ sky130_fd_sc_hd__inv_2
X_4500_ _1296_ _1554_ _1555_ VGND VGND VPWR VPWR _1556_ sky130_fd_sc_hd__a21o_1
XFILLER_0_53_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_5_349 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_26_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3782__B1 _0624_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4431_ _1296_ _1487_ _1490_ VGND VGND VPWR VPWR _1491_ sky130_fd_sc_hd__a21o_1
XANTENNA_1 _0560_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_67_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4362_ cu.reg_file.reg_a\[5\] _1276_ _1287_ cu.reg_file.reg_sp\[5\] VGND VGND VPWR
+ VPWR _1425_ sky130_fd_sc_hd__a22o_1
X_6101_ clknet_leaf_26_clk _0135_ net195 VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__dfrtp_4
X_4293_ cu.reg_file.reg_e\[2\] _1283_ _1285_ cu.reg_file.reg_l\[2\] _1358_ VGND VGND
+ VPWR VPWR _1359_ sky130_fd_sc_hd__a221o_1
XTAP_322 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3313_ _0374_ cu.id.cb_opcode_x\[1\] cu.id.cb_opcode_x\[0\] VGND VGND VPWR VPWR _0389_
+ sky130_fd_sc_hd__or3_1
XTAP_300 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3244_ _2884_ net150 _2934_ VGND VGND VPWR VPWR _0320_ sky130_fd_sc_hd__and3b_2
XTAP_355 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6032_ clknet_leaf_3_clk _0070_ net156 VGND VGND VPWR VPWR cu.reg_file.reg_e\[6\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_377 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3175_ _2911_ VGND VGND VPWR VPWR _2912_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_49_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_28 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_88_171 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XPHY_39 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_355 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5211__A0 _0619_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_29_271 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5816_ cu.reg_file.reg_sp\[10\] _2536_ VGND VGND VPWR VPWR _2598_ sky130_fd_sc_hd__nand2_1
X_2959_ mc.rw.state\[0\] mc.rw.state\[2\] _2695_ VGND VGND VPWR VPWR _2700_ sky130_fd_sc_hd__and3b_1
XFILLER_0_8_187 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5762__A1 cu.reg_file.reg_sp\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5747_ _0740_ _2116_ _2537_ _2948_ VGND VGND VPWR VPWR _2538_ sky130_fd_sc_hd__o31a_2
X_5678_ _1489_ _1631_ _1661_ VGND VGND VPWR VPWR _2490_ sky130_fd_sc_hd__or3_2
XANTENNA__5514__A1 net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_32_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4629_ _1669_ VGND VGND VPWR VPWR _1670_ sky130_fd_sc_hd__clkbuf_4
XANTENNA__5514__B2 net62 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3706__A _0545_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5132__S _2066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4971__S _1798_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_63_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3764__B1 _0429_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_211 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_23_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3616__A cu.id.cb_opcode_y\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_277 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput60 net60 VGND VGND VPWR VPWR programmable_gpio_out[0] sky130_fd_sc_hd__buf_2
Xoutput82 net82 VGND VGND VPWR VPWR ss0[6] sky130_fd_sc_hd__clkbuf_4
Xoutput93 net93 VGND VGND VPWR VPWR ss2[1] sky130_fd_sc_hd__clkbuf_4
Xoutput71 net71 VGND VGND VPWR VPWR programmable_gpio_wr[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_37_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5831__A cu.reg_file.reg_sp\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3819__A1 cu.reg_file.reg_mem\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5441__A0 _2022_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4980_ _1943_ _1955_ _1967_ VGND VGND VPWR VPWR _1968_ sky130_fd_sc_hd__or3_1
XFILLER_0_85_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_377 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3931_ _0976_ VGND VGND VPWR VPWR _1007_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_325 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3862_ _0923_ _0937_ VGND VGND VPWR VPWR _0938_ sky130_fd_sc_hd__nand2_1
X_5601_ net80 _1633_ _2413_ _2416_ VGND VGND VPWR VPWR _2417_ sky130_fd_sc_hd__o22a_1
XFILLER_0_5_124 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5532_ cu.reg_file.reg_mem\[0\] _2350_ _2351_ VGND VGND VPWR VPWR _2352_ sky130_fd_sc_hd__mux2_1
XANTENNA__3755__B1 _0429_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3793_ cu.pc.pc_o\[11\] _0740_ _0868_ VGND VGND VPWR VPWR _0869_ sky130_fd_sc_hd__a21o_1
XFILLER_0_81_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_14_425 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_26_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5463_ _2289_ VGND VGND VPWR VPWR _0191_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_41_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4414_ _1463_ _1474_ VGND VGND VPWR VPWR _1475_ sky130_fd_sc_hd__or2_1
X_5394_ _1190_ net128 _2237_ VGND VGND VPWR VPWR _2242_ sky130_fd_sc_hd__mux2_1
X_4345_ _1271_ _1408_ VGND VGND VPWR VPWR _1409_ sky130_fd_sc_hd__nor2_1
XFILLER_0_22_491 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4276_ _0295_ _1318_ VGND VGND VPWR VPWR _1343_ sky130_fd_sc_hd__nor2_2
XANTENNA__4483__A1 _1296_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6015_ clknet_leaf_4_clk _0053_ net173 VGND VGND VPWR VPWR cu.reg_file.reg_c\[5\]
+ sky130_fd_sc_hd__dfrtp_4
X_3227_ _2916_ _2917_ _2919_ VGND VGND VPWR VPWR _0303_ sky130_fd_sc_hd__and3b_2
XTAP_196 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5680__B1 cu.reg_file.reg_mem\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3158_ cu.id.opcode\[2\] cu.id.opcode\[6\] cu.id.opcode\[7\] cu.id.opcode\[1\] VGND
+ VGND VPWR VPWR _2895_ sky130_fd_sc_hd__nor4b_1
XFILLER_0_96_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3089_ _2751_ _2825_ ih.t.count\[8\] VGND VGND VPWR VPWR _2827_ sky130_fd_sc_hd__a21oi_1
XANTENNA__5432__A0 _2022_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5188__A _1646_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_64_303 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_241 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5127__S _2069_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5423__A0 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_95_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5726__A1 net19 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_43_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5037__S _2002_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4130_ _0777_ _0949_ _1197_ _1199_ VGND VGND VPWR VPWR _1200_ sky130_fd_sc_hd__a22o_1
XFILLER_0_48_89 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4465__A1 cu.reg_file.reg_b\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4061_ _1131_ _1134_ _0517_ VGND VGND VPWR VPWR _1135_ sky130_fd_sc_hd__o21a_1
X_3012_ ih.t.timer_max\[5\] ih.t.timer_max\[6\] _2749_ VGND VGND VPWR VPWR _2750_
+ sky130_fd_sc_hd__or3_2
XANTENNA__4465__B2 cu.reg_file.reg_h\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_64_88 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4905__A cu.id.cb_opcode_x\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4963_ _1952_ VGND VGND VPWR VPWR _0028_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_86_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3914_ _2936_ _0386_ _0312_ _0323_ _0984_ VGND VGND VPWR VPWR _0990_ sky130_fd_sc_hd__a2111o_1
X_4894_ _1887_ _1888_ VGND VGND VPWR VPWR _1889_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_46_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_336 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3845_ _0895_ _0892_ VGND VGND VPWR VPWR _0921_ sky130_fd_sc_hd__and2b_1
XFILLER_0_6_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_14_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3776_ cu.reg_file.reg_b\[5\] _0426_ _0429_ cu.reg_file.reg_d\[5\] VGND VGND VPWR
+ VPWR _0852_ sky130_fd_sc_hd__a22o_1
X_5515_ _1374_ _2333_ _2334_ VGND VGND VPWR VPWR _2335_ sky130_fd_sc_hd__or3_1
XFILLER_0_73_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5446_ _1640_ VGND VGND VPWR VPWR _2274_ sky130_fd_sc_hd__buf_2
XFILLER_0_14_277 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5377_ _1192_ net121 _2226_ VGND VGND VPWR VPWR _2232_ sky130_fd_sc_hd__mux2_1
XFILLER_0_1_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_4328_ _1387_ _1388_ _1392_ VGND VGND VPWR VPWR _1393_ sky130_fd_sc_hd__o21a_2
Xfanout179 net180 VGND VGND VPWR VPWR net179 sky130_fd_sc_hd__clkbuf_4
Xfanout168 net169 VGND VGND VPWR VPWR net168 sky130_fd_sc_hd__clkbuf_4
Xfanout157 net163 VGND VGND VPWR VPWR net157 sky130_fd_sc_hd__clkbuf_2
XANTENNA__3703__B _0528_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4087__A _1144_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4259_ cu.reg_file.reg_e\[0\] _1315_ _1317_ cu.reg_file.reg_l\[0\] _1326_ VGND VGND
+ VPWR VPWR _1327_ sky130_fd_sc_hd__a221o_1
XFILLER_0_96_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XTAP_1104 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5405__A0 _0619_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1137 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1126 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1115 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5956__A1 _2372_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_1159 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1148 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_461 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_92_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5708__B2 _1646_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_33_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_542 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_33_564 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5892__A0 _1260_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_clkbuf_leaf_8_clk_A clknet_2_2__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4447__B2 cu.pc.pc_o\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4447__A1 cu.id.imm_i\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_87_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5320__S _2195_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_409 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_314 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_291 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_208 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3630_ cu.alu_f\[2\] _0498_ _0628_ cu.reg_file.reg_mem\[2\] _0705_ VGND VGND VPWR
+ VPWR _0706_ sky130_fd_sc_hd__a221o_1
X_3561_ cu.reg_file.reg_d\[6\] _0415_ _0432_ cu.reg_file.reg_b\[6\] VGND VGND VPWR
+ VPWR _0637_ sky130_fd_sc_hd__a22o_1
XANTENNA__3076__A ih.t.timer_max\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5300_ _2187_ VGND VGND VPWR VPWR _0130_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_51_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6280_ clknet_leaf_13_clk _0262_ net180 VGND VGND VPWR VPWR ih.t.timer_max\[20\]
+ sky130_fd_sc_hd__dfrtp_1
XFILLER_0_11_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3492_ net142 _0532_ _0545_ _0558_ _0567_ VGND VGND VPWR VPWR _0568_ sky130_fd_sc_hd__a221o_1
X_5231_ _1367_ _1625_ _2139_ VGND VGND VPWR VPWR _2140_ sky130_fd_sc_hd__or3_2
X_5162_ _2094_ VGND VGND VPWR VPWR _0085_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5992__RESET_B net161 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5093_ cu.reg_file.reg_d\[5\] _2049_ _2039_ VGND VGND VPWR VPWR _2050_ sky130_fd_sc_hd__mux2_1
X_4113_ _2946_ _2947_ VGND VGND VPWR VPWR _1186_ sky130_fd_sc_hd__or2_2
X_4044_ _1113_ _1117_ VGND VGND VPWR VPWR _1118_ sky130_fd_sc_hd__nor2_1
XANTENNA__4635__A _1672_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5938__A1 _2372_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_59_461 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_46_100 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3949__B1 alu.Cin VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5995_ clknet_leaf_0_clk _0033_ net154 VGND VGND VPWR VPWR cu.reg_file.reg_a\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_74_442 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_59_494 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4946_ _1931_ _1936_ _1808_ VGND VGND VPWR VPWR _1937_ sky130_fd_sc_hd__mux2_1
X_4877_ cu.pc.pc_o\[6\] _1860_ VGND VGND VPWR VPWR _1873_ sky130_fd_sc_hd__nor2_1
X_3828_ _0887_ _0901_ _0903_ VGND VGND VPWR VPWR _0904_ sky130_fd_sc_hd__a21o_1
X_3759_ cu.reg_file.reg_b\[6\] _0743_ _0624_ cu.reg_file.reg_sp\[14\] VGND VGND VPWR
+ VPWR _0835_ sky130_fd_sc_hd__a22o_1
XFILLER_0_42_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5405__S _2248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5429_ _2022_ net70 _2262_ VGND VGND VPWR VPWR _2263_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_280 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3101__A1 ih.t.timer_max\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_84_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4601__A1 _1364_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_464 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3168__A1 _2893_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_40_309 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_33_361 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_406 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_707 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_25 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_729 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3340__A1 cu.reg_file.reg_sp\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3340__B2 cu.reg_file.reg_d\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_501 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_output40_A net40 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5050__S _2006_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_75_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4800_ _2932_ _0330_ VGND VGND VPWR VPWR _1802_ sky130_fd_sc_hd__or2_1
XFILLER_0_0_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_37 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2992_ _2729_ ih.ih.ih.prev_data\[7\] _2730_ ih.ih.ih.prev_data\[8\] VGND VGND VPWR
+ VPWR _2731_ sky130_fd_sc_hd__o22a_1
X_5780_ _1144_ _2566_ _2545_ VGND VGND VPWR VPWR _2567_ sky130_fd_sc_hd__mux2_1
XFILLER_0_83_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_56_475 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4731_ _2946_ _1301_ _1300_ VGND VGND VPWR VPWR _1740_ sky130_fd_sc_hd__a21oi_1
XFILLER_0_8_539 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4662_ net225 _1691_ _1687_ VGND VGND VPWR VPWR _1694_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_71_412 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3613_ cu.alu_f\[3\] _0498_ _0494_ cu.reg_file.reg_mem\[3\] _0688_ VGND VGND VPWR
+ VPWR _0689_ sky130_fd_sc_hd__a221o_1
X_4593_ _1434_ _1635_ VGND VGND VPWR VPWR _1637_ sky130_fd_sc_hd__nand2_1
XFILLER_0_12_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_43_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_51_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3544_ _0377_ _0393_ VGND VGND VPWR VPWR _0620_ sky130_fd_sc_hd__nor2_1
XANTENNA__5733__B mc.cl.next_data\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6263_ clknet_leaf_15_clk _0245_ net179 VGND VGND VPWR VPWR ih.t.timer_max\[11\]
+ sky130_fd_sc_hd__dfrtp_2
XFILLER_0_10_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3475_ _0399_ _0550_ VGND VGND VPWR VPWR _0551_ sky130_fd_sc_hd__nand2_1
X_5214_ _2129_ VGND VGND VPWR VPWR _0102_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5856__A0 _1263_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6194_ clknet_leaf_34_clk net1 net162 VGND VGND VPWR VPWR ih.ip_ed.prev_data sky130_fd_sc_hd__dfrtp_1
XANTENNA__3331__B2 _2877_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout194_A net195 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_36_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5145_ _2083_ cu.reg_file.reg_h\[7\] _2069_ VGND VGND VPWR VPWR _2084_ sky130_fd_sc_hd__mux2_1
X_5076_ _0367_ _2037_ VGND VGND VPWR VPWR _2038_ sky130_fd_sc_hd__and2_1
X_4027_ _1100_ VGND VGND VPWR VPWR _1101_ sky130_fd_sc_hd__inv_2
XFILLER_0_79_545 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5978_ clknet_leaf_29_clk _0016_ net188 VGND VGND VPWR VPWR cu.pc.pc_o\[0\] sky130_fd_sc_hd__dfrtp_1
X_4929_ cu.pc.pc_o\[9\] cu.pc.pc_o\[8\] _1233_ VGND VGND VPWR VPWR _1921_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_34_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5544__C1 _1661_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_353 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5135__S _2066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3322__A1 _0361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4275__A cu.reg_file.reg_l\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_206 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_53_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire141 _2324_ VGND VGND VPWR VPWR net141 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_25_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_25_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_40_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_203 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_40_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output88_A net88 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3561__B2 cu.reg_file.reg_b\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3561__A1 cu.reg_file.reg_d\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_247 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_504 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_515 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3260_ _0335_ VGND VGND VPWR VPWR _0336_ sky130_fd_sc_hd__clkbuf_4
XTAP_526 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3191_ _2888_ _2889_ _2927_ VGND VGND VPWR VPWR _2928_ sky130_fd_sc_hd__and3_1
XTAP_559 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5066__A1 _1191_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_22_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4185__A _0387_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5901_ ih.t.timer_max\[19\] _1187_ _2654_ VGND VGND VPWR VPWR _2658_ sky130_fd_sc_hd__mux2_1
XANTENNA__3589__C_N _0374_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_72_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_76_537 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_29_420 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3845__A_N _0895_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5832_ cu.reg_file.reg_sp\[12\] _2536_ VGND VGND VPWR VPWR _2612_ sky130_fd_sc_hd__nand2_1
X_5763_ _2550_ _2551_ VGND VGND VPWR VPWR _2552_ sky130_fd_sc_hd__xor2_1
XANTENNA__4577__B1 _1209_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4714_ _1728_ VGND VGND VPWR VPWR ih.t.next_count\[26\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_91_529 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2975_ _2709_ ih.ih.ih.prev_data\[1\] _2710_ ih.ih.ih.prev_data\[11\] _2713_ VGND
+ VGND VPWR VPWR _2714_ sky130_fd_sc_hd__o221a_1
XFILLER_0_29_497 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5694_ ih.t.timer_max\[28\] _2151_ _2320_ ih.t.timer_max\[12\] VGND VGND VPWR VPWR
+ _2502_ sky130_fd_sc_hd__a22oi_1
XFILLER_0_44_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4645_ ih.t.count\[4\] _1679_ _1670_ VGND VGND VPWR VPWR _1682_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_71_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_21_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_320 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_128 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4576_ _2702_ _1190_ _1213_ _2697_ VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__a22o_1
X_3527_ _0548_ _0602_ VGND VGND VPWR VPWR _0603_ sky130_fd_sc_hd__nor2_4
X_6315_ clknet_leaf_36_clk _0003_ net158 VGND VGND VPWR VPWR cu.id.starting_int_service
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_12_375 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_397 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5829__A0 cu.reg_file.reg_sp\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6246_ clknet_leaf_42_clk _0228_ net155 VGND VGND VPWR VPWR cu.reg_file.reg_sp\[2\]
+ sky130_fd_sc_hd__dfrtp_4
X_3458_ cu.pc.pc_o\[1\] _0501_ VGND VGND VPWR VPWR _0534_ sky130_fd_sc_hd__and2_1
XANTENNA_clkbuf_leaf_33_clk_A clknet_2_1__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6177_ clknet_leaf_19_clk _0211_ net183 VGND VGND VPWR VPWR cu.reg_file.reg_mem\[13\]
+ sky130_fd_sc_hd__dfrtp_2
X_3389_ _2892_ _2897_ net150 VGND VGND VPWR VPWR _0465_ sky130_fd_sc_hd__and3_1
X_5128_ _2072_ VGND VGND VPWR VPWR _0073_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4095__A _0566_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5059_ _2027_ VGND VGND VPWR VPWR _0049_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5638__B _1330_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_35_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_242 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_445 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__3791__B2 cu.reg_file.reg_sp\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3791__A1 cu.reg_file.reg_b\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2997__B net27 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_15_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_30_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5599__A2 _2205_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output126_A net126 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_58_526 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_504 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_312 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4733__A _2893_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3349__A _0405_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_275 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_106 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3782__B2 cu.reg_file.reg_sp\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3782__A1 cu.reg_file.reg_b\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_2 _0617_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4430_ cu.id.imm_i\[8\] _1294_ _1297_ cu.pc.pc_o\[8\] _1489_ VGND VGND VPWR VPWR
+ _1490_ sky130_fd_sc_hd__a221o_1
XFILLER_0_1_501 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_41_459 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3084__A ih.t.timer_max\[9\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4361_ _1415_ _1416_ _1418_ _1424_ VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__a211o_1
X_6100_ clknet_leaf_20_clk _0134_ net189 VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__dfrtp_4
XFILLER_0_1_556 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_150 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4292_ cu.reg_file.reg_a\[2\] _1276_ _1286_ cu.reg_file.reg_sp\[2\] VGND VGND VPWR
+ VPWR _1358_ sky130_fd_sc_hd__a22o_1
XTAP_323 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3312_ cu.id.cb_opcode_x\[1\] _0387_ VGND VGND VPWR VPWR _0388_ sky130_fd_sc_hd__nand2_1
XTAP_312 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_301 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_21_194 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_3243_ _2892_ _2884_ net150 _2897_ VGND VGND VPWR VPWR _0319_ sky130_fd_sc_hd__o211a_1
XTAP_334 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6031_ clknet_leaf_1_clk _0069_ net154 VGND VGND VPWR VPWR cu.reg_file.reg_e\[5\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_378 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3174_ _2909_ _2910_ VGND VGND VPWR VPWR _2911_ sky130_fd_sc_hd__or2_2
XFILLER_0_83_76 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_83_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_49_559 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5739__A cu.reg_file.reg_sp\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_fanout157_A net163 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5815_ cu.reg_file.reg_sp\[10\] _2536_ VGND VGND VPWR VPWR _2597_ sky130_fd_sc_hd__or2_1
XFILLER_0_76_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_401 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2958_ _2695_ mc.rw.state\[0\] VGND VGND VPWR VPWR _2699_ sky130_fd_sc_hd__nor2_2
XFILLER_0_29_294 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5746_ _0986_ _2532_ _2536_ VGND VGND VPWR VPWR _2537_ sky130_fd_sc_hd__o21ai_1
X_5677_ ih.t.timer_max\[24\] _2151_ _2320_ ih.t.timer_max\[8\] VGND VGND VPWR VPWR
+ _2489_ sky130_fd_sc_hd__a22oi_1
XANTENNA__4970__A0 _1209_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_44_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3773__A1 cu.reg_file.reg_a\[5\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3773__B2 cu.reg_file.reg_mem\[13\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4628_ ih.t.enable _2869_ VGND VGND VPWR VPWR _1669_ sky130_fd_sc_hd__and2_1
XFILLER_0_4_350 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_448 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4559_ cu.pc.pc_o\[15\] _1321_ _1314_ cu.reg_file.reg_d\[7\] _1611_ VGND VGND VPWR
+ VPWR _1612_ sky130_fd_sc_hd__a221o_1
X_6229_ clknet_leaf_14_clk ih.t.next_count\[17\] net177 VGND VGND VPWR VPWR ih.t.count\[17\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__4818__A _0343_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5413__S _2248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_890 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3441__B _0516_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_86_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_334 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5450__A1 net68 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5450__B2 net69 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3764__B2 cu.reg_file.reg_d\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3764__A1 cu.reg_file.reg_b\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_35_297 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__3516__A1 cu.reg_file.reg_b\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_289 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3516__B2 cu.reg_file.reg_a\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
Xoutput61 net61 VGND VGND VPWR VPWR programmable_gpio_out[1] sky130_fd_sc_hd__clkbuf_4
Xoutput50 net50 VGND VGND VPWR VPWR memory_address_out[9] sky130_fd_sc_hd__clkbuf_4
Xoutput94 net94 VGND VGND VPWR VPWR ss2[2] sky130_fd_sc_hd__clkbuf_4
Xoutput72 net72 VGND VGND VPWR VPWR programmable_gpio_wr[4] sky130_fd_sc_hd__buf_2
Xoutput83 net83 VGND VGND VPWR VPWR ss0[7] sky130_fd_sc_hd__buf_2
XANTENNA__4728__A _1672_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5550__C _1661_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3819__A2 _0640_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_37_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4492__A2 _1530_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5441__A1 net74 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3930_ _0999_ _0997_ _1005_ VGND VGND VPWR VPWR _1006_ sky130_fd_sc_hd__o21ai_1
XFILLER_0_58_389 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_529 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3861_ _0887_ _0922_ VGND VGND VPWR VPWR _0937_ sky130_fd_sc_hd__nand2_1
XFILLER_0_73_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5600_ net112 _2147_ _2225_ net120 _2415_ VGND VGND VPWR VPWR _2416_ sky130_fd_sc_hd__a221o_1
X_3792_ cu.reg_file.reg_d\[3\] _0488_ _0741_ cu.reg_file.reg_h\[3\] _0867_ VGND VGND
+ VPWR VPWR _0868_ sky130_fd_sc_hd__a221o_1
XFILLER_0_54_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4952__A0 _1213_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_253 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__3755__B2 cu.reg_file.reg_d\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5531_ _1739_ VGND VGND VPWR VPWR _2351_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_5_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_14_437 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_41_201 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5462_ net61 _2085_ _2288_ VGND VGND VPWR VPWR _2289_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_43 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4413_ _1332_ _1473_ VGND VGND VPWR VPWR _1474_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_68_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5393_ _2241_ VGND VGND VPWR VPWR _0169_ sky130_fd_sc_hd__clkbuf_1
X_4344_ cu.reg_file.reg_c\[4\] _1281_ _1407_ VGND VGND VPWR VPWR _1408_ sky130_fd_sc_hd__a21oi_1
XANTENNA__3542__A _0617_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4275_ cu.reg_file.reg_l\[1\] _1317_ VGND VGND VPWR VPWR _1342_ sky130_fd_sc_hd__and2_1
X_6014_ clknet_leaf_3_clk _0052_ net156 VGND VGND VPWR VPWR cu.reg_file.reg_c\[4\]
+ sky130_fd_sc_hd__dfrtp_4
XTAP_197 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3226_ _0300_ _0301_ VGND VGND VPWR VPWR _0302_ sky130_fd_sc_hd__nor2_1
X_3157_ cu.id.opcode\[0\] VGND VGND VPWR VPWR _2894_ sky130_fd_sc_hd__buf_4
XFILLER_0_27_80 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_96_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3088_ ih.t.count\[8\] _2751_ _2825_ VGND VGND VPWR VPWR _2826_ sky130_fd_sc_hd__and3_1
XANTENNA__5432__A1 net71 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_323 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_301 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_367 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_345 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_64_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_220 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5729_ _2518_ mc.cl.next_data\[3\] _2111_ VGND VGND VPWR VPWR _2525_ sky130_fd_sc_hd__and3_1
XFILLER_0_91_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_72_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_17_286 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_32_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_60_554 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_32_267 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5671__B2 net8 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5671__A1 net15 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5423__A1 _2085_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4283__A _1335_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_142 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_67_175 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_67_186 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_82_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_70_318 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_36_562 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5318__S _2195_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_63_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_23_256 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_11_418 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_output70_A net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_48_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4060_ _1120_ _0773_ _1132_ _1133_ VGND VGND VPWR VPWR _1134_ sky130_fd_sc_hd__a31o_1
X_3011_ _2748_ VGND VGND VPWR VPWR _2749_ sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__5662__B2 ih.t.timer_max\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_407 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3673__B1 _0748_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5289__A _1364_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4905__B cu.pc.pc_o\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4962_ cu.pc.pc_o\[12\] _1951_ _1814_ VGND VGND VPWR VPWR _1952_ sky130_fd_sc_hd__mux2_1
X_4893_ _1875_ _1878_ _1876_ VGND VGND VPWR VPWR _1888_ sky130_fd_sc_hd__o21a_1
XFILLER_0_46_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_46_304 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3913_ _0966_ _0971_ _0987_ _0988_ _0296_ VGND VGND VPWR VPWR _0989_ sky130_fd_sc_hd__a41o_2
XFILLER_0_46_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3844_ _0747_ _0751_ VGND VGND VPWR VPWR _0920_ sky130_fd_sc_hd__or2b_1
XFILLER_0_73_178 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_434 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3775_ cu.reg_file.reg_sp\[13\] _0636_ _0748_ cu.reg_file.reg_h\[5\] VGND VGND VPWR
+ VPWR _0851_ sky130_fd_sc_hd__a22o_1
XFILLER_0_89_75 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5514_ net63 _1638_ _2279_ net62 VGND VGND VPWR VPWR _2334_ sky130_fd_sc_hd__a22o_1
XFILLER_0_54_392 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_489 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_565 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_89_86 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5445_ _2273_ VGND VGND VPWR VPWR _0189_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__5350__A0 _1052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_66_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5752__A cu.reg_file.reg_sp\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5376_ _2231_ VGND VGND VPWR VPWR _0162_ sky130_fd_sc_hd__clkbuf_1
X_4327_ cu.reg_file.reg_c\[3\] _1313_ _1389_ _1391_ VGND VGND VPWR VPWR _1392_ sky130_fd_sc_hd__a211o_1
Xfanout169 net182 VGND VGND VPWR VPWR net169 sky130_fd_sc_hd__clkbuf_2
Xfanout158 net160 VGND VGND VPWR VPWR net158 sky130_fd_sc_hd__clkbuf_4
XANTENNA__4087__B _1160_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5102__B1 _2951_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4258_ cu.reg_file.reg_sp\[0\] _0993_ _1322_ _1299_ _1325_ VGND VGND VPWR VPWR _1326_
+ sky130_fd_sc_hd__a221o_1
X_3209_ cu.id.state\[2\] VGND VGND VPWR VPWR _2946_ sky130_fd_sc_hd__inv_2
X_4189_ _1194_ _1258_ _1027_ VGND VGND VPWR VPWR _1259_ sky130_fd_sc_hd__mux2_1
XTAP_1105 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__5405__A1 net132 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_96_259 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_1138 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1127 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1116 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1149 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_77_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_315 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_37_337 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4550__B _1598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5138__S _2066_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3447__A _0373_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4392__A1 cu.reg_file.reg_c\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5341__A0 _1192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_18_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_87_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_68_440 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_95_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_476 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_55_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_28_359 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_83_498 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5580__B1 _2225_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3560_ _0413_ VGND VGND VPWR VPWR _0636_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_51_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_215 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5230_ _2138_ VGND VGND VPWR VPWR _2139_ sky130_fd_sc_hd__buf_2
XANTENNA__5572__A _1649_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3491_ _0566_ _0547_ _0550_ VGND VGND VPWR VPWR _0567_ sky130_fd_sc_hd__and3_1
X_5161_ cu.reg_file.reg_l\[5\] _1191_ _2088_ VGND VGND VPWR VPWR _2094_ sky130_fd_sc_hd__mux2_1
XANTENNA__3477__B_N _0528_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5092_ _1191_ _1209_ _2035_ VGND VGND VPWR VPWR _2049_ sky130_fd_sc_hd__mux2_1
X_4112_ _1027_ _1075_ _1183_ _1185_ VGND VGND VPWR VPWR _0009_ sky130_fd_sc_hd__o22a_1
XFILLER_0_75_66 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4043_ _0588_ _1059_ VGND VGND VPWR VPWR _1117_ sky130_fd_sc_hd__or2_1
XANTENNA__3820__A _0892_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_78_204 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_91_54 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_78_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5994_ clknet_leaf_0_clk _0032_ net154 VGND VGND VPWR VPWR cu.reg_file.reg_a\[0\]
+ sky130_fd_sc_hd__dfrtp_4
XFILLER_0_93_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_91_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4354__C _1417_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_473 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4945_ _1934_ _1935_ _1798_ VGND VGND VPWR VPWR _1936_ sky130_fd_sc_hd__mux2_1
XFILLER_0_74_421 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4876_ cu.pc.pc_o\[6\] _1860_ VGND VGND VPWR VPWR _1872_ sky130_fd_sc_hd__and2_1
XFILLER_0_61_104 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_253 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_27_381 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3827_ _0902_ _0885_ VGND VGND VPWR VPWR _0903_ sky130_fd_sc_hd__nor2_1
XFILLER_0_61_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3758_ cu.reg_file.reg_d\[6\] _0488_ _0741_ cu.reg_file.reg_h\[6\] VGND VGND VPWR
+ VPWR _0834_ sky130_fd_sc_hd__a22o_1
X_3689_ _0761_ _0764_ VGND VGND VPWR VPWR _0765_ sky130_fd_sc_hd__nor2_1
X_5428_ _2139_ _2194_ VGND VGND VPWR VPWR _2262_ sky130_fd_sc_hd__nand2_1
XFILLER_0_30_568 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5359_ _2221_ VGND VGND VPWR VPWR _0155_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3885__B1 _0773_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5626__A1 _1666_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4826__A _1299_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3101__A2 ih.t.timer_max\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4545__B _1598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_69_248 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_77_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4601__A2 _1489_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_402 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_25_307 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_80_435 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_52_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5562__B1 _2204_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_468 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__5314__A0 _1052_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3905__A _0350_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_0_429 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5865__A1 ih.t.timer_max\[10\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_719 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_708 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_37 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__3340__A2 _0413_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__2999__A_N net70 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5617__A1 net97 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5331__S _2206_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_88_513 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_557 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_61_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_2991_ net16 VGND VGND VPWR VPWR _2730_ sky130_fd_sc_hd__inv_2
XFILLER_0_28_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4730_ _1364_ _1489_ _1644_ VGND VGND VPWR VPWR _1739_ sky130_fd_sc_hd__a21oi_4
X_4661_ ih.t.count\[8\] ih.t.count\[9\] _1689_ VGND VGND VPWR VPWR _1693_ sky130_fd_sc_hd__and3_1
XFILLER_0_83_262 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_71_424 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3612_ cu.reg_file.reg_h\[3\] _0495_ _0499_ cu.reg_file.reg_a\[3\] VGND VGND VPWR
+ VPWR _0688_ sky130_fd_sc_hd__a22o_1
X_4592_ _1434_ _1629_ _1635_ VGND VGND VPWR VPWR _1636_ sky130_fd_sc_hd__or3b_2
XFILLER_0_3_212 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_362 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3543_ _0618_ VGND VGND VPWR VPWR _0619_ sky130_fd_sc_hd__buf_4
X_6262_ clknet_leaf_15_clk _0244_ net179 VGND VGND VPWR VPWR ih.t.timer_max\[10\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__5305__A0 _1261_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3474_ _0392_ _0384_ VGND VGND VPWR VPWR _0550_ sky130_fd_sc_hd__and2b_1
XANTENNA__4101__A1_N _0918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6193_ clknet_leaf_20_clk _0226_ net190 VGND VGND VPWR VPWR mc.cl.next_data\[7\]
+ sky130_fd_sc_hd__dfrtp_1
X_5213_ _1052_ ih.gpio_interrupt_mask\[1\] _2127_ VGND VGND VPWR VPWR _2129_ sky130_fd_sc_hd__mux2_1
XFILLER_0_86_98 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5144_ _1263_ _1110_ _2066_ VGND VGND VPWR VPWR _2083_ sky130_fd_sc_hd__mux2_1
XFILLER_0_19_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_fanout187_A net188 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5075_ _0352_ _1790_ VGND VGND VPWR VPWR _2037_ sky130_fd_sc_hd__and2b_1
X_4026_ _1060_ _0588_ VGND VGND VPWR VPWR _1100_ sky130_fd_sc_hd__or2_1
XFILLER_0_79_557 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4292__B1 _1286_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_281 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_47_432 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_19_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5977_ clknet_leaf_35_clk _0014_ net159 VGND VGND VPWR VPWR cu.alu_f\[7\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_74_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4928_ _1918_ _1919_ VGND VGND VPWR VPWR _1920_ sky130_fd_sc_hd__nand2_1
XFILLER_0_47_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3398__A2 _2878_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_19_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_34_115 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_4859_ _1855_ _1856_ _1799_ VGND VGND VPWR VPWR _1857_ sky130_fd_sc_hd__mux2_1
XANTENNA_clkbuf_leaf_7_clk_A clknet_2_2__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_343 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_30_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_42_192 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_30_398 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_15_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_505 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_57_218 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_38_410 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_38_443 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_38_465 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_446 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5326__S _2195_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3635__A _0587_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3561__A2 _0415_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_505 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_516 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_527 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3190_ _2902_ cu.id.alu_opcode\[3\] VGND VGND VPWR VPWR _2927_ sky130_fd_sc_hd__nor2_1
X_5900_ _2657_ VGND VGND VPWR VPWR _0260_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_72_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_76_549 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_5831_ cu.reg_file.reg_sp\[12\] _2536_ VGND VGND VPWR VPWR _2611_ sky130_fd_sc_hd__or2_1
X_2974_ _2711_ ih.ih.ih.prev_data\[2\] _2712_ ih.ih.ih.prev_data\[3\] VGND VGND VPWR
+ VPWR _2713_ sky130_fd_sc_hd__o22a_1
XFILLER_0_8_326 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_5762_ cu.reg_file.reg_sp\[1\] _2543_ _2541_ VGND VGND VPWR VPWR _2551_ sky130_fd_sc_hd__a21bo_1
XANTENNA__4577__B2 _2697_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4577__A1 _2702_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4713_ _1726_ _1727_ _1669_ VGND VGND VPWR VPWR _1728_ sky130_fd_sc_hd__and3b_1
XFILLER_0_44_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5693_ net4 _1650_ _2488_ _2501_ VGND VGND VPWR VPWR _0209_ sky130_fd_sc_hd__a31o_1
X_4644_ _1681_ VGND VGND VPWR VPWR ih.t.next_count\[3\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_71_287 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_21_93 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_24_170 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_4575_ _2702_ _1188_ _1222_ _2697_ VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__a22o_1
XANTENNA__5236__S _1667_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_332 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3526_ _0519_ _0555_ VGND VGND VPWR VPWR _0602_ sky130_fd_sc_hd__or2b_2
X_6314_ clknet_leaf_36_clk net200 net160 VGND VGND VPWR VPWR cu.id.is_halted sky130_fd_sc_hd__dfrtp_1
XFILLER_0_12_365 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_6245_ clknet_leaf_2_clk _0227_ net155 VGND VGND VPWR VPWR cu.reg_file.reg_sp\[1\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__5760__A cu.reg_file.reg_sp\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3457_ _0464_ _0487_ _0482_ cu.reg_file.reg_l\[1\] VGND VGND VPWR VPWR _0533_ sky130_fd_sc_hd__o211a_1
X_6176_ clknet_leaf_19_clk _0210_ net185 VGND VGND VPWR VPWR cu.reg_file.reg_mem\[12\]
+ sky130_fd_sc_hd__dfrtp_4
XANTENNA__4501__A1 cu.pc.pc_o\[12\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3388_ _0458_ _0463_ VGND VGND VPWR VPWR _0464_ sky130_fd_sc_hd__nor2_2
X_5127_ _2071_ cu.reg_file.reg_h\[1\] _2069_ VGND VGND VPWR VPWR _2072_ sky130_fd_sc_hd__mux2_1
X_5058_ cu.reg_file.reg_c\[1\] _1051_ _2025_ VGND VGND VPWR VPWR _2027_ sky130_fd_sc_hd__mux2_1
X_4009_ _0600_ _1041_ VGND VGND VPWR VPWR _1083_ sky130_fd_sc_hd__nor2_1
XANTENNA__4095__B _1110_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_376 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_79_354 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_207 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_79_387 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4568__B2 _1614_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_47_240 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5765__A0 cu.reg_file.reg_sp\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_35_413 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_62_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_50_416 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3791__A2 _0743_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4740__A1 _2908_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4985__S _1808_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_89_118 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_107 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA_output119_A net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_85_324 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_42_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4559__A1 cu.pc.pc_o\[15\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4559__B2 cu.reg_file.reg_d\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5756__A0 _1073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_541 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_53_243 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3782__A2 _0743_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_405 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA_3 _1188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4360_ _1351_ _1422_ _1423_ VGND VGND VPWR VPWR _1424_ sky130_fd_sc_hd__and3_1
XFILLER_0_6_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3311_ cu.id.cb_opcode_x\[0\] VGND VGND VPWR VPWR _0387_ sky130_fd_sc_hd__buf_4
X_4291_ _1350_ _1352_ _1353_ _1354_ _1357_ VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__a221o_4
XTAP_324 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_302 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6030_ clknet_leaf_1_clk _0068_ net153 VGND VGND VPWR VPWR cu.reg_file.reg_e\[4\]
+ sky130_fd_sc_hd__dfrtp_4
X_3242_ _2938_ _2931_ VGND VGND VPWR VPWR _0318_ sky130_fd_sc_hd__nor2_1
XTAP_335 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3173_ _2900_ _2899_ VGND VGND VPWR VPWR _2910_ sky130_fd_sc_hd__or2b_1
XTAP_368 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_83_33 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_49_505 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_88_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__5747__B1 _2948_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5814_ _2596_ VGND VGND VPWR VPWR _0235_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_64_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_123 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_91_349 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_2957_ mc.rw.state\[2\] VGND VGND VPWR VPWR _2698_ sky130_fd_sc_hd__inv_2
XFILLER_0_32_81 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5745_ _2535_ VGND VGND VPWR VPWR _2536_ sky130_fd_sc_hd__buf_2
XFILLER_0_44_210 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_44_221 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5676_ _1641_ _2344_ VGND VGND VPWR VPWR _2488_ sky130_fd_sc_hd__nor2_2
XFILLER_0_17_479 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_44_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4627_ _2706_ _1664_ _1668_ _1647_ _1371_ VGND VGND VPWR VPWR mc.rw.next_state\[2\]
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_44_276 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4558_ cu.reg_file.reg_sp\[15\] _0992_ _1343_ cu.id.imm_i\[15\] _1323_ VGND VGND
+ VPWR VPWR _1611_ sky130_fd_sc_hd__a221o_1
X_4489_ _1333_ _1545_ VGND VGND VPWR VPWR _1546_ sky130_fd_sc_hd__or2_1
XFILLER_0_12_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3509_ _0582_ _0584_ VGND VGND VPWR VPWR _0585_ sky130_fd_sc_hd__nand2_1
X_6228_ clknet_leaf_11_clk ih.t.next_count\[16\] net177 VGND VGND VPWR VPWR ih.t.count\[16\]
+ sky130_fd_sc_hd__dfrtp_2
XTAP_880 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_6159_ clknet_leaf_18_clk _0193_ net172 VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__dfrtp_4
XANTENNA__4818__B _1299_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_891 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_79_140 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xclkbuf_leaf_37_clk clknet_2_1__leaf_clk VGND VGND VPWR VPWR clknet_leaf_37_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__3461__A1 cu.reg_file.reg_c\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_327 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_82_338 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_12_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_23_405 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3764__A2 _0426_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3185__A _2920_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_23_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_31_460 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput51 net51 VGND VGND VPWR VPWR memory_data_out[0] sky130_fd_sc_hd__clkbuf_4
Xoutput40 net40 VGND VGND VPWR VPWR memory_address_out[14] sky130_fd_sc_hd__buf_2
Xoutput84 net84 VGND VGND VPWR VPWR ss1[0] sky130_fd_sc_hd__clkbuf_4
Xoutput73 net73 VGND VGND VPWR VPWR programmable_gpio_wr[5] sky130_fd_sc_hd__buf_2
Xoutput62 net62 VGND VGND VPWR VPWR programmable_gpio_out[2] sky130_fd_sc_hd__clkbuf_4
Xoutput95 net95 VGND VGND VPWR VPWR ss2[3] sky130_fd_sc_hd__clkbuf_4
Xclkbuf_leaf_28_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_28_clk sky130_fd_sc_hd__clkbuf_16
XFILLER_0_58_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_85_176 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_3860_ _0813_ _0935_ VGND VGND VPWR VPWR _0936_ sky130_fd_sc_hd__or2b_1
XFILLER_0_54_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_clkbuf_leaf_32_clk_A clknet_2_1__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3791_ cu.reg_file.reg_b\[3\] _0743_ _0624_ cu.reg_file.reg_sp\[11\] VGND VGND VPWR
+ VPWR _0867_ sky130_fd_sc_hd__a22o_1
XPHY_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5530_ _2329_ _2330_ _2343_ _2349_ VGND VGND VPWR VPWR _2350_ sky130_fd_sc_hd__o31a_4
XFILLER_0_54_541 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3755__A2 _0426_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_81_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5461_ _2287_ _2284_ VGND VGND VPWR VPWR _2288_ sky130_fd_sc_hd__nor2_1
X_4412_ _1467_ _1468_ _1472_ VGND VGND VPWR VPWR _1473_ sky130_fd_sc_hd__o21ai_4
XFILLER_0_41_246 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_78_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5392_ _1188_ net127 _2237_ VGND VGND VPWR VPWR _2241_ sky130_fd_sc_hd__mux2_1
XFILLER_0_78_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4343_ cu.reg_file.reg_e\[4\] _1283_ _1285_ cu.reg_file.reg_l\[4\] _1406_ VGND VGND
+ VPWR VPWR _1407_ sky130_fd_sc_hd__a221o_1
X_4274_ _0340_ _1295_ _1298_ cu.pc.pc_o\[1\] _1305_ VGND VGND VPWR VPWR _1341_ sky130_fd_sc_hd__a221o_1
XANTENNA__5665__C1 _1660_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6013_ clknet_leaf_4_clk _0051_ net170 VGND VGND VPWR VPWR cu.reg_file.reg_c\[3\]
+ sky130_fd_sc_hd__dfrtp_4
X_3225_ _2876_ _2875_ VGND VGND VPWR VPWR _0301_ sky130_fd_sc_hd__nand2b_4
XTAP_198 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_3156_ _2892_ VGND VGND VPWR VPWR _2893_ sky130_fd_sc_hd__clkbuf_4
X_3087_ ih.t.timer_max\[7\] _2750_ ih.t.timer_max\[8\] VGND VGND VPWR VPWR _2825_
+ sky130_fd_sc_hd__o21ai_1
Xclkbuf_leaf_19_clk clknet_2_3__leaf_clk VGND VGND VPWR VPWR clknet_leaf_19_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__5469__B _2284_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4373__B _1434_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_335 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_91_102 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_76_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3708__A_N _0710_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5728_ net20 _2519_ _2524_ VGND VGND VPWR VPWR _0221_ sky130_fd_sc_hd__a21o_1
X_3989_ _0558_ _0694_ _0822_ _0545_ _1062_ VGND VGND VPWR VPWR _1063_ sky130_fd_sc_hd__a221o_1
XFILLER_0_17_254 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_60_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3717__B _0663_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5659_ net107 _2204_ _2471_ _1401_ VGND VGND VPWR VPWR _2472_ sky130_fd_sc_hd__a22o_1
XFILLER_0_20_408 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4829__A _0341_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_67_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_67_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_23_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_28_508 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_36_530 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3908__A _2918_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_51_522 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_63_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4698__B1 _1687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3643__A _0652_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_31_290 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__4458__B _1511_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output63_A net63 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_3_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5111__A1 _1189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3010_ ih.t.timer_max\[4\] _2747_ VGND VGND VPWR VPWR _2748_ sky130_fd_sc_hd__or2_1
XANTENNA__3673__A1 cu.reg_file.reg_sp\[8\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3673__B2 cu.reg_file.reg_h\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4961_ _1941_ _1950_ _1808_ VGND VGND VPWR VPWR _1951_ sky130_fd_sc_hd__mux2_1
X_4892_ _1885_ _1886_ VGND VGND VPWR VPWR _1887_ sky130_fd_sc_hd__and2b_1
X_3912_ _2936_ _2881_ _0469_ VGND VGND VPWR VPWR _0988_ sky130_fd_sc_hd__o21a_1
XFILLER_0_19_519 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_3843_ _0832_ VGND VGND VPWR VPWR _0919_ sky130_fd_sc_hd__inv_2
XFILLER_0_73_157 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_89_32 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_13_94 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_3774_ cu.id.imm_i\[13\] _0739_ _0849_ _0653_ VGND VGND VPWR VPWR _0850_ sky130_fd_sc_hd__a22oi_4
XFILLER_0_81_190 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5513_ net60 _2277_ _2179_ net61 VGND VGND VPWR VPWR _2333_ sky130_fd_sc_hd__a22o_1
XFILLER_0_14_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_42_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5444_ _2022_ net75 _2272_ VGND VGND VPWR VPWR _2273_ sky130_fd_sc_hd__mux2_1
Xclkbuf_leaf_8_clk clknet_2_2__leaf_clk VGND VGND VPWR VPWR clknet_leaf_8_clk sky130_fd_sc_hd__clkbuf_16
XANTENNA__4689__B1 _1687_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5375_ _1190_ net120 _2226_ VGND VGND VPWR VPWR _2231_ sky130_fd_sc_hd__mux2_1
X_4326_ cu.pc.pc_o\[3\] _1322_ _1315_ cu.reg_file.reg_e\[3\] _1390_ VGND VGND VPWR
+ VPWR _1391_ sky130_fd_sc_hd__a221o_1
Xfanout159 net160 VGND VGND VPWR VPWR net159 sky130_fd_sc_hd__clkbuf_4
XANTENNA__5102__A1 _2035_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4257_ _0343_ _2950_ _1319_ _1324_ VGND VGND VPWR VPWR _1325_ sky130_fd_sc_hd__a31o_1
X_3208_ _2907_ _2915_ _2930_ _2944_ VGND VGND VPWR VPWR _2945_ sky130_fd_sc_hd__o211ai_1
X_4188_ cu.alu_f\[6\] _1256_ _1257_ VGND VGND VPWR VPWR _1258_ sky130_fd_sc_hd__mux2_1
XFILLER_0_38_91 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4861__A0 cu.pc.pc_o\[4\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3139_ cu.id.opcode\[7\] VGND VGND VPWR VPWR _2876_ sky130_fd_sc_hd__clkbuf_4
XFILLER_0_96_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_96_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_1128 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1117 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_1106 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_89_290 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_1139 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_49_154 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_37_305 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_92_477 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__5419__S _2248_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_52_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_382 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_45_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3447__B cu.id.cb_opcode_y\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5341__A1 net105 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_216 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__6196__D net9 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4993__S _1798_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_68_452 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_output101_A net101 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_55_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_55_146 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XANTENNA__4368__C1 _1364_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5580__B2 net119 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5580__A1 net111 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_24_533 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__3357__B _0405_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_449 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3490_ _0560_ _0562_ _0564_ _0565_ VGND VGND VPWR VPWR _0566_ sky130_fd_sc_hd__o31a_4
XANTENNA__5853__A cu.reg_file.reg_sp\[14\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_59_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5160_ _2093_ VGND VGND VPWR VPWR _0084_ sky130_fd_sc_hd__clkbuf_1
X_5091_ _2048_ VGND VGND VPWR VPWR _0060_ sky130_fd_sc_hd__clkbuf_1
X_4111_ cu.alu_f\[2\] _1184_ _0370_ VGND VGND VPWR VPWR _1185_ sky130_fd_sc_hd__a21o_1
XANTENNA__5096__A0 cu.reg_file.reg_d\[6\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4042_ _0531_ _0632_ _0566_ _0558_ VGND VGND VPWR VPWR _1116_ sky130_fd_sc_hd__a2bb2o_1
XANTENNA__3646__A1 _0652_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_91_44 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_59_441 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5993_ clknet_leaf_33_clk _0031_ net161 VGND VGND VPWR VPWR cu.pc.pc_o\[15\] sky130_fd_sc_hd__dfrtp_4
X_4944_ _1222_ _1931_ _1794_ VGND VGND VPWR VPWR _1935_ sky130_fd_sc_hd__mux2_1
XFILLER_0_46_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_74_455 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4875_ _1871_ VGND VGND VPWR VPWR _0021_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_74_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3826_ _0882_ VGND VGND VPWR VPWR _0902_ sky130_fd_sc_hd__inv_2
XANTENNA__5020__A0 _1260_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_34_319 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5571__B2 net3 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5571__A1 net10 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_265 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_27_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3757_ _0829_ _0832_ VGND VGND VPWR VPWR _0833_ sky130_fd_sc_hd__xnor2_4
XANTENNA__3582__B1 _0499_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3688_ _0716_ _0763_ VGND VGND VPWR VPWR _0764_ sky130_fd_sc_hd__xnor2_1
XFILLER_0_30_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
X_5427_ _2261_ VGND VGND VPWR VPWR _0183_ sky130_fd_sc_hd__clkbuf_1
X_5358_ _1192_ net113 _2215_ VGND VGND VPWR VPWR _2221_ sky130_fd_sc_hd__mux2_1
XFILLER_0_10_260 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4309_ _1371_ _1372_ _1374_ VGND VGND VPWR VPWR _1375_ sky130_fd_sc_hd__a21o_1
XANTENNA__5087__A0 cu.reg_file.reg_d\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5289_ _1364_ _2169_ VGND VGND VPWR VPWR _2181_ sky130_fd_sc_hd__nor2_8
XANTENNA__4826__B cu.pc.pc_o\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4834__A0 _1073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__6036__RESET_B net188 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4842__A cu.id.cb_opcode_y\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_77_293 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3458__A cu.pc.pc_o\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_499 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_18_360 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5011__A0 _1189_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_20_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_33_385 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4565__C_N _1598_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5314__A1 net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_709 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_29_49 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5078__A0 cu.reg_file.reg_d\[0\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5617__A2 _2194_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_45_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_88_525 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_88_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_61_36 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_2990_ net15 VGND VGND VPWR VPWR _2729_ sky130_fd_sc_hd__inv_2
XFILLER_0_61_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4660_ _1691_ _1692_ VGND VGND VPWR VPWR ih.t.next_count\[8\] sky130_fd_sc_hd__nor2_1
XFILLER_0_83_274 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_56_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5002__A0 _1051_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_9_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_3611_ cu.reg_file.reg_c\[3\] _0485_ _0489_ cu.reg_file.reg_e\[3\] _0686_ VGND VGND
+ VPWR VPWR _0687_ sky130_fd_sc_hd__a221o_1
X_4591_ _1455_ _1473_ VGND VGND VPWR VPWR _1635_ sky130_fd_sc_hd__nor2_1
X_3542_ _0617_ VGND VGND VPWR VPWR _0618_ sky130_fd_sc_hd__buf_4
XANTENNA__3919__A_N _0986_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_12_547 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_24_374 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
X_6261_ clknet_leaf_15_clk _0243_ net179 VGND VGND VPWR VPWR ih.t.timer_max\[9\] sky130_fd_sc_hd__dfstp_1
XANTENNA__4583__D_N _1614_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__5305__A1 net91 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3473_ _0548_ _0393_ VGND VGND VPWR VPWR _0549_ sky130_fd_sc_hd__nor2_1
X_6192_ clknet_leaf_22_clk _0225_ net191 VGND VGND VPWR VPWR mc.cl.next_data\[6\]
+ sky130_fd_sc_hd__dfrtp_1
X_5212_ _2128_ VGND VGND VPWR VPWR _0101_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__3316__B1 _2950_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5143_ _2082_ VGND VGND VPWR VPWR _0078_ sky130_fd_sc_hd__clkbuf_1
XANTENNA__4927__A _2920_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5074_ _0617_ _1622_ _2035_ VGND VGND VPWR VPWR _2036_ sky130_fd_sc_hd__mux2_1
XFILLER_0_79_503 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__4292__A1 cu.reg_file.reg_a\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4025_ _1092_ _1098_ _1069_ VGND VGND VPWR VPWR _1099_ sky130_fd_sc_hd__a21oi_1
XANTENNA__4292__B2 cu.reg_file.reg_sp\[2\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_79_569 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_47_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5976_ clknet_leaf_35_clk _0013_ net159 VGND VGND VPWR VPWR cu.alu_f\[6\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_19_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5477__B _2284_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4927_ _2920_ _1521_ VGND VGND VPWR VPWR _1919_ sky130_fd_sc_hd__nand2_1
XANTENNA__3278__A _2883_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_62_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4858_ _1160_ _1850_ _1795_ VGND VGND VPWR VPWR _1856_ sky130_fd_sc_hd__mux2_1
X_3809_ cu.reg_file.reg_mem\[10\] _0640_ _0883_ _0884_ VGND VGND VPWR VPWR _0885_
+ sky130_fd_sc_hd__a211oi_2
XANTENNA__5544__B2 ih.t.timer_max\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3555__B1 _0536_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4789_ _0350_ _0358_ VGND VGND VPWR VPWR _1791_ sky130_fd_sc_hd__nor2_1
XFILLER_0_30_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_85_517 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XANTENNA__4572__A _0516_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_93_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_31_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_38_477 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4338__A2 _1401_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_80_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5535__A1 net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_65_296 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_65_285 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_53_458 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xwire143 _1280_ VGND VGND VPWR VPWR net143 sky130_fd_sc_hd__clkbuf_2
XFILLER_0_33_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5299__A0 _1190_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__3635__B _0710_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_21_333 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_506 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_56_58 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_72_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4274__B2 cu.pc.pc_o\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4274__A1 _0340_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_72_35 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5223__A0 _1194_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_29_400 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5830_ _2610_ VGND VGND VPWR VPWR _0237_ sky130_fd_sc_hd__clkbuf_1
X_2973_ net11 VGND VGND VPWR VPWR _2712_ sky130_fd_sc_hd__inv_2
X_5761_ _2548_ _2549_ VGND VGND VPWR VPWR _2550_ sky130_fd_sc_hd__nor2_1
XANTENNA__4577__A2 _1192_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4712_ ih.t.count\[24\] ih.t.count\[25\] _1720_ ih.t.count\[26\] VGND VGND VPWR VPWR
+ _1727_ sky130_fd_sc_hd__a31o_1
XANTENNA__3098__A ih.t.timer_max\[1\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_71_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5692_ _2500_ _1643_ cu.reg_file.reg_mem\[11\] _1646_ VGND VGND VPWR VPWR _2501_
+ sky130_fd_sc_hd__a2bb2o_1
XFILLER_0_44_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_4643_ _1679_ _1680_ _1672_ VGND VGND VPWR VPWR _1681_ sky130_fd_sc_hd__and3b_1
XFILLER_0_71_266 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XANTENNA__5526__A1 net16 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_4_533 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_24_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4574_ _2702_ _1075_ _1226_ _2697_ VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__a22o_1
XFILLER_0_12_344 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3525_ _0575_ _0588_ _0600_ VGND VGND VPWR VPWR _0601_ sky130_fd_sc_hd__and3_1
X_6313_ clknet_leaf_36_clk _0006_ net158 VGND VGND VPWR VPWR cu.id.state\[2\] sky130_fd_sc_hd__dfrtp_1
XFILLER_0_24_182 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
X_6244_ clknet_leaf_36_clk _0015_ net158 VGND VGND VPWR VPWR cu.id.interrupt_requested
+ sky130_fd_sc_hd__dfrtp_1
X_3456_ _0531_ VGND VGND VPWR VPWR _0532_ sky130_fd_sc_hd__inv_2
X_6175_ clknet_leaf_19_clk _0209_ net184 VGND VGND VPWR VPWR cu.reg_file.reg_mem\[11\]
+ sky130_fd_sc_hd__dfrtp_2
X_3387_ _0336_ _0460_ _0462_ VGND VGND VPWR VPWR _0463_ sky130_fd_sc_hd__a21o_2
X_5126_ _1623_ _1050_ _2066_ VGND VGND VPWR VPWR _2071_ sky130_fd_sc_hd__mux2_1
X_5057_ _2026_ VGND VGND VPWR VPWR _0048_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_79_311 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA__5462__A0 net61 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_4008_ _0570_ _0763_ VGND VGND VPWR VPWR _1082_ sky130_fd_sc_hd__nor2_1
XFILLER_0_39_219 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_5959_ _2689_ VGND VGND VPWR VPWR _0287_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_75_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__3776__B1 _0429_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_90_531 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_35_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_7_393 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_371 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_50_439 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4740__A2 _0361_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_30_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XANTENNA__4559__A2 _1321_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_38_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_42_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_66_550 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_26_414 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_93_391 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_26_447 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_81_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XANTENNA__5337__S _2206_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_26_469 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_53_299 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_41_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_41_428 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA_4 _1188_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output93_A net93 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
X_3310_ _2877_ _2880_ VGND VGND VPWR VPWR _0386_ sky130_fd_sc_hd__nand2_2
X_4290_ _1356_ _1354_ VGND VGND VPWR VPWR _1357_ sky130_fd_sc_hd__nor2_1
XTAP_314 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_303 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_67_68 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_325 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__3381__A cu.id.starting_int_service VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3241_ _2943_ _0316_ VGND VGND VPWR VPWR _0317_ sky130_fd_sc_hd__nand2_1
XANTENNA__5692__B1 cu.reg_file.reg_mem\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3172_ cu.id.opcode\[6\] cu.id.opcode\[7\] VGND VGND VPWR VPWR _2909_ sky130_fd_sc_hd__or2_1
XTAP_369 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4196__B _1027_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_clkbuf_leaf_6_clk_A clknet_2_2__leaf_clk VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_83_67 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5444__A0 _2022_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_49_517 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4643__C _1672_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_76_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_76_347 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5747__A1 _0740_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_5813_ cu.reg_file.reg_sp\[9\] _2595_ _2539_ VGND VGND VPWR VPWR _2596_ sky130_fd_sc_hd__mux2_1
XANTENNA__3758__B1 _0741_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_2956_ _2696_ VGND VGND VPWR VPWR _2697_ sky130_fd_sc_hd__clkbuf_8
XFILLER_0_17_425 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_17_436 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
X_5744_ _2534_ VGND VGND VPWR VPWR _2535_ sky130_fd_sc_hd__clkbuf_2
X_5675_ _2487_ VGND VGND VPWR VPWR _0205_ sky130_fd_sc_hd__clkbuf_1
XFILLER_0_89_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_4626_ _1651_ _1667_ _1657_ _1351_ VGND VGND VPWR VPWR _1668_ sky130_fd_sc_hd__a31o_1
XFILLER_0_32_417 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
X_4557_ cu.pc.pc_o\[15\] _1485_ _1609_ VGND VGND VPWR VPWR _1610_ sky130_fd_sc_hd__o21a_1
X_4488_ _1305_ _1541_ _1544_ VGND VGND VPWR VPWR _1545_ sky130_fd_sc_hd__o21ai_4
X_3508_ cu.id.cb_opcode_y\[2\] _0361_ _0437_ _0341_ _0583_ VGND VGND VPWR VPWR _0584_
+ sky130_fd_sc_hd__a221o_1
X_6227_ clknet_leaf_12_clk ih.t.next_count\[15\] net177 VGND VGND VPWR VPWR ih.t.count\[15\]
+ sky130_fd_sc_hd__dfrtp_1
XANTENNA__4486__A1 cu.pc.pc_o\[11\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_3439_ _0514_ _0400_ VGND VGND VPWR VPWR _0515_ sky130_fd_sc_hd__or2b_1
X_6158_ clknet_leaf_16_clk _0192_ net181 VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__dfrtp_4
XTAP_870 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__4486__B2 cu.reg_file.reg_d\[3\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XTAP_892 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_881 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
X_5109_ cu.reg_file.reg_e\[3\] _1187_ _2056_ VGND VGND VPWR VPWR _2060_ sky130_fd_sc_hd__mux2_1
XANTENNA__5435__A0 _2022_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6089_ clknet_leaf_8_clk _0123_ net168 VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__dfrtp_4
XANTENNA__5738__A1 net25 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_82_306 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_55_509 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_48_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__3749__B1 _0741_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_380 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_63_520 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4410__B2 cu.reg_file.reg_e\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4410__A1 cu.pc.pc_o\[7\] VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__6199__D net12 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_50_236 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_16_480 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_31_472 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput41 net41 VGND VGND VPWR VPWR memory_address_out[15] sky130_fd_sc_hd__clkbuf_4
Xoutput52 net52 VGND VGND VPWR VPWR memory_data_out[1] sky130_fd_sc_hd__clkbuf_4
Xoutput85 net85 VGND VGND VPWR VPWR ss1[1] sky130_fd_sc_hd__clkbuf_4
Xoutput74 net74 VGND VGND VPWR VPWR programmable_gpio_wr[6] sky130_fd_sc_hd__buf_2
Xoutput63 net63 VGND VGND VPWR VPWR programmable_gpio_out[3] sky130_fd_sc_hd__clkbuf_4
Xoutput96 net96 VGND VGND VPWR VPWR ss2[4] sky130_fd_sc_hd__clkbuf_4
XANTENNA__5426__A0 _2022_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA_output131_A net131 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_53_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_85_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_58_369 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_39_561 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_3790_ _0865_ VGND VGND VPWR VPWR _0866_ sky130_fd_sc_hd__inv_2
XPHY_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_180 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_54_553 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_81_383 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5460_ _1369_ _2179_ VGND VGND VPWR VPWR _2287_ sky130_fd_sc_hd__nand2_1
X_4411_ cu.reg_file.reg_c\[7\] _1313_ _1469_ _1471_ VGND VGND VPWR VPWR _1472_ sky130_fd_sc_hd__a211o_1
XANTENNA__4165__B1 _0824_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_41_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_41_236 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__5901__A1 _1187_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XFILLER_0_75_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
X_5391_ _2240_ VGND VGND VPWR VPWR _0168_ sky130_fd_sc_hd__clkbuf_1
X_4342_ cu.reg_file.reg_a\[4\] _1276_ _1287_ cu.reg_file.reg_sp\[4\] VGND VGND VPWR
+ VPWR _1406_ sky130_fd_sc_hd__a22o_1
X_4273_ _1271_ _1339_ VGND VGND VPWR VPWR _1340_ sky130_fd_sc_hd__nor2_1
XFILLER_0_1_388 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XANTENNA__4468__A1 _1521_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XANTENNA__4000__A _1073_ VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
X_6012_ clknet_leaf_4_clk _0050_ net170 VGND VGND VPWR VPWR cu.reg_file.reg_c\[2\]
+ sky130_fd_sc_hd__dfrtp_2
X_3224_ _0298_ _0299_ VGND VGND VPWR VPWR _0300_ sky130_fd_sc_hd__nand2_1
.ends

