VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO Eighty_Twos
  CLASS BLOCK ;
  FOREIGN Eighty_Twos ;
  ORIGIN 0.000 0.000 ;
  SIZE 197.090 BY 207.810 ;
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 24.340 10.640 25.940 196.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 177.940 10.640 179.540 196.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 30.030 191.600 31.630 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 183.210 191.600 184.810 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 196.080 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 196.080 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 26.730 191.600 28.330 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.280 179.910 191.600 181.510 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END clk
  PIN cs
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.247500 ;
    PORT
      LAYER met3 ;
        RECT 193.090 44.240 197.090 44.840 ;
    END
  END cs
  PIN gpi[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END gpi[0]
  PIN gpi[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 193.090 146.240 197.090 146.840 ;
    END
  END gpi[10]
  PIN gpi[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END gpi[11]
  PIN gpi[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 193.090 68.040 197.090 68.640 ;
    END
  END gpi[12]
  PIN gpi[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 203.810 10.030 207.810 ;
    END
  END gpi[13]
  PIN gpi[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 0.000 142.050 4.000 ;
    END
  END gpi[14]
  PIN gpi[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 193.090 125.840 197.090 126.440 ;
    END
  END gpi[15]
  PIN gpi[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 115.640 4.000 116.240 ;
    END
  END gpi[16]
  PIN gpi[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 193.090 20.440 197.090 21.040 ;
    END
  END gpi[17]
  PIN gpi[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END gpi[18]
  PIN gpi[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 119.230 0.000 119.510 4.000 ;
    END
  END gpi[19]
  PIN gpi[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END gpi[1]
  PIN gpi[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END gpi[20]
  PIN gpi[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 193.090 30.640 197.090 31.240 ;
    END
  END gpi[21]
  PIN gpi[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END gpi[22]
  PIN gpi[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 154.650 203.810 154.930 207.810 ;
    END
  END gpi[23]
  PIN gpi[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 141.770 203.810 142.050 207.810 ;
    END
  END gpi[24]
  PIN gpi[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 149.640 4.000 150.240 ;
    END
  END gpi[25]
  PIN gpi[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 193.090 136.040 197.090 136.640 ;
    END
  END gpi[26]
  PIN gpi[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 193.090 159.840 197.090 160.440 ;
    END
  END gpi[27]
  PIN gpi[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 173.440 4.000 174.040 ;
    END
  END gpi[28]
  PIN gpi[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 0.000 109.850 4.000 ;
    END
  END gpi[29]
  PIN gpi[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END gpi[2]
  PIN gpi[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 197.240 4.000 197.840 ;
    END
  END gpi[30]
  PIN gpi[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END gpi[31]
  PIN gpi[32]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 203.810 122.730 207.810 ;
    END
  END gpi[32]
  PIN gpi[33]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 203.810 32.570 207.810 ;
    END
  END gpi[33]
  PIN gpi[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.196500 ;
    PORT
      LAYER met2 ;
        RECT 41.950 0.000 42.230 4.000 ;
    END
  END gpi[3]
  PIN gpi[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met2 ;
        RECT 77.370 203.810 77.650 207.810 ;
    END
  END gpi[4]
  PIN gpi[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 186.850 203.810 187.130 207.810 ;
    END
  END gpi[5]
  PIN gpi[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.159000 ;
    PORT
      LAYER met2 ;
        RECT 186.850 0.000 187.130 4.000 ;
    END
  END gpi[6]
  PIN gpi[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.126000 ;
    PORT
      LAYER met2 ;
        RECT 99.910 203.810 100.190 207.810 ;
    END
  END gpi[7]
  PIN gpi[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 203.810 196.790 207.810 ;
    END
  END gpi[8]
  PIN gpi[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 164.310 0.000 164.590 4.000 ;
    END
  END gpi[9]
  PIN gpo[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 87.030 203.810 87.310 207.810 ;
    END
  END gpo[0]
  PIN gpo[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 20.440 4.000 21.040 ;
    END
  END gpo[10]
  PIN gpo[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 193.090 54.440 197.090 55.040 ;
    END
  END gpo[11]
  PIN gpo[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.240 4.000 44.840 ;
    END
  END gpo[12]
  PIN gpo[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 193.090 78.240 197.090 78.840 ;
    END
  END gpo[13]
  PIN gpo[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 0.090 203.810 0.370 207.810 ;
    END
  END gpo[14]
  PIN gpo[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 132.110 203.810 132.390 207.810 ;
    END
  END gpo[15]
  PIN gpo[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END gpo[16]
  PIN gpo[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END gpo[17]
  PIN gpo[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 125.840 4.000 126.440 ;
    END
  END gpo[18]
  PIN gpo[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 109.570 203.810 109.850 207.810 ;
    END
  END gpo[19]
  PIN gpo[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 78.240 4.000 78.840 ;
    END
  END gpo[1]
  PIN gpo[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 193.090 193.840 197.090 194.440 ;
    END
  END gpo[20]
  PIN gpo[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 64.490 203.810 64.770 207.810 ;
    END
  END gpo[21]
  PIN gpo[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END gpo[22]
  PIN gpo[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END gpo[23]
  PIN gpo[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 193.090 183.640 197.090 184.240 ;
    END
  END gpo[24]
  PIN gpo[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.840 4.000 92.440 ;
    END
  END gpo[25]
  PIN gpo[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 74.150 0.000 74.430 4.000 ;
    END
  END gpo[26]
  PIN gpo[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 193.090 170.040 197.090 170.640 ;
    END
  END gpo[27]
  PIN gpo[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 193.090 6.840 197.090 7.440 ;
    END
  END gpo[28]
  PIN gpo[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 45.170 203.810 45.450 207.810 ;
    END
  END gpo[29]
  PIN gpo[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 193.090 102.040 197.090 102.640 ;
    END
  END gpo[2]
  PIN gpo[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END gpo[30]
  PIN gpo[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 64.490 0.000 64.770 4.000 ;
    END
  END gpo[31]
  PIN gpo[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END gpo[32]
  PIN gpo[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met3 ;
        RECT 193.090 112.240 197.090 112.840 ;
    END
  END gpo[33]
  PIN gpo[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 96.690 0.000 96.970 4.000 ;
    END
  END gpo[3]
  PIN gpo[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 177.190 203.810 177.470 207.810 ;
    END
  END gpo[4]
  PIN gpo[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 164.310 203.810 164.590 207.810 ;
    END
  END gpo[5]
  PIN gpo[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.445500 ;
    PORT
      LAYER met2 ;
        RECT 22.630 203.810 22.910 207.810 ;
    END
  END gpo[6]
  PIN gpo[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 54.830 203.810 55.110 207.810 ;
    END
  END gpo[7]
  PIN gpo[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met2 ;
        RECT 132.110 0.000 132.390 4.000 ;
    END
  END gpo[8]
  PIN gpo[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 0.000 68.040 4.000 68.640 ;
    END
  END gpo[9]
  PIN nrst
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213000 ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END nrst
  PIN store_en
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.795200 ;
    PORT
      LAYER met3 ;
        RECT 193.090 88.440 197.090 89.040 ;
    END
  END store_en
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 191.360 195.925 ;
      LAYER met1 ;
        RECT 0.070 10.640 192.210 196.080 ;
      LAYER met2 ;
        RECT 0.650 203.530 9.470 204.410 ;
        RECT 10.310 203.530 22.350 204.410 ;
        RECT 23.190 203.530 32.010 204.410 ;
        RECT 32.850 203.530 44.890 204.410 ;
        RECT 45.730 203.530 54.550 204.410 ;
        RECT 55.390 203.530 64.210 204.410 ;
        RECT 65.050 203.530 77.090 204.410 ;
        RECT 77.930 203.530 86.750 204.410 ;
        RECT 87.590 203.530 99.630 204.410 ;
        RECT 100.470 203.530 109.290 204.410 ;
        RECT 110.130 203.530 122.170 204.410 ;
        RECT 123.010 203.530 131.830 204.410 ;
        RECT 132.670 203.530 141.490 204.410 ;
        RECT 142.330 203.530 154.370 204.410 ;
        RECT 155.210 203.530 164.030 204.410 ;
        RECT 164.870 203.530 176.910 204.410 ;
        RECT 177.750 203.530 186.570 204.410 ;
        RECT 187.410 203.530 192.190 204.410 ;
        RECT 0.100 4.280 192.190 203.530 ;
        RECT 0.650 4.000 9.470 4.280 ;
        RECT 10.310 4.000 19.130 4.280 ;
        RECT 19.970 4.000 32.010 4.280 ;
        RECT 32.850 4.000 41.670 4.280 ;
        RECT 42.510 4.000 54.550 4.280 ;
        RECT 55.390 4.000 64.210 4.280 ;
        RECT 65.050 4.000 73.870 4.280 ;
        RECT 74.710 4.000 86.750 4.280 ;
        RECT 87.590 4.000 96.410 4.280 ;
        RECT 97.250 4.000 109.290 4.280 ;
        RECT 110.130 4.000 118.950 4.280 ;
        RECT 119.790 4.000 131.830 4.280 ;
        RECT 132.670 4.000 141.490 4.280 ;
        RECT 142.330 4.000 151.150 4.280 ;
        RECT 151.990 4.000 164.030 4.280 ;
        RECT 164.870 4.000 173.690 4.280 ;
        RECT 174.530 4.000 186.570 4.280 ;
        RECT 187.410 4.000 192.190 4.280 ;
      LAYER met3 ;
        RECT 3.990 194.840 193.090 196.005 ;
        RECT 3.990 193.440 192.690 194.840 ;
        RECT 3.990 184.640 193.090 193.440 ;
        RECT 4.400 183.240 192.690 184.640 ;
        RECT 3.990 174.440 193.090 183.240 ;
        RECT 4.400 173.040 193.090 174.440 ;
        RECT 3.990 171.040 193.090 173.040 ;
        RECT 3.990 169.640 192.690 171.040 ;
        RECT 3.990 160.840 193.090 169.640 ;
        RECT 4.400 159.440 192.690 160.840 ;
        RECT 3.990 150.640 193.090 159.440 ;
        RECT 4.400 149.240 193.090 150.640 ;
        RECT 3.990 147.240 193.090 149.240 ;
        RECT 3.990 145.840 192.690 147.240 ;
        RECT 3.990 137.040 193.090 145.840 ;
        RECT 4.400 135.640 192.690 137.040 ;
        RECT 3.990 126.840 193.090 135.640 ;
        RECT 4.400 125.440 192.690 126.840 ;
        RECT 3.990 116.640 193.090 125.440 ;
        RECT 4.400 115.240 193.090 116.640 ;
        RECT 3.990 113.240 193.090 115.240 ;
        RECT 3.990 111.840 192.690 113.240 ;
        RECT 3.990 103.040 193.090 111.840 ;
        RECT 4.400 101.640 192.690 103.040 ;
        RECT 3.990 92.840 193.090 101.640 ;
        RECT 4.400 91.440 193.090 92.840 ;
        RECT 3.990 89.440 193.090 91.440 ;
        RECT 3.990 88.040 192.690 89.440 ;
        RECT 3.990 79.240 193.090 88.040 ;
        RECT 4.400 77.840 192.690 79.240 ;
        RECT 3.990 69.040 193.090 77.840 ;
        RECT 4.400 67.640 192.690 69.040 ;
        RECT 3.990 58.840 193.090 67.640 ;
        RECT 4.400 57.440 193.090 58.840 ;
        RECT 3.990 55.440 193.090 57.440 ;
        RECT 3.990 54.040 192.690 55.440 ;
        RECT 3.990 45.240 193.090 54.040 ;
        RECT 4.400 43.840 192.690 45.240 ;
        RECT 3.990 35.040 193.090 43.840 ;
        RECT 4.400 33.640 193.090 35.040 ;
        RECT 3.990 31.640 193.090 33.640 ;
        RECT 3.990 30.240 192.690 31.640 ;
        RECT 3.990 21.440 193.090 30.240 ;
        RECT 4.400 20.040 192.690 21.440 ;
        RECT 3.990 11.240 193.090 20.040 ;
        RECT 4.400 9.840 193.090 11.240 ;
        RECT 3.990 7.840 193.090 9.840 ;
        RECT 3.990 6.975 192.690 7.840 ;
      LAYER met4 ;
        RECT 48.135 19.895 145.065 194.305 ;
  END
END Eighty_Twos
END LIBRARY

